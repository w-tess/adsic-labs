**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [26 16 160] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_14_PCB_wire_2p0inch_highloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 -1.3077575657901009e-02
GC_1_2 b_1 NI_1 NS_2 0 1.3851810838323535e-03
GC_1_3 b_1 NI_1 NS_3 0 -2.6206809722674823e-07
GC_1_4 b_1 NI_1 NS_4 0 -3.7495376870490346e-06
GC_1_5 b_1 NI_1 NS_5 0 -2.7819412649520358e-04
GC_1_6 b_1 NI_1 NS_6 0 4.6297784662633300e-04
GC_1_7 b_1 NI_1 NS_7 0 1.3195316947854435e-03
GC_1_8 b_1 NI_1 NS_8 0 5.4935810838291593e-04
GC_1_9 b_1 NI_1 NS_9 0 -2.7628707830369883e-03
GC_1_10 b_1 NI_1 NS_10 0 -8.1702960577214928e-04
GC_1_11 b_1 NI_1 NS_11 0 3.5326194217735240e-03
GC_1_12 b_1 NI_1 NS_12 0 2.5338003494739768e-03
GC_1_13 b_1 NI_1 NS_13 0 1.1824215167209342e-03
GC_1_14 b_1 NI_1 NS_14 0 -4.1997919360091483e-03
GC_1_15 b_1 NI_1 NS_15 0 -1.7498497484580156e-03
GC_1_16 b_1 NI_1 NS_16 0 2.6968875331490551e-03
GC_1_17 b_1 NI_1 NS_17 0 -3.1387253129775311e-04
GC_1_18 b_1 NI_1 NS_18 0 -1.8984355421804193e-04
GC_1_19 b_1 NI_1 NS_19 0 3.9674908773077461e-03
GC_1_20 b_1 NI_1 NS_20 0 2.9857924899115109e-04
GC_1_21 b_1 NI_1 NS_21 0 -7.4413898752019921e-03
GC_1_22 b_1 NI_1 NS_22 0 -1.3618331607426655e-02
GC_1_23 b_1 NI_1 NS_23 0 4.4052529700013528e-03
GC_1_24 b_1 NI_1 NS_24 0 1.3511450566459538e-02
GC_1_25 b_1 NI_1 NS_25 0 6.7110134907060288e-03
GC_1_26 b_1 NI_1 NS_26 0 -3.9862641894755184e-03
GC_1_27 b_1 NI_1 NS_27 0 -1.3390053159841231e-02
GC_1_28 b_1 NI_1 NS_28 0 6.9023312149961967e-04
GC_1_29 b_1 NI_1 NS_29 0 7.8426027215748491e-03
GC_1_30 b_1 NI_1 NS_30 0 1.8947657846528946e-03
GC_1_31 b_1 NI_1 NS_31 0 1.0544114974705733e-02
GC_1_32 b_1 NI_1 NS_32 0 -1.9595452275828550e-02
GC_1_33 b_1 NI_1 NS_33 0 -1.7809618055612247e-02
GC_1_34 b_1 NI_1 NS_34 0 1.9141982754547052e-02
GC_1_35 b_1 NI_1 NS_35 0 7.6787743766726299e-03
GC_1_36 b_1 NI_1 NS_36 0 -1.4142911445394878e-03
GC_1_37 b_1 NI_1 NS_37 0 -1.5647917037334789e-02
GC_1_38 b_1 NI_1 NS_38 0 -4.7614903566561839e-03
GC_1_39 b_1 NI_1 NS_39 0 8.0618568963727790e-03
GC_1_40 b_1 NI_1 NS_40 0 7.2869895044589588e-03
GC_1_41 b_1 NI_1 NS_41 0 8.1170040783415231e-03
GC_1_42 b_1 NI_1 NS_42 0 -5.9990842974454173e-03
GC_1_43 b_1 NI_1 NS_43 0 -1.3980589235184478e-02
GC_1_44 b_1 NI_1 NS_44 0 4.5682738336424028e-03
GC_1_45 b_1 NI_1 NS_45 0 6.2307821482152246e-03
GC_1_46 b_1 NI_1 NS_46 0 2.4081616521146897e-03
GC_1_47 b_1 NI_1 NS_47 0 -6.2859259532728950e-03
GC_1_48 b_1 NI_1 NS_48 0 -1.1107051215958732e-02
GC_1_49 b_1 NI_1 NS_49 0 2.1280730654035310e-03
GC_1_50 b_1 NI_1 NS_50 0 1.1947396614296972e-02
GC_1_51 b_1 NI_1 NS_51 0 4.2092181380885456e-03
GC_1_52 b_1 NI_1 NS_52 0 -1.1609525185983017e-03
GC_1_53 b_1 NI_1 NS_53 0 -4.9313047700377541e-03
GC_1_54 b_1 NI_1 NS_54 0 1.0532426449717895e-03
GC_1_55 b_1 NI_1 NS_55 0 3.0238805602791304e-03
GC_1_56 b_1 NI_1 NS_56 0 6.9985668908831983e-04
GC_1_57 b_1 NI_1 NS_57 0 -2.2205265102976553e-03
GC_1_58 b_1 NI_1 NS_58 0 4.9428523590553297e-04
GC_1_59 b_1 NI_1 NS_59 0 3.0655101856454977e-03
GC_1_60 b_1 NI_1 NS_60 0 2.3037295682999523e-03
GC_1_61 b_1 NI_1 NS_61 0 -1.5339095928932412e-03
GC_1_62 b_1 NI_1 NS_62 0 -6.6977523797265954e-04
GC_1_63 b_1 NI_1 NS_63 0 1.8873377871796466e-03
GC_1_64 b_1 NI_1 NS_64 0 6.8441611640669437e-04
GC_1_65 b_1 NI_1 NS_65 0 -1.5620994940070121e-03
GC_1_66 b_1 NI_1 NS_66 0 1.2263485505595833e-03
GC_1_67 b_1 NI_1 NS_67 0 3.9751899193916440e-03
GC_1_68 b_1 NI_1 NS_68 0 1.4060873640009222e-03
GC_1_69 b_1 NI_1 NS_69 0 -1.5528113430304227e-03
GC_1_70 b_1 NI_1 NS_70 0 7.4659511700874819e-05
GC_1_71 b_1 NI_1 NS_71 0 2.8290376322292333e-03
GC_1_72 b_1 NI_1 NS_72 0 -6.8617020675090182e-04
GC_1_73 b_1 NI_1 NS_73 0 -1.8781842572438718e-03
GC_1_74 b_1 NI_1 NS_74 0 2.0100714537211613e-03
GC_1_75 b_1 NI_1 NS_75 0 4.9079326878394038e-03
GC_1_76 b_1 NI_1 NS_76 0 -1.8215468359406971e-04
GC_1_77 b_1 NI_1 NS_77 0 -1.6564605115434354e-03
GC_1_78 b_1 NI_1 NS_78 0 9.3019010342196620e-04
GC_1_79 b_1 NI_1 NS_79 0 3.0643001553695101e-03
GC_1_80 b_1 NI_1 NS_80 0 -2.8465122061003948e-03
GC_1_81 b_1 NI_1 NS_81 0 -1.4568575903714243e-03
GC_1_82 b_1 NI_1 NS_82 0 3.2233585197213922e-03
GC_1_83 b_1 NI_1 NS_83 0 3.8009943564278437e-03
GC_1_84 b_1 NI_1 NS_84 0 -2.9784231906301497e-03
GC_1_85 b_1 NI_1 NS_85 0 -1.8786945472106229e-03
GC_1_86 b_1 NI_1 NS_86 0 -3.8879223983061492e-03
GC_1_87 b_1 NI_1 NS_87 0 -4.0380170454161907e-04
GC_1_88 b_1 NI_1 NS_88 0 2.3675226288496134e-03
GC_1_89 b_1 NI_1 NS_89 0 -1.0556794297925798e-05
GC_1_90 b_1 NI_1 NS_90 0 -2.1452512941284554e-05
GC_1_91 b_1 NI_1 NS_91 0 8.4229612476062325e-04
GC_1_92 b_1 NI_1 NS_92 0 -3.7965172925199099e-03
GC_1_93 b_1 NI_1 NS_93 0 3.4279131023536144e-04
GC_1_94 b_1 NI_1 NS_94 0 3.3487732415310350e-03
GC_1_95 b_1 NI_1 NS_95 0 1.3577072327638348e-03
GC_1_96 b_1 NI_1 NS_96 0 -2.3752473045804577e-03
GC_1_97 b_1 NI_1 NS_97 0 2.1858950999851176e-03
GC_1_98 b_1 NI_1 NS_98 0 3.3360403257720718e-03
GC_1_99 b_1 NI_1 NS_99 0 1.1689683902370773e-03
GC_1_100 b_1 NI_1 NS_100 0 2.4033203960212926e-03
GC_1_101 b_1 NI_1 NS_101 0 -8.1092242504170577e-04
GC_1_102 b_1 NI_1 NS_102 0 -1.9781509790563197e-03
GC_1_103 b_1 NI_1 NS_103 0 3.9749449703226731e-04
GC_1_104 b_1 NI_1 NS_104 0 -2.6833646704893972e-03
GC_1_105 b_1 NI_1 NS_105 0 9.8234519887786787e-04
GC_1_106 b_1 NI_1 NS_106 0 2.7459694004676187e-03
GC_1_107 b_1 NI_1 NS_107 0 1.0390528567683220e-03
GC_1_108 b_1 NI_1 NS_108 0 -2.4207680352576542e-03
GC_1_109 b_1 NI_1 NS_109 0 -1.0837521621894820e-03
GC_1_110 b_1 NI_1 NS_110 0 1.5920956224601483e-03
GC_1_111 b_1 NI_1 NS_111 0 -1.1067857241654118e-08
GC_1_112 b_1 NI_1 NS_112 0 -2.8131625101367103e-09
GC_1_113 b_1 NI_1 NS_113 0 2.2673375171328769e-06
GC_1_114 b_1 NI_1 NS_114 0 5.3151463752614834e-07
GC_1_115 b_1 NI_1 NS_115 0 1.8229768971867504e-02
GC_1_116 b_1 NI_1 NS_116 0 6.7517747779893599e-03
GC_1_117 b_1 NI_1 NS_117 0 4.8176237406255103e-07
GC_1_118 b_1 NI_1 NS_118 0 1.4329614168124728e-06
GC_1_119 b_1 NI_1 NS_119 0 6.0824999945254567e-03
GC_1_120 b_1 NI_1 NS_120 0 1.8254880323254384e-03
GC_1_121 b_1 NI_1 NS_121 0 -6.0663216004818426e-03
GC_1_122 b_1 NI_1 NS_122 0 -6.4127997028286623e-04
GC_1_123 b_1 NI_1 NS_123 0 7.3353149342791132e-03
GC_1_124 b_1 NI_1 NS_124 0 -1.2858414056027881e-02
GC_1_125 b_1 NI_1 NS_125 0 8.4354710028741661e-03
GC_1_126 b_1 NI_1 NS_126 0 -2.1165010913373427e-04
GC_1_127 b_1 NI_1 NS_127 0 -9.6680547443697556e-03
GC_1_128 b_1 NI_1 NS_128 0 2.5853966643882521e-03
GC_1_129 b_1 NI_1 NS_129 0 -8.8080249442280528e-03
GC_1_130 b_1 NI_1 NS_130 0 -2.4394897882313686e-02
GC_1_131 b_1 NI_1 NS_131 0 -8.6848124533620106e-04
GC_1_132 b_1 NI_1 NS_132 0 4.1758872051821262e-03
GC_1_133 b_1 NI_1 NS_133 0 7.1854582274890168e-03
GC_1_134 b_1 NI_1 NS_134 0 -9.9750178948579122e-04
GC_1_135 b_1 NI_1 NS_135 0 -2.5219943873861370e-02
GC_1_136 b_1 NI_1 NS_136 0 4.8141538601170946e-03
GC_1_137 b_1 NI_1 NS_137 0 -1.9618485114991212e-02
GC_1_138 b_1 NI_1 NS_138 0 8.5369576203501074e-04
GC_1_139 b_1 NI_1 NS_139 0 1.0773090203853511e-02
GC_1_140 b_1 NI_1 NS_140 0 -2.7350692474235059e-03
GC_1_141 b_1 NI_1 NS_141 0 -4.8270291391232191e-03
GC_1_142 b_1 NI_1 NS_142 0 4.5019523413195837e-02
GC_1_143 b_1 NI_1 NS_143 0 -1.2641866833814196e-02
GC_1_144 b_1 NI_1 NS_144 0 -3.2184671887946923e-04
GC_1_145 b_1 NI_1 NS_145 0 1.5975293983663728e-02
GC_1_146 b_1 NI_1 NS_146 0 -3.9759266204381317e-03
GC_1_147 b_1 NI_1 NS_147 0 3.2145903249934778e-02
GC_1_148 b_1 NI_1 NS_148 0 1.8555230541492759e-02
GC_1_149 b_1 NI_1 NS_149 0 -1.2594982553996055e-02
GC_1_150 b_1 NI_1 NS_150 0 1.1569141782556884e-04
GC_1_151 b_1 NI_1 NS_151 0 1.7251925944377657e-02
GC_1_152 b_1 NI_1 NS_152 0 -3.5175897355458369e-02
GC_1_153 b_1 NI_1 NS_153 0 1.3984016088098796e-02
GC_1_154 b_1 NI_1 NS_154 0 4.8235365206254167e-03
GC_1_155 b_1 NI_1 NS_155 0 -1.4410945404248027e-02
GC_1_156 b_1 NI_1 NS_156 0 1.9244703412420953e-04
GC_1_157 b_1 NI_1 NS_157 0 -2.0124185788695650e-02
GC_1_158 b_1 NI_1 NS_158 0 -3.0196941856939684e-02
GC_1_159 b_1 NI_1 NS_159 0 1.0516052223712267e-02
GC_1_160 b_1 NI_1 NS_160 0 3.6210369250344078e-03
GC_1_161 b_1 NI_1 NS_161 0 -2.6839334853586368e-02
GC_1_162 b_1 NI_1 NS_162 0 1.1127464824650563e-02
GC_1_163 b_1 NI_1 NS_163 0 -1.4106856955881358e-02
GC_1_164 b_1 NI_1 NS_164 0 -2.5292733643898220e-03
GC_1_165 b_1 NI_1 NS_165 0 7.5511384056998112e-03
GC_1_166 b_1 NI_1 NS_166 0 1.6110670303257110e-03
GC_1_167 b_1 NI_1 NS_167 0 -8.7782798416482534e-04
GC_1_168 b_1 NI_1 NS_168 0 2.4406473856554225e-02
GC_1_169 b_1 NI_1 NS_169 0 -7.6159538818854700e-03
GC_1_170 b_1 NI_1 NS_170 0 2.7280778895468388e-04
GC_1_171 b_1 NI_1 NS_171 0 -5.5398018609179478e-04
GC_1_172 b_1 NI_1 NS_172 0 -5.5347552424719285e-03
GC_1_173 b_1 NI_1 NS_173 0 8.2549295156051430e-03
GC_1_174 b_1 NI_1 NS_174 0 7.0291658244709954e-03
GC_1_175 b_1 NI_1 NS_175 0 -7.2657828553996566e-04
GC_1_176 b_1 NI_1 NS_176 0 1.2096249880014608e-02
GC_1_177 b_1 NI_1 NS_177 0 -5.1449933010362511e-03
GC_1_178 b_1 NI_1 NS_178 0 -1.3736740083024836e-04
GC_1_179 b_1 NI_1 NS_179 0 -1.8277917732876198e-03
GC_1_180 b_1 NI_1 NS_180 0 -5.1663778979150433e-03
GC_1_181 b_1 NI_1 NS_181 0 9.2806004053513236e-03
GC_1_182 b_1 NI_1 NS_182 0 5.4201888408802312e-03
GC_1_183 b_1 NI_1 NS_183 0 3.5139970262974187e-03
GC_1_184 b_1 NI_1 NS_184 0 1.1696927542125219e-02
GC_1_185 b_1 NI_1 NS_185 0 -6.1352204731379822e-03
GC_1_186 b_1 NI_1 NS_186 0 1.4322934935951789e-03
GC_1_187 b_1 NI_1 NS_187 0 -2.8179422592280799e-03
GC_1_188 b_1 NI_1 NS_188 0 -7.3386927850469762e-03
GC_1_189 b_1 NI_1 NS_189 0 9.9491567342893401e-03
GC_1_190 b_1 NI_1 NS_190 0 3.3701752947640738e-03
GC_1_191 b_1 NI_1 NS_191 0 8.1727436024223044e-03
GC_1_192 b_1 NI_1 NS_192 0 1.0256343564889170e-02
GC_1_193 b_1 NI_1 NS_193 0 -6.9843105263184737e-03
GC_1_194 b_1 NI_1 NS_194 0 2.9455097438636558e-03
GC_1_195 b_1 NI_1 NS_195 0 -5.6339149178409494e-03
GC_1_196 b_1 NI_1 NS_196 0 -8.0804968512090750e-03
GC_1_197 b_1 NI_1 NS_197 0 9.8431594290583572e-03
GC_1_198 b_1 NI_1 NS_198 0 5.5952313827845469e-04
GC_1_199 b_1 NI_1 NS_199 0 -1.0789843398086163e-02
GC_1_200 b_1 NI_1 NS_200 0 1.2190784534326305e-02
GC_1_201 b_1 NI_1 NS_201 0 9.6746160643738470e-03
GC_1_202 b_1 NI_1 NS_202 0 5.0623913848552912e-03
GC_1_203 b_1 NI_1 NS_203 0 -1.9022005986450378e-05
GC_1_204 b_1 NI_1 NS_204 0 3.1756644648914916e-05
GC_1_205 b_1 NI_1 NS_205 0 -7.1157907395909608e-03
GC_1_206 b_1 NI_1 NS_206 0 4.4965754708824780e-03
GC_1_207 b_1 NI_1 NS_207 0 -7.6591575737087105e-03
GC_1_208 b_1 NI_1 NS_208 0 -5.3141664589059579e-03
GC_1_209 b_1 NI_1 NS_209 0 9.4991951729312511e-03
GC_1_210 b_1 NI_1 NS_210 0 -1.7114737154242047e-03
GC_1_211 b_1 NI_1 NS_211 0 1.2463031433085886e-02
GC_1_212 b_1 NI_1 NS_212 0 -1.3561705396320832e-03
GC_1_213 b_1 NI_1 NS_213 0 -5.0733887030775717e-03
GC_1_214 b_1 NI_1 NS_214 0 -2.7549337256449640e-03
GC_1_215 b_1 NI_1 NS_215 0 -2.2333207468812765e-03
GC_1_216 b_1 NI_1 NS_216 0 6.5928668697620351e-03
GC_1_217 b_1 NI_1 NS_217 0 8.9636625837498565e-03
GC_1_218 b_1 NI_1 NS_218 0 1.2895545396009276e-04
GC_1_219 b_1 NI_1 NS_219 0 1.2489930355578899e-02
GC_1_220 b_1 NI_1 NS_220 0 1.7708869693264513e-03
GC_1_221 b_1 NI_1 NS_221 0 -5.3741342131808697e-03
GC_1_222 b_1 NI_1 NS_222 0 4.1561547985190144e-03
GC_1_223 b_1 NI_1 NS_223 0 -1.8427481189287522e-03
GC_1_224 b_1 NI_1 NS_224 0 -5.6872752486660854e-03
GC_1_225 b_1 NI_1 NS_225 0 2.0875930792225757e-07
GC_1_226 b_1 NI_1 NS_226 0 -2.4399571741935520e-07
GC_1_227 b_1 NI_1 NS_227 0 -1.1437014872363319e-05
GC_1_228 b_1 NI_1 NS_228 0 1.8295056856632399e-05
GC_1_229 b_1 NI_1 NS_229 0 7.7623631688390335e-03
GC_1_230 b_1 NI_1 NS_230 0 -1.6012429819179362e-03
GC_1_231 b_1 NI_1 NS_231 0 -1.2109163074623930e-08
GC_1_232 b_1 NI_1 NS_232 0 -8.8417590504038885e-07
GC_1_233 b_1 NI_1 NS_233 0 1.0417924324583035e-04
GC_1_234 b_1 NI_1 NS_234 0 -5.1170037850179048e-04
GC_1_235 b_1 NI_1 NS_235 0 -1.9362887985344141e-03
GC_1_236 b_1 NI_1 NS_236 0 -5.9765172108607869e-04
GC_1_237 b_1 NI_1 NS_237 0 2.9418128645628651e-03
GC_1_238 b_1 NI_1 NS_238 0 2.2635993047207740e-03
GC_1_239 b_1 NI_1 NS_239 0 -3.5704327589455988e-03
GC_1_240 b_1 NI_1 NS_240 0 -3.0490673763287723e-03
GC_1_241 b_1 NI_1 NS_241 0 -1.7073725775933386e-03
GC_1_242 b_1 NI_1 NS_242 0 5.8427846669151491e-03
GC_1_243 b_1 NI_1 NS_243 0 4.3666970100778874e-03
GC_1_244 b_1 NI_1 NS_244 0 -2.4750965249272935e-03
GC_1_245 b_1 NI_1 NS_245 0 -1.1000888430814992e-04
GC_1_246 b_1 NI_1 NS_246 0 -1.0334512903076414e-04
GC_1_247 b_1 NI_1 NS_247 0 -4.4523052984915398e-03
GC_1_248 b_1 NI_1 NS_248 0 -9.2440307396499523e-04
GC_1_249 b_1 NI_1 NS_249 0 9.1241543833800072e-03
GC_1_250 b_1 NI_1 NS_250 0 1.7784746375459161e-02
GC_1_251 b_1 NI_1 NS_251 0 -4.0272971001455160e-03
GC_1_252 b_1 NI_1 NS_252 0 -1.7846771806168733e-02
GC_1_253 b_1 NI_1 NS_253 0 -8.2177715191523674e-03
GC_1_254 b_1 NI_1 NS_254 0 4.1736008749562710e-03
GC_1_255 b_1 NI_1 NS_255 0 1.7063484687004131e-02
GC_1_256 b_1 NI_1 NS_256 0 -4.3909977322205846e-04
GC_1_257 b_1 NI_1 NS_257 0 -9.2787160081823604e-03
GC_1_258 b_1 NI_1 NS_258 0 -3.2069945516728523e-03
GC_1_259 b_1 NI_1 NS_259 0 -1.3713361965228434e-02
GC_1_260 b_1 NI_1 NS_260 0 2.2836239953980878e-02
GC_1_261 b_1 NI_1 NS_261 0 2.2839552393961387e-02
GC_1_262 b_1 NI_1 NS_262 0 -2.2669171312948658e-02
GC_1_263 b_1 NI_1 NS_263 0 -9.2392853314757009e-03
GC_1_264 b_1 NI_1 NS_264 0 9.0811376155357714e-04
GC_1_265 b_1 NI_1 NS_265 0 1.8480132532803027e-02
GC_1_266 b_1 NI_1 NS_266 0 6.2442241030503587e-03
GC_1_267 b_1 NI_1 NS_267 0 -9.1760808825051936e-03
GC_1_268 b_1 NI_1 NS_268 0 -9.4609794905343974e-03
GC_1_269 b_1 NI_1 NS_269 0 -9.9743264482213233e-03
GC_1_270 b_1 NI_1 NS_270 0 6.3961885386635232e-03
GC_1_271 b_1 NI_1 NS_271 0 1.6838481102741960e-02
GC_1_272 b_1 NI_1 NS_272 0 -4.8501205084066678e-03
GC_1_273 b_1 NI_1 NS_273 0 -7.2149225369889970e-03
GC_1_274 b_1 NI_1 NS_274 0 -3.4092354578978581e-03
GC_1_275 b_1 NI_1 NS_275 0 6.8281954719585725e-03
GC_1_276 b_1 NI_1 NS_276 0 1.3297053324820403e-02
GC_1_277 b_1 NI_1 NS_277 0 -1.8195824534275376e-03
GC_1_278 b_1 NI_1 NS_278 0 -1.4401720113390958e-02
GC_1_279 b_1 NI_1 NS_279 0 -4.9860069971232350e-03
GC_1_280 b_1 NI_1 NS_280 0 1.0394629019308838e-03
GC_1_281 b_1 NI_1 NS_281 0 6.0026097697297269e-03
GC_1_282 b_1 NI_1 NS_282 0 -1.1030574878201705e-03
GC_1_283 b_1 NI_1 NS_283 0 -3.4642734364388871e-03
GC_1_284 b_1 NI_1 NS_284 0 -1.0876297929212997e-03
GC_1_285 b_1 NI_1 NS_285 0 2.7180517521761057e-03
GC_1_286 b_1 NI_1 NS_286 0 -5.0782105589906596e-04
GC_1_287 b_1 NI_1 NS_287 0 -3.2964856509136663e-03
GC_1_288 b_1 NI_1 NS_288 0 -2.8951315922092122e-03
GC_1_289 b_1 NI_1 NS_289 0 2.0159621881281299e-03
GC_1_290 b_1 NI_1 NS_290 0 7.7577849499497304e-04
GC_1_291 b_1 NI_1 NS_291 0 -2.0162760630027293e-03
GC_1_292 b_1 NI_1 NS_292 0 -9.6646512749078411e-04
GC_1_293 b_1 NI_1 NS_293 0 2.1216220343160054e-03
GC_1_294 b_1 NI_1 NS_294 0 -1.4709118335084631e-03
GC_1_295 b_1 NI_1 NS_295 0 -4.1847944562909073e-03
GC_1_296 b_1 NI_1 NS_296 0 -1.8129441562875206e-03
GC_1_297 b_1 NI_1 NS_297 0 2.3697817652576854e-03
GC_1_298 b_1 NI_1 NS_298 0 -3.7075719352222894e-04
GC_1_299 b_1 NI_1 NS_299 0 -3.0172215283848949e-03
GC_1_300 b_1 NI_1 NS_300 0 4.6233692493955180e-04
GC_1_301 b_1 NI_1 NS_301 0 2.7064446320338620e-03
GC_1_302 b_1 NI_1 NS_302 0 -2.7282256796825862e-03
GC_1_303 b_1 NI_1 NS_303 0 -5.0393282341897163e-03
GC_1_304 b_1 NI_1 NS_304 0 -1.2783040351664764e-04
GC_1_305 b_1 NI_1 NS_305 0 2.4346778108484020e-03
GC_1_306 b_1 NI_1 NS_306 0 -2.1719821015994140e-03
GC_1_307 b_1 NI_1 NS_307 0 -3.2449804044284189e-03
GC_1_308 b_1 NI_1 NS_308 0 2.6005310513265993e-03
GC_1_309 b_1 NI_1 NS_309 0 1.7436680446217688e-03
GC_1_310 b_1 NI_1 NS_310 0 -4.7503555602780865e-03
GC_1_311 b_1 NI_1 NS_311 0 -3.6339959509242947e-03
GC_1_312 b_1 NI_1 NS_312 0 2.5967283187350904e-03
GC_1_313 b_1 NI_1 NS_313 0 -2.8319057300553504e-03
GC_1_314 b_1 NI_1 NS_314 0 3.9895611145249052e-03
GC_1_315 b_1 NI_1 NS_315 0 -2.2141465854295827e-04
GC_1_316 b_1 NI_1 NS_316 0 -4.2135156478468007e-03
GC_1_317 b_1 NI_1 NS_317 0 -9.8958396334079424e-06
GC_1_318 b_1 NI_1 NS_318 0 7.5257580410616705e-06
GC_1_319 b_1 NI_1 NS_319 0 -1.3539532717406016e-03
GC_1_320 b_1 NI_1 NS_320 0 3.3754867364988645e-03
GC_1_321 b_1 NI_1 NS_321 0 -9.6985114955971832e-04
GC_1_322 b_1 NI_1 NS_322 0 -4.3479519128989457e-03
GC_1_323 b_1 NI_1 NS_323 0 -1.0009104611191882e-03
GC_1_324 b_1 NI_1 NS_324 0 2.2213067654239531e-03
GC_1_325 b_1 NI_1 NS_325 0 -1.6517261451508955e-03
GC_1_326 b_1 NI_1 NS_326 0 -4.4093120919419665e-03
GC_1_327 b_1 NI_1 NS_327 0 -1.4483164113443176e-03
GC_1_328 b_1 NI_1 NS_328 0 -2.4971461095301159e-03
GC_1_329 b_1 NI_1 NS_329 0 7.8219531514154260e-04
GC_1_330 b_1 NI_1 NS_330 0 2.5933467042053913e-03
GC_1_331 b_1 NI_1 NS_331 0 -6.9628504516090653e-04
GC_1_332 b_1 NI_1 NS_332 0 2.8792034901541472e-03
GC_1_333 b_1 NI_1 NS_333 0 -1.4353710703639581e-03
GC_1_334 b_1 NI_1 NS_334 0 -2.7718619392427786e-03
GC_1_335 b_1 NI_1 NS_335 0 -1.1678495857965199e-03
GC_1_336 b_1 NI_1 NS_336 0 2.6661993124953787e-03
GC_1_337 b_1 NI_1 NS_337 0 7.8075943466351103e-04
GC_1_338 b_1 NI_1 NS_338 0 -1.8746156136009921e-03
GC_1_339 b_1 NI_1 NS_339 0 2.3789690379687181e-08
GC_1_340 b_1 NI_1 NS_340 0 -6.0253482765046754e-08
GC_1_341 b_1 NI_1 NS_341 0 -9.0373275433935194e-07
GC_1_342 b_1 NI_1 NS_342 0 3.2031385932357687e-06
GC_1_343 b_1 NI_1 NS_343 0 2.9495781541059697e-03
GC_1_344 b_1 NI_1 NS_344 0 -6.1234119963752014e-04
GC_1_345 b_1 NI_1 NS_345 0 2.7949880247010815e-08
GC_1_346 b_1 NI_1 NS_346 0 -3.1702432499492385e-08
GC_1_347 b_1 NI_1 NS_347 0 2.0347278449610806e-04
GC_1_348 b_1 NI_1 NS_348 0 1.3799473859673318e-04
GC_1_349 b_1 NI_1 NS_349 0 5.6259278867111235e-04
GC_1_350 b_1 NI_1 NS_350 0 2.6570817171653430e-04
GC_1_351 b_1 NI_1 NS_351 0 3.1064667357130222e-03
GC_1_352 b_1 NI_1 NS_352 0 -2.2048923971853063e-03
GC_1_353 b_1 NI_1 NS_353 0 -1.5822543810086924e-03
GC_1_354 b_1 NI_1 NS_354 0 -2.6870784552691352e-03
GC_1_355 b_1 NI_1 NS_355 0 -2.0496562077166047e-03
GC_1_356 b_1 NI_1 NS_356 0 -3.7885102902007685e-03
GC_1_357 b_1 NI_1 NS_357 0 -4.9745615347427307e-03
GC_1_358 b_1 NI_1 NS_358 0 -1.5415295611829773e-03
GC_1_359 b_1 NI_1 NS_359 0 2.9290598381321984e-04
GC_1_360 b_1 NI_1 NS_360 0 1.9565108914326823e-04
GC_1_361 b_1 NI_1 NS_361 0 -2.8663286944718754e-03
GC_1_362 b_1 NI_1 NS_362 0 -9.5746369397000915e-04
GC_1_363 b_1 NI_1 NS_363 0 -2.2151869990957460e-02
GC_1_364 b_1 NI_1 NS_364 0 -1.0226316050092915e-02
GC_1_365 b_1 NI_1 NS_365 0 1.1324964778460372e-03
GC_1_366 b_1 NI_1 NS_366 0 2.0395319713006642e-02
GC_1_367 b_1 NI_1 NS_367 0 -5.8416210173243572e-03
GC_1_368 b_1 NI_1 NS_368 0 4.6116288232749443e-03
GC_1_369 b_1 NI_1 NS_369 0 5.7171498002332498e-03
GC_1_370 b_1 NI_1 NS_370 0 3.4516070764761521e-02
GC_1_371 b_1 NI_1 NS_371 0 8.0342761959906299e-03
GC_1_372 b_1 NI_1 NS_372 0 2.7930240306842185e-03
GC_1_373 b_1 NI_1 NS_373 0 -7.7724214964439604e-03
GC_1_374 b_1 NI_1 NS_374 0 2.9556754323995484e-02
GC_1_375 b_1 NI_1 NS_375 0 5.0768430142714455e-02
GC_1_376 b_1 NI_1 NS_376 0 -2.0072961102686377e-02
GC_1_377 b_1 NI_1 NS_377 0 7.9195785261018965e-03
GC_1_378 b_1 NI_1 NS_378 0 -1.6364409984739659e-03
GC_1_379 b_1 NI_1 NS_379 0 2.9084860001785985e-02
GC_1_380 b_1 NI_1 NS_380 0 -2.6464736593899429e-02
GC_1_381 b_1 NI_1 NS_381 0 -6.7250677010260501e-03
GC_1_382 b_1 NI_1 NS_382 0 -9.8822057179754775e-03
GC_1_383 b_1 NI_1 NS_383 0 8.4630826882353544e-03
GC_1_384 b_1 NI_1 NS_384 0 -8.0277980858305328e-03
GC_1_385 b_1 NI_1 NS_385 0 -1.8994952670628965e-02
GC_1_386 b_1 NI_1 NS_386 0 -2.5238422123919302e-02
GC_1_387 b_1 NI_1 NS_387 0 -5.4717850937434408e-03
GC_1_388 b_1 NI_1 NS_388 0 -2.8547841795536744e-03
GC_1_389 b_1 NI_1 NS_389 0 -1.7741074142562405e-02
GC_1_390 b_1 NI_1 NS_390 0 -1.3132230479676280e-02
GC_1_391 b_1 NI_1 NS_391 0 -4.8178007911030656e-03
GC_1_392 b_1 NI_1 NS_392 0 1.2541404259819212e-02
GC_1_393 b_1 NI_1 NS_393 0 -3.4590901728862159e-03
GC_1_394 b_1 NI_1 NS_394 0 1.5412380194080328e-03
GC_1_395 b_1 NI_1 NS_395 0 -7.1865218186604280e-04
GC_1_396 b_1 NI_1 NS_396 0 7.0058606429342285e-03
GC_1_397 b_1 NI_1 NS_397 0 1.8820411281323356e-03
GC_1_398 b_1 NI_1 NS_398 0 8.5748803355927306e-05
GC_1_399 b_1 NI_1 NS_399 0 3.1400256685555324e-04
GC_1_400 b_1 NI_1 NS_400 0 -1.9467011484858314e-03
GC_1_401 b_1 NI_1 NS_401 0 -1.8563356155217418e-03
GC_1_402 b_1 NI_1 NS_402 0 -1.6182086453746134e-03
GC_1_403 b_1 NI_1 NS_403 0 -2.1290963631129846e-03
GC_1_404 b_1 NI_1 NS_404 0 1.6850438918243513e-03
GC_1_405 b_1 NI_1 NS_405 0 7.6361034722424140e-04
GC_1_406 b_1 NI_1 NS_406 0 1.8527544762886151e-04
GC_1_407 b_1 NI_1 NS_407 0 -6.9730352436409211e-04
GC_1_408 b_1 NI_1 NS_408 0 -1.6780698211294270e-03
GC_1_409 b_1 NI_1 NS_409 0 -2.6815283771762172e-03
GC_1_410 b_1 NI_1 NS_410 0 -8.2749104579960128e-04
GC_1_411 b_1 NI_1 NS_411 0 -4.9989643564299965e-04
GC_1_412 b_1 NI_1 NS_412 0 2.9288646769845515e-03
GC_1_413 b_1 NI_1 NS_413 0 1.3533577789987892e-03
GC_1_414 b_1 NI_1 NS_414 0 -8.5805557051073830e-04
GC_1_415 b_1 NI_1 NS_415 0 -2.4189241805641268e-03
GC_1_416 b_1 NI_1 NS_416 0 -2.2676207872691064e-03
GC_1_417 b_1 NI_1 NS_417 0 -3.5540452699943975e-03
GC_1_418 b_1 NI_1 NS_418 0 7.4852702206970926e-04
GC_1_419 b_1 NI_1 NS_419 0 2.4633835839580295e-03
GC_1_420 b_1 NI_1 NS_420 0 3.0182798439779661e-03
GC_1_421 b_1 NI_1 NS_421 0 9.8455418912004960e-04
GC_1_422 b_1 NI_1 NS_422 0 -2.9418100609102447e-03
GC_1_423 b_1 NI_1 NS_423 0 -4.7678000310426042e-03
GC_1_424 b_1 NI_1 NS_424 0 5.4340225271683148e-05
GC_1_425 b_1 NI_1 NS_425 0 -1.7083703564014403e-03
GC_1_426 b_1 NI_1 NS_426 0 3.7124270138559094e-03
GC_1_427 b_1 NI_1 NS_427 0 -7.6587643484793497e-04
GC_1_428 b_1 NI_1 NS_428 0 1.5006814834019342e-03
GC_1_429 b_1 NI_1 NS_429 0 3.2213016671005456e-03
GC_1_430 b_1 NI_1 NS_430 0 -1.3508683621748624e-03
GC_1_431 b_1 NI_1 NS_431 0 -2.9326074906924854e-06
GC_1_432 b_1 NI_1 NS_432 0 8.7469702082612298e-06
GC_1_433 b_1 NI_1 NS_433 0 -1.8200418648386203e-03
GC_1_434 b_1 NI_1 NS_434 0 -2.5277363336050690e-03
GC_1_435 b_1 NI_1 NS_435 0 -2.4072534073868333e-03
GC_1_436 b_1 NI_1 NS_436 0 2.4886635241563376e-03
GC_1_437 b_1 NI_1 NS_437 0 1.0142619049036408e-03
GC_1_438 b_1 NI_1 NS_438 0 2.4256812017993280e-03
GC_1_439 b_1 NI_1 NS_439 0 8.5775930065578384e-04
GC_1_440 b_1 NI_1 NS_440 0 -2.6994852973402559e-03
GC_1_441 b_1 NI_1 NS_441 0 -3.0644787207095847e-04
GC_1_442 b_1 NI_1 NS_442 0 1.6741356690644210e-03
GC_1_443 b_1 NI_1 NS_443 0 -1.7840540679053948e-03
GC_1_444 b_1 NI_1 NS_444 0 -3.1181081247855653e-04
GC_1_445 b_1 NI_1 NS_445 0 1.4004539637538394e-03
GC_1_446 b_1 NI_1 NS_446 0 1.9709615797124020e-03
GC_1_447 b_1 NI_1 NS_447 0 1.0449287362756718e-03
GC_1_448 b_1 NI_1 NS_448 0 -2.2998045682780664e-03
GC_1_449 b_1 NI_1 NS_449 0 -6.9799494563789184e-04
GC_1_450 b_1 NI_1 NS_450 0 -1.4668898799569078e-03
GC_1_451 b_1 NI_1 NS_451 0 -1.3735491330375937e-03
GC_1_452 b_1 NI_1 NS_452 0 -3.1252861563721321e-04
GC_1_453 b_1 NI_1 NS_453 0 7.1030065532240196e-09
GC_1_454 b_1 NI_1 NS_454 0 -2.4710001485461635e-08
GC_1_455 b_1 NI_1 NS_455 0 -4.5275410590251481e-07
GC_1_456 b_1 NI_1 NS_456 0 1.6341839063988990e-06
GC_1_457 b_1 NI_1 NS_457 0 -1.1990417494770154e-04
GC_1_458 b_1 NI_1 NS_458 0 -2.1506583650043852e-06
GC_1_459 b_1 NI_1 NS_459 0 -2.4444181869517410e-10
GC_1_460 b_1 NI_1 NS_460 0 2.5345872105997169e-09
GC_1_461 b_1 NI_1 NS_461 0 1.5459797321879491e-06
GC_1_462 b_1 NI_1 NS_462 0 -1.4954279553507424e-06
GC_1_463 b_1 NI_1 NS_463 0 -2.6328536416109721e-08
GC_1_464 b_1 NI_1 NS_464 0 -6.1347873549544356e-06
GC_1_465 b_1 NI_1 NS_465 0 -7.5890813287154378e-06
GC_1_466 b_1 NI_1 NS_466 0 6.3141454132102551e-07
GC_1_467 b_1 NI_1 NS_467 0 -9.4093710326879636e-07
GC_1_468 b_1 NI_1 NS_468 0 -4.4034014664471327e-06
GC_1_469 b_1 NI_1 NS_469 0 -1.5515996091878922e-05
GC_1_470 b_1 NI_1 NS_470 0 -1.2262226854320398e-06
GC_1_471 b_1 NI_1 NS_471 0 -5.1272331084723988e-06
GC_1_472 b_1 NI_1 NS_472 0 1.9057488954927098e-05
GC_1_473 b_1 NI_1 NS_473 0 4.3659579714125282e-06
GC_1_474 b_1 NI_1 NS_474 0 -3.1091685775347459e-06
GC_1_475 b_1 NI_1 NS_475 0 1.2739373771324426e-07
GC_1_476 b_1 NI_1 NS_476 0 -2.6189011077477678e-06
GC_1_477 b_1 NI_1 NS_477 0 -2.4695118996629760e-05
GC_1_478 b_1 NI_1 NS_478 0 2.8214913375080709e-05
GC_1_479 b_1 NI_1 NS_479 0 2.7678010939608789e-05
GC_1_480 b_1 NI_1 NS_480 0 -8.8491167123092485e-06
GC_1_481 b_1 NI_1 NS_481 0 -7.7786901490916476e-06
GC_1_482 b_1 NI_1 NS_482 0 -4.1717376937000054e-06
GC_1_483 b_1 NI_1 NS_483 0 1.2852721310710080e-05
GC_1_484 b_1 NI_1 NS_484 0 2.5989432197929272e-05
GC_1_485 b_1 NI_1 NS_485 0 1.3965873953305457e-06
GC_1_486 b_1 NI_1 NS_486 0 -8.8467713497858762e-06
GC_1_487 b_1 NI_1 NS_487 0 -2.7274070196427769e-05
GC_1_488 b_1 NI_1 NS_488 0 5.0518926545830929e-06
GC_1_489 b_1 NI_1 NS_489 0 4.0358168245698754e-05
GC_1_490 b_1 NI_1 NS_490 0 9.5136818803633682e-06
GC_1_491 b_1 NI_1 NS_491 0 -2.8939298143949531e-06
GC_1_492 b_1 NI_1 NS_492 0 -4.3230654360941788e-06
GC_1_493 b_1 NI_1 NS_493 0 1.3068135383984228e-05
GC_1_494 b_1 NI_1 NS_494 0 1.8039409445944825e-05
GC_1_495 b_1 NI_1 NS_495 0 3.4806889754966687e-06
GC_1_496 b_1 NI_1 NS_496 0 -1.0690735109510123e-05
GC_1_497 b_1 NI_1 NS_497 0 -6.1534218532278669e-06
GC_1_498 b_1 NI_1 NS_498 0 1.0246667669107377e-06
GC_1_499 b_1 NI_1 NS_499 0 1.8579425134837087e-05
GC_1_500 b_1 NI_1 NS_500 0 4.7194965170093430e-06
GC_1_501 b_1 NI_1 NS_501 0 -1.7163671058541620e-07
GC_1_502 b_1 NI_1 NS_502 0 -4.0410338239184102e-06
GC_1_503 b_1 NI_1 NS_503 0 5.3110690603834932e-06
GC_1_504 b_1 NI_1 NS_504 0 1.3887857538476306e-05
GC_1_505 b_1 NI_1 NS_505 0 7.3444730001178477e-06
GC_1_506 b_1 NI_1 NS_506 0 -1.1159205118327633e-05
GC_1_507 b_1 NI_1 NS_507 0 -1.3421715236458289e-06
GC_1_508 b_1 NI_1 NS_508 0 1.0174183386021314e-06
GC_1_509 b_1 NI_1 NS_509 0 1.0876590979840572e-05
GC_1_510 b_1 NI_1 NS_510 0 3.8402785230580925e-06
GC_1_511 b_1 NI_1 NS_511 0 1.6848231938441983e-06
GC_1_512 b_1 NI_1 NS_512 0 -6.0383775016051198e-07
GC_1_513 b_1 NI_1 NS_513 0 5.6746775701362120e-06
GC_1_514 b_1 NI_1 NS_514 0 1.5928962077412817e-06
GC_1_515 b_1 NI_1 NS_515 0 3.3876857670137650e-06
GC_1_516 b_1 NI_1 NS_516 0 2.0447826012803304e-06
GC_1_517 b_1 NI_1 NS_517 0 1.1009150564419416e-05
GC_1_518 b_1 NI_1 NS_518 0 3.6665169529882541e-06
GC_1_519 b_1 NI_1 NS_519 0 4.8524824080097361e-06
GC_1_520 b_1 NI_1 NS_520 0 -9.3154851253556022e-08
GC_1_521 b_1 NI_1 NS_521 0 9.9846404485454234e-06
GC_1_522 b_1 NI_1 NS_522 0 -1.1688006959200438e-06
GC_1_523 b_1 NI_1 NS_523 0 8.2907545265570333e-06
GC_1_524 b_1 NI_1 NS_524 0 2.9619522292149753e-06
GC_1_525 b_1 NI_1 NS_525 0 1.9135356772703823e-05
GC_1_526 b_1 NI_1 NS_526 0 -5.6872192956509124e-06
GC_1_527 b_1 NI_1 NS_527 0 7.2561492281017364e-06
GC_1_528 b_1 NI_1 NS_528 0 -4.0375690947185186e-06
GC_1_529 b_1 NI_1 NS_529 0 1.3814375078115959e-05
GC_1_530 b_1 NI_1 NS_530 0 -1.2017012207963864e-05
GC_1_531 b_1 NI_1 NS_531 0 1.2524732497661204e-05
GC_1_532 b_1 NI_1 NS_532 0 -3.9196656912671611e-06
GC_1_533 b_1 NI_1 NS_533 0 9.3874027572219420e-06
GC_1_534 b_1 NI_1 NS_534 0 -2.7008491502144383e-05
GC_1_535 b_1 NI_1 NS_535 0 2.5340514268338131e-06
GC_1_536 b_1 NI_1 NS_536 0 -1.2433576141289434e-05
GC_1_537 b_1 NI_1 NS_537 0 -8.1011417799400451e-06
GC_1_538 b_1 NI_1 NS_538 0 -1.8935730184699154e-05
GC_1_539 b_1 NI_1 NS_539 0 -4.4539202387794539e-06
GC_1_540 b_1 NI_1 NS_540 0 -1.2056803182112205e-05
GC_1_541 b_1 NI_1 NS_541 0 5.2729053246588910e-05
GC_1_542 b_1 NI_1 NS_542 0 -8.9465544133772773e-05
GC_1_543 b_1 NI_1 NS_543 0 -9.8695738088673526e-06
GC_1_544 b_1 NI_1 NS_544 0 5.5951776949728550e-07
GC_1_545 b_1 NI_1 NS_545 0 3.8236082281730305e-07
GC_1_546 b_1 NI_1 NS_546 0 -1.3957348952537372e-07
GC_1_547 b_1 NI_1 NS_547 0 -2.6066256150927539e-06
GC_1_548 b_1 NI_1 NS_548 0 -2.3472560403143718e-06
GC_1_549 b_1 NI_1 NS_549 0 -4.4561577908256142e-06
GC_1_550 b_1 NI_1 NS_550 0 2.3602450172532859e-07
GC_1_551 b_1 NI_1 NS_551 0 -1.7027355507051956e-05
GC_1_552 b_1 NI_1 NS_552 0 9.6526753420072147e-06
GC_1_553 b_1 NI_1 NS_553 0 -8.5113172944890925e-06
GC_1_554 b_1 NI_1 NS_554 0 3.7251828213227478e-05
GC_1_555 b_1 NI_1 NS_555 0 -7.2790849411971916e-06
GC_1_556 b_1 NI_1 NS_556 0 3.7957320119752530e-07
GC_1_557 b_1 NI_1 NS_557 0 -1.3447171408941609e-05
GC_1_558 b_1 NI_1 NS_558 0 1.9992894790493110e-06
GC_1_559 b_1 NI_1 NS_559 0 -4.6778654391756952e-06
GC_1_560 b_1 NI_1 NS_560 0 -3.4374763006582938e-06
GC_1_561 b_1 NI_1 NS_561 0 -6.4554994626799839e-06
GC_1_562 b_1 NI_1 NS_562 0 1.0434673332689180e-06
GC_1_563 b_1 NI_1 NS_563 0 -3.0715773663287049e-06
GC_1_564 b_1 NI_1 NS_564 0 8.7380281211515957e-07
GC_1_565 b_1 NI_1 NS_565 0 -1.8084091449414782e-06
GC_1_566 b_1 NI_1 NS_566 0 -9.3492553452635466e-07
GC_1_567 b_1 NI_1 NS_567 0 -2.5769931072136170e-10
GC_1_568 b_1 NI_1 NS_568 0 4.1862387056011173e-10
GC_1_569 b_1 NI_1 NS_569 0 2.1402119757677950e-09
GC_1_570 b_1 NI_1 NS_570 0 -2.6513264309540877e-08
GC_1_571 b_1 NI_1 NS_571 0 -3.8127618243054336e-05
GC_1_572 b_1 NI_1 NS_572 0 2.2429770296472153e-06
GC_1_573 b_1 NI_1 NS_573 0 5.7510756613961427e-11
GC_1_574 b_1 NI_1 NS_574 0 3.0676920984028503e-09
GC_1_575 b_1 NI_1 NS_575 0 -1.9281110935481452e-06
GC_1_576 b_1 NI_1 NS_576 0 -1.7008096195617562e-06
GC_1_577 b_1 NI_1 NS_577 0 -5.6014742201550229e-06
GC_1_578 b_1 NI_1 NS_578 0 2.8809782733150529e-06
GC_1_579 b_1 NI_1 NS_579 0 -1.6609396165968357e-05
GC_1_580 b_1 NI_1 NS_580 0 1.9115783992859909e-05
GC_1_581 b_1 NI_1 NS_581 0 1.5381277700843868e-05
GC_1_582 b_1 NI_1 NS_582 0 1.0271581209289325e-05
GC_1_583 b_1 NI_1 NS_583 0 1.7283130657142685e-05
GC_1_584 b_1 NI_1 NS_584 0 2.3212263410403662e-05
GC_1_585 b_1 NI_1 NS_585 0 3.0965021174760464e-05
GC_1_586 b_1 NI_1 NS_586 0 5.3090203270968456e-06
GC_1_587 b_1 NI_1 NS_587 0 -3.3865846603746305e-06
GC_1_588 b_1 NI_1 NS_588 0 -2.1456123687085187e-06
GC_1_589 b_1 NI_1 NS_589 0 1.7199398202451132e-05
GC_1_590 b_1 NI_1 NS_590 0 -2.1238079077130038e-06
GC_1_591 b_1 NI_1 NS_591 0 1.2959165088019967e-04
GC_1_592 b_1 NI_1 NS_592 0 3.5268879846131514e-05
GC_1_593 b_1 NI_1 NS_593 0 -2.8361254280399520e-05
GC_1_594 b_1 NI_1 NS_594 0 -1.0001870928486552e-04
GC_1_595 b_1 NI_1 NS_595 0 2.5325861958929697e-05
GC_1_596 b_1 NI_1 NS_596 0 -3.1108754036155923e-05
GC_1_597 b_1 NI_1 NS_597 0 -4.1100399421461918e-05
GC_1_598 b_1 NI_1 NS_598 0 -1.6753409185215682e-04
GC_1_599 b_1 NI_1 NS_599 0 -4.1818796508857966e-05
GC_1_600 b_1 NI_1 NS_600 0 -5.5999251305126259e-06
GC_1_601 b_1 NI_1 NS_601 0 2.2902358278411213e-05
GC_1_602 b_1 NI_1 NS_602 0 -1.5132347450534878e-04
GC_1_603 b_1 NI_1 NS_603 0 -2.3194036291446376e-04
GC_1_604 b_1 NI_1 NS_604 0 1.1299732194006234e-04
GC_1_605 b_1 NI_1 NS_605 0 -3.7469245066163350e-05
GC_1_606 b_1 NI_1 NS_606 0 1.3726671842994912e-05
GC_1_607 b_1 NI_1 NS_607 0 -1.3772298261734381e-04
GC_1_608 b_1 NI_1 NS_608 0 1.2973732668858273e-04
GC_1_609 b_1 NI_1 NS_609 0 3.6014580459039122e-05
GC_1_610 b_1 NI_1 NS_610 0 4.1758562882016404e-05
GC_1_611 b_1 NI_1 NS_611 0 -3.8325643077279527e-05
GC_1_612 b_1 NI_1 NS_612 0 4.2732816956013462e-05
GC_1_613 b_1 NI_1 NS_613 0 8.7551061748031848e-05
GC_1_614 b_1 NI_1 NS_614 0 1.1830579977033164e-04
GC_1_615 b_1 NI_1 NS_615 0 2.7199706151306579e-05
GC_1_616 b_1 NI_1 NS_616 0 1.0487347513925878e-05
GC_1_617 b_1 NI_1 NS_617 0 8.6918390797216294e-05
GC_1_618 b_1 NI_1 NS_618 0 6.5387623415457402e-05
GC_1_619 b_1 NI_1 NS_619 0 2.0649678663307343e-05
GC_1_620 b_1 NI_1 NS_620 0 -5.7329129905617912e-05
GC_1_621 b_1 NI_1 NS_621 0 1.7010777862364386e-05
GC_1_622 b_1 NI_1 NS_622 0 -8.6980471918995415e-06
GC_1_623 b_1 NI_1 NS_623 0 8.3266740916594054e-06
GC_1_624 b_1 NI_1 NS_624 0 -3.3101616471253901e-05
GC_1_625 b_1 NI_1 NS_625 0 -8.8261838370693839e-06
GC_1_626 b_1 NI_1 NS_626 0 3.3237480204381289e-07
GC_1_627 b_1 NI_1 NS_627 0 -2.3513350115789503e-06
GC_1_628 b_1 NI_1 NS_628 0 8.4561590396524091e-06
GC_1_629 b_1 NI_1 NS_629 0 1.0134444151928945e-05
GC_1_630 b_1 NI_1 NS_630 0 6.1702244373529140e-06
GC_1_631 b_1 NI_1 NS_631 0 1.2106296708449743e-05
GC_1_632 b_1 NI_1 NS_632 0 -7.8948444101772782e-06
GC_1_633 b_1 NI_1 NS_633 0 -3.4457719645756991e-06
GC_1_634 b_1 NI_1 NS_634 0 -5.4105727583616130e-07
GC_1_635 b_1 NI_1 NS_635 0 2.5534795467902545e-06
GC_1_636 b_1 NI_1 NS_636 0 7.3550292759749945e-06
GC_1_637 b_1 NI_1 NS_637 0 1.3648108139347366e-05
GC_1_638 b_1 NI_1 NS_638 0 2.7056951847831875e-06
GC_1_639 b_1 NI_1 NS_639 0 4.5460332843596275e-06
GC_1_640 b_1 NI_1 NS_640 0 -1.4254844430092434e-05
GC_1_641 b_1 NI_1 NS_641 0 -5.8809758975686397e-06
GC_1_642 b_1 NI_1 NS_642 0 4.1779280557322787e-06
GC_1_643 b_1 NI_1 NS_643 0 1.0407133900258957e-05
GC_1_644 b_1 NI_1 NS_644 0 9.8673482856852675e-06
GC_1_645 b_1 NI_1 NS_645 0 1.7371587674168731e-05
GC_1_646 b_1 NI_1 NS_646 0 -4.2134163554901156e-06
GC_1_647 b_1 NI_1 NS_647 0 -9.1860362040983230e-06
GC_1_648 b_1 NI_1 NS_648 0 -1.5417459336232890e-05
GC_1_649 b_1 NI_1 NS_649 0 -3.9937462921714397e-06
GC_1_650 b_1 NI_1 NS_650 0 1.3459827800278997e-05
GC_1_651 b_1 NI_1 NS_651 0 2.1061339055209568e-05
GC_1_652 b_1 NI_1 NS_652 0 -6.9754286162137272e-07
GC_1_653 b_1 NI_1 NS_653 0 9.0885522481808230e-06
GC_1_654 b_1 NI_1 NS_654 0 -1.7352306203978696e-05
GC_1_655 b_1 NI_1 NS_655 0 1.8901171594397829e-06
GC_1_656 b_1 NI_1 NS_656 0 -1.4898997365206833e-05
GC_1_657 b_1 NI_1 NS_657 0 -1.3643855850568576e-05
GC_1_658 b_1 NI_1 NS_658 0 4.0672393101359127e-06
GC_1_659 b_1 NI_1 NS_659 0 1.3198585075412352e-08
GC_1_660 b_1 NI_1 NS_660 0 -4.9292708817307030e-08
GC_1_661 b_1 NI_1 NS_661 0 8.7094375253196080e-06
GC_1_662 b_1 NI_1 NS_662 0 1.1413291482407200e-05
GC_1_663 b_1 NI_1 NS_663 0 1.0949792347002537e-05
GC_1_664 b_1 NI_1 NS_664 0 -1.1467445742355033e-05
GC_1_665 b_1 NI_1 NS_665 0 -3.5677400524012549e-06
GC_1_666 b_1 NI_1 NS_666 0 -1.0053466146405010e-05
GC_1_667 b_1 NI_1 NS_667 0 -2.0108126116167848e-06
GC_1_668 b_1 NI_1 NS_668 0 1.3050038459178061e-05
GC_1_669 b_1 NI_1 NS_669 0 9.7275560318863426e-07
GC_1_670 b_1 NI_1 NS_670 0 -7.2791644972848783e-06
GC_1_671 b_1 NI_1 NS_671 0 7.4349154440459069e-06
GC_1_672 b_1 NI_1 NS_672 0 1.7180971658735462e-06
GC_1_673 b_1 NI_1 NS_673 0 -6.1040294984975425e-06
GC_1_674 b_1 NI_1 NS_674 0 -8.8986487325647160e-06
GC_1_675 b_1 NI_1 NS_675 0 -4.1281685758378263e-06
GC_1_676 b_1 NI_1 NS_676 0 9.6390248418877161e-06
GC_1_677 b_1 NI_1 NS_677 0 3.3246453370566033e-06
GC_1_678 b_1 NI_1 NS_678 0 6.0744663520002685e-06
GC_1_679 b_1 NI_1 NS_679 0 5.7495181646459397e-06
GC_1_680 b_1 NI_1 NS_680 0 5.2304198756832159e-07
GC_1_681 b_1 NI_1 NS_681 0 5.7043206283872192e-11
GC_1_682 b_1 NI_1 NS_682 0 1.4838853948537982e-10
GC_1_683 b_1 NI_1 NS_683 0 6.0313697961434863e-09
GC_1_684 b_1 NI_1 NS_684 0 -8.4056175185868739e-09
GC_1_685 b_1 NI_1 NS_685 0 6.6701490246950346e-05
GC_1_686 b_1 NI_1 NS_686 0 2.1487593113722078e-07
GC_1_687 b_1 NI_1 NS_687 0 2.2380668209054809e-11
GC_1_688 b_1 NI_1 NS_688 0 -9.9152092431020436e-10
GC_1_689 b_1 NI_1 NS_689 0 4.3114279902238446e-07
GC_1_690 b_1 NI_1 NS_690 0 1.8615289531319374e-07
GC_1_691 b_1 NI_1 NS_691 0 6.0533473004313551e-07
GC_1_692 b_1 NI_1 NS_692 0 5.0362668621704696e-07
GC_1_693 b_1 NI_1 NS_693 0 2.9724324468424571e-06
GC_1_694 b_1 NI_1 NS_694 0 -1.5630087690921464e-06
GC_1_695 b_1 NI_1 NS_695 0 -1.1990738041424137e-06
GC_1_696 b_1 NI_1 NS_696 0 -1.1274223172713372e-06
GC_1_697 b_1 NI_1 NS_697 0 2.3740973804667618e-06
GC_1_698 b_1 NI_1 NS_698 0 -8.7014361544288491e-07
GC_1_699 b_1 NI_1 NS_699 0 -2.5791855801999536e-06
GC_1_700 b_1 NI_1 NS_700 0 -6.4188239898857804e-06
GC_1_701 b_1 NI_1 NS_701 0 1.1120405169811142e-07
GC_1_702 b_1 NI_1 NS_702 0 1.6980772037795315e-06
GC_1_703 b_1 NI_1 NS_703 0 -1.7225276156704670e-06
GC_1_704 b_1 NI_1 NS_704 0 5.0765299801755539e-07
GC_1_705 b_1 NI_1 NS_705 0 3.1223283398785453e-06
GC_1_706 b_1 NI_1 NS_706 0 -4.3467334270915486e-06
GC_1_707 b_1 NI_1 NS_707 0 -6.6651234546803577e-06
GC_1_708 b_1 NI_1 NS_708 0 1.1614607025116634e-06
GC_1_709 b_1 NI_1 NS_709 0 -4.7510515756048819e-07
GC_1_710 b_1 NI_1 NS_710 0 1.6872439520213062e-06
GC_1_711 b_1 NI_1 NS_711 0 -2.1293716842352186e-06
GC_1_712 b_1 NI_1 NS_712 0 -4.2560152914789083e-06
GC_1_713 b_1 NI_1 NS_713 0 -2.2153029186094944e-06
GC_1_714 b_1 NI_1 NS_714 0 2.1659200625242935e-06
GC_1_715 b_1 NI_1 NS_715 0 3.1593370700088968e-06
GC_1_716 b_1 NI_1 NS_716 0 3.0711637056328444e-06
GC_1_717 b_1 NI_1 NS_717 0 -6.0923082511330965e-06
GC_1_718 b_1 NI_1 NS_718 0 -4.4508802780496267e-06
GC_1_719 b_1 NI_1 NS_719 0 -1.2975249857838159e-06
GC_1_720 b_1 NI_1 NS_720 0 2.1675952668669274e-06
GC_1_721 b_1 NI_1 NS_721 0 2.8169568021362270e-07
GC_1_722 b_1 NI_1 NS_722 0 -2.8035795586186740e-06
GC_1_723 b_1 NI_1 NS_723 0 -3.1939610604328982e-06
GC_1_724 b_1 NI_1 NS_724 0 1.8340042060102757e-06
GC_1_725 b_1 NI_1 NS_725 0 -3.1234118303491942e-07
GC_1_726 b_1 NI_1 NS_726 0 2.3430253997579803e-06
GC_1_727 b_1 NI_1 NS_727 0 -1.4637172335766488e-06
GC_1_728 b_1 NI_1 NS_728 0 -2.6210648393144875e-06
GC_1_729 b_1 NI_1 NS_729 0 -1.8974252865670412e-06
GC_1_730 b_1 NI_1 NS_730 0 1.3687529716579467e-06
GC_1_731 b_1 NI_1 NS_731 0 1.1585925632264011e-06
GC_1_732 b_1 NI_1 NS_732 0 -6.4540652719473749e-07
GC_1_733 b_1 NI_1 NS_733 0 -3.5960772126802328e-06
GC_1_734 b_1 NI_1 NS_734 0 2.8645391862162086e-07
GC_1_735 b_1 NI_1 NS_735 0 -8.2546538260808026e-07
GC_1_736 b_1 NI_1 NS_736 0 7.2322604869650604e-07
GC_1_737 b_1 NI_1 NS_737 0 -1.8925809065824413e-06
GC_1_738 b_1 NI_1 NS_738 0 -1.3277323206558993e-06
GC_1_739 b_1 NI_1 NS_739 0 -1.4489409937888748e-06
GC_1_740 b_1 NI_1 NS_740 0 5.5829974849458577e-07
GC_1_741 b_1 NI_1 NS_741 0 -1.0698697004329278e-06
GC_1_742 b_1 NI_1 NS_742 0 -5.9277137671907856e-07
GC_1_743 b_1 NI_1 NS_743 0 -2.3266422409217864e-06
GC_1_744 b_1 NI_1 NS_744 0 -6.7325042795127172e-07
GC_1_745 b_1 NI_1 NS_745 0 -2.8005575822005168e-06
GC_1_746 b_1 NI_1 NS_746 0 -5.7579604098330063e-07
GC_1_747 b_1 NI_1 NS_747 0 -2.0701486110218062e-06
GC_1_748 b_1 NI_1 NS_748 0 2.3474597420323596e-07
GC_1_749 b_1 NI_1 NS_749 0 -2.5970654227936913e-06
GC_1_750 b_1 NI_1 NS_750 0 1.0366584562903118e-07
GC_1_751 b_1 NI_1 NS_751 0 -3.9148792414820219e-06
GC_1_752 b_1 NI_1 NS_752 0 -7.2842823073807339e-07
GC_1_753 b_1 NI_1 NS_753 0 -5.2762864252069513e-06
GC_1_754 b_1 NI_1 NS_754 0 1.8897604776495205e-06
GC_1_755 b_1 NI_1 NS_755 0 -2.9592146633652752e-06
GC_1_756 b_1 NI_1 NS_756 0 1.7284778153242393e-06
GC_1_757 b_1 NI_1 NS_757 0 -3.7956743303695738e-06
GC_1_758 b_1 NI_1 NS_758 0 2.9627451811167990e-06
GC_1_759 b_1 NI_1 NS_759 0 -5.2520803366240319e-06
GC_1_760 b_1 NI_1 NS_760 0 1.3679661614965092e-06
GC_1_761 b_1 NI_1 NS_761 0 -2.9739722128864600e-06
GC_1_762 b_1 NI_1 NS_762 0 7.6177906559748348e-06
GC_1_763 b_1 NI_1 NS_763 0 -1.9309243732355516e-06
GC_1_764 b_1 NI_1 NS_764 0 4.3923521136705281e-06
GC_1_765 b_1 NI_1 NS_765 0 1.5636688114064320e-06
GC_1_766 b_1 NI_1 NS_766 0 4.8436709892747677e-06
GC_1_767 b_1 NI_1 NS_767 0 -9.8795309155149944e-07
GC_1_768 b_1 NI_1 NS_768 0 3.6442588135305073e-06
GC_1_769 b_1 NI_1 NS_769 0 -1.0320720134545872e-05
GC_1_770 b_1 NI_1 NS_770 0 3.3102413321429392e-05
GC_1_771 b_1 NI_1 NS_771 0 1.3164909029001369e-06
GC_1_772 b_1 NI_1 NS_772 0 1.2184828977595657e-06
GC_1_773 b_1 NI_1 NS_773 0 -9.3710917921602539e-08
GC_1_774 b_1 NI_1 NS_774 0 8.7634007816137938e-08
GC_1_775 b_1 NI_1 NS_775 0 -3.3515352414707102e-07
GC_1_776 b_1 NI_1 NS_776 0 2.6717607234162035e-06
GC_1_777 b_1 NI_1 NS_777 0 7.2368311131835902e-07
GC_1_778 b_1 NI_1 NS_778 0 1.5966554211957487e-07
GC_1_779 b_1 NI_1 NS_779 0 3.0760805100985005e-06
GC_1_780 b_1 NI_1 NS_780 0 -2.7795582289444609e-06
GC_1_781 b_1 NI_1 NS_781 0 -1.9947497444675968e-07
GC_1_782 b_1 NI_1 NS_782 0 -1.1674120378683225e-05
GC_1_783 b_1 NI_1 NS_783 0 1.9433167553049848e-06
GC_1_784 b_1 NI_1 NS_784 0 -6.7943780134503402e-07
GC_1_785 b_1 NI_1 NS_785 0 4.3063510962476958e-06
GC_1_786 b_1 NI_1 NS_786 0 -1.7890105539125543e-07
GC_1_787 b_1 NI_1 NS_787 0 1.2121026772739589e-06
GC_1_788 b_1 NI_1 NS_788 0 1.8711460744924319e-06
GC_1_789 b_1 NI_1 NS_789 0 1.6466082677821691e-06
GC_1_790 b_1 NI_1 NS_790 0 -7.9762638984555255e-07
GC_1_791 b_1 NI_1 NS_791 0 5.9154016731862128e-07
GC_1_792 b_1 NI_1 NS_792 0 4.7824094466641006e-07
GC_1_793 b_1 NI_1 NS_793 0 6.8251371407376970e-07
GC_1_794 b_1 NI_1 NS_794 0 -9.6216799664748684e-08
GC_1_795 b_1 NI_1 NS_795 0 2.5753539695459647e-11
GC_1_796 b_1 NI_1 NS_796 0 -9.7279566208026095e-11
GC_1_797 b_1 NI_1 NS_797 0 -1.9600538533723910e-09
GC_1_798 b_1 NI_1 NS_798 0 4.2972470809647094e-09
GC_1_799 b_1 NI_1 NS_799 0 -6.1954754676191002e-05
GC_1_800 b_1 NI_1 NS_800 0 3.1010306822547913e-07
GC_1_801 b_1 NI_1 NS_801 0 1.6335222240018869e-11
GC_1_802 b_1 NI_1 NS_802 0 -8.7577506511756706e-11
GC_1_803 b_1 NI_1 NS_803 0 -1.1069944223560813e-06
GC_1_804 b_1 NI_1 NS_804 0 -1.7649936582932537e-06
GC_1_805 b_1 NI_1 NS_805 0 -1.9904438820119717e-06
GC_1_806 b_1 NI_1 NS_806 0 1.9660066780424967e-06
GC_1_807 b_1 NI_1 NS_807 0 -9.5690915150157322e-06
GC_1_808 b_1 NI_1 NS_808 0 6.6947451932457139e-07
GC_1_809 b_1 NI_1 NS_809 0 -2.0966142220717011e-07
GC_1_810 b_1 NI_1 NS_810 0 3.5162866639762272e-06
GC_1_811 b_1 NI_1 NS_811 0 -2.1093973898424736e-06
GC_1_812 b_1 NI_1 NS_812 0 1.1709183041963191e-05
GC_1_813 b_1 NI_1 NS_813 0 6.8681820516804274e-06
GC_1_814 b_1 NI_1 NS_814 0 1.2213099662179149e-05
GC_1_815 b_1 NI_1 NS_815 0 -2.0257219219094535e-06
GC_1_816 b_1 NI_1 NS_816 0 -2.2559685047026348e-06
GC_1_817 b_1 NI_1 NS_817 0 1.6633461102023282e-06
GC_1_818 b_1 NI_1 NS_818 0 1.0211518333581011e-06
GC_1_819 b_1 NI_1 NS_819 0 7.4141103416645533e-06
GC_1_820 b_1 NI_1 NS_820 0 3.8490357317088379e-05
GC_1_821 b_1 NI_1 NS_821 0 2.2911888642951947e-05
GC_1_822 b_1 NI_1 NS_822 0 -1.2059859990209158e-05
GC_1_823 b_1 NI_1 NS_823 0 8.4232956953175023e-06
GC_1_824 b_1 NI_1 NS_824 0 1.7608848895286437e-06
GC_1_825 b_1 NI_1 NS_825 0 4.7761689953949868e-05
GC_1_826 b_1 NI_1 NS_826 0 -2.5200272790429622e-05
GC_1_827 b_1 NI_1 NS_827 0 -9.4026341041243322e-07
GC_1_828 b_1 NI_1 NS_828 0 -8.0488290835822408e-06
GC_1_829 b_1 NI_1 NS_829 0 3.4272857740911033e-05
GC_1_830 b_1 NI_1 NS_830 0 -7.7701605693957179e-06
GC_1_831 b_1 NI_1 NS_831 0 -3.8695799316197772e-05
GC_1_832 b_1 NI_1 NS_832 0 -5.1800869353347996e-05
GC_1_833 b_1 NI_1 NS_833 0 -4.5827305730402849e-06
GC_1_834 b_1 NI_1 NS_834 0 -4.5466890848144618e-06
GC_1_835 b_1 NI_1 NS_835 0 -3.9429359182428298e-05
GC_1_836 b_1 NI_1 NS_836 0 -1.9669239802882115e-05
GC_1_837 b_1 NI_1 NS_837 0 -4.8828626132733461e-06
GC_1_838 b_1 NI_1 NS_838 0 6.5890060003302604e-06
GC_1_839 b_1 NI_1 NS_839 0 -8.6504783459213907e-06
GC_1_840 b_1 NI_1 NS_840 0 -6.8353885908475828e-07
GC_1_841 b_1 NI_1 NS_841 0 -1.4941086012048991e-05
GC_1_842 b_1 NI_1 NS_842 0 2.4266070306498082e-05
GC_1_843 b_1 NI_1 NS_843 0 1.0803054147931686e-06
GC_1_844 b_1 NI_1 NS_844 0 2.6351381273034198e-06
GC_1_845 b_1 NI_1 NS_845 0 3.0586506151893946e-06
GC_1_846 b_1 NI_1 NS_846 0 1.8296340852320316e-05
GC_1_847 b_1 NI_1 NS_847 0 7.7541133254390095e-06
GC_1_848 b_1 NI_1 NS_848 0 -1.6862230106078220e-06
GC_1_849 b_1 NI_1 NS_849 0 2.9848518227932247e-06
GC_1_850 b_1 NI_1 NS_850 0 -3.4525580208383781e-07
GC_1_851 b_1 NI_1 NS_851 0 7.3238433162841771e-06
GC_1_852 b_1 NI_1 NS_852 0 -4.5245347822424613e-06
GC_1_853 b_1 NI_1 NS_853 0 -8.5067556456567978e-07
GC_1_854 b_1 NI_1 NS_854 0 -5.4051529114568876e-07
GC_1_855 b_1 NI_1 NS_855 0 -1.6424460013381049e-06
GC_1_856 b_1 NI_1 NS_856 0 2.2866377948124080e-07
GC_1_857 b_1 NI_1 NS_857 0 1.5096012088851366e-06
GC_1_858 b_1 NI_1 NS_858 0 1.1390136992916757e-07
GC_1_859 b_1 NI_1 NS_859 0 3.6033424970138488e-06
GC_1_860 b_1 NI_1 NS_860 0 -8.9568557468048640e-07
GC_1_861 b_1 NI_1 NS_861 0 -7.2227980088304346e-08
GC_1_862 b_1 NI_1 NS_862 0 -3.6299696741049643e-07
GC_1_863 b_1 NI_1 NS_863 0 -5.1726377129253901e-07
GC_1_864 b_1 NI_1 NS_864 0 5.5090656374660594e-07
GC_1_865 b_1 NI_1 NS_865 0 2.4011118302071183e-06
GC_1_866 b_1 NI_1 NS_866 0 2.0003029243194903e-07
GC_1_867 b_1 NI_1 NS_867 0 3.3592408410955226e-06
GC_1_868 b_1 NI_1 NS_868 0 -2.8048532574468143e-06
GC_1_869 b_1 NI_1 NS_869 0 -2.6349799223930938e-07
GC_1_870 b_1 NI_1 NS_870 0 -4.2644315289323677e-08
GC_1_871 b_1 NI_1 NS_871 0 7.5184377004930060e-07
GC_1_872 b_1 NI_1 NS_872 0 1.0635517219827041e-06
GC_1_873 b_1 NI_1 NS_873 0 3.5136225677402775e-06
GC_1_874 b_1 NI_1 NS_874 0 7.3949840095078865e-08
GC_1_875 b_1 NI_1 NS_875 0 2.4236023780556246e-06
GC_1_876 b_1 NI_1 NS_876 0 -4.5985037418008654e-06
GC_1_877 b_1 NI_1 NS_877 0 4.5788589767699476e-07
GC_1_878 b_1 NI_1 NS_878 0 1.1656972745797443e-06
GC_1_879 b_1 NI_1 NS_879 0 3.6840101181412070e-06
GC_1_880 b_1 NI_1 NS_880 0 -6.3709724081119493e-07
GC_1_881 b_1 NI_1 NS_881 0 5.5747486870316607e-06
GC_1_882 b_1 NI_1 NS_882 0 -9.4415504632486433e-07
GC_1_883 b_1 NI_1 NS_883 0 -1.6037184436263482e-05
GC_1_884 b_1 NI_1 NS_884 0 -1.0587186233726855e-05
GC_1_885 b_1 NI_1 NS_885 0 9.9725411741341356e-07
GC_1_886 b_1 NI_1 NS_886 0 -7.4331373304826086e-06
GC_1_887 b_1 NI_1 NS_887 0 -6.5807512805485100e-08
GC_1_888 b_1 NI_1 NS_888 0 -1.4868637282113048e-07
GC_1_889 b_1 NI_1 NS_889 0 1.8274069908192643e-06
GC_1_890 b_1 NI_1 NS_890 0 -1.8611960233675400e-06
GC_1_891 b_1 NI_1 NS_891 0 5.4345063871437239e-07
GC_1_892 b_1 NI_1 NS_892 0 -3.3780317887553656e-06
GC_1_893 b_1 NI_1 NS_893 0 3.3863496998023347e-06
GC_1_894 b_1 NI_1 NS_894 0 -1.3093449499728824e-06
GC_1_895 b_1 NI_1 NS_895 0 4.5638629755796472e-06
GC_1_896 b_1 NI_1 NS_896 0 -7.9243940648845461e-07
GC_1_897 b_1 NI_1 NS_897 0 -2.0240625991196655e-07
GC_1_898 b_1 NI_1 NS_898 0 -2.0622476842503352e-07
GC_1_899 b_1 NI_1 NS_899 0 7.0565393377887776e-07
GC_1_900 b_1 NI_1 NS_900 0 1.3955201855801988e-06
GC_1_901 b_1 NI_1 NS_901 0 -7.0553621634654420e-07
GC_1_902 b_1 NI_1 NS_902 0 -1.4723673487529553e-06
GC_1_903 b_1 NI_1 NS_903 0 -6.2774372062465125e-07
GC_1_904 b_1 NI_1 NS_904 0 8.2971958479122943e-07
GC_1_905 b_1 NI_1 NS_905 0 2.2261796398987170e-07
GC_1_906 b_1 NI_1 NS_906 0 6.5380890399128053e-07
GC_1_907 b_1 NI_1 NS_907 0 5.9764946882790926e-07
GC_1_908 b_1 NI_1 NS_908 0 2.1145311927392387e-08
GC_1_909 b_1 NI_1 NS_909 0 1.4034065087524767e-11
GC_1_910 b_1 NI_1 NS_910 0 1.0178152774509873e-12
GC_1_911 b_1 NI_1 NS_911 0 4.3186487448021170e-10
GC_1_912 b_1 NI_1 NS_912 0 1.6518485973502456e-09
GC_1_913 b_1 NI_1 NS_913 0 1.3439637471726088e-05
GC_1_914 b_1 NI_1 NS_914 0 -5.8811639067700940e-08
GC_1_915 b_1 NI_1 NS_915 0 -1.4973651109209550e-11
GC_1_916 b_1 NI_1 NS_916 0 1.3623467904103493e-10
GC_1_917 b_1 NI_1 NS_917 0 3.6109501594648911e-07
GC_1_918 b_1 NI_1 NS_918 0 -1.7974057119663528e-07
GC_1_919 b_1 NI_1 NS_919 0 2.8426232599836713e-07
GC_1_920 b_1 NI_1 NS_920 0 -3.5218292675242587e-07
GC_1_921 b_1 NI_1 NS_921 0 5.0389371682057103e-07
GC_1_922 b_1 NI_1 NS_922 0 -1.4258623372861138e-06
GC_1_923 b_1 NI_1 NS_923 0 -1.1608910122242875e-06
GC_1_924 b_1 NI_1 NS_924 0 -4.7429564324690532e-07
GC_1_925 b_1 NI_1 NS_925 0 -3.4574756200746869e-07
GC_1_926 b_1 NI_1 NS_926 0 -6.3124048701464298e-07
GC_1_927 b_1 NI_1 NS_927 0 -2.5929912189319981e-06
GC_1_928 b_1 NI_1 NS_928 0 -6.5714230444093196e-07
GC_1_929 b_1 NI_1 NS_929 0 7.1939754171038316e-07
GC_1_930 b_1 NI_1 NS_930 0 3.6304573578050671e-07
GC_1_931 b_1 NI_1 NS_931 0 -7.3971065377502899e-07
GC_1_932 b_1 NI_1 NS_932 0 3.6642636660124864e-07
GC_1_933 b_1 NI_1 NS_933 0 -1.0222420098565529e-06
GC_1_934 b_1 NI_1 NS_934 0 5.8988384921640021e-07
GC_1_935 b_1 NI_1 NS_935 0 -4.1600465611074540e-07
GC_1_936 b_1 NI_1 NS_936 0 2.6264354001885697e-07
GC_1_937 b_1 NI_1 NS_937 0 -8.5727219522009608e-07
GC_1_938 b_1 NI_1 NS_938 0 4.4631304796778164e-07
GC_1_939 b_1 NI_1 NS_939 0 1.5253915617366407e-07
GC_1_940 b_1 NI_1 NS_940 0 1.1341010866690232e-06
GC_1_941 b_1 NI_1 NS_941 0 -5.9583494646991186e-07
GC_1_942 b_1 NI_1 NS_942 0 1.1918712108249603e-07
GC_1_943 b_1 NI_1 NS_943 0 -1.9185660306496886e-06
GC_1_944 b_1 NI_1 NS_944 0 1.2734571457808126e-06
GC_1_945 b_1 NI_1 NS_945 0 2.0855889527150006e-06
GC_1_946 b_1 NI_1 NS_946 0 2.8031309403767581e-07
GC_1_947 b_1 NI_1 NS_947 0 -6.8889828372355174e-07
GC_1_948 b_1 NI_1 NS_948 0 1.8836134764747142e-07
GC_1_949 b_1 NI_1 NS_949 0 9.8343422441323734e-07
GC_1_950 b_1 NI_1 NS_950 0 1.7053682618962538e-06
GC_1_951 b_1 NI_1 NS_951 0 -2.2785245808326664e-07
GC_1_952 b_1 NI_1 NS_952 0 -5.8892789080117272e-07
GC_1_953 b_1 NI_1 NS_953 0 -9.2869865517955615e-07
GC_1_954 b_1 NI_1 NS_954 0 4.1600975204450351e-07
GC_1_955 b_1 NI_1 NS_955 0 1.4319962513667778e-06
GC_1_956 b_1 NI_1 NS_956 0 7.1444759469523358e-07
GC_1_957 b_1 NI_1 NS_957 0 -3.3565453908114355e-07
GC_1_958 b_1 NI_1 NS_958 0 -2.2026683155327463e-07
GC_1_959 b_1 NI_1 NS_959 0 -5.3855027329264775e-08
GC_1_960 b_1 NI_1 NS_960 0 1.4317868402542614e-06
GC_1_961 b_1 NI_1 NS_961 0 4.8359320521918686e-07
GC_1_962 b_1 NI_1 NS_962 0 -7.6448870025528634e-07
GC_1_963 b_1 NI_1 NS_963 0 -3.5361624168478885e-07
GC_1_964 b_1 NI_1 NS_964 0 4.2725036325638248e-08
GC_1_965 b_1 NI_1 NS_965 0 3.2259204678572204e-07
GC_1_966 b_1 NI_1 NS_966 0 3.9012931760579889e-07
GC_1_967 b_1 NI_1 NS_967 0 -1.4407256124595710e-07
GC_1_968 b_1 NI_1 NS_968 0 -1.1227657715674928e-08
GC_1_969 b_1 NI_1 NS_969 0 1.4059238094774264e-07
GC_1_970 b_1 NI_1 NS_970 0 1.2582111777466113e-07
GC_1_971 b_1 NI_1 NS_971 0 -1.9006704547673381e-07
GC_1_972 b_1 NI_1 NS_972 0 -6.9875918603160823e-08
GC_1_973 b_1 NI_1 NS_973 0 3.8836561742552791e-08
GC_1_974 b_1 NI_1 NS_974 0 1.9898314876185474e-07
GC_1_975 b_1 NI_1 NS_975 0 -1.1133965462397343e-07
GC_1_976 b_1 NI_1 NS_976 0 9.3792321961629411e-09
GC_1_977 b_1 NI_1 NS_977 0 4.6150751308462358e-08
GC_1_978 b_1 NI_1 NS_978 0 7.8744506028674841e-09
GC_1_979 b_1 NI_1 NS_979 0 -2.9781812341170399e-07
GC_1_980 b_1 NI_1 NS_980 0 -5.3926537220122785e-08
GC_1_981 b_1 NI_1 NS_981 0 -9.1414023886036529e-08
GC_1_982 b_1 NI_1 NS_982 0 6.3222389103798743e-08
GC_1_983 b_1 NI_1 NS_983 0 -2.3130298366943066e-07
GC_1_984 b_1 NI_1 NS_984 0 7.8668917297580387e-08
GC_1_985 b_1 NI_1 NS_985 0 -1.3284201847162289e-07
GC_1_986 b_1 NI_1 NS_986 0 -6.8245269144299801e-08
GC_1_987 b_1 NI_1 NS_987 0 -4.3126488636912351e-07
GC_1_988 b_1 NI_1 NS_988 0 -5.7483646955421057e-08
GC_1_989 b_1 NI_1 NS_989 0 -4.2237555782447771e-07
GC_1_990 b_1 NI_1 NS_990 0 6.4399203327046516e-08
GC_1_991 b_1 NI_1 NS_991 0 -4.4356281923081705e-07
GC_1_992 b_1 NI_1 NS_992 0 1.4475419366082026e-07
GC_1_993 b_1 NI_1 NS_993 0 -5.1284985608864835e-07
GC_1_994 b_1 NI_1 NS_994 0 1.0392226392216272e-07
GC_1_995 b_1 NI_1 NS_995 0 -9.6728434400121380e-07
GC_1_996 b_1 NI_1 NS_996 0 -1.0044880874691566e-07
GC_1_997 b_1 NI_1 NS_997 0 2.6364149412660422e-06
GC_1_998 b_1 NI_1 NS_998 0 3.0037205276037852e-06
GC_1_999 b_1 NI_1 NS_999 0 -6.1832919260756550e-07
GC_1_1000 b_1 NI_1 NS_1000 0 1.0424218587488890e-06
GC_1_1001 b_1 NI_1 NS_1001 0 9.1726242603909509e-09
GC_1_1002 b_1 NI_1 NS_1002 0 2.5504718174527994e-08
GC_1_1003 b_1 NI_1 NS_1003 0 -4.7322550825853925e-07
GC_1_1004 b_1 NI_1 NS_1004 0 8.3082223239234102e-07
GC_1_1005 b_1 NI_1 NS_1005 0 9.3290629157831377e-09
GC_1_1006 b_1 NI_1 NS_1006 0 3.8802042225248755e-07
GC_1_1007 b_1 NI_1 NS_1007 0 -8.7284245953432691e-07
GC_1_1008 b_1 NI_1 NS_1008 0 -7.3755133695306748e-08
GC_1_1009 b_1 NI_1 NS_1009 0 -9.8359148890076430e-07
GC_1_1010 b_1 NI_1 NS_1010 0 -1.8073755521871289e-07
GC_1_1011 b_1 NI_1 NS_1011 0 1.0888652741678155e-07
GC_1_1012 b_1 NI_1 NS_1012 0 -1.4767569188511779e-07
GC_1_1013 b_1 NI_1 NS_1013 0 6.7378564383500656e-08
GC_1_1014 b_1 NI_1 NS_1014 0 1.3250443864128178e-08
GC_1_1015 b_1 NI_1 NS_1015 0 -6.9949612618207880e-08
GC_1_1016 b_1 NI_1 NS_1016 0 1.6113303619873345e-07
GC_1_1017 b_1 NI_1 NS_1017 0 2.9099302997449126e-08
GC_1_1018 b_1 NI_1 NS_1018 0 -4.0233291011964655e-08
GC_1_1019 b_1 NI_1 NS_1019 0 -8.1240446495969615e-08
GC_1_1020 b_1 NI_1 NS_1020 0 1.6008186830063477e-07
GC_1_1021 b_1 NI_1 NS_1021 0 5.6406813854015007e-08
GC_1_1022 b_1 NI_1 NS_1022 0 -1.6261378089410085e-08
GC_1_1023 b_1 NI_1 NS_1023 0 -1.1764356489354584e-11
GC_1_1024 b_1 NI_1 NS_1024 0 5.1442654168098170e-12
GC_1_1025 b_1 NI_1 NS_1025 0 -3.3968959700383056e-10
GC_1_1026 b_1 NI_1 NS_1026 0 -9.7415117878258192e-10
GC_1_1027 b_1 NI_1 NS_1027 0 -2.7508945777840313e-05
GC_1_1028 b_1 NI_1 NS_1028 0 -1.0597555891506710e-08
GC_1_1029 b_1 NI_1 NS_1029 0 1.0238602241791736e-11
GC_1_1030 b_1 NI_1 NS_1030 0 -5.9556851229906745e-11
GC_1_1031 b_1 NI_1 NS_1031 0 -6.3653660479131467e-07
GC_1_1032 b_1 NI_1 NS_1032 0 -1.0748115441599618e-06
GC_1_1033 b_1 NI_1 NS_1033 0 -1.4323563797717064e-06
GC_1_1034 b_1 NI_1 NS_1034 0 2.3248327185690436e-06
GC_1_1035 b_1 NI_1 NS_1035 0 -3.8131152001132450e-06
GC_1_1036 b_1 NI_1 NS_1036 0 2.1795942028616508e-06
GC_1_1037 b_1 NI_1 NS_1037 0 1.9255558595379840e-06
GC_1_1038 b_1 NI_1 NS_1038 0 -2.3466180970278790e-07
GC_1_1039 b_1 NI_1 NS_1039 0 1.4104623108568041e-06
GC_1_1040 b_1 NI_1 NS_1040 0 5.7203933500303993e-06
GC_1_1041 b_1 NI_1 NS_1041 0 3.7051999369784538e-06
GC_1_1042 b_1 NI_1 NS_1042 0 3.2538169624462978e-06
GC_1_1043 b_1 NI_1 NS_1043 0 -1.4742151996485657e-06
GC_1_1044 b_1 NI_1 NS_1044 0 -9.4918334590915179e-07
GC_1_1045 b_1 NI_1 NS_1045 0 9.7320356791067220e-07
GC_1_1046 b_1 NI_1 NS_1046 0 -2.1860338939620328e-06
GC_1_1047 b_1 NI_1 NS_1047 0 6.4354295070577751e-06
GC_1_1048 b_1 NI_1 NS_1048 0 8.5306920824907914e-06
GC_1_1049 b_1 NI_1 NS_1049 0 1.3303316379626706e-06
GC_1_1050 b_1 NI_1 NS_1050 0 -9.3979889626311533e-07
GC_1_1051 b_1 NI_1 NS_1051 0 1.0706358364326949e-06
GC_1_1052 b_1 NI_1 NS_1052 0 -1.9034724561710593e-06
GC_1_1053 b_1 NI_1 NS_1053 0 1.4528584448675629e-05
GC_1_1054 b_1 NI_1 NS_1054 0 -4.1922129564045466e-06
GC_1_1055 b_1 NI_1 NS_1055 0 -2.0125599398982585e-07
GC_1_1056 b_1 NI_1 NS_1056 0 6.7953454945009254e-07
GC_1_1057 b_1 NI_1 NS_1057 0 4.9185731740301409e-06
GC_1_1058 b_1 NI_1 NS_1058 0 -2.1983552566062362e-06
GC_1_1059 b_1 NI_1 NS_1059 0 -7.4680117793014575e-07
GC_1_1060 b_1 NI_1 NS_1060 0 -1.4996612953607686e-05
GC_1_1061 b_1 NI_1 NS_1061 0 -7.6214299920028800e-08
GC_1_1062 b_1 NI_1 NS_1062 0 9.7377272691973808e-07
GC_1_1063 b_1 NI_1 NS_1063 0 -7.9309470845856223e-06
GC_1_1064 b_1 NI_1 NS_1064 0 -8.5785661254947106e-06
GC_1_1065 b_1 NI_1 NS_1065 0 -6.2159288755519954e-07
GC_1_1066 b_1 NI_1 NS_1066 0 -2.1586647565540568e-06
GC_1_1067 b_1 NI_1 NS_1067 0 -8.3452604308228820e-09
GC_1_1068 b_1 NI_1 NS_1068 0 1.2073960960205957e-06
GC_1_1069 b_1 NI_1 NS_1069 0 -7.7192758971547030e-06
GC_1_1070 b_1 NI_1 NS_1070 0 1.9618085179197188e-06
GC_1_1071 b_1 NI_1 NS_1071 0 2.4500474071729283e-07
GC_1_1072 b_1 NI_1 NS_1072 0 -1.6819730219654643e-06
GC_1_1073 b_1 NI_1 NS_1073 0 1.1608984849320913e-06
GC_1_1074 b_1 NI_1 NS_1074 0 3.0678682796291355e-06
GC_1_1075 b_1 NI_1 NS_1075 0 -9.7673335589809980e-07
GC_1_1076 b_1 NI_1 NS_1076 0 2.0311471355105232e-06
GC_1_1077 b_1 NI_1 NS_1077 0 4.5640899366946350e-07
GC_1_1078 b_1 NI_1 NS_1078 0 -1.2309827319597460e-06
GC_1_1079 b_1 NI_1 NS_1079 0 3.2453575023360024e-06
GC_1_1080 b_1 NI_1 NS_1080 0 -8.8264335797575143e-07
GC_1_1081 b_1 NI_1 NS_1081 0 -1.6148480230007144e-07
GC_1_1082 b_1 NI_1 NS_1082 0 5.1316752860974584e-07
GC_1_1083 b_1 NI_1 NS_1083 0 -8.4629646814944673e-07
GC_1_1084 b_1 NI_1 NS_1084 0 -4.1984284719566242e-07
GC_1_1085 b_1 NI_1 NS_1085 0 9.9341967893318775e-07
GC_1_1086 b_1 NI_1 NS_1086 0 -1.2690036826535599e-06
GC_1_1087 b_1 NI_1 NS_1087 0 1.4441137191261077e-06
GC_1_1088 b_1 NI_1 NS_1088 0 -5.7046350091479201e-07
GC_1_1089 b_1 NI_1 NS_1089 0 -3.4131937899494509e-08
GC_1_1090 b_1 NI_1 NS_1090 0 9.6986038599166660e-08
GC_1_1091 b_1 NI_1 NS_1091 0 -5.9769572083376677e-07
GC_1_1092 b_1 NI_1 NS_1092 0 -3.4061585818694250e-07
GC_1_1093 b_1 NI_1 NS_1093 0 9.6764809538452811e-07
GC_1_1094 b_1 NI_1 NS_1094 0 -1.0810604950279121e-06
GC_1_1095 b_1 NI_1 NS_1095 0 1.3955285728348506e-06
GC_1_1096 b_1 NI_1 NS_1096 0 -1.2449209242943618e-06
GC_1_1097 b_1 NI_1 NS_1097 0 1.6144271052288160e-07
GC_1_1098 b_1 NI_1 NS_1098 0 -4.3250410688902463e-08
GC_1_1099 b_1 NI_1 NS_1099 0 -4.8925181850679352e-07
GC_1_1100 b_1 NI_1 NS_1100 0 -5.0362502674259778e-07
GC_1_1101 b_1 NI_1 NS_1101 0 1.0632934744194061e-06
GC_1_1102 b_1 NI_1 NS_1102 0 -8.0455379898035858e-07
GC_1_1103 b_1 NI_1 NS_1103 0 1.2280565465868681e-06
GC_1_1104 b_1 NI_1 NS_1104 0 -2.1206267084338879e-06
GC_1_1105 b_1 NI_1 NS_1105 0 4.9661462222739672e-07
GC_1_1106 b_1 NI_1 NS_1106 0 -2.5357229450726540e-07
GC_1_1107 b_1 NI_1 NS_1107 0 -2.4769332259669225e-07
GC_1_1108 b_1 NI_1 NS_1108 0 -9.1984635275966867e-07
GC_1_1109 b_1 NI_1 NS_1109 0 1.9186317111693919e-06
GC_1_1110 b_1 NI_1 NS_1110 0 -1.0012987231731998e-06
GC_1_1111 b_1 NI_1 NS_1111 0 -8.0998302409131586e-06
GC_1_1112 b_1 NI_1 NS_1112 0 -9.1470443203761767e-07
GC_1_1113 b_1 NI_1 NS_1113 0 -3.1608301656091077e-07
GC_1_1114 b_1 NI_1 NS_1114 0 -3.6264850965385275e-06
GC_1_1115 b_1 NI_1 NS_1115 0 -4.9018272969275402e-08
GC_1_1116 b_1 NI_1 NS_1116 0 -3.3202810865230287e-08
GC_1_1117 b_1 NI_1 NS_1117 0 -1.0294207779192870e-07
GC_1_1118 b_1 NI_1 NS_1118 0 -1.2361446890951357e-06
GC_1_1119 b_1 NI_1 NS_1119 0 -1.0227371138756875e-06
GC_1_1120 b_1 NI_1 NS_1120 0 -6.6783097908288506e-07
GC_1_1121 b_1 NI_1 NS_1121 0 1.4569217195397530e-06
GC_1_1122 b_1 NI_1 NS_1122 0 -7.6152643169874754e-07
GC_1_1123 b_1 NI_1 NS_1123 0 1.9436911686863176e-06
GC_1_1124 b_1 NI_1 NS_1124 0 -1.8722481408128170e-06
GC_1_1125 b_1 NI_1 NS_1125 0 -2.2230806034672048e-07
GC_1_1126 b_1 NI_1 NS_1126 0 3.2515854106087799e-07
GC_1_1127 b_1 NI_1 NS_1127 0 2.1538544104732469e-07
GC_1_1128 b_1 NI_1 NS_1128 0 5.2991274333894390e-07
GC_1_1129 b_1 NI_1 NS_1129 0 -1.0774256416695313e-07
GC_1_1130 b_1 NI_1 NS_1130 0 -2.8383025954633880e-07
GC_1_1131 b_1 NI_1 NS_1131 0 8.1703886129939581e-09
GC_1_1132 b_1 NI_1 NS_1132 0 -9.6163704087025897e-08
GC_1_1133 b_1 NI_1 NS_1133 0 -8.8650245271560952e-08
GC_1_1134 b_1 NI_1 NS_1134 0 4.2005512054087013e-08
GC_1_1135 b_1 NI_1 NS_1135 0 -1.2200395410459134e-07
GC_1_1136 b_1 NI_1 NS_1136 0 -5.3538704787285406e-08
GC_1_1137 b_1 NI_1 NS_1137 0 6.1368284736184142e-12
GC_1_1138 b_1 NI_1 NS_1138 0 -1.6270949392971857e-12
GC_1_1139 b_1 NI_1 NS_1139 0 3.5453293829172617e-10
GC_1_1140 b_1 NI_1 NS_1140 0 6.9229622217861102e-10
GC_1_1141 b_1 NI_1 NS_1141 0 5.5770362728948789e-06
GC_1_1142 b_1 NI_1 NS_1142 0 -6.0661703531600921e-08
GC_1_1143 b_1 NI_1 NS_1143 0 -3.1618767091057349e-11
GC_1_1144 b_1 NI_1 NS_1144 0 4.1808051847100716e-10
GC_1_1145 b_1 NI_1 NS_1145 0 8.7028958035008214e-08
GC_1_1146 b_1 NI_1 NS_1146 0 -7.3629563344290221e-08
GC_1_1147 b_1 NI_1 NS_1147 0 3.8985453958308887e-09
GC_1_1148 b_1 NI_1 NS_1148 0 8.3796046559543148e-08
GC_1_1149 b_1 NI_1 NS_1149 0 6.3125370447641811e-07
GC_1_1150 b_1 NI_1 NS_1150 0 -8.3251284196113968e-07
GC_1_1151 b_1 NI_1 NS_1151 0 -9.1906436841819005e-07
GC_1_1152 b_1 NI_1 NS_1152 0 7.4744386054534755e-08
GC_1_1153 b_1 NI_1 NS_1153 0 5.4098495399094928e-07
GC_1_1154 b_1 NI_1 NS_1154 0 4.5916135147898073e-08
GC_1_1155 b_1 NI_1 NS_1155 0 -1.3830487557748705e-06
GC_1_1156 b_1 NI_1 NS_1156 0 -9.7965322224859343e-07
GC_1_1157 b_1 NI_1 NS_1157 0 3.0645728312439700e-07
GC_1_1158 b_1 NI_1 NS_1158 0 2.0540827079896341e-07
GC_1_1159 b_1 NI_1 NS_1159 0 -5.6263412791054066e-07
GC_1_1160 b_1 NI_1 NS_1160 0 7.1032653167075279e-07
GC_1_1161 b_1 NI_1 NS_1161 0 1.9975475391551389e-06
GC_1_1162 b_1 NI_1 NS_1162 0 -6.2826557627466827e-07
GC_1_1163 b_1 NI_1 NS_1163 0 -2.6418463540165651e-06
GC_1_1164 b_1 NI_1 NS_1164 0 3.8240853108779037e-07
GC_1_1165 b_1 NI_1 NS_1165 0 4.1242829606835476e-08
GC_1_1166 b_1 NI_1 NS_1166 0 1.4294320017982218e-06
GC_1_1167 b_1 NI_1 NS_1167 0 2.3346803223060024e-07
GC_1_1168 b_1 NI_1 NS_1168 0 -1.8326922251824578e-06
GC_1_1169 b_1 NI_1 NS_1169 0 -8.6531545887579878e-07
GC_1_1170 b_1 NI_1 NS_1170 0 1.3761787872450734e-06
GC_1_1171 b_1 NI_1 NS_1171 0 2.2851557004760655e-06
GC_1_1172 b_1 NI_1 NS_1172 0 2.9656045764094944e-06
GC_1_1173 b_1 NI_1 NS_1173 0 -2.0507148844792816e-06
GC_1_1174 b_1 NI_1 NS_1174 0 -3.4923365980902166e-06
GC_1_1175 b_1 NI_1 NS_1175 0 -2.8720388861340612e-07
GC_1_1176 b_1 NI_1 NS_1176 0 1.5382510729207017e-06
GC_1_1177 b_1 NI_1 NS_1177 0 1.7081739067506851e-06
GC_1_1178 b_1 NI_1 NS_1178 0 -1.8792223133430614e-06
GC_1_1179 b_1 NI_1 NS_1179 0 -1.6427703125683742e-06
GC_1_1180 b_1 NI_1 NS_1180 0 1.0311220252027908e-06
GC_1_1181 b_1 NI_1 NS_1181 0 4.2908079030846074e-07
GC_1_1182 b_1 NI_1 NS_1182 0 1.8543841340277980e-06
GC_1_1183 b_1 NI_1 NS_1183 0 2.5930379535056047e-07
GC_1_1184 b_1 NI_1 NS_1184 0 -2.2598887483401473e-06
GC_1_1185 b_1 NI_1 NS_1185 0 -7.4201414028607817e-07
GC_1_1186 b_1 NI_1 NS_1186 0 9.6146792327830604e-07
GC_1_1187 b_1 NI_1 NS_1187 0 2.0833923213325708e-06
GC_1_1188 b_1 NI_1 NS_1188 0 -1.8848775709928121e-08
GC_1_1189 b_1 NI_1 NS_1189 0 -1.8132679243074056e-06
GC_1_1190 b_1 NI_1 NS_1190 0 -3.2980086345427977e-07
GC_1_1191 b_1 NI_1 NS_1191 0 -9.5362714945672343e-08
GC_1_1192 b_1 NI_1 NS_1192 0 7.6458380674783890e-07
GC_1_1193 b_1 NI_1 NS_1193 0 2.1964075308747233e-07
GC_1_1194 b_1 NI_1 NS_1194 0 -5.5285408377651080e-07
GC_1_1195 b_1 NI_1 NS_1195 0 -2.4027915193345908e-07
GC_1_1196 b_1 NI_1 NS_1196 0 4.2925615253186780e-07
GC_1_1197 b_1 NI_1 NS_1197 0 1.0687531703890824e-07
GC_1_1198 b_1 NI_1 NS_1198 0 -2.2410637597473001e-07
GC_1_1199 b_1 NI_1 NS_1199 0 -4.5515340082244786e-07
GC_1_1200 b_1 NI_1 NS_1200 0 3.0526517919262870e-07
GC_1_1201 b_1 NI_1 NS_1201 0 2.0651295333710467e-07
GC_1_1202 b_1 NI_1 NS_1202 0 1.6780208929117503e-08
GC_1_1203 b_1 NI_1 NS_1203 0 -1.4742983152109624e-07
GC_1_1204 b_1 NI_1 NS_1204 0 1.9351597761662741e-07
GC_1_1205 b_1 NI_1 NS_1205 0 2.4897442194225535e-08
GC_1_1206 b_1 NI_1 NS_1206 0 -1.4136273492701904e-07
GC_1_1207 b_1 NI_1 NS_1207 0 -3.4516562564858358e-07
GC_1_1208 b_1 NI_1 NS_1208 0 2.7933039674541865e-07
GC_1_1209 b_1 NI_1 NS_1209 0 1.1041828230171893e-07
GC_1_1210 b_1 NI_1 NS_1210 0 -2.3166559256339420e-08
GC_1_1211 b_1 NI_1 NS_1211 0 -1.1146422843207088e-07
GC_1_1212 b_1 NI_1 NS_1212 0 2.2575710090691902e-07
GC_1_1213 b_1 NI_1 NS_1213 0 -1.8955337482132207e-08
GC_1_1214 b_1 NI_1 NS_1214 0 -1.6880170076561466e-07
GC_1_1215 b_1 NI_1 NS_1215 0 -2.8643069097839047e-07
GC_1_1216 b_1 NI_1 NS_1216 0 1.8674637275506719e-07
GC_1_1217 b_1 NI_1 NS_1217 0 -1.1166126888900960e-07
GC_1_1218 b_1 NI_1 NS_1218 0 -5.9934119337634844e-08
GC_1_1219 b_1 NI_1 NS_1219 0 -1.7481578475826626e-07
GC_1_1220 b_1 NI_1 NS_1220 0 2.0346164717057045e-07
GC_1_1221 b_1 NI_1 NS_1221 0 -2.9232296964884173e-07
GC_1_1222 b_1 NI_1 NS_1222 0 -3.9929749188308510e-08
GC_1_1223 b_1 NI_1 NS_1223 0 -4.9681227135799169e-07
GC_1_1224 b_1 NI_1 NS_1224 0 5.7772029539622710e-08
GC_1_1225 b_1 NI_1 NS_1225 0 2.7719568818716643e-06
GC_1_1226 b_1 NI_1 NS_1226 0 4.3304257297998862e-07
GC_1_1227 b_1 NI_1 NS_1227 0 -3.2409812184842252e-07
GC_1_1228 b_1 NI_1 NS_1228 0 6.7640696814948879e-07
GC_1_1229 b_1 NI_1 NS_1229 0 1.2398649645977117e-08
GC_1_1230 b_1 NI_1 NS_1230 0 1.2812502572687916e-08
GC_1_1231 b_1 NI_1 NS_1231 0 -6.7518772978340081e-09
GC_1_1232 b_1 NI_1 NS_1232 0 4.6496685133454310e-07
GC_1_1233 b_1 NI_1 NS_1233 0 -1.2602595943226098e-07
GC_1_1234 b_1 NI_1 NS_1234 0 2.6654242296891681e-07
GC_1_1235 b_1 NI_1 NS_1235 0 -4.8112943550968628e-07
GC_1_1236 b_1 NI_1 NS_1236 0 9.8550137207964495e-08
GC_1_1237 b_1 NI_1 NS_1237 0 -9.4591670889202899e-07
GC_1_1238 b_1 NI_1 NS_1238 0 4.8604653450201114e-07
GC_1_1239 b_1 NI_1 NS_1239 0 -1.8710246440725365e-07
GC_1_1240 b_1 NI_1 NS_1240 0 -7.9281357130715413e-08
GC_1_1241 b_1 NI_1 NS_1241 0 1.6412110459388455e-08
GC_1_1242 b_1 NI_1 NS_1242 0 -1.4793960472081853e-07
GC_1_1243 b_1 NI_1 NS_1243 0 8.6145547433575407e-08
GC_1_1244 b_1 NI_1 NS_1244 0 1.0231862764690105e-07
GC_1_1245 b_1 NI_1 NS_1245 0 -1.1791419285479237e-07
GC_1_1246 b_1 NI_1 NS_1246 0 -1.5795355077707331e-07
GC_1_1247 b_1 NI_1 NS_1247 0 -7.0288333582887699e-08
GC_1_1248 b_1 NI_1 NS_1248 0 8.1122645825886532e-08
GC_1_1249 b_1 NI_1 NS_1249 0 -4.4816947122412782e-10
GC_1_1250 b_1 NI_1 NS_1250 0 -3.7626805442986324e-08
GC_1_1251 b_1 NI_1 NS_1251 0 -8.0397622846783845e-12
GC_1_1252 b_1 NI_1 NS_1252 0 7.1579129726139311e-12
GC_1_1253 b_1 NI_1 NS_1253 0 9.6679308890493451e-10
GC_1_1254 b_1 NI_1 NS_1254 0 -3.3561978645393174e-10
GC_1_1255 b_1 NI_1 NS_1255 0 -1.2624774919759490e-05
GC_1_1256 b_1 NI_1 NS_1256 0 1.6614498917458670e-08
GC_1_1257 b_1 NI_1 NS_1257 0 2.1156791733859395e-11
GC_1_1258 b_1 NI_1 NS_1258 0 -3.0722763271680945e-10
GC_1_1259 b_1 NI_1 NS_1259 0 -3.4980938929532835e-07
GC_1_1260 b_1 NI_1 NS_1260 0 -9.9927065582844404e-07
GC_1_1261 b_1 NI_1 NS_1261 0 -9.3440149864286681e-07
GC_1_1262 b_1 NI_1 NS_1262 0 1.7812981889050790e-06
GC_1_1263 b_1 NI_1 NS_1263 0 -3.3145705061615105e-06
GC_1_1264 b_1 NI_1 NS_1264 0 8.1232046624510609e-07
GC_1_1265 b_1 NI_1 NS_1265 0 9.4647152482036973e-07
GC_1_1266 b_1 NI_1 NS_1266 0 -2.3710222534920450e-07
GC_1_1267 b_1 NI_1 NS_1267 0 5.4137163190697463e-07
GC_1_1268 b_1 NI_1 NS_1268 0 4.5112145834752356e-06
GC_1_1269 b_1 NI_1 NS_1269 0 1.6155112262548026e-06
GC_1_1270 b_1 NI_1 NS_1270 0 3.0375444094245314e-06
GC_1_1271 b_1 NI_1 NS_1271 0 -8.7084008683706689e-07
GC_1_1272 b_1 NI_1 NS_1272 0 -5.9646298363486803e-07
GC_1_1273 b_1 NI_1 NS_1273 0 4.7061514660394062e-07
GC_1_1274 b_1 NI_1 NS_1274 0 -1.1586884354833402e-06
GC_1_1275 b_1 NI_1 NS_1275 0 2.8699782659822701e-06
GC_1_1276 b_1 NI_1 NS_1276 0 1.0313952861481981e-05
GC_1_1277 b_1 NI_1 NS_1277 0 4.5228581560728192e-06
GC_1_1278 b_1 NI_1 NS_1278 0 -7.5297937495991424e-07
GC_1_1279 b_1 NI_1 NS_1279 0 1.6523542132837095e-06
GC_1_1280 b_1 NI_1 NS_1280 0 -4.2608573490463162e-07
GC_1_1281 b_1 NI_1 NS_1281 0 1.6706021651728678e-05
GC_1_1282 b_1 NI_1 NS_1282 0 -4.4199325781548106e-06
GC_1_1283 b_1 NI_1 NS_1283 0 2.2368611257723632e-07
GC_1_1284 b_1 NI_1 NS_1284 0 -1.0416399298374731e-06
GC_1_1285 b_1 NI_1 NS_1285 0 9.3469223821362583e-06
GC_1_1286 b_1 NI_1 NS_1286 0 -7.0992943368862869e-07
GC_1_1287 b_1 NI_1 NS_1287 0 -5.5727601009676410e-06
GC_1_1288 b_1 NI_1 NS_1288 0 -1.9751240852650745e-05
GC_1_1289 b_1 NI_1 NS_1289 0 -6.0103078718306195e-07
GC_1_1290 b_1 NI_1 NS_1290 0 -8.9964383671354777e-07
GC_1_1291 b_1 NI_1 NS_1291 0 -1.1428658574247873e-05
GC_1_1292 b_1 NI_1 NS_1292 0 -1.0988290649535122e-05
GC_1_1293 b_1 NI_1 NS_1293 0 -2.2555822882514152e-06
GC_1_1294 b_1 NI_1 NS_1294 0 2.5926792138208369e-07
GC_1_1295 b_1 NI_1 NS_1295 0 -1.9214226527668540e-06
GC_1_1296 b_1 NI_1 NS_1296 0 -7.8273434043320070e-07
GC_1_1297 b_1 NI_1 NS_1297 0 -9.6694382758991426e-06
GC_1_1298 b_1 NI_1 NS_1298 0 5.8238608399825813e-06
GC_1_1299 b_1 NI_1 NS_1299 0 -3.0070379455774259e-07
GC_1_1300 b_1 NI_1 NS_1300 0 1.6096116546284328e-07
GC_1_1301 b_1 NI_1 NS_1301 0 -1.6035958833777506e-06
GC_1_1302 b_1 NI_1 NS_1302 0 5.7948443022033633e-06
GC_1_1303 b_1 NI_1 NS_1303 0 2.0456008827918957e-06
GC_1_1304 b_1 NI_1 NS_1304 0 1.9760439166860847e-06
GC_1_1305 b_1 NI_1 NS_1305 0 6.0757046210884015e-07
GC_1_1306 b_1 NI_1 NS_1306 0 -8.9292419185837336e-08
GC_1_1307 b_1 NI_1 NS_1307 0 3.3238970100988191e-06
GC_1_1308 b_1 NI_1 NS_1308 0 -4.3020817764518419e-07
GC_1_1309 b_1 NI_1 NS_1309 0 -5.1720331664259144e-08
GC_1_1310 b_1 NI_1 NS_1310 0 3.3333385138378275e-08
GC_1_1311 b_1 NI_1 NS_1311 0 -8.0692554517263397e-07
GC_1_1312 b_1 NI_1 NS_1312 0 -2.3783518975845425e-07
GC_1_1313 b_1 NI_1 NS_1313 0 3.8090018835305686e-07
GC_1_1314 b_1 NI_1 NS_1314 0 -5.1763393886864828e-07
GC_1_1315 b_1 NI_1 NS_1315 0 1.1838650259703670e-06
GC_1_1316 b_1 NI_1 NS_1316 0 -3.2905040350187232e-08
GC_1_1317 b_1 NI_1 NS_1317 0 2.3909378165552666e-08
GC_1_1318 b_1 NI_1 NS_1318 0 4.9139863410260330e-08
GC_1_1319 b_1 NI_1 NS_1319 0 -5.6752164826798390e-07
GC_1_1320 b_1 NI_1 NS_1320 0 -5.4511895121540461e-08
GC_1_1321 b_1 NI_1 NS_1321 0 4.9423749436177013e-07
GC_1_1322 b_1 NI_1 NS_1322 0 -5.0922585893968493e-07
GC_1_1323 b_1 NI_1 NS_1323 0 1.1633692376335517e-06
GC_1_1324 b_1 NI_1 NS_1324 0 -6.8915176154383945e-07
GC_1_1325 b_1 NI_1 NS_1325 0 5.6878914422873829e-08
GC_1_1326 b_1 NI_1 NS_1326 0 -7.3032406744999975e-12
GC_1_1327 b_1 NI_1 NS_1327 0 -5.7572917232830658e-07
GC_1_1328 b_1 NI_1 NS_1328 0 -6.5420228901857981e-08
GC_1_1329 b_1 NI_1 NS_1329 0 6.3198136249246717e-07
GC_1_1330 b_1 NI_1 NS_1330 0 -5.0017555707981110e-07
GC_1_1331 b_1 NI_1 NS_1331 0 8.4908653166779729e-07
GC_1_1332 b_1 NI_1 NS_1332 0 -1.3993603292584332e-06
GC_1_1333 b_1 NI_1 NS_1333 0 1.0851464920796851e-07
GC_1_1334 b_1 NI_1 NS_1334 0 -6.0235381620259452e-08
GC_1_1335 b_1 NI_1 NS_1335 0 -3.9931200571413556e-07
GC_1_1336 b_1 NI_1 NS_1336 0 -2.0520897951652222e-07
GC_1_1337 b_1 NI_1 NS_1337 0 1.1352398591482740e-06
GC_1_1338 b_1 NI_1 NS_1338 0 -8.8090186619465855e-07
GC_1_1339 b_1 NI_1 NS_1339 0 -4.1524217160468467e-06
GC_1_1340 b_1 NI_1 NS_1340 0 6.0076417930567948e-07
GC_1_1341 b_1 NI_1 NS_1341 0 -5.6337449373852473e-07
GC_1_1342 b_1 NI_1 NS_1342 0 -1.9350557577504503e-06
GC_1_1343 b_1 NI_1 NS_1343 0 -2.9192658064150436e-08
GC_1_1344 b_1 NI_1 NS_1344 0 -9.6995575247984301e-09
GC_1_1345 b_1 NI_1 NS_1345 0 -3.5869169467994532e-07
GC_1_1346 b_1 NI_1 NS_1346 0 -2.9247555264357250e-07
GC_1_1347 b_1 NI_1 NS_1347 0 -4.7717727604781798e-07
GC_1_1348 b_1 NI_1 NS_1348 0 -1.7395719069175722e-07
GC_1_1349 b_1 NI_1 NS_1349 0 8.5945807319976419e-07
GC_1_1350 b_1 NI_1 NS_1350 0 -7.5659574809881944e-07
GC_1_1351 b_1 NI_1 NS_1351 0 6.0934982376939002e-07
GC_1_1352 b_1 NI_1 NS_1352 0 -1.0778282438870586e-06
GC_1_1353 b_1 NI_1 NS_1353 0 9.0828870702236679e-08
GC_1_1354 b_1 NI_1 NS_1354 0 1.4507020224151880e-07
GC_1_1355 b_1 NI_1 NS_1355 0 1.5780207422438009e-07
GC_1_1356 b_1 NI_1 NS_1356 0 4.4524739614981855e-07
GC_1_1357 b_1 NI_1 NS_1357 0 2.3130304379866481e-08
GC_1_1358 b_1 NI_1 NS_1358 0 -1.6507878054137226e-07
GC_1_1359 b_1 NI_1 NS_1359 0 -3.7596769907357745e-08
GC_1_1360 b_1 NI_1 NS_1360 0 -1.2378262361303168e-07
GC_1_1361 b_1 NI_1 NS_1361 0 -8.6474604705123461e-08
GC_1_1362 b_1 NI_1 NS_1362 0 1.2324407763772904e-07
GC_1_1363 b_1 NI_1 NS_1363 0 -9.0133036593611958e-09
GC_1_1364 b_1 NI_1 NS_1364 0 -3.7917691596676893e-09
GC_1_1365 b_1 NI_1 NS_1365 0 2.2956463436555228e-12
GC_1_1366 b_1 NI_1 NS_1366 0 -3.3975543871863607e-12
GC_1_1367 b_1 NI_1 NS_1367 0 -7.3117264020247804e-10
GC_1_1368 b_1 NI_1 NS_1368 0 -8.2654847221324910e-11
GD_1_1 b_1 NI_1 NA_1 0 -8.8592633367533483e-03
GD_1_2 b_1 NI_1 NA_2 0 -4.2259674030547542e-03
GD_1_3 b_1 NI_1 NA_3 0 1.3004902192097227e-02
GD_1_4 b_1 NI_1 NA_4 0 5.9084065482663012e-04
GD_1_5 b_1 NI_1 NA_5 0 5.6585682801942395e-06
GD_1_6 b_1 NI_1 NA_6 0 2.4210595786006727e-06
GD_1_7 b_1 NI_1 NA_7 0 -3.6554696157799598e-06
GD_1_8 b_1 NI_1 NA_8 0 1.0039627760117894e-05
GD_1_9 b_1 NI_1 NA_9 0 -1.8680218656177269e-06
GD_1_10 b_1 NI_1 NA_10 0 5.6280493176681220e-06
GD_1_11 b_1 NI_1 NA_11 0 -6.4899006105884963e-07
GD_1_12 b_1 NI_1 NA_12 0 3.5859754888125554e-06
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 1.8230039061899118e-02
GC_2_2 b_2 NI_2 NS_2 0 6.7517748588041661e-03
GC_2_3 b_2 NI_2 NS_3 0 4.8176235412146930e-07
GC_2_4 b_2 NI_2 NS_4 0 1.4329617485962278e-06
GC_2_5 b_2 NI_2 NS_5 0 6.0825248487266885e-03
GC_2_6 b_2 NI_2 NS_6 0 1.8254985159630479e-03
GC_2_7 b_2 NI_2 NS_7 0 -6.0663489091265961e-03
GC_2_8 b_2 NI_2 NS_8 0 -6.4127978922103165e-04
GC_2_9 b_2 NI_2 NS_9 0 7.3353526262885781e-03
GC_2_10 b_2 NI_2 NS_10 0 -1.2858434177101818e-02
GC_2_11 b_2 NI_2 NS_11 0 8.4355295081309355e-03
GC_2_12 b_2 NI_2 NS_12 0 -2.1165104320126709e-04
GC_2_13 b_2 NI_2 NS_13 0 -9.6680534989310001e-03
GC_2_14 b_2 NI_2 NS_14 0 2.5854036631835406e-03
GC_2_15 b_2 NI_2 NS_15 0 -8.8080269224896299e-03
GC_2_16 b_2 NI_2 NS_16 0 -2.4395023146212697e-02
GC_2_17 b_2 NI_2 NS_17 0 -8.6848627101713735e-04
GC_2_18 b_2 NI_2 NS_18 0 4.1759068882033156e-03
GC_2_19 b_2 NI_2 NS_19 0 7.1854996224088932e-03
GC_2_20 b_2 NI_2 NS_20 0 -9.9751747952556060e-04
GC_2_21 b_2 NI_2 NS_21 0 -2.5219867220426000e-02
GC_2_22 b_2 NI_2 NS_22 0 4.8140735355620386e-03
GC_2_23 b_2 NI_2 NS_23 0 -1.9618673441073656e-02
GC_2_24 b_2 NI_2 NS_24 0 8.5360791904722964e-04
GC_2_25 b_2 NI_2 NS_25 0 1.0773125157927606e-02
GC_2_26 b_2 NI_2 NS_26 0 -2.7351328804441585e-03
GC_2_27 b_2 NI_2 NS_27 0 -4.8272985082159128e-03
GC_2_28 b_2 NI_2 NS_28 0 4.5019507995646163e-02
GC_2_29 b_2 NI_2 NS_29 0 -1.2641959584080568e-02
GC_2_30 b_2 NI_2 NS_30 0 -3.2181137565287277e-04
GC_2_31 b_2 NI_2 NS_31 0 1.5975179694205862e-02
GC_2_32 b_2 NI_2 NS_32 0 -3.9761003575212416e-03
GC_2_33 b_2 NI_2 NS_33 0 3.2145894844490770e-02
GC_2_34 b_2 NI_2 NS_34 0 1.8555664776058883e-02
GC_2_35 b_2 NI_2 NS_35 0 -1.2595027817914458e-02
GC_2_36 b_2 NI_2 NS_36 0 1.1573529122424000e-04
GC_2_37 b_2 NI_2 NS_37 0 1.7251990989723499e-02
GC_2_38 b_2 NI_2 NS_38 0 -3.5175740088199958e-02
GC_2_39 b_2 NI_2 NS_39 0 1.3984105281888428e-02
GC_2_40 b_2 NI_2 NS_40 0 4.8235505429299729e-03
GC_2_41 b_2 NI_2 NS_41 0 -1.4410964269810112e-02
GC_2_42 b_2 NI_2 NS_42 0 1.9249748290731244e-04
GC_2_43 b_2 NI_2 NS_43 0 -2.0124073649327872e-02
GC_2_44 b_2 NI_2 NS_44 0 -3.0196986780034719e-02
GC_2_45 b_2 NI_2 NS_45 0 1.0516088412861276e-02
GC_2_46 b_2 NI_2 NS_46 0 3.6210340231066056e-03
GC_2_47 b_2 NI_2 NS_47 0 -2.6839303910668966e-02
GC_2_48 b_2 NI_2 NS_48 0 1.1127446656882185e-02
GC_2_49 b_2 NI_2 NS_49 0 -1.4106901817026965e-02
GC_2_50 b_2 NI_2 NS_50 0 -2.5293090443954357e-03
GC_2_51 b_2 NI_2 NS_51 0 7.5511422011574937e-03
GC_2_52 b_2 NI_2 NS_52 0 1.6110587602041755e-03
GC_2_53 b_2 NI_2 NS_53 0 -8.7786011049233875e-04
GC_2_54 b_2 NI_2 NS_54 0 2.4406497512945189e-02
GC_2_55 b_2 NI_2 NS_55 0 -7.6159627408168519e-03
GC_2_56 b_2 NI_2 NS_56 0 2.7281640949137305e-04
GC_2_57 b_2 NI_2 NS_57 0 -5.5397748036337916e-04
GC_2_58 b_2 NI_2 NS_58 0 -5.5347504684661649e-03
GC_2_59 b_2 NI_2 NS_59 0 8.2549319693739926e-03
GC_2_60 b_2 NI_2 NS_60 0 7.0291735461128612e-03
GC_2_61 b_2 NI_2 NS_61 0 -7.2658614181994618e-04
GC_2_62 b_2 NI_2 NS_62 0 1.2096258797943465e-02
GC_2_63 b_2 NI_2 NS_63 0 -5.1449971133258592e-03
GC_2_64 b_2 NI_2 NS_64 0 -1.3736254715227184e-04
GC_2_65 b_2 NI_2 NS_65 0 -1.8277901983705202e-03
GC_2_66 b_2 NI_2 NS_66 0 -5.1663735910053221e-03
GC_2_67 b_2 NI_2 NS_67 0 9.2805974918669671e-03
GC_2_68 b_2 NI_2 NS_68 0 5.4201891255769071e-03
GC_2_69 b_2 NI_2 NS_69 0 3.5139830703434082e-03
GC_2_70 b_2 NI_2 NS_70 0 1.1696931131325933e-02
GC_2_71 b_2 NI_2 NS_71 0 -6.1352297753534341e-03
GC_2_72 b_2 NI_2 NS_72 0 1.4322953320917383e-03
GC_2_73 b_2 NI_2 NS_73 0 -2.8179573100192527e-03
GC_2_74 b_2 NI_2 NS_74 0 -7.3386810051825069e-03
GC_2_75 b_2 NI_2 NS_75 0 9.9491352723307096e-03
GC_2_76 b_2 NI_2 NS_76 0 3.3701742004156000e-03
GC_2_77 b_2 NI_2 NS_77 0 8.1727144660940863e-03
GC_2_78 b_2 NI_2 NS_78 0 1.0256376601752959e-02
GC_2_79 b_2 NI_2 NS_79 0 -6.9843353386215773e-03
GC_2_80 b_2 NI_2 NS_80 0 2.9455291783147390e-03
GC_2_81 b_2 NI_2 NS_81 0 -5.6339165862952702e-03
GC_2_82 b_2 NI_2 NS_82 0 -8.0804392929484017e-03
GC_2_83 b_2 NI_2 NS_83 0 9.8431188819430165e-03
GC_2_84 b_2 NI_2 NS_84 0 5.5956605507856069e-04
GC_2_85 b_2 NI_2 NS_85 0 -1.0789780644149208e-02
GC_2_86 b_2 NI_2 NS_86 0 1.2190659140759598e-02
GC_2_87 b_2 NI_2 NS_87 0 9.6746764539523480e-03
GC_2_88 b_2 NI_2 NS_88 0 5.0624616423630584e-03
GC_2_89 b_2 NI_2 NS_89 0 -1.9019902556747380e-05
GC_2_90 b_2 NI_2 NS_90 0 3.1757032473048231e-05
GC_2_91 b_2 NI_2 NS_91 0 -7.1157513096728325e-03
GC_2_92 b_2 NI_2 NS_92 0 4.4966089266802308e-03
GC_2_93 b_2 NI_2 NS_93 0 -7.6591177680452116e-03
GC_2_94 b_2 NI_2 NS_94 0 -5.3141664629227352e-03
GC_2_95 b_2 NI_2 NS_95 0 9.4991996307270052e-03
GC_2_96 b_2 NI_2 NS_96 0 -1.7114390495441764e-03
GC_2_97 b_2 NI_2 NS_97 0 1.2463051630688823e-02
GC_2_98 b_2 NI_2 NS_98 0 -1.3561359797575044e-03
GC_2_99 b_2 NI_2 NS_99 0 -5.0733906037891321e-03
GC_2_100 b_2 NI_2 NS_100 0 -2.7549348882787046e-03
GC_2_101 b_2 NI_2 NS_101 0 -2.2333264439641873e-03
GC_2_102 b_2 NI_2 NS_102 0 6.5928662730748468e-03
GC_2_103 b_2 NI_2 NS_103 0 8.9636634146078326e-03
GC_2_104 b_2 NI_2 NS_104 0 1.2895392433878640e-04
GC_2_105 b_2 NI_2 NS_105 0 1.2489929382331589e-02
GC_2_106 b_2 NI_2 NS_106 0 1.7708857219725759e-03
GC_2_107 b_2 NI_2 NS_107 0 -5.3741340359903609e-03
GC_2_108 b_2 NI_2 NS_108 0 4.1561546109872838e-03
GC_2_109 b_2 NI_2 NS_109 0 -1.8427479441608344e-03
GC_2_110 b_2 NI_2 NS_110 0 -5.6872754356419300e-03
GC_2_111 b_2 NI_2 NS_111 0 2.0875928785291602e-07
GC_2_112 b_2 NI_2 NS_112 0 -2.4399578241098077e-07
GC_2_113 b_2 NI_2 NS_113 0 -1.1437013034868182e-05
GC_2_114 b_2 NI_2 NS_114 0 1.8295056790630626e-05
GC_2_115 b_2 NI_2 NS_115 0 -1.3077575657918679e-02
GC_2_116 b_2 NI_2 NS_116 0 1.3851810838321856e-03
GC_2_117 b_2 NI_2 NS_117 0 -2.6206809722675156e-07
GC_2_118 b_2 NI_2 NS_118 0 -3.7495376870487568e-06
GC_2_119 b_2 NI_2 NS_119 0 -2.7819412649494803e-04
GC_2_120 b_2 NI_2 NS_120 0 4.6297784662617064e-04
GC_2_121 b_2 NI_2 NS_121 0 1.3195316947856943e-03
GC_2_122 b_2 NI_2 NS_122 0 5.4935810838243357e-04
GC_2_123 b_2 NI_2 NS_123 0 -2.7628707830373894e-03
GC_2_124 b_2 NI_2 NS_124 0 -8.1702960577355950e-04
GC_2_125 b_2 NI_2 NS_125 0 3.5326194217725386e-03
GC_2_126 b_2 NI_2 NS_126 0 2.5338003494739798e-03
GC_2_127 b_2 NI_2 NS_127 0 1.1824215167199710e-03
GC_2_128 b_2 NI_2 NS_128 0 -4.1997919360099636e-03
GC_2_129 b_2 NI_2 NS_129 0 -1.7498497484614815e-03
GC_2_130 b_2 NI_2 NS_130 0 2.6968875331504728e-03
GC_2_131 b_2 NI_2 NS_131 0 -3.1387253129655729e-04
GC_2_132 b_2 NI_2 NS_132 0 -1.8984355421809357e-04
GC_2_133 b_2 NI_2 NS_133 0 3.9674908773075310e-03
GC_2_134 b_2 NI_2 NS_134 0 2.9857924899183446e-04
GC_2_135 b_2 NI_2 NS_135 0 -7.4413898752046107e-03
GC_2_136 b_2 NI_2 NS_136 0 -1.3618331607425224e-02
GC_2_137 b_2 NI_2 NS_137 0 4.4052529700029704e-03
GC_2_138 b_2 NI_2 NS_138 0 1.3511450566460931e-02
GC_2_139 b_2 NI_2 NS_139 0 6.7110134907057556e-03
GC_2_140 b_2 NI_2 NS_140 0 -3.9862641894750596e-03
GC_2_141 b_2 NI_2 NS_141 0 -1.3390053159840857e-02
GC_2_142 b_2 NI_2 NS_142 0 6.9023312150232735e-04
GC_2_143 b_2 NI_2 NS_143 0 7.8426027215753348e-03
GC_2_144 b_2 NI_2 NS_144 0 1.8947657846531943e-03
GC_2_145 b_2 NI_2 NS_145 0 1.0544114974704123e-02
GC_2_146 b_2 NI_2 NS_146 0 -1.9595452275827405e-02
GC_2_147 b_2 NI_2 NS_147 0 -1.7809618055608809e-02
GC_2_148 b_2 NI_2 NS_148 0 1.9141982754548405e-02
GC_2_149 b_2 NI_2 NS_149 0 7.6787743766728632e-03
GC_2_150 b_2 NI_2 NS_150 0 -1.4142911445391127e-03
GC_2_151 b_2 NI_2 NS_151 0 -1.5647917037332763e-02
GC_2_152 b_2 NI_2 NS_152 0 -4.7614903566545602e-03
GC_2_153 b_2 NI_2 NS_153 0 8.0618568963733775e-03
GC_2_154 b_2 NI_2 NS_154 0 7.2869895044586014e-03
GC_2_155 b_2 NI_2 NS_155 0 8.1170040783417000e-03
GC_2_156 b_2 NI_2 NS_156 0 -5.9990842974447268e-03
GC_2_157 b_2 NI_2 NS_157 0 -1.3980589235182254e-02
GC_2_158 b_2 NI_2 NS_158 0 4.5682738336424696e-03
GC_2_159 b_2 NI_2 NS_159 0 6.2307821482156427e-03
GC_2_160 b_2 NI_2 NS_160 0 2.4081616521147032e-03
GC_2_161 b_2 NI_2 NS_161 0 -6.2859259532714257e-03
GC_2_162 b_2 NI_2 NS_162 0 -1.1107051215957600e-02
GC_2_163 b_2 NI_2 NS_163 0 2.1280730654042379e-03
GC_2_164 b_2 NI_2 NS_164 0 1.1947396614296037e-02
GC_2_165 b_2 NI_2 NS_165 0 4.2092181380888397e-03
GC_2_166 b_2 NI_2 NS_166 0 -1.1609525185980215e-03
GC_2_167 b_2 NI_2 NS_167 0 -4.9313047700363872e-03
GC_2_168 b_2 NI_2 NS_168 0 1.0532426449720680e-03
GC_2_169 b_2 NI_2 NS_169 0 3.0238805602796071e-03
GC_2_170 b_2 NI_2 NS_170 0 6.9985668908834455e-04
GC_2_171 b_2 NI_2 NS_171 0 -2.2205265102970529e-03
GC_2_172 b_2 NI_2 NS_172 0 4.9428523590564378e-04
GC_2_173 b_2 NI_2 NS_173 0 3.0655101856460502e-03
GC_2_174 b_2 NI_2 NS_174 0 2.3037295683004588e-03
GC_2_175 b_2 NI_2 NS_175 0 -1.5339095928920683e-03
GC_2_176 b_2 NI_2 NS_176 0 -6.6977523797219041e-04
GC_2_177 b_2 NI_2 NS_177 0 1.8873377871802353e-03
GC_2_178 b_2 NI_2 NS_178 0 6.8441611640691869e-04
GC_2_179 b_2 NI_2 NS_179 0 -1.5620994940060511e-03
GC_2_180 b_2 NI_2 NS_180 0 1.2263485505598489e-03
GC_2_181 b_2 NI_2 NS_181 0 3.9751899193924134e-03
GC_2_182 b_2 NI_2 NS_182 0 1.4060873640020085e-03
GC_2_183 b_2 NI_2 NS_183 0 -1.5528113430281333e-03
GC_2_184 b_2 NI_2 NS_184 0 7.4659511701641120e-05
GC_2_185 b_2 NI_2 NS_185 0 2.8290376322304173e-03
GC_2_186 b_2 NI_2 NS_186 0 -6.8617020675040699e-04
GC_2_187 b_2 NI_2 NS_187 0 -1.8781842572414289e-03
GC_2_188 b_2 NI_2 NS_188 0 2.0100714537215946e-03
GC_2_189 b_2 NI_2 NS_189 0 4.9079326878410335e-03
GC_2_190 b_2 NI_2 NS_190 0 -1.8215468359191909e-04
GC_2_191 b_2 NI_2 NS_191 0 -1.6564605115377425e-03
GC_2_192 b_2 NI_2 NS_192 0 9.3019010342163780e-04
GC_2_193 b_2 NI_2 NS_193 0 3.0643001553729990e-03
GC_2_194 b_2 NI_2 NS_194 0 -2.8465122060995188e-03
GC_2_195 b_2 NI_2 NS_195 0 -1.4568575903653339e-03
GC_2_196 b_2 NI_2 NS_196 0 3.2233585197185195e-03
GC_2_197 b_2 NI_2 NS_197 0 3.8009943564368182e-03
GC_2_198 b_2 NI_2 NS_198 0 -2.9784231906263728e-03
GC_2_199 b_2 NI_2 NS_199 0 -1.8786945472682136e-03
GC_2_200 b_2 NI_2 NS_200 0 -3.8879223982944745e-03
GC_2_201 b_2 NI_2 NS_201 0 -4.0380170453442566e-04
GC_2_202 b_2 NI_2 NS_202 0 2.3675226288339046e-03
GC_2_203 b_2 NI_2 NS_203 0 -1.0556794298080710e-05
GC_2_204 b_2 NI_2 NS_204 0 -2.1452512941681735e-05
GC_2_205 b_2 NI_2 NS_205 0 8.4229612476317383e-04
GC_2_206 b_2 NI_2 NS_206 0 -3.7965172925296773e-03
GC_2_207 b_2 NI_2 NS_207 0 3.4279131023208281e-04
GC_2_208 b_2 NI_2 NS_208 0 3.3487732415227699e-03
GC_2_209 b_2 NI_2 NS_209 0 1.3577072327752384e-03
GC_2_210 b_2 NI_2 NS_210 0 -2.3752473045855495e-03
GC_2_211 b_2 NI_2 NS_211 0 2.1858950999962133e-03
GC_2_212 b_2 NI_2 NS_212 0 3.3360403257568518e-03
GC_2_213 b_2 NI_2 NS_213 0 1.1689683902379984e-03
GC_2_214 b_2 NI_2 NS_214 0 2.4033203960224323e-03
GC_2_215 b_2 NI_2 NS_215 0 -8.1092242503903495e-04
GC_2_216 b_2 NI_2 NS_216 0 -1.9781509790535220e-03
GC_2_217 b_2 NI_2 NS_217 0 3.9749449703149785e-04
GC_2_218 b_2 NI_2 NS_218 0 -2.6833646704886027e-03
GC_2_219 b_2 NI_2 NS_219 0 9.8234519887813675e-04
GC_2_220 b_2 NI_2 NS_220 0 2.7459694004685455e-03
GC_2_221 b_2 NI_2 NS_221 0 1.0390528567681089e-03
GC_2_222 b_2 NI_2 NS_222 0 -2.4207680352574222e-03
GC_2_223 b_2 NI_2 NS_223 0 -1.0837521621897010e-03
GC_2_224 b_2 NI_2 NS_224 0 1.5920956224602810e-03
GC_2_225 b_2 NI_2 NS_225 0 -1.1067857241680959e-08
GC_2_226 b_2 NI_2 NS_226 0 -2.8131625100977339e-09
GC_2_227 b_2 NI_2 NS_227 0 2.2673375171341543e-06
GC_2_228 b_2 NI_2 NS_228 0 5.3151463752411419e-07
GC_2_229 b_2 NI_2 NS_229 0 2.9495792726215112e-03
GC_2_230 b_2 NI_2 NS_230 0 -6.1234121947676594e-04
GC_2_231 b_2 NI_2 NS_231 0 2.7949878385541875e-08
GC_2_232 b_2 NI_2 NS_232 0 -3.1702388072309191e-08
GC_2_233 b_2 NI_2 NS_233 0 2.0347269598136963e-04
GC_2_234 b_2 NI_2 NS_234 0 1.3799469331437654e-04
GC_2_235 b_2 NI_2 NS_235 0 5.6259274490763882e-04
GC_2_236 b_2 NI_2 NS_236 0 2.6570823306473382e-04
GC_2_237 b_2 NI_2 NS_237 0 3.1064666446457114e-03
GC_2_238 b_2 NI_2 NS_238 0 -2.2048919772135835e-03
GC_2_239 b_2 NI_2 NS_239 0 -1.5822541432357643e-03
GC_2_240 b_2 NI_2 NS_240 0 -2.6870784023858398e-03
GC_2_241 b_2 NI_2 NS_241 0 -2.0496554889941404e-03
GC_2_242 b_2 NI_2 NS_242 0 -3.7885102412030594e-03
GC_2_243 b_2 NI_2 NS_243 0 -4.9745613666760703e-03
GC_2_244 b_2 NI_2 NS_244 0 -1.5415311521883974e-03
GC_2_245 b_2 NI_2 NS_245 0 2.9290574614371099e-04
GC_2_246 b_2 NI_2 NS_246 0 1.9565159619311094e-04
GC_2_247 b_2 NI_2 NS_247 0 -2.8663291474148754e-03
GC_2_248 b_2 NI_2 NS_248 0 -9.5746385504127127e-04
GC_2_249 b_2 NI_2 NS_249 0 -2.2151871586076614e-02
GC_2_250 b_2 NI_2 NS_250 0 -1.0226316681949583e-02
GC_2_251 b_2 NI_2 NS_251 0 1.1324969792815148e-03
GC_2_252 b_2 NI_2 NS_252 0 2.0395321144443517e-02
GC_2_253 b_2 NI_2 NS_253 0 -5.8416211634823769e-03
GC_2_254 b_2 NI_2 NS_254 0 4.6116292304264608e-03
GC_2_255 b_2 NI_2 NS_255 0 5.7171509182161982e-03
GC_2_256 b_2 NI_2 NS_256 0 3.4516071258136272e-02
GC_2_257 b_2 NI_2 NS_257 0 8.0342763886237564e-03
GC_2_258 b_2 NI_2 NS_258 0 2.7930238789601485e-03
GC_2_259 b_2 NI_2 NS_259 0 -7.7724209649965492e-03
GC_2_260 b_2 NI_2 NS_260 0 2.9556754670022767e-02
GC_2_261 b_2 NI_2 NS_261 0 5.0768429824633934e-02
GC_2_262 b_2 NI_2 NS_262 0 -2.0072962242951624e-02
GC_2_263 b_2 NI_2 NS_263 0 7.9195784236485416e-03
GC_2_264 b_2 NI_2 NS_264 0 -1.6364410949631948e-03
GC_2_265 b_2 NI_2 NS_265 0 2.9084859400548325e-02
GC_2_266 b_2 NI_2 NS_266 0 -2.6464736335252596e-02
GC_2_267 b_2 NI_2 NS_267 0 -6.7250676030620833e-03
GC_2_268 b_2 NI_2 NS_268 0 -9.8822055521542926e-03
GC_2_269 b_2 NI_2 NS_269 0 8.4630825888769388e-03
GC_2_270 b_2 NI_2 NS_270 0 -8.0277978687476846e-03
GC_2_271 b_2 NI_2 NS_271 0 -1.8994952145513517e-02
GC_2_272 b_2 NI_2 NS_272 0 -2.5238421805226313e-02
GC_2_273 b_2 NI_2 NS_273 0 -5.4717849959770434e-03
GC_2_274 b_2 NI_2 NS_274 0 -2.8547841827361725e-03
GC_2_275 b_2 NI_2 NS_275 0 -1.7741073806988972e-02
GC_2_276 b_2 NI_2 NS_276 0 -1.3132230207121672e-02
GC_2_277 b_2 NI_2 NS_277 0 -4.8178006004423943e-03
GC_2_278 b_2 NI_2 NS_278 0 1.2541404095801793e-02
GC_2_279 b_2 NI_2 NS_279 0 -3.4590900613967199e-03
GC_2_280 b_2 NI_2 NS_280 0 1.5412381719795960e-03
GC_2_281 b_2 NI_2 NS_281 0 -7.1865144567420972e-04
GC_2_282 b_2 NI_2 NS_282 0 7.0058605784199604e-03
GC_2_283 b_2 NI_2 NS_283 0 1.8820413841029871e-03
GC_2_284 b_2 NI_2 NS_284 0 8.5748619143940320e-05
GC_2_285 b_2 NI_2 NS_285 0 3.1400281534097173e-04
GC_2_286 b_2 NI_2 NS_286 0 -1.9467014119337795e-03
GC_2_287 b_2 NI_2 NS_287 0 -1.8563352640916424e-03
GC_2_288 b_2 NI_2 NS_288 0 -1.6182088771356617e-03
GC_2_289 b_2 NI_2 NS_289 0 -2.1290960700133888e-03
GC_2_290 b_2 NI_2 NS_290 0 1.6850433455973452e-03
GC_2_291 b_2 NI_2 NS_291 0 7.6361045370997754e-04
GC_2_292 b_2 NI_2 NS_292 0 1.8527513037901096e-04
GC_2_293 b_2 NI_2 NS_293 0 -6.9730354411923852e-04
GC_2_294 b_2 NI_2 NS_294 0 -1.6780703341174393e-03
GC_2_295 b_2 NI_2 NS_295 0 -2.6815282169833188e-03
GC_2_296 b_2 NI_2 NS_296 0 -8.2749160397336142e-04
GC_2_297 b_2 NI_2 NS_297 0 -4.9989688575079769e-04
GC_2_298 b_2 NI_2 NS_298 0 2.9288639063664744e-03
GC_2_299 b_2 NI_2 NS_299 0 1.3533574670609901e-03
GC_2_300 b_2 NI_2 NS_300 0 -8.5805587459256930e-04
GC_2_301 b_2 NI_2 NS_301 0 -2.4189247508466386e-03
GC_2_302 b_2 NI_2 NS_302 0 -2.2676209709430206e-03
GC_2_303 b_2 NI_2 NS_303 0 -3.5540455364462798e-03
GC_2_304 b_2 NI_2 NS_304 0 7.4852673501159446e-04
GC_2_305 b_2 NI_2 NS_305 0 2.4633829778002731e-03
GC_2_306 b_2 NI_2 NS_306 0 3.0182799552168531e-03
GC_2_307 b_2 NI_2 NS_307 0 9.8455399410401438e-04
GC_2_308 b_2 NI_2 NS_308 0 -2.9418100018954773e-03
GC_2_309 b_2 NI_2 NS_309 0 -4.7678001582966423e-03
GC_2_310 b_2 NI_2 NS_310 0 5.4340316487482121e-05
GC_2_311 b_2 NI_2 NS_311 0 -1.7083702925141939e-03
GC_2_312 b_2 NI_2 NS_312 0 3.7124268853424409e-03
GC_2_313 b_2 NI_2 NS_313 0 -7.6587734480741752e-04
GC_2_314 b_2 NI_2 NS_314 0 1.5006835278413978e-03
GC_2_315 b_2 NI_2 NS_315 0 3.2213013460885538e-03
GC_2_316 b_2 NI_2 NS_316 0 -1.3508686582678691e-03
GC_2_317 b_2 NI_2 NS_317 0 -2.9326239923893263e-06
GC_2_318 b_2 NI_2 NS_318 0 8.7469591660207792e-06
GC_2_319 b_2 NI_2 NS_319 0 -1.8200422844684423e-03
GC_2_320 b_2 NI_2 NS_320 0 -2.5277365468768342e-03
GC_2_321 b_2 NI_2 NS_321 0 -2.4072537648056622e-03
GC_2_322 b_2 NI_2 NS_322 0 2.4886636555887360e-03
GC_2_323 b_2 NI_2 NS_323 0 1.0142618788330706e-03
GC_2_324 b_2 NI_2 NS_324 0 2.4256808521002662e-03
GC_2_325 b_2 NI_2 NS_325 0 8.5775914702243918e-04
GC_2_326 b_2 NI_2 NS_326 0 -2.6994858348549748e-03
GC_2_327 b_2 NI_2 NS_327 0 -3.0644780738181370e-04
GC_2_328 b_2 NI_2 NS_328 0 1.6741356978676677e-03
GC_2_329 b_2 NI_2 NS_329 0 -1.7840539158117958e-03
GC_2_330 b_2 NI_2 NS_330 0 -3.1181076893642602e-04
GC_2_331 b_2 NI_2 NS_331 0 1.4004539382215157e-03
GC_2_332 b_2 NI_2 NS_332 0 1.9709616317316867e-03
GC_2_333 b_2 NI_2 NS_333 0 1.0449287577521927e-03
GC_2_334 b_2 NI_2 NS_334 0 -2.2998045192744393e-03
GC_2_335 b_2 NI_2 NS_335 0 -6.9799496653780678e-04
GC_2_336 b_2 NI_2 NS_336 0 -1.4668898647731416e-03
GC_2_337 b_2 NI_2 NS_337 0 -1.3735491585586416e-03
GC_2_338 b_2 NI_2 NS_338 0 -3.1252860516914880e-04
GC_2_339 b_2 NI_2 NS_339 0 7.1030028256060112e-09
GC_2_340 b_2 NI_2 NS_340 0 -2.4709996242732650e-08
GC_2_341 b_2 NI_2 NS_341 0 -4.5275393918210935e-07
GC_2_342 b_2 NI_2 NS_342 0 1.6341836566458982e-06
GC_2_343 b_2 NI_2 NS_343 0 7.7517773778853728e-03
GC_2_344 b_2 NI_2 NS_344 0 -1.6012310594381263e-03
GC_2_345 b_2 NI_2 NS_345 0 -1.2107575666080743e-08
GC_2_346 b_2 NI_2 NS_346 0 -8.8419586430203635e-07
GC_2_347 b_2 NI_2 NS_347 0 1.0389377947345378e-04
GC_2_348 b_2 NI_2 NS_348 0 -5.1165589632056981e-04
GC_2_349 b_2 NI_2 NS_349 0 -1.9366724880200566e-03
GC_2_350 b_2 NI_2 NS_350 0 -5.9740804149900466e-04
GC_2_351 b_2 NI_2 NS_351 0 2.9415452896669123e-03
GC_2_352 b_2 NI_2 NS_352 0 2.2646130278170971e-03
GC_2_353 b_2 NI_2 NS_353 0 -3.5699577149257669e-03
GC_2_354 b_2 NI_2 NS_354 0 -3.0486836838590102e-03
GC_2_355 b_2 NI_2 NS_355 0 -1.7071501568238681e-03
GC_2_356 b_2 NI_2 NS_356 0 5.8436838666205398e-03
GC_2_357 b_2 NI_2 NS_357 0 4.3687530436905065e-03
GC_2_358 b_2 NI_2 NS_358 0 -2.4745967049057682e-03
GC_2_359 b_2 NI_2 NS_359 0 -1.1051197485519853e-04
GC_2_360 b_2 NI_2 NS_360 0 -1.0369084873499772e-04
GC_2_361 b_2 NI_2 NS_361 0 -4.4520053128230506e-03
GC_2_362 b_2 NI_2 NS_362 0 -9.2458240841154066e-04
GC_2_363 b_2 NI_2 NS_363 0 9.1257593927417772e-03
GC_2_364 b_2 NI_2 NS_364 0 1.7785327687101470e-02
GC_2_365 b_2 NI_2 NS_365 0 -4.0274380463636390e-03
GC_2_366 b_2 NI_2 NS_366 0 -1.7847943499154681e-02
GC_2_367 b_2 NI_2 NS_367 0 -8.2175435813232091e-03
GC_2_368 b_2 NI_2 NS_368 0 4.1736391799597570e-03
GC_2_369 b_2 NI_2 NS_369 0 1.7064439428660535e-02
GC_2_370 b_2 NI_2 NS_370 0 -4.4005705420395371e-04
GC_2_371 b_2 NI_2 NS_371 0 -9.2787949621601987e-03
GC_2_372 b_2 NI_2 NS_372 0 -3.2071945428810782e-03
GC_2_373 b_2 NI_2 NS_373 0 -1.3712651090382026e-02
GC_2_374 b_2 NI_2 NS_374 0 2.2836662053447115e-02
GC_2_375 b_2 NI_2 NS_375 0 2.2839357165334383e-02
GC_2_376 b_2 NI_2 NS_376 0 -2.2670702905947613e-02
GC_2_377 b_2 NI_2 NS_377 0 -9.2392572685181598e-03
GC_2_378 b_2 NI_2 NS_378 0 9.0801440054633206e-04
GC_2_379 b_2 NI_2 NS_379 0 1.8480442543301921e-02
GC_2_380 b_2 NI_2 NS_380 0 6.2433937813125770e-03
GC_2_381 b_2 NI_2 NS_381 0 -9.1763268352659504e-03
GC_2_382 b_2 NI_2 NS_382 0 -9.4611046174689975e-03
GC_2_383 b_2 NI_2 NS_383 0 -9.9741852673505774e-03
GC_2_384 b_2 NI_2 NS_384 0 6.3961382701889277e-03
GC_2_385 b_2 NI_2 NS_385 0 1.6838377576843935e-02
GC_2_386 b_2 NI_2 NS_386 0 -4.8507523614030818e-03
GC_2_387 b_2 NI_2 NS_387 0 -7.2149762239858695e-03
GC_2_388 b_2 NI_2 NS_388 0 -3.4093174612818793e-03
GC_2_389 b_2 NI_2 NS_389 0 6.8284576463739219e-03
GC_2_390 b_2 NI_2 NS_390 0 1.3296720248934787e-02
GC_2_391 b_2 NI_2 NS_391 0 -1.8198397290107380e-03
GC_2_392 b_2 NI_2 NS_392 0 -1.4401884725728122e-02
GC_2_393 b_2 NI_2 NS_393 0 -4.9859625706528358e-03
GC_2_394 b_2 NI_2 NS_394 0 1.0394190570049459e-03
GC_2_395 b_2 NI_2 NS_395 0 6.0026878584690897e-03
GC_2_396 b_2 NI_2 NS_396 0 -1.1033368423158797e-03
GC_2_397 b_2 NI_2 NS_397 0 -3.4642734771405405e-03
GC_2_398 b_2 NI_2 NS_398 0 -1.0877136295650300e-03
GC_2_399 b_2 NI_2 NS_399 0 2.7180843192213962e-03
GC_2_400 b_2 NI_2 NS_400 0 -5.0793037241864884e-04
GC_2_401 b_2 NI_2 NS_401 0 -3.2964042742944203e-03
GC_2_402 b_2 NI_2 NS_402 0 -2.8952144423371596e-03
GC_2_403 b_2 NI_2 NS_403 0 2.0160578131157123e-03
GC_2_404 b_2 NI_2 NS_404 0 7.7561498992574326e-04
GC_2_405 b_2 NI_2 NS_405 0 -2.0162392358003601e-03
GC_2_406 b_2 NI_2 NS_406 0 -9.6653808865190881e-04
GC_2_407 b_2 NI_2 NS_407 0 2.1216790410996246e-03
GC_2_408 b_2 NI_2 NS_408 0 -1.4710183113699846e-03
GC_2_409 b_2 NI_2 NS_409 0 -4.1846676197283455e-03
GC_2_410 b_2 NI_2 NS_410 0 -1.8129776339244359e-03
GC_2_411 b_2 NI_2 NS_411 0 2.3699534346868795e-03
GC_2_412 b_2 NI_2 NS_412 0 -3.7091486379361028e-04
GC_2_413 b_2 NI_2 NS_413 0 -3.0171271284337611e-03
GC_2_414 b_2 NI_2 NS_414 0 4.6227949902273986e-04
GC_2_415 b_2 NI_2 NS_415 0 2.7066174204063327e-03
GC_2_416 b_2 NI_2 NS_416 0 -2.7283516400600154e-03
GC_2_417 b_2 NI_2 NS_417 0 -5.0391209614568267e-03
GC_2_418 b_2 NI_2 NS_418 0 -1.2777720509594227e-04
GC_2_419 b_2 NI_2 NS_419 0 2.4350415202187030e-03
GC_2_420 b_2 NI_2 NS_420 0 -2.1722385743882301e-03
GC_2_421 b_2 NI_2 NS_421 0 -3.2447311674065238e-03
GC_2_422 b_2 NI_2 NS_422 0 2.6004814944434384e-03
GC_2_423 b_2 NI_2 NS_423 0 1.7440028190431509e-03
GC_2_424 b_2 NI_2 NS_424 0 -4.7506654664725241e-03
GC_2_425 b_2 NI_2 NS_425 0 -3.6334488908336023e-03
GC_2_426 b_2 NI_2 NS_426 0 2.5968949548931513e-03
GC_2_427 b_2 NI_2 NS_427 0 -2.8337755503635518e-03
GC_2_428 b_2 NI_2 NS_428 0 3.9869976680980898e-03
GC_2_429 b_2 NI_2 NS_429 0 -2.2097291659768591e-04
GC_2_430 b_2 NI_2 NS_430 0 -4.2143931767534559e-03
GC_2_431 b_2 NI_2 NS_431 0 -9.9004930717312887e-06
GC_2_432 b_2 NI_2 NS_432 0 7.5068431570776734e-06
GC_2_433 b_2 NI_2 NS_433 0 -1.3536752221605566e-03
GC_2_434 b_2 NI_2 NS_434 0 3.3750369352797730e-03
GC_2_435 b_2 NI_2 NS_435 0 -9.6981082599738549e-04
GC_2_436 b_2 NI_2 NS_436 0 -4.3483886339256966e-03
GC_2_437 b_2 NI_2 NS_437 0 -1.0004295426337179e-03
GC_2_438 b_2 NI_2 NS_438 0 2.2215356041265775e-03
GC_2_439 b_2 NI_2 NS_439 0 -1.6509349865853028e-03
GC_2_440 b_2 NI_2 NS_440 0 -4.4091720150585424e-03
GC_2_441 b_2 NI_2 NS_441 0 -1.4483889308222768e-03
GC_2_442 b_2 NI_2 NS_442 0 -2.4971171259750482e-03
GC_2_443 b_2 NI_2 NS_443 0 7.8206440214795671e-04
GC_2_444 b_2 NI_2 NS_444 0 2.5934686425242003e-03
GC_2_445 b_2 NI_2 NS_445 0 -6.9629932558045945e-04
GC_2_446 b_2 NI_2 NS_446 0 2.8791308451955001e-03
GC_2_447 b_2 NI_2 NS_447 0 -1.4354331597146233e-03
GC_2_448 b_2 NI_2 NS_448 0 -2.7718926043723271e-03
GC_2_449 b_2 NI_2 NS_449 0 -1.1678459034003472e-03
GC_2_450 b_2 NI_2 NS_450 0 2.6661739427565573e-03
GC_2_451 b_2 NI_2 NS_451 0 7.8077002249662888e-04
GC_2_452 b_2 NI_2 NS_452 0 -1.8746307425867408e-03
GC_2_453 b_2 NI_2 NS_453 0 2.3791410613138728e-08
GC_2_454 b_2 NI_2 NS_454 0 -6.0255378988179937e-08
GC_2_455 b_2 NI_2 NS_455 0 -9.0379195589119467e-07
GC_2_456 b_2 NI_2 NS_456 0 3.2032331613926917e-06
GC_2_457 b_2 NI_2 NS_457 0 -3.8126145421109555e-05
GC_2_458 b_2 NI_2 NS_458 0 2.2429780013294595e-06
GC_2_459 b_2 NI_2 NS_459 0 5.7510315309722728e-11
GC_2_460 b_2 NI_2 NS_460 0 3.0677000352002756e-09
GC_2_461 b_2 NI_2 NS_461 0 -1.9278399077390812e-06
GC_2_462 b_2 NI_2 NS_462 0 -1.7007509566656212e-06
GC_2_463 b_2 NI_2 NS_463 0 -5.6017352409557403e-06
GC_2_464 b_2 NI_2 NS_464 0 2.8809340764108912e-06
GC_2_465 b_2 NI_2 NS_465 0 -1.6609148419360369e-05
GC_2_466 b_2 NI_2 NS_466 0 1.9115494014770666e-05
GC_2_467 b_2 NI_2 NS_467 0 1.5381838597530011e-05
GC_2_468 b_2 NI_2 NS_468 0 1.0271588431257469e-05
GC_2_469 b_2 NI_2 NS_469 0 1.7283121532183457e-05
GC_2_470 b_2 NI_2 NS_470 0 2.3212332368670635e-05
GC_2_471 b_2 NI_2 NS_471 0 3.0964746108475604e-05
GC_2_472 b_2 NI_2 NS_472 0 5.3078390946276810e-06
GC_2_473 b_2 NI_2 NS_473 0 -3.3865371779836663e-06
GC_2_474 b_2 NI_2 NS_474 0 -2.1454163663258833e-06
GC_2_475 b_2 NI_2 NS_475 0 1.7199892457945204e-05
GC_2_476 b_2 NI_2 NS_476 0 -2.1239549379839019e-06
GC_2_477 b_2 NI_2 NS_477 0 1.2959268469623852e-04
GC_2_478 b_2 NI_2 NS_478 0 3.5267997551867905e-05
GC_2_479 b_2 NI_2 NS_479 0 -2.8363536859844153e-05
GC_2_480 b_2 NI_2 NS_480 0 -1.0001971518228863e-04
GC_2_481 b_2 NI_2 NS_481 0 2.5326198621965190e-05
GC_2_482 b_2 NI_2 NS_482 0 -3.1109552973910961e-05
GC_2_483 b_2 NI_2 NS_483 0 -4.1103625530690115e-05
GC_2_484 b_2 NI_2 NS_484 0 -1.6753401710173658e-04
GC_2_485 b_2 NI_2 NS_485 0 -4.1819867668073262e-05
GC_2_486 b_2 NI_2 NS_486 0 -5.5994630457197798e-06
GC_2_487 b_2 NI_2 NS_487 0 2.2900988024227043e-05
GC_2_488 b_2 NI_2 NS_488 0 -1.5132579087555076e-04
GC_2_489 b_2 NI_2 NS_489 0 -2.3194062423213379e-04
GC_2_490 b_2 NI_2 NS_490 0 1.1300294384142839e-04
GC_2_491 b_2 NI_2 NS_491 0 -3.7469906456433307e-05
GC_2_492 b_2 NI_2 NS_492 0 1.3727346467279548e-05
GC_2_493 b_2 NI_2 NS_493 0 -1.3772206140927795e-04
GC_2_494 b_2 NI_2 NS_494 0 1.2973991904714015e-04
GC_2_495 b_2 NI_2 NS_495 0 3.6015990846596232e-05
GC_2_496 b_2 NI_2 NS_496 0 4.1758736164586717e-05
GC_2_497 b_2 NI_2 NS_497 0 -3.8325873675016681e-05
GC_2_498 b_2 NI_2 NS_498 0 4.2733754681994854e-05
GC_2_499 b_2 NI_2 NS_499 0 8.7553203531928582e-05
GC_2_500 b_2 NI_2 NS_500 0 1.1830509384616555e-04
GC_2_501 b_2 NI_2 NS_501 0 2.7200342385980316e-05
GC_2_502 b_2 NI_2 NS_502 0 1.0487248115855233e-05
GC_2_503 b_2 NI_2 NS_503 0 8.6919301602754177e-05
GC_2_504 b_2 NI_2 NS_504 0 6.5387413420267844e-05
GC_2_505 b_2 NI_2 NS_505 0 2.0648990354311142e-05
GC_2_506 b_2 NI_2 NS_506 0 -5.7329958705323692e-05
GC_2_507 b_2 NI_2 NS_507 0 1.7010943409808137e-05
GC_2_508 b_2 NI_2 NS_508 0 -8.6982096013409108e-06
GC_2_509 b_2 NI_2 NS_509 0 8.3263451945088089e-06
GC_2_510 b_2 NI_2 NS_510 0 -3.3101469207872683e-05
GC_2_511 b_2 NI_2 NS_511 0 -8.8263224347399455e-06
GC_2_512 b_2 NI_2 NS_512 0 3.3245522078929201e-07
GC_2_513 b_2 NI_2 NS_513 0 -2.3512434032311600e-06
GC_2_514 b_2 NI_2 NS_514 0 8.4561785160927535e-06
GC_2_515 b_2 NI_2 NS_515 0 1.0134608853512476e-05
GC_2_516 b_2 NI_2 NS_516 0 6.1703155359101972e-06
GC_2_517 b_2 NI_2 NS_517 0 1.2106283434026199e-05
GC_2_518 b_2 NI_2 NS_518 0 -7.8948002966209239e-06
GC_2_519 b_2 NI_2 NS_519 0 -3.4458125858481598e-06
GC_2_520 b_2 NI_2 NS_520 0 -5.4102916634246623e-07
GC_2_521 b_2 NI_2 NS_521 0 2.5535447627906504e-06
GC_2_522 b_2 NI_2 NS_522 0 7.3550393086767715e-06
GC_2_523 b_2 NI_2 NS_523 0 1.3648180774188222e-05
GC_2_524 b_2 NI_2 NS_524 0 2.7057424102060667e-06
GC_2_525 b_2 NI_2 NS_525 0 4.5460289824291641e-06
GC_2_526 b_2 NI_2 NS_526 0 -1.4254776148381142e-05
GC_2_527 b_2 NI_2 NS_527 0 -5.8809806720570141e-06
GC_2_528 b_2 NI_2 NS_528 0 4.1779762857959373e-06
GC_2_529 b_2 NI_2 NS_529 0 1.0407199106658150e-05
GC_2_530 b_2 NI_2 NS_530 0 9.8673809492871069e-06
GC_2_531 b_2 NI_2 NS_531 0 1.7371591512955435e-05
GC_2_532 b_2 NI_2 NS_532 0 -4.2133739970412172e-06
GC_2_533 b_2 NI_2 NS_533 0 -9.1859982607328866e-06
GC_2_534 b_2 NI_2 NS_534 0 -1.5417369730909773e-05
GC_2_535 b_2 NI_2 NS_535 0 -3.9937420604051080e-06
GC_2_536 b_2 NI_2 NS_536 0 1.3459879586596607e-05
GC_2_537 b_2 NI_2 NS_537 0 2.1061386147212581e-05
GC_2_538 b_2 NI_2 NS_538 0 -6.9747259698229141e-07
GC_2_539 b_2 NI_2 NS_539 0 9.0884856063751424e-06
GC_2_540 b_2 NI_2 NS_540 0 -1.7352201611856742e-05
GC_2_541 b_2 NI_2 NS_541 0 1.8906919983534022e-06
GC_2_542 b_2 NI_2 NS_542 0 -1.4899317806407173e-05
GC_2_543 b_2 NI_2 NS_543 0 -1.3643680222395739e-05
GC_2_544 b_2 NI_2 NS_544 0 4.0673710546740363e-06
GC_2_545 b_2 NI_2 NS_545 0 1.3202617770948745e-08
GC_2_546 b_2 NI_2 NS_546 0 -4.9292960769132304e-08
GC_2_547 b_2 NI_2 NS_547 0 8.7095219841643637e-06
GC_2_548 b_2 NI_2 NS_548 0 1.1413355381623932e-05
GC_2_549 b_2 NI_2 NS_549 0 1.0949854761009922e-05
GC_2_550 b_2 NI_2 NS_550 0 -1.1467430611896881e-05
GC_2_551 b_2 NI_2 NS_551 0 -3.5678216235840095e-06
GC_2_552 b_2 NI_2 NS_552 0 -1.0053365341892320e-05
GC_2_553 b_2 NI_2 NS_553 0 -2.0108394133224388e-06
GC_2_554 b_2 NI_2 NS_554 0 1.3050215603618248e-05
GC_2_555 b_2 NI_2 NS_555 0 9.7274307634934138e-07
GC_2_556 b_2 NI_2 NS_556 0 -7.2791931750609059e-06
GC_2_557 b_2 NI_2 NS_557 0 7.4348965660094463e-06
GC_2_558 b_2 NI_2 NS_558 0 1.7180574063960692e-06
GC_2_559 b_2 NI_2 NS_559 0 -6.1040138549410502e-06
GC_2_560 b_2 NI_2 NS_560 0 -8.8986588134885606e-06
GC_2_561 b_2 NI_2 NS_561 0 -4.1281705341514484e-06
GC_2_562 b_2 NI_2 NS_562 0 9.6390058961427223e-06
GC_2_563 b_2 NI_2 NS_563 0 3.3246533001382367e-06
GC_2_564 b_2 NI_2 NS_564 0 6.0744636677885924e-06
GC_2_565 b_2 NI_2 NS_565 0 5.7495240499624785e-06
GC_2_566 b_2 NI_2 NS_566 0 5.2303417392620955e-07
GC_2_567 b_2 NI_2 NS_567 0 5.7042482092918390e-11
GC_2_568 b_2 NI_2 NS_568 0 1.4838925086350135e-10
GC_2_569 b_2 NI_2 NS_569 0 6.0314121284059970e-09
GC_2_570 b_2 NI_2 NS_570 0 -8.4056564596109882e-09
GC_2_571 b_2 NI_2 NS_571 0 -1.1889665190136687e-04
GC_2_572 b_2 NI_2 NS_572 0 -2.1515751052027916e-06
GC_2_573 b_2 NI_2 NS_573 0 -2.4447828841623735e-10
GC_2_574 b_2 NI_2 NS_574 0 2.5353387457701169e-09
GC_2_575 b_2 NI_2 NS_575 0 1.5643085700313063e-06
GC_2_576 b_2 NI_2 NS_576 0 -1.5218359475695793e-06
GC_2_577 b_2 NI_2 NS_577 0 -8.9297830737699720e-09
GC_2_578 b_2 NI_2 NS_578 0 -6.1820522471670406e-06
GC_2_579 b_2 NI_2 NS_579 0 -7.6539314483315976e-06
GC_2_580 b_2 NI_2 NS_580 0 5.3261378272329129e-07
GC_2_581 b_2 NI_2 NS_581 0 -9.8452203377515357e-07
GC_2_582 b_2 NI_2 NS_582 0 -4.3923453456296181e-06
GC_2_583 b_2 NI_2 NS_583 0 -1.5585557096571115e-05
GC_2_584 b_2 NI_2 NS_584 0 -1.3013886552039649e-06
GC_2_585 b_2 NI_2 NS_585 0 -5.3235186219972581e-06
GC_2_586 b_2 NI_2 NS_586 0 1.9150005299466030e-05
GC_2_587 b_2 NI_2 NS_587 0 4.4241060801470735e-06
GC_2_588 b_2 NI_2 NS_588 0 -3.1123180198401221e-06
GC_2_589 b_2 NI_2 NS_589 0 1.2804786107827318e-07
GC_2_590 b_2 NI_2 NS_590 0 -2.5891790723550555e-06
GC_2_591 b_2 NI_2 NS_591 0 -2.4876404743375842e-05
GC_2_592 b_2 NI_2 NS_592 0 2.8210753953300287e-05
GC_2_593 b_2 NI_2 NS_593 0 2.7762971664200824e-05
GC_2_594 b_2 NI_2 NS_594 0 -8.7259229447981464e-06
GC_2_595 b_2 NI_2 NS_595 0 -7.7819273879627227e-06
GC_2_596 b_2 NI_2 NS_596 0 -4.1753176951320778e-06
GC_2_597 b_2 NI_2 NS_597 0 1.2787917415274856e-05
GC_2_598 b_2 NI_2 NS_598 0 2.6107424771221397e-05
GC_2_599 b_2 NI_2 NS_599 0 1.4270067896338161e-06
GC_2_600 b_2 NI_2 NS_600 0 -8.8305599645571942e-06
GC_2_601 b_2 NI_2 NS_601 0 -2.7324696858414378e-05
GC_2_602 b_2 NI_2 NS_602 0 5.0137308266355514e-06
GC_2_603 b_2 NI_2 NS_603 0 4.0396636126122139e-05
GC_2_604 b_2 NI_2 NS_604 0 9.6550503763662491e-06
GC_2_605 b_2 NI_2 NS_605 0 -2.8820962081267942e-06
GC_2_606 b_2 NI_2 NS_606 0 -4.3143669172992278e-06
GC_2_607 b_2 NI_2 NS_607 0 1.3053639094992278e-05
GC_2_608 b_2 NI_2 NS_608 0 1.8104097724720489e-05
GC_2_609 b_2 NI_2 NS_609 0 3.5097808089726455e-06
GC_2_610 b_2 NI_2 NS_610 0 -1.0678067842191033e-05
GC_2_611 b_2 NI_2 NS_611 0 -6.1544161233581069e-06
GC_2_612 b_2 NI_2 NS_612 0 1.0310052394207302e-06
GC_2_613 b_2 NI_2 NS_613 0 1.8592830052407238e-05
GC_2_614 b_2 NI_2 NS_614 0 4.7647994636989809e-06
GC_2_615 b_2 NI_2 NS_615 0 -1.6257204329740137e-07
GC_2_616 b_2 NI_2 NS_616 0 -4.0317312744565410e-06
GC_2_617 b_2 NI_2 NS_617 0 5.3001344430040513e-06
GC_2_618 b_2 NI_2 NS_618 0 1.3913341154526265e-05
GC_2_619 b_2 NI_2 NS_619 0 7.3647531479878706e-06
GC_2_620 b_2 NI_2 NS_620 0 -1.1146120799689468e-05
GC_2_621 b_2 NI_2 NS_621 0 -1.3430338836535959e-06
GC_2_622 b_2 NI_2 NS_622 0 1.0232544103023052e-06
GC_2_623 b_2 NI_2 NS_623 0 1.0874239562731582e-05
GC_2_624 b_2 NI_2 NS_624 0 3.8626541644343327e-06
GC_2_625 b_2 NI_2 NS_625 0 1.6867603292858436e-06
GC_2_626 b_2 NI_2 NS_626 0 -5.9600513575350683e-07
GC_2_627 b_2 NI_2 NS_627 0 5.6731245568656106e-06
GC_2_628 b_2 NI_2 NS_628 0 1.6014341794102558e-06
GC_2_629 b_2 NI_2 NS_629 0 3.3818685123247231e-06
GC_2_630 b_2 NI_2 NS_630 0 2.0535677158039071e-06
GC_2_631 b_2 NI_2 NS_631 0 1.1002372514272964e-05
GC_2_632 b_2 NI_2 NS_632 0 3.6804860206141826e-06
GC_2_633 b_2 NI_2 NS_633 0 4.8497229807595525e-06
GC_2_634 b_2 NI_2 NS_634 0 -8.6121374771457664e-08
GC_2_635 b_2 NI_2 NS_635 0 9.9794195515369079e-06
GC_2_636 b_2 NI_2 NS_636 0 -1.1587618576747175e-06
GC_2_637 b_2 NI_2 NS_637 0 8.2788150445617330e-06
GC_2_638 b_2 NI_2 NS_638 0 2.9673088558733744e-06
GC_2_639 b_2 NI_2 NS_639 0 1.9120276973391630e-05
GC_2_640 b_2 NI_2 NS_640 0 -5.6689228093488515e-06
GC_2_641 b_2 NI_2 NS_641 0 7.2485954099759134e-06
GC_2_642 b_2 NI_2 NS_642 0 -4.0295064560293275e-06
GC_2_643 b_2 NI_2 NS_643 0 1.3800813643098931e-05
GC_2_644 b_2 NI_2 NS_644 0 -1.2000538269531615e-05
GC_2_645 b_2 NI_2 NS_645 0 1.2506358506717436e-05
GC_2_646 b_2 NI_2 NS_646 0 -3.9183446889610967e-06
GC_2_647 b_2 NI_2 NS_647 0 9.3634143384864689e-06
GC_2_648 b_2 NI_2 NS_648 0 -2.6978357460782655e-05
GC_2_649 b_2 NI_2 NS_649 0 2.5168592268940938e-06
GC_2_650 b_2 NI_2 NS_650 0 -1.2425235333244613e-05
GC_2_651 b_2 NI_2 NS_651 0 -8.1224251343218550e-06
GC_2_652 b_2 NI_2 NS_652 0 -1.8906424102071361e-05
GC_2_653 b_2 NI_2 NS_653 0 -4.4970473668116960e-06
GC_2_654 b_2 NI_2 NS_654 0 -1.2065329369989343e-05
GC_2_655 b_2 NI_2 NS_655 0 5.2902141876645946e-05
GC_2_656 b_2 NI_2 NS_656 0 -8.9264416266488785e-05
GC_2_657 b_2 NI_2 NS_657 0 -9.8974227905403725e-06
GC_2_658 b_2 NI_2 NS_658 0 6.3392400347989702e-07
GC_2_659 b_2 NI_2 NS_659 0 3.8297080116946243e-07
GC_2_660 b_2 NI_2 NS_660 0 -1.3807140751481266e-07
GC_2_661 b_2 NI_2 NS_661 0 -2.6243895052963541e-06
GC_2_662 b_2 NI_2 NS_662 0 -2.3105603753959717e-06
GC_2_663 b_2 NI_2 NS_663 0 -4.4577508265747636e-06
GC_2_664 b_2 NI_2 NS_664 0 2.7145411372357149e-07
GC_2_665 b_2 NI_2 NS_665 0 -1.7068913101714160e-05
GC_2_666 b_2 NI_2 NS_666 0 9.6343682918614459e-06
GC_2_667 b_2 NI_2 NS_667 0 -8.5804544315371991e-06
GC_2_668 b_2 NI_2 NS_668 0 3.7246477444496816e-05
GC_2_669 b_2 NI_2 NS_669 0 -7.2739652247995409e-06
GC_2_670 b_2 NI_2 NS_670 0 3.7766515731380429e-07
GC_2_671 b_2 NI_2 NS_671 0 -1.3438136112483517e-05
GC_2_672 b_2 NI_2 NS_672 0 1.9879390826485144e-06
GC_2_673 b_2 NI_2 NS_673 0 -4.6768386269797029e-06
GC_2_674 b_2 NI_2 NS_674 0 -3.4323461850717753e-06
GC_2_675 b_2 NI_2 NS_675 0 -6.4511240799349945e-06
GC_2_676 b_2 NI_2 NS_676 0 1.0470457215021574e-06
GC_2_677 b_2 NI_2 NS_677 0 -3.0717703405032320e-06
GC_2_678 b_2 NI_2 NS_678 0 8.7596277011058588e-07
GC_2_679 b_2 NI_2 NS_679 0 -1.8095974103547490e-06
GC_2_680 b_2 NI_2 NS_680 0 -9.3346424913158260e-07
GC_2_681 b_2 NI_2 NS_681 0 -2.5782249015160393e-10
GC_2_682 b_2 NI_2 NS_682 0 4.1882528775927913e-10
GC_2_683 b_2 NI_2 NS_683 0 2.1382058932723421e-09
GC_2_684 b_2 NI_2 NS_684 0 -2.6515544213761256e-08
GC_2_685 b_2 NI_2 NS_685 0 -6.2021626709423257e-05
GC_2_686 b_2 NI_2 NS_686 0 3.1006124253686665e-07
GC_2_687 b_2 NI_2 NS_687 0 1.6341689521018586e-11
GC_2_688 b_2 NI_2 NS_688 0 -8.7701220840072195e-11
GC_2_689 b_2 NI_2 NS_689 0 -1.1181529415063307e-06
GC_2_690 b_2 NI_2 NS_690 0 -1.7690614888983087e-06
GC_2_691 b_2 NI_2 NS_691 0 -1.9757200225012559e-06
GC_2_692 b_2 NI_2 NS_692 0 1.9724312780572612e-06
GC_2_693 b_2 NI_2 NS_693 0 -9.5765593063874671e-06
GC_2_694 b_2 NI_2 NS_694 0 6.8034136613391432e-07
GC_2_695 b_2 NI_2 NS_695 0 -2.2987481038458849e-07
GC_2_696 b_2 NI_2 NS_696 0 3.5063290314872800e-06
GC_2_697 b_2 NI_2 NS_697 0 -2.0994415670304274e-06
GC_2_698 b_2 NI_2 NS_698 0 1.1705852359787371e-05
GC_2_699 b_2 NI_2 NS_699 0 6.8703457329792806e-06
GC_2_700 b_2 NI_2 NS_700 0 1.2241242737182216e-05
GC_2_701 b_2 NI_2 NS_701 0 -2.0277601157354628e-06
GC_2_702 b_2 NI_2 NS_702 0 -2.2588482069851019e-06
GC_2_703 b_2 NI_2 NS_703 0 1.6453776754194627e-06
GC_2_704 b_2 NI_2 NS_704 0 1.0187566512107025e-06
GC_2_705 b_2 NI_2 NS_705 0 7.3910975614293019e-06
GC_2_706 b_2 NI_2 NS_706 0 3.8498707711955123e-05
GC_2_707 b_2 NI_2 NS_707 0 2.2957037801936800e-05
GC_2_708 b_2 NI_2 NS_708 0 -1.2018263828446583e-05
GC_2_709 b_2 NI_2 NS_709 0 8.4099953827387901e-06
GC_2_710 b_2 NI_2 NS_710 0 1.7737176793971525e-06
GC_2_711 b_2 NI_2 NS_711 0 4.7831240784761748e-05
GC_2_712 b_2 NI_2 NS_712 0 -2.5191947081810410e-05
GC_2_713 b_2 NI_2 NS_713 0 -9.1802611209784247e-07
GC_2_714 b_2 NI_2 NS_714 0 -8.0507038261386457e-06
GC_2_715 b_2 NI_2 NS_715 0 3.4285634382887531e-05
GC_2_716 b_2 NI_2 NS_716 0 -7.7290034913422946e-06
GC_2_717 b_2 NI_2 NS_717 0 -3.8666328320067861e-05
GC_2_718 b_2 NI_2 NS_718 0 -5.1897463357019726e-05
GC_2_719 b_2 NI_2 NS_719 0 -4.5703072675549051e-06
GC_2_720 b_2 NI_2 NS_720 0 -4.5524722373524250e-06
GC_2_721 b_2 NI_2 NS_721 0 -3.9431764743747368e-05
GC_2_722 b_2 NI_2 NS_722 0 -1.9713947869860132e-05
GC_2_723 b_2 NI_2 NS_723 0 -4.8992954662857712e-06
GC_2_724 b_2 NI_2 NS_724 0 6.5785889776379930e-06
GC_2_725 b_2 NI_2 NS_725 0 -8.6427728546088723e-06
GC_2_726 b_2 NI_2 NS_726 0 -6.9219581670300355e-07
GC_2_727 b_2 NI_2 NS_727 0 -1.4971145567403596e-05
GC_2_728 b_2 NI_2 NS_728 0 2.4256383700411538e-05
GC_2_729 b_2 NI_2 NS_729 0 1.0744564743488149e-06
GC_2_730 b_2 NI_2 NS_730 0 2.6313448247121744e-06
GC_2_731 b_2 NI_2 NS_731 0 3.0498313594826664e-06
GC_2_732 b_2 NI_2 NS_732 0 1.8288499585978226e-05
GC_2_733 b_2 NI_2 NS_733 0 7.7498869528168542e-06
GC_2_734 b_2 NI_2 NS_734 0 -1.6761099826007991e-06
GC_2_735 b_2 NI_2 NS_735 0 2.9830302135466017e-06
GC_2_736 b_2 NI_2 NS_736 0 -3.4643355292559714e-07
GC_2_737 b_2 NI_2 NS_737 0 7.3243737586906262e-06
GC_2_738 b_2 NI_2 NS_738 0 -4.5247748967194984e-06
GC_2_739 b_2 NI_2 NS_739 0 -8.5040071629311501e-07
GC_2_740 b_2 NI_2 NS_740 0 -5.4040893319202232e-07
GC_2_741 b_2 NI_2 NS_741 0 -1.6433403296149142e-06
GC_2_742 b_2 NI_2 NS_742 0 2.2712868141613826e-07
GC_2_743 b_2 NI_2 NS_743 0 1.5096355901412225e-06
GC_2_744 b_2 NI_2 NS_744 0 1.1119823339675059e-07
GC_2_745 b_2 NI_2 NS_745 0 3.6029706071552695e-06
GC_2_746 b_2 NI_2 NS_746 0 -8.9726882061888266e-07
GC_2_747 b_2 NI_2 NS_747 0 -7.2239132190555617e-08
GC_2_748 b_2 NI_2 NS_748 0 -3.6343486233547505e-07
GC_2_749 b_2 NI_2 NS_749 0 -5.1807472322338076e-07
GC_2_750 b_2 NI_2 NS_750 0 5.4927178351110710e-07
GC_2_751 b_2 NI_2 NS_751 0 2.4014210242824821e-06
GC_2_752 b_2 NI_2 NS_752 0 1.9776803630927372e-07
GC_2_753 b_2 NI_2 NS_753 0 3.3593916205523121e-06
GC_2_754 b_2 NI_2 NS_754 0 -2.8068110404911311e-06
GC_2_755 b_2 NI_2 NS_755 0 -2.6296997882578301e-07
GC_2_756 b_2 NI_2 NS_756 0 -4.3648794398174012e-08
GC_2_757 b_2 NI_2 NS_757 0 7.5093165882650579e-07
GC_2_758 b_2 NI_2 NS_758 0 1.0609989104410428e-06
GC_2_759 b_2 NI_2 NS_759 0 3.5142752808073165e-06
GC_2_760 b_2 NI_2 NS_760 0 7.2317541997660593e-08
GC_2_761 b_2 NI_2 NS_761 0 2.4243670763603613e-06
GC_2_762 b_2 NI_2 NS_762 0 -4.6016436103198682e-06
GC_2_763 b_2 NI_2 NS_763 0 4.5912225370370790e-07
GC_2_764 b_2 NI_2 NS_764 0 1.1635549418280078e-06
GC_2_765 b_2 NI_2 NS_765 0 3.6822517975380021e-06
GC_2_766 b_2 NI_2 NS_766 0 -6.4052937860993710e-07
GC_2_767 b_2 NI_2 NS_767 0 5.5776230227320351e-06
GC_2_768 b_2 NI_2 NS_768 0 -9.4618306718035505e-07
GC_2_769 b_2 NI_2 NS_769 0 -1.6056020974324721e-05
GC_2_770 b_2 NI_2 NS_770 0 -1.0583731514723755e-05
GC_2_771 b_2 NI_2 NS_771 0 9.9491805291303825e-07
GC_2_772 b_2 NI_2 NS_772 0 -7.4396870851722032e-06
GC_2_773 b_2 NI_2 NS_773 0 -6.5942377748439504e-08
GC_2_774 b_2 NI_2 NS_774 0 -1.4872747827613943e-07
GC_2_775 b_2 NI_2 NS_775 0 1.8258042147572597e-06
GC_2_776 b_2 NI_2 NS_776 0 -1.8648513345069797e-06
GC_2_777 b_2 NI_2 NS_777 0 5.4044241914556100e-07
GC_2_778 b_2 NI_2 NS_778 0 -3.3794477374817534e-06
GC_2_779 b_2 NI_2 NS_779 0 3.3892700434864533e-06
GC_2_780 b_2 NI_2 NS_780 0 -1.3110593117844272e-06
GC_2_781 b_2 NI_2 NS_781 0 4.5672059294476322e-06
GC_2_782 b_2 NI_2 NS_782 0 -7.9721498384081721e-07
GC_2_783 b_2 NI_2 NS_783 0 -2.0258037870048441e-07
GC_2_784 b_2 NI_2 NS_784 0 -2.0551945713702369e-07
GC_2_785 b_2 NI_2 NS_785 0 7.0588802684820616e-07
GC_2_786 b_2 NI_2 NS_786 0 1.3963566889670417e-06
GC_2_787 b_2 NI_2 NS_787 0 -7.0583199464074040e-07
GC_2_788 b_2 NI_2 NS_788 0 -1.4718784159130441e-06
GC_2_789 b_2 NI_2 NS_789 0 -6.2725011510701891e-07
GC_2_790 b_2 NI_2 NS_790 0 8.2981048051161381e-07
GC_2_791 b_2 NI_2 NS_791 0 2.2262537396722139e-07
GC_2_792 b_2 NI_2 NS_792 0 6.5365093461954275e-07
GC_2_793 b_2 NI_2 NS_793 0 5.9754305938926936e-07
GC_2_794 b_2 NI_2 NS_794 0 2.1049137021780889e-08
GC_2_795 b_2 NI_2 NS_795 0 1.4042999542042702e-11
GC_2_796 b_2 NI_2 NS_796 0 1.0067811068084359e-12
GC_2_797 b_2 NI_2 NS_797 0 4.3083016999081001e-10
GC_2_798 b_2 NI_2 NS_798 0 1.6517095706668085e-09
GC_2_799 b_2 NI_2 NS_799 0 6.6651390091120995e-05
GC_2_800 b_2 NI_2 NS_800 0 2.1491735470289441e-07
GC_2_801 b_2 NI_2 NS_801 0 2.2385582314026420e-11
GC_2_802 b_2 NI_2 NS_802 0 -9.9158411192619067e-10
GC_2_803 b_2 NI_2 NS_803 0 4.2970867777043392e-07
GC_2_804 b_2 NI_2 NS_804 0 1.8577071549275925e-07
GC_2_805 b_2 NI_2 NS_805 0 6.0303231364804118e-07
GC_2_806 b_2 NI_2 NS_806 0 5.0409507908008327e-07
GC_2_807 b_2 NI_2 NS_807 0 2.9694845315045038e-06
GC_2_808 b_2 NI_2 NS_808 0 -1.5587272831873766e-06
GC_2_809 b_2 NI_2 NS_809 0 -1.1975759032880572e-06
GC_2_810 b_2 NI_2 NS_810 0 -1.1247595618262901e-06
GC_2_811 b_2 NI_2 NS_811 0 2.3738782294223852e-06
GC_2_812 b_2 NI_2 NS_812 0 -8.6541707036134626e-07
GC_2_813 b_2 NI_2 NS_813 0 -2.5702159196746251e-06
GC_2_814 b_2 NI_2 NS_814 0 -6.4135429900295284e-06
GC_2_815 b_2 NI_2 NS_815 0 1.0932674577371273e-07
GC_2_816 b_2 NI_2 NS_816 0 1.6956899255649889e-06
GC_2_817 b_2 NI_2 NS_817 0 -1.7209484409897409e-06
GC_2_818 b_2 NI_2 NS_818 0 5.0733426177017622e-07
GC_2_819 b_2 NI_2 NS_819 0 3.1297098754843176e-06
GC_2_820 b_2 NI_2 NS_820 0 -4.3417947524309823e-06
GC_2_821 b_2 NI_2 NS_821 0 -6.6647729736885000e-06
GC_2_822 b_2 NI_2 NS_822 0 1.1555774680286786e-06
GC_2_823 b_2 NI_2 NS_823 0 -4.7409986507306165e-07
GC_2_824 b_2 NI_2 NS_824 0 1.6879960103636680e-06
GC_2_825 b_2 NI_2 NS_825 0 -2.1234785306110889e-06
GC_2_826 b_2 NI_2 NS_826 0 -4.2598558797826172e-06
GC_2_827 b_2 NI_2 NS_827 0 -2.2157159838621164e-06
GC_2_828 b_2 NI_2 NS_828 0 2.1650792338535210e-06
GC_2_829 b_2 NI_2 NS_829 0 3.1625503122525481e-06
GC_2_830 b_2 NI_2 NS_830 0 3.0747064988599888e-06
GC_2_831 b_2 NI_2 NS_831 0 -6.0917990908137832e-06
GC_2_832 b_2 NI_2 NS_832 0 -4.4592812667806961e-06
GC_2_833 b_2 NI_2 NS_833 0 -1.2974854790708514e-06
GC_2_834 b_2 NI_2 NS_834 0 2.1674364101038580e-06
GC_2_835 b_2 NI_2 NS_835 0 2.8446441055612250e-07
GC_2_836 b_2 NI_2 NS_836 0 -2.8074512685806640e-06
GC_2_837 b_2 NI_2 NS_837 0 -3.1954507512292324e-06
GC_2_838 b_2 NI_2 NS_838 0 1.8332574996962073e-06
GC_2_839 b_2 NI_2 NS_839 0 -3.1171932357648657e-07
GC_2_840 b_2 NI_2 NS_840 0 2.3433548072648849e-06
GC_2_841 b_2 NI_2 NS_841 0 -1.4634078054773629e-06
GC_2_842 b_2 NI_2 NS_842 0 -2.6245703186603722e-06
GC_2_843 b_2 NI_2 NS_843 0 -1.8978822214254370e-06
GC_2_844 b_2 NI_2 NS_844 0 1.3684811477005939e-06
GC_2_845 b_2 NI_2 NS_845 0 1.1604802834171357e-06
GC_2_846 b_2 NI_2 NS_846 0 -6.4651733091833623e-07
GC_2_847 b_2 NI_2 NS_847 0 -3.5975082791493297e-06
GC_2_848 b_2 NI_2 NS_848 0 2.8531232213316487e-07
GC_2_849 b_2 NI_2 NS_849 0 -8.2535291876990135e-07
GC_2_850 b_2 NI_2 NS_850 0 7.2325707151211299e-07
GC_2_851 b_2 NI_2 NS_851 0 -1.8919625459763084e-06
GC_2_852 b_2 NI_2 NS_852 0 -1.3288984113246450e-06
GC_2_853 b_2 NI_2 NS_853 0 -1.4489680149472238e-06
GC_2_854 b_2 NI_2 NS_854 0 5.5809484210612648e-07
GC_2_855 b_2 NI_2 NS_855 0 -1.0695911213046222e-06
GC_2_856 b_2 NI_2 NS_856 0 -5.9316168121813291e-07
GC_2_857 b_2 NI_2 NS_857 0 -2.3263765400405105e-06
GC_2_858 b_2 NI_2 NS_858 0 -6.7330250580343929e-07
GC_2_859 b_2 NI_2 NS_859 0 -2.7997954353571166e-06
GC_2_860 b_2 NI_2 NS_860 0 -5.7610636960952808e-07
GC_2_861 b_2 NI_2 NS_861 0 -2.0698222997692857e-06
GC_2_862 b_2 NI_2 NS_862 0 2.3466868171903605e-07
GC_2_863 b_2 NI_2 NS_863 0 -2.5964214982585391e-06
GC_2_864 b_2 NI_2 NS_864 0 1.0337946502357992e-07
GC_2_865 b_2 NI_2 NS_865 0 -3.9140716066031654e-06
GC_2_866 b_2 NI_2 NS_866 0 -7.2803030927597530e-07
GC_2_867 b_2 NI_2 NS_867 0 -5.2745676303496874e-06
GC_2_868 b_2 NI_2 NS_868 0 1.8892502784242825e-06
GC_2_869 b_2 NI_2 NS_869 0 -2.9583279846254258e-06
GC_2_870 b_2 NI_2 NS_870 0 1.7283196473432765e-06
GC_2_871 b_2 NI_2 NS_871 0 -3.7941645853739669e-06
GC_2_872 b_2 NI_2 NS_872 0 2.9619616956216754e-06
GC_2_873 b_2 NI_2 NS_873 0 -5.2505210474322237e-06
GC_2_874 b_2 NI_2 NS_874 0 1.3684591221162666e-06
GC_2_875 b_2 NI_2 NS_875 0 -2.9715069794637034e-06
GC_2_876 b_2 NI_2 NS_876 0 7.6158265118010663e-06
GC_2_877 b_2 NI_2 NS_877 0 -1.9293754537941810e-06
GC_2_878 b_2 NI_2 NS_878 0 4.3918274340375839e-06
GC_2_879 b_2 NI_2 NS_879 0 1.5652483429145344e-06
GC_2_880 b_2 NI_2 NS_880 0 4.8415894279686688e-06
GC_2_881 b_2 NI_2 NS_881 0 -9.8516279710853324e-07
GC_2_882 b_2 NI_2 NS_882 0 3.6448224555297086e-06
GC_2_883 b_2 NI_2 NS_883 0 -1.0328822506933486e-05
GC_2_884 b_2 NI_2 NS_884 0 3.3088910168695070e-05
GC_2_885 b_2 NI_2 NS_885 0 1.3184333882808799e-06
GC_2_886 b_2 NI_2 NS_886 0 1.2141105086765114e-06
GC_2_887 b_2 NI_2 NS_887 0 -9.3725708105693050e-08
GC_2_888 b_2 NI_2 NS_888 0 8.7540955283798467e-08
GC_2_889 b_2 NI_2 NS_889 0 -3.3374167491612421e-07
GC_2_890 b_2 NI_2 NS_890 0 2.6694957532224243e-06
GC_2_891 b_2 NI_2 NS_891 0 7.2381473657441745e-07
GC_2_892 b_2 NI_2 NS_892 0 1.5751253119483511e-07
GC_2_893 b_2 NI_2 NS_893 0 3.0782505594516152e-06
GC_2_894 b_2 NI_2 NS_894 0 -2.7783591944957311e-06
GC_2_895 b_2 NI_2 NS_895 0 -1.9583439496015484e-07
GC_2_896 b_2 NI_2 NS_896 0 -1.1673003655431016e-05
GC_2_897 b_2 NI_2 NS_897 0 1.9428742222391279e-06
GC_2_898 b_2 NI_2 NS_898 0 -6.7931500062307902e-07
GC_2_899 b_2 NI_2 NS_899 0 4.3055689052218414e-06
GC_2_900 b_2 NI_2 NS_900 0 -1.7836180993988445e-07
GC_2_901 b_2 NI_2 NS_901 0 1.2120141523623256e-06
GC_2_902 b_2 NI_2 NS_902 0 1.8707237607204383e-06
GC_2_903 b_2 NI_2 NS_903 0 1.6462418732088611e-06
GC_2_904 b_2 NI_2 NS_904 0 -7.9777745354164259e-07
GC_2_905 b_2 NI_2 NS_905 0 5.9154556168255298e-07
GC_2_906 b_2 NI_2 NS_906 0 4.7809425097655395e-07
GC_2_907 b_2 NI_2 NS_907 0 6.8253534297053343e-07
GC_2_908 b_2 NI_2 NS_908 0 -9.6305430277920707e-08
GC_2_909 b_2 NI_2 NS_909 0 2.5759382143566203e-11
GC_2_910 b_2 NI_2 NS_910 0 -9.7284717954239938e-11
GC_2_911 b_2 NI_2 NS_911 0 -1.9602989061836594e-09
GC_2_912 b_2 NI_2 NS_912 0 4.2975237764717973e-09
GC_2_913 b_2 NI_2 NS_913 0 -2.7508922052763034e-05
GC_2_914 b_2 NI_2 NS_914 0 -1.0597458287312382e-08
GC_2_915 b_2 NI_2 NS_915 0 1.0238646407598247e-11
GC_2_916 b_2 NI_2 NS_916 0 -5.9557464810675279e-11
GC_2_917 b_2 NI_2 NS_917 0 -6.3653704589666123e-07
GC_2_918 b_2 NI_2 NS_918 0 -1.0748177356444395e-06
GC_2_919 b_2 NI_2 NS_919 0 -1.4323565688762948e-06
GC_2_920 b_2 NI_2 NS_920 0 2.3248382014099810e-06
GC_2_921 b_2 NI_2 NS_921 0 -3.8131237734988199e-06
GC_2_922 b_2 NI_2 NS_922 0 2.1795998807068459e-06
GC_2_923 b_2 NI_2 NS_923 0 1.9255579806869868e-06
GC_2_924 b_2 NI_2 NS_924 0 -2.3466645414956548e-07
GC_2_925 b_2 NI_2 NS_925 0 1.4104719736434773e-06
GC_2_926 b_2 NI_2 NS_926 0 5.7203978535943588e-06
GC_2_927 b_2 NI_2 NS_927 0 3.7052046287584900e-06
GC_2_928 b_2 NI_2 NS_928 0 3.2538242839706593e-06
GC_2_929 b_2 NI_2 NS_929 0 -1.4742156889951279e-06
GC_2_930 b_2 NI_2 NS_930 0 -9.4918496675115681e-07
GC_2_931 b_2 NI_2 NS_931 0 9.7320375229584416e-07
GC_2_932 b_2 NI_2 NS_932 0 -2.1860386396217035e-06
GC_2_933 b_2 NI_2 NS_933 0 6.4354679623061415e-06
GC_2_934 b_2 NI_2 NS_934 0 8.5306761737827501e-06
GC_2_935 b_2 NI_2 NS_935 0 1.3303141618421924e-06
GC_2_936 b_2 NI_2 NS_936 0 -9.3980790802304171e-07
GC_2_937 b_2 NI_2 NS_937 0 1.0706268758807727e-06
GC_2_938 b_2 NI_2 NS_938 0 -1.9034799825205395e-06
GC_2_939 b_2 NI_2 NS_939 0 1.4528565928154613e-05
GC_2_940 b_2 NI_2 NS_940 0 -4.1922350032154194e-06
GC_2_941 b_2 NI_2 NS_941 0 -2.0125078470442396e-07
GC_2_942 b_2 NI_2 NS_942 0 6.7953922563270037e-07
GC_2_943 b_2 NI_2 NS_943 0 4.9185689211490024e-06
GC_2_944 b_2 NI_2 NS_944 0 -2.1983531229219365e-06
GC_2_945 b_2 NI_2 NS_945 0 -7.4682447092262442e-07
GC_2_946 b_2 NI_2 NS_946 0 -1.4996633867449370e-05
GC_2_947 b_2 NI_2 NS_947 0 -7.6209581413551377e-08
GC_2_948 b_2 NI_2 NS_948 0 9.7376823371865617e-07
GC_2_949 b_2 NI_2 NS_949 0 -7.9309861629249349e-06
GC_2_950 b_2 NI_2 NS_950 0 -8.5785743389528530e-06
GC_2_951 b_2 NI_2 NS_951 0 -6.2161152900106812e-07
GC_2_952 b_2 NI_2 NS_952 0 -2.1586599844064495e-06
GC_2_953 b_2 NI_2 NS_953 0 -8.3539927817447303e-09
GC_2_954 b_2 NI_2 NS_954 0 1.2073829248621493e-06
GC_2_955 b_2 NI_2 NS_955 0 -7.7193087237810621e-06
GC_2_956 b_2 NI_2 NS_956 0 1.9618656783549399e-06
GC_2_957 b_2 NI_2 NS_957 0 2.4499709127524057e-07
GC_2_958 b_2 NI_2 NS_958 0 -1.6819644954938615e-06
GC_2_959 b_2 NI_2 NS_959 0 1.1608825696966975e-06
GC_2_960 b_2 NI_2 NS_960 0 3.0678971503349163e-06
GC_2_961 b_2 NI_2 NS_961 0 -9.7670739390748371e-07
GC_2_962 b_2 NI_2 NS_962 0 2.0311639889408109e-06
GC_2_963 b_2 NI_2 NS_963 0 4.5640379539990658e-07
GC_2_964 b_2 NI_2 NS_964 0 -1.2309758687970394e-06
GC_2_965 b_2 NI_2 NS_965 0 3.2453682011166394e-06
GC_2_966 b_2 NI_2 NS_966 0 -8.8263120207557856e-07
GC_2_967 b_2 NI_2 NS_967 0 -1.6147957172388211e-07
GC_2_968 b_2 NI_2 NS_968 0 5.1317112704051707e-07
GC_2_969 b_2 NI_2 NS_969 0 -8.4629639191842616e-07
GC_2_970 b_2 NI_2 NS_970 0 -4.1983599429020138e-07
GC_2_971 b_2 NI_2 NS_971 0 9.9341481865769933e-07
GC_2_972 b_2 NI_2 NS_972 0 -1.2689965157976694e-06
GC_2_973 b_2 NI_2 NS_973 0 1.4441204397436968e-06
GC_2_974 b_2 NI_2 NS_974 0 -5.7045136988017212e-07
GC_2_975 b_2 NI_2 NS_975 0 -3.4126546784858690e-08
GC_2_976 b_2 NI_2 NS_976 0 9.6990932247128628e-08
GC_2_977 b_2 NI_2 NS_977 0 -5.9769069420404148e-07
GC_2_978 b_2 NI_2 NS_978 0 -3.4060902663865262e-07
GC_2_979 b_2 NI_2 NS_979 0 9.6764876660693377e-07
GC_2_980 b_2 NI_2 NS_980 0 -1.0810511075610741e-06
GC_2_981 b_2 NI_2 NS_981 0 1.3955425404753142e-06
GC_2_982 b_2 NI_2 NS_982 0 -1.2449166718245761e-06
GC_2_983 b_2 NI_2 NS_983 0 1.6144774289636528e-07
GC_2_984 b_2 NI_2 NS_984 0 -4.3250650603336581e-08
GC_2_985 b_2 NI_2 NS_985 0 -4.8924862890199979e-07
GC_2_986 b_2 NI_2 NS_986 0 -5.0362145214746667e-07
GC_2_987 b_2 NI_2 NS_987 0 1.0632923605108969e-06
GC_2_988 b_2 NI_2 NS_988 0 -8.0454766664028744e-07
GC_2_989 b_2 NI_2 NS_989 0 1.2280651786767847e-06
GC_2_990 b_2 NI_2 NS_990 0 -2.1206220131127492e-06
GC_2_991 b_2 NI_2 NS_991 0 4.9661651558734029e-07
GC_2_992 b_2 NI_2 NS_992 0 -2.5356650205116670e-07
GC_2_993 b_2 NI_2 NS_993 0 -2.4767997685841302e-07
GC_2_994 b_2 NI_2 NS_994 0 -9.1983803127624398e-07
GC_2_995 b_2 NI_2 NS_995 0 1.9186433827364441e-06
GC_2_996 b_2 NI_2 NS_996 0 -1.0012864395638282e-06
GC_2_997 b_2 NI_2 NS_997 0 -8.0998212494302278e-06
GC_2_998 b_2 NI_2 NS_998 0 -9.1473985001352207e-07
GC_2_999 b_2 NI_2 NS_999 0 -3.1606968397067282e-07
GC_2_1000 b_2 NI_2 NS_1000 0 -3.6265001157662142e-06
GC_2_1001 b_2 NI_2 NS_1001 0 -4.9018415219799729e-08
GC_2_1002 b_2 NI_2 NS_1002 0 -3.3203002681491843e-08
GC_2_1003 b_2 NI_2 NS_1003 0 -1.0293810003620717e-07
GC_2_1004 b_2 NI_2 NS_1004 0 -1.2361463220473070e-06
GC_2_1005 b_2 NI_2 NS_1005 0 -1.0227317970889141e-06
GC_2_1006 b_2 NI_2 NS_1006 0 -6.6783220411544225e-07
GC_2_1007 b_2 NI_2 NS_1007 0 1.4569246945511633e-06
GC_2_1008 b_2 NI_2 NS_1008 0 -7.6152077873564570e-07
GC_2_1009 b_2 NI_2 NS_1009 0 1.9436944987371934e-06
GC_2_1010 b_2 NI_2 NS_1010 0 -1.8722415279397244e-06
GC_2_1011 b_2 NI_2 NS_1011 0 -2.2230874970804511e-07
GC_2_1012 b_2 NI_2 NS_1012 0 3.2515815368862006e-07
GC_2_1013 b_2 NI_2 NS_1013 0 2.1538305907720173e-07
GC_2_1014 b_2 NI_2 NS_1014 0 5.2991254226998600e-07
GC_2_1015 b_2 NI_2 NS_1015 0 -1.0774198666067165e-07
GC_2_1016 b_2 NI_2 NS_1016 0 -2.8383169422512264e-07
GC_2_1017 b_2 NI_2 NS_1017 0 8.1692111392639076e-09
GC_2_1018 b_2 NI_2 NS_1018 0 -9.6164747548183296e-08
GC_2_1019 b_2 NI_2 NS_1019 0 -8.8650340815797607e-08
GC_2_1020 b_2 NI_2 NS_1020 0 4.2005206235258952e-08
GC_2_1021 b_2 NI_2 NS_1021 0 -1.2200393278080286e-07
GC_2_1022 b_2 NI_2 NS_1022 0 -5.3538817591796084e-08
GC_2_1023 b_2 NI_2 NS_1023 0 6.1368478177311984e-12
GC_2_1024 b_2 NI_2 NS_1024 0 -1.6271206019768649e-12
GC_2_1025 b_2 NI_2 NS_1025 0 3.5453162714959252e-10
GC_2_1026 b_2 NI_2 NS_1026 0 6.9229676089785939e-10
GC_2_1027 b_2 NI_2 NS_1027 0 1.3443286591066164e-05
GC_2_1028 b_2 NI_2 NS_1028 0 -5.8799810368818040e-08
GC_2_1029 b_2 NI_2 NS_1029 0 -1.4953926555597338e-11
GC_2_1030 b_2 NI_2 NS_1030 0 1.3605168213287575e-10
GC_2_1031 b_2 NI_2 NS_1031 0 3.6053358753150889e-07
GC_2_1032 b_2 NI_2 NS_1032 0 -1.8115038164155767e-07
GC_2_1033 b_2 NI_2 NS_1033 0 2.8267810900599002e-07
GC_2_1034 b_2 NI_2 NS_1034 0 -3.5350018278176721e-07
GC_2_1035 b_2 NI_2 NS_1035 0 4.9947347174824239e-07
GC_2_1036 b_2 NI_2 NS_1036 0 -1.4260701463557728e-06
GC_2_1037 b_2 NI_2 NS_1037 0 -1.1620830946740480e-06
GC_2_1038 b_2 NI_2 NS_1038 0 -4.7166461198678293e-07
GC_2_1039 b_2 NI_2 NS_1039 0 -3.4835192819467737e-07
GC_2_1040 b_2 NI_2 NS_1040 0 -6.2923206251864981e-07
GC_2_1041 b_2 NI_2 NS_1041 0 -2.5926063427104733e-06
GC_2_1042 b_2 NI_2 NS_1042 0 -6.4982329396946384e-07
GC_2_1043 b_2 NI_2 NS_1043 0 7.1999384734597792e-07
GC_2_1044 b_2 NI_2 NS_1044 0 3.6092312426302965e-07
GC_2_1045 b_2 NI_2 NS_1045 0 -7.3896662075199212e-07
GC_2_1046 b_2 NI_2 NS_1046 0 3.6755301329171026e-07
GC_2_1047 b_2 NI_2 NS_1047 0 -1.0208056756980538e-06
GC_2_1048 b_2 NI_2 NS_1048 0 5.9502488779393783e-07
GC_2_1049 b_2 NI_2 NS_1049 0 -4.1423519585251237e-07
GC_2_1050 b_2 NI_2 NS_1050 0 2.6100158170502966e-07
GC_2_1051 b_2 NI_2 NS_1051 0 -8.5708675784622281e-07
GC_2_1052 b_2 NI_2 NS_1052 0 4.4785383997809174e-07
GC_2_1053 b_2 NI_2 NS_1053 0 1.5654094656157338e-07
GC_2_1054 b_2 NI_2 NS_1054 0 1.1343652134545988e-06
GC_2_1055 b_2 NI_2 NS_1055 0 -5.9604691290274052e-07
GC_2_1056 b_2 NI_2 NS_1056 0 1.1950655657052493e-07
GC_2_1057 b_2 NI_2 NS_1057 0 -1.9175642419314803e-06
GC_2_1058 b_2 NI_2 NS_1058 0 1.2778547598152152e-06
GC_2_1059 b_2 NI_2 NS_1059 0 2.0881303467389491e-06
GC_2_1060 b_2 NI_2 NS_1060 0 2.7546847854629766e-07
GC_2_1061 b_2 NI_2 NS_1061 0 -6.8903156918258435e-07
GC_2_1062 b_2 NI_2 NS_1062 0 1.8923875877891653e-07
GC_2_1063 b_2 NI_2 NS_1063 0 9.8702499774833262e-07
GC_2_1064 b_2 NI_2 NS_1064 0 1.7040544033339144e-06
GC_2_1065 b_2 NI_2 NS_1065 0 -2.2913286719671584e-07
GC_2_1066 b_2 NI_2 NS_1066 0 -5.8920974110383955e-07
GC_2_1067 b_2 NI_2 NS_1067 0 -9.2846695334972176e-07
GC_2_1068 b_2 NI_2 NS_1068 0 4.1750094643629186e-07
GC_2_1069 b_2 NI_2 NS_1069 0 1.4336540955649042e-06
GC_2_1070 b_2 NI_2 NS_1070 0 7.1202858588146108e-07
GC_2_1071 b_2 NI_2 NS_1071 0 -3.3623679245679884e-07
GC_2_1072 b_2 NI_2 NS_1072 0 -2.1999175018858330e-07
GC_2_1073 b_2 NI_2 NS_1073 0 -5.1611380891488108e-08
GC_2_1074 b_2 NI_2 NS_1074 0 1.4321515299777107e-06
GC_2_1075 b_2 NI_2 NS_1075 0 4.8239743516439178e-07
GC_2_1076 b_2 NI_2 NS_1076 0 -7.6567470990908646e-07
GC_2_1077 b_2 NI_2 NS_1077 0 -3.5368866033713721e-07
GC_2_1078 b_2 NI_2 NS_1078 0 4.3186405387376900e-08
GC_2_1079 b_2 NI_2 NS_1079 0 3.2325001434396593e-07
GC_2_1080 b_2 NI_2 NS_1080 0 3.8951617691011563e-07
GC_2_1081 b_2 NI_2 NS_1081 0 -1.4421297378298842e-07
GC_2_1082 b_2 NI_2 NS_1082 0 -1.1106747421118052e-08
GC_2_1083 b_2 NI_2 NS_1083 0 1.4081964288717094e-07
GC_2_1084 b_2 NI_2 NS_1084 0 1.2556229657107889e-07
GC_2_1085 b_2 NI_2 NS_1085 0 -1.9026600156880872e-07
GC_2_1086 b_2 NI_2 NS_1086 0 -6.9780300476069068e-08
GC_2_1087 b_2 NI_2 NS_1087 0 3.9138826974970751e-08
GC_2_1088 b_2 NI_2 NS_1088 0 1.9887773433200087e-07
GC_2_1089 b_2 NI_2 NS_1089 0 -1.1141304676930686e-07
GC_2_1090 b_2 NI_2 NS_1090 0 9.4557682827556229e-09
GC_2_1091 b_2 NI_2 NS_1091 0 4.6234666905744456e-08
GC_2_1092 b_2 NI_2 NS_1092 0 7.7274118748349035e-09
GC_2_1093 b_2 NI_2 NS_1093 0 -2.9801165218328529e-07
GC_2_1094 b_2 NI_2 NS_1094 0 -5.3663208643793118e-08
GC_2_1095 b_2 NI_2 NS_1095 0 -9.1173315554246913e-08
GC_2_1096 b_2 NI_2 NS_1096 0 6.3261914073962288e-08
GC_2_1097 b_2 NI_2 NS_1097 0 -2.3127810893288200e-07
GC_2_1098 b_2 NI_2 NS_1098 0 7.8911622205050031e-08
GC_2_1099 b_2 NI_2 NS_1099 0 -1.3267302404789674e-07
GC_2_1100 b_2 NI_2 NS_1100 0 -6.8277668600850482e-08
GC_2_1101 b_2 NI_2 NS_1101 0 -4.3132410261711414e-07
GC_2_1102 b_2 NI_2 NS_1102 0 -5.7064342384234027e-08
GC_2_1103 b_2 NI_2 NS_1103 0 -4.2194785476566187e-07
GC_2_1104 b_2 NI_2 NS_1104 0 6.4455266595139592e-08
GC_2_1105 b_2 NI_2 NS_1105 0 -4.4334323077985314e-07
GC_2_1106 b_2 NI_2 NS_1106 0 1.4505114094508527e-07
GC_2_1107 b_2 NI_2 NS_1107 0 -5.1253876122343317e-07
GC_2_1108 b_2 NI_2 NS_1108 0 1.0382042858051606e-07
GC_2_1109 b_2 NI_2 NS_1109 0 -9.6705480163560004e-07
GC_2_1110 b_2 NI_2 NS_1110 0 -9.9958288592050460e-08
GC_2_1111 b_2 NI_2 NS_1111 0 2.6356996757142701e-06
GC_2_1112 b_2 NI_2 NS_1112 0 3.0027959200091508e-06
GC_2_1113 b_2 NI_2 NS_1113 0 -6.1775117154675484e-07
GC_2_1114 b_2 NI_2 NS_1114 0 1.0421154476472191e-06
GC_2_1115 b_2 NI_2 NS_1115 0 9.1780980548871867e-09
GC_2_1116 b_2 NI_2 NS_1116 0 2.5495408937644127e-08
GC_2_1117 b_2 NI_2 NS_1117 0 -4.7283643637877157e-07
GC_2_1118 b_2 NI_2 NS_1118 0 8.3077585890271831e-07
GC_2_1119 b_2 NI_2 NS_1119 0 9.5163104834931166e-09
GC_2_1120 b_2 NI_2 NS_1120 0 3.8773674643880595e-07
GC_2_1121 b_2 NI_2 NS_1121 0 -8.7248176210624591e-07
GC_2_1122 b_2 NI_2 NS_1122 0 -7.3605725682289776e-08
GC_2_1123 b_2 NI_2 NS_1123 0 -9.8320735408307547e-07
GC_2_1124 b_2 NI_2 NS_1124 0 -1.8084314256228258e-07
GC_2_1125 b_2 NI_2 NS_1125 0 1.0885127022959826e-07
GC_2_1126 b_2 NI_2 NS_1126 0 -1.4767353714400131e-07
GC_2_1127 b_2 NI_2 NS_1127 0 6.7365673416575397e-08
GC_2_1128 b_2 NI_2 NS_1128 0 1.3222899505792587e-08
GC_2_1129 b_2 NI_2 NS_1129 0 -6.9919532120965149e-08
GC_2_1130 b_2 NI_2 NS_1130 0 1.6104204130988646e-07
GC_2_1131 b_2 NI_2 NS_1131 0 2.8981756188290599e-08
GC_2_1132 b_2 NI_2 NS_1132 0 -4.0222916000207849e-08
GC_2_1133 b_2 NI_2 NS_1133 0 -8.1261213848560592e-08
GC_2_1134 b_2 NI_2 NS_1134 0 1.6009599317785755e-07
GC_2_1135 b_2 NI_2 NS_1135 0 5.6392897117972219e-08
GC_2_1136 b_2 NI_2 NS_1136 0 -1.6240574341618343e-08
GC_2_1137 b_2 NI_2 NS_1137 0 -1.1754894037699271e-11
GC_2_1138 b_2 NI_2 NS_1138 0 5.1377865769960826e-12
GC_2_1139 b_2 NI_2 NS_1139 0 -3.4035926148512298e-10
GC_2_1140 b_2 NI_2 NS_1140 0 -9.7344879290884305e-10
GC_2_1141 b_2 NI_2 NS_1141 0 -1.2624301388947050e-05
GC_2_1142 b_2 NI_2 NS_1142 0 1.6605035165257951e-08
GC_2_1143 b_2 NI_2 NS_1143 0 2.1156629577664854e-11
GC_2_1144 b_2 NI_2 NS_1144 0 -3.0722398633290562e-10
GC_2_1145 b_2 NI_2 NS_1145 0 -3.4970532593843347e-07
GC_2_1146 b_2 NI_2 NS_1146 0 -9.9914995439939111e-07
GC_2_1147 b_2 NI_2 NS_1147 0 -9.3464108741122802e-07
GC_2_1148 b_2 NI_2 NS_1148 0 1.7814211585069677e-06
GC_2_1149 b_2 NI_2 NS_1149 0 -3.3141586806292383e-06
GC_2_1150 b_2 NI_2 NS_1150 0 8.1245822586061759e-07
GC_2_1151 b_2 NI_2 NS_1151 0 9.4712103063257263e-07
GC_2_1152 b_2 NI_2 NS_1152 0 -2.3716196159424203e-07
GC_2_1153 b_2 NI_2 NS_1153 0 5.4159301521075016e-07
GC_2_1154 b_2 NI_2 NS_1154 0 4.5114361135140793e-06
GC_2_1155 b_2 NI_2 NS_1155 0 1.6161387651133794e-06
GC_2_1156 b_2 NI_2 NS_1156 0 3.0361302588018449e-06
GC_2_1157 b_2 NI_2 NS_1157 0 -8.7111953036492395e-07
GC_2_1158 b_2 NI_2 NS_1158 0 -5.9629273272493845e-07
GC_2_1159 b_2 NI_2 NS_1159 0 4.7104036759173226e-07
GC_2_1160 b_2 NI_2 NS_1160 0 -1.1590520673606388e-06
GC_2_1161 b_2 NI_2 NS_1161 0 2.8710413221612542e-06
GC_2_1162 b_2 NI_2 NS_1162 0 1.0312480713973841e-05
GC_2_1163 b_2 NI_2 NS_1163 0 4.5202385033562908e-06
GC_2_1164 b_2 NI_2 NS_1164 0 -7.5372068953807139e-07
GC_2_1165 b_2 NI_2 NS_1165 0 1.6526201801225566e-06
GC_2_1166 b_2 NI_2 NS_1166 0 -4.2690991953935434e-07
GC_2_1167 b_2 NI_2 NS_1167 0 1.6702708240733496e-05
GC_2_1168 b_2 NI_2 NS_1168 0 -4.4193880617204907e-06
GC_2_1169 b_2 NI_2 NS_1169 0 2.2260104326354222e-07
GC_2_1170 b_2 NI_2 NS_1170 0 -1.0410952305169067e-06
GC_2_1171 b_2 NI_2 NS_1171 0 9.3453497632000322e-06
GC_2_1172 b_2 NI_2 NS_1172 0 -7.1207921816839812e-07
GC_2_1173 b_2 NI_2 NS_1173 0 -5.5720390445561965e-06
GC_2_1174 b_2 NI_2 NS_1174 0 -1.9745305001164619e-05
GC_2_1175 b_2 NI_2 NS_1175 0 -6.0170096527701270e-07
GC_2_1176 b_2 NI_2 NS_1176 0 -8.9886614529680733e-07
GC_2_1177 b_2 NI_2 NS_1177 0 -1.1426759357460531e-05
GC_2_1178 b_2 NI_2 NS_1178 0 -1.0985922130551234e-05
GC_2_1179 b_2 NI_2 NS_1179 0 -2.2538843134633765e-06
GC_2_1180 b_2 NI_2 NS_1180 0 2.5922546928373163e-07
GC_2_1181 b_2 NI_2 NS_1181 0 -1.9214949855249674e-06
GC_2_1182 b_2 NI_2 NS_1182 0 -7.8162596592877525e-07
GC_2_1183 b_2 NI_2 NS_1183 0 -9.6669571219765965e-06
GC_2_1184 b_2 NI_2 NS_1184 0 5.8218554538991858e-06
GC_2_1185 b_2 NI_2 NS_1185 0 -2.9987017248958069e-07
GC_2_1186 b_2 NI_2 NS_1186 0 1.6066091324819642e-07
GC_2_1187 b_2 NI_2 NS_1187 0 -1.6024799068673516e-06
GC_2_1188 b_2 NI_2 NS_1188 0 5.7938318339637000e-06
GC_2_1189 b_2 NI_2 NS_1189 0 2.0440915534265262e-06
GC_2_1190 b_2 NI_2 NS_1190 0 1.9749665009256539e-06
GC_2_1191 b_2 NI_2 NS_1191 0 6.0777021516361615e-07
GC_2_1192 b_2 NI_2 NS_1192 0 -8.9639870154055870e-08
GC_2_1193 b_2 NI_2 NS_1193 0 3.3231634983171416e-06
GC_2_1194 b_2 NI_2 NS_1194 0 -4.3001366775514505e-07
GC_2_1195 b_2 NI_2 NS_1195 0 -5.2001361801033780e-08
GC_2_1196 b_2 NI_2 NS_1196 0 3.3450964365307643e-08
GC_2_1197 b_2 NI_2 NS_1197 0 -8.0680299794069427e-07
GC_2_1198 b_2 NI_2 NS_1198 0 -2.3790136138170533e-07
GC_2_1199 b_2 NI_2 NS_1199 0 3.8122934985385072e-07
GC_2_1200 b_2 NI_2 NS_1200 0 -5.1760987527687322e-07
GC_2_1201 b_2 NI_2 NS_1201 0 1.1837436132921259e-06
GC_2_1202 b_2 NI_2 NS_1202 0 -3.2959682556131892e-08
GC_2_1203 b_2 NI_2 NS_1203 0 2.3779791579680737e-08
GC_2_1204 b_2 NI_2 NS_1204 0 4.9143009376544571e-08
GC_2_1205 b_2 NI_2 NS_1205 0 -5.6742768077024496e-07
GC_2_1206 b_2 NI_2 NS_1206 0 -5.4636635665052227e-08
GC_2_1207 b_2 NI_2 NS_1207 0 4.9448331416561021e-07
GC_2_1208 b_2 NI_2 NS_1208 0 -5.0932364531909706e-07
GC_2_1209 b_2 NI_2 NS_1209 0 1.1632153447629343e-06
GC_2_1210 b_2 NI_2 NS_1210 0 -6.8919926909943468e-07
GC_2_1211 b_2 NI_2 NS_1211 0 5.6824274420254855e-08
GC_2_1212 b_2 NI_2 NS_1212 0 3.4948802964509609e-11
GC_2_1213 b_2 NI_2 NS_1213 0 -5.7560681132535920e-07
GC_2_1214 b_2 NI_2 NS_1214 0 -6.5638698022343762e-08
GC_2_1215 b_2 NI_2 NS_1215 0 6.3212230611493758e-07
GC_2_1216 b_2 NI_2 NS_1216 0 -5.0035747673175157e-07
GC_2_1217 b_2 NI_2 NS_1217 0 8.4891803007304569e-07
GC_2_1218 b_2 NI_2 NS_1218 0 -1.3993919976931137e-06
GC_2_1219 b_2 NI_2 NS_1219 0 1.0856745839993926e-07
GC_2_1220 b_2 NI_2 NS_1220 0 -6.0253282435149129e-08
GC_2_1221 b_2 NI_2 NS_1221 0 -3.9935569883638671e-07
GC_2_1222 b_2 NI_2 NS_1222 0 -2.0554161137891716e-07
GC_2_1223 b_2 NI_2 NS_1223 0 1.1352888975133143e-06
GC_2_1224 b_2 NI_2 NS_1224 0 -8.8116737631473315e-07
GC_2_1225 b_2 NI_2 NS_1225 0 -4.1532553362216341e-06
GC_2_1226 b_2 NI_2 NS_1226 0 6.0164525716014825e-07
GC_2_1227 b_2 NI_2 NS_1227 0 -5.6369531774946773e-07
GC_2_1228 b_2 NI_2 NS_1228 0 -1.9351405050868588e-06
GC_2_1229 b_2 NI_2 NS_1229 0 -2.9200051328004840e-08
GC_2_1230 b_2 NI_2 NS_1230 0 -9.6976426056041127e-09
GC_2_1231 b_2 NI_2 NS_1231 0 -3.5883455771398271e-07
GC_2_1232 b_2 NI_2 NS_1232 0 -2.9257611229552754e-07
GC_2_1233 b_2 NI_2 NS_1233 0 -4.7734292842816864e-07
GC_2_1234 b_2 NI_2 NS_1234 0 -1.7399166003996378e-07
GC_2_1235 b_2 NI_2 NS_1235 0 8.5953398371234001e-07
GC_2_1236 b_2 NI_2 NS_1236 0 -7.5679554158193093e-07
GC_2_1237 b_2 NI_2 NS_1237 0 6.0934348841617696e-07
GC_2_1238 b_2 NI_2 NS_1238 0 -1.0781668824622172e-06
GC_2_1239 b_2 NI_2 NS_1239 0 9.0839675592967979e-08
GC_2_1240 b_2 NI_2 NS_1240 0 1.4512025909803173e-07
GC_2_1241 b_2 NI_2 NS_1241 0 1.5784771070563888e-07
GC_2_1242 b_2 NI_2 NS_1242 0 4.4529267731877747e-07
GC_2_1243 b_2 NI_2 NS_1243 0 2.3088285653824172e-08
GC_2_1244 b_2 NI_2 NS_1244 0 -1.6503927986311406e-07
GC_2_1245 b_2 NI_2 NS_1245 0 -3.7569017275980923e-08
GC_2_1246 b_2 NI_2 NS_1246 0 -1.2372632954783143e-07
GC_2_1247 b_2 NI_2 NS_1247 0 -8.6481926392337842e-08
GC_2_1248 b_2 NI_2 NS_1248 0 1.2325197059870009e-07
GC_2_1249 b_2 NI_2 NS_1249 0 -9.0267394135875301e-09
GC_2_1250 b_2 NI_2 NS_1250 0 -3.7854347783692081e-09
GC_2_1251 b_2 NI_2 NS_1251 0 2.2963634837077365e-12
GC_2_1252 b_2 NI_2 NS_1252 0 -3.3972979845764074e-12
GC_2_1253 b_2 NI_2 NS_1253 0 -7.3122637319264288e-10
GC_2_1254 b_2 NI_2 NS_1254 0 -8.2737041404112543e-11
GC_2_1255 b_2 NI_2 NS_1255 0 5.5755233249049324e-06
GC_2_1256 b_2 NI_2 NS_1256 0 -6.0659995502399974e-08
GC_2_1257 b_2 NI_2 NS_1257 0 -3.1618552896067530e-11
GC_2_1258 b_2 NI_2 NS_1258 0 4.1807644493839025e-10
GC_2_1259 b_2 NI_2 NS_1259 0 8.6995342826697660e-08
GC_2_1260 b_2 NI_2 NS_1260 0 -7.3605856807355659e-08
GC_2_1261 b_2 NI_2 NS_1261 0 3.8660217678375328e-09
GC_2_1262 b_2 NI_2 NS_1262 0 8.3839956210091608e-08
GC_2_1263 b_2 NI_2 NS_1263 0 6.3124894410310040e-07
GC_2_1264 b_2 NI_2 NS_1264 0 -8.3236113913339872e-07
GC_2_1265 b_2 NI_2 NS_1265 0 -9.1896948938193899e-07
GC_2_1266 b_2 NI_2 NS_1266 0 7.4767600830941548e-08
GC_2_1267 b_2 NI_2 NS_1267 0 5.4102910042275900e-07
GC_2_1268 b_2 NI_2 NS_1268 0 4.6009580349822230e-08
GC_2_1269 b_2 NI_2 NS_1269 0 -1.3827626199935668e-06
GC_2_1270 b_2 NI_2 NS_1270 0 -9.7963500739675335e-07
GC_2_1271 b_2 NI_2 NS_1271 0 3.0638153973673792e-07
GC_2_1272 b_2 NI_2 NS_1272 0 2.0537911092863431e-07
GC_2_1273 b_2 NI_2 NS_1273 0 -5.6258821460563622e-07
GC_2_1274 b_2 NI_2 NS_1274 0 7.1028200868542315e-07
GC_2_1275 b_2 NI_2 NS_1275 0 1.9977094694063597e-06
GC_2_1276 b_2 NI_2 NS_1276 0 -6.2823252667733160e-07
GC_2_1277 b_2 NI_2 NS_1277 0 -2.6418325397511948e-06
GC_2_1278 b_2 NI_2 NS_1278 0 3.8227294567619549e-07
GC_2_1279 b_2 NI_2 NS_1279 0 4.1279216098346333e-08
GC_2_1280 b_2 NI_2 NS_1280 0 1.4294009844376045e-06
GC_2_1281 b_2 NI_2 NS_1281 0 2.3354973587487856e-07
GC_2_1282 b_2 NI_2 NS_1282 0 -1.8328018888726209e-06
GC_2_1283 b_2 NI_2 NS_1283 0 -8.6530550596159443e-07
GC_2_1284 b_2 NI_2 NS_1284 0 1.3761334683490092e-06
GC_2_1285 b_2 NI_2 NS_1285 0 2.2852342363416874e-06
GC_2_1286 b_2 NI_2 NS_1286 0 2.9655735738289613e-06
GC_2_1287 b_2 NI_2 NS_1287 0 -2.0507619370379609e-06
GC_2_1288 b_2 NI_2 NS_1288 0 -3.4924529704201600e-06
GC_2_1289 b_2 NI_2 NS_1289 0 -2.8718749731831979e-07
GC_2_1290 b_2 NI_2 NS_1290 0 1.5382141646105776e-06
GC_2_1291 b_2 NI_2 NS_1291 0 1.7081594516816934e-06
GC_2_1292 b_2 NI_2 NS_1292 0 -1.8793184495793729e-06
GC_2_1293 b_2 NI_2 NS_1293 0 -1.6427719821182413e-06
GC_2_1294 b_2 NI_2 NS_1294 0 1.0311044448704443e-06
GC_2_1295 b_2 NI_2 NS_1295 0 4.2910644183948357e-07
GC_2_1296 b_2 NI_2 NS_1296 0 1.8543445156432694e-06
GC_2_1297 b_2 NI_2 NS_1297 0 2.5925872988293640e-07
GC_2_1298 b_2 NI_2 NS_1298 0 -2.2599443564932194e-06
GC_2_1299 b_2 NI_2 NS_1299 0 -7.4200626671807644e-07
GC_2_1300 b_2 NI_2 NS_1300 0 9.6144879720118187e-07
GC_2_1301 b_2 NI_2 NS_1301 0 2.0833942470600015e-06
GC_2_1302 b_2 NI_2 NS_1302 0 -1.8913984094096332e-08
GC_2_1303 b_2 NI_2 NS_1303 0 -1.8132846643543070e-06
GC_2_1304 b_2 NI_2 NS_1304 0 -3.2980298542881406e-07
GC_2_1305 b_2 NI_2 NS_1305 0 -9.5351350444908930e-08
GC_2_1306 b_2 NI_2 NS_1306 0 7.6456726018225267e-07
GC_2_1307 b_2 NI_2 NS_1307 0 2.1964087934885977e-07
GC_2_1308 b_2 NI_2 NS_1308 0 -5.5288913064722348e-07
GC_2_1309 b_2 NI_2 NS_1309 0 -2.4027522741763492e-07
GC_2_1310 b_2 NI_2 NS_1310 0 4.2923991682513514e-07
GC_2_1311 b_2 NI_2 NS_1311 0 1.0687595538810058e-07
GC_2_1312 b_2 NI_2 NS_1312 0 -2.2412005325287203e-07
GC_2_1313 b_2 NI_2 NS_1313 0 -4.5513544762560777e-07
GC_2_1314 b_2 NI_2 NS_1314 0 3.0524944485674127e-07
GC_2_1315 b_2 NI_2 NS_1315 0 2.0652151452208203e-07
GC_2_1316 b_2 NI_2 NS_1316 0 1.6753144264659561e-08
GC_2_1317 b_2 NI_2 NS_1317 0 -1.4742341202148027e-07
GC_2_1318 b_2 NI_2 NS_1318 0 1.9350205783788473e-07
GC_2_1319 b_2 NI_2 NS_1319 0 2.4902970825114813e-08
GC_2_1320 b_2 NI_2 NS_1320 0 -1.4137812783569027e-07
GC_2_1321 b_2 NI_2 NS_1321 0 -3.4514292767197126e-07
GC_2_1322 b_2 NI_2 NS_1322 0 2.7931866718646379e-07
GC_2_1323 b_2 NI_2 NS_1323 0 1.1043774217858132e-07
GC_2_1324 b_2 NI_2 NS_1324 0 -2.3194593463466130e-08
GC_2_1325 b_2 NI_2 NS_1325 0 -1.1145133026085654e-07
GC_2_1326 b_2 NI_2 NS_1326 0 2.2574248495932455e-07
GC_2_1327 b_2 NI_2 NS_1327 0 -1.8935198294873309e-08
GC_2_1328 b_2 NI_2 NS_1328 0 -1.6882368292556763e-07
GC_2_1329 b_2 NI_2 NS_1329 0 -2.8639917305756959e-07
GC_2_1330 b_2 NI_2 NS_1330 0 1.8674261379016836e-07
GC_2_1331 b_2 NI_2 NS_1331 0 -1.1162273286388968e-07
GC_2_1332 b_2 NI_2 NS_1332 0 -5.9977948880440899e-08
GC_2_1333 b_2 NI_2 NS_1333 0 -1.7478663285066386e-07
GC_2_1334 b_2 NI_2 NS_1334 0 2.0344659536992369e-07
GC_2_1335 b_2 NI_2 NS_1335 0 -2.9228607105152202e-07
GC_2_1336 b_2 NI_2 NS_1336 0 -3.9974519212994674e-08
GC_2_1337 b_2 NI_2 NS_1337 0 -4.9673892409098923e-07
GC_2_1338 b_2 NI_2 NS_1338 0 5.7782125303590741e-08
GC_2_1339 b_2 NI_2 NS_1339 0 2.7716646177908911e-06
GC_2_1340 b_2 NI_2 NS_1340 0 4.3275028998124637e-07
GC_2_1341 b_2 NI_2 NS_1341 0 -3.2405514259860497e-07
GC_2_1342 b_2 NI_2 NS_1342 0 6.7628446925409451e-07
GC_2_1343 b_2 NI_2 NS_1343 0 1.2397616163885931e-08
GC_2_1344 b_2 NI_2 NS_1344 0 1.2810103880696708e-08
GC_2_1345 b_2 NI_2 NS_1345 0 -6.7256860606633889e-09
GC_2_1346 b_2 NI_2 NS_1346 0 4.6490300825517555e-07
GC_2_1347 b_2 NI_2 NS_1347 0 -1.2602629599951513e-07
GC_2_1348 b_2 NI_2 NS_1348 0 2.6648573241699668e-07
GC_2_1349 b_2 NI_2 NS_1349 0 -4.8106150041836877e-07
GC_2_1350 b_2 NI_2 NS_1350 0 9.8571602757997863e-08
GC_2_1351 b_2 NI_2 NS_1351 0 -9.4580799769025161e-07
GC_2_1352 b_2 NI_2 NS_1352 0 4.8604632934928411e-07
GC_2_1353 b_2 NI_2 NS_1353 0 -1.8710927637909151e-07
GC_2_1354 b_2 NI_2 NS_1354 0 -7.9276884371400712e-08
GC_2_1355 b_2 NI_2 NS_1355 0 1.6398868717794845e-08
GC_2_1356 b_2 NI_2 NS_1356 0 -1.4792164204296224e-07
GC_2_1357 b_2 NI_2 NS_1357 0 8.6143360211949760e-08
GC_2_1358 b_2 NI_2 NS_1358 0 1.0231039009664216e-07
GC_2_1359 b_2 NI_2 NS_1359 0 -1.1792082971010515e-07
GC_2_1360 b_2 NI_2 NS_1360 0 -1.5795717957238686e-07
GC_2_1361 b_2 NI_2 NS_1361 0 -7.0287850399368265e-08
GC_2_1362 b_2 NI_2 NS_1362 0 8.1119490193013362e-08
GC_2_1363 b_2 NI_2 NS_1363 0 -4.4652726918279637e-10
GC_2_1364 b_2 NI_2 NS_1364 0 -3.7628560061260789e-08
GC_2_1365 b_2 NI_2 NS_1365 0 -8.0395725235290242e-12
GC_2_1366 b_2 NI_2 NS_1366 0 7.1577536593994342e-12
GC_2_1367 b_2 NI_2 NS_1367 0 9.6678219865435842e-10
GC_2_1368 b_2 NI_2 NS_1368 0 -3.3560578106431397e-10
GD_2_1 b_2 NI_2 NA_1 0 -4.2260012133238578e-03
GD_2_2 b_2 NI_2 NA_2 0 -8.8592633367534403e-03
GD_2_3 b_2 NI_2 NA_3 0 5.9084076902141743e-04
GD_2_4 b_2 NI_2 NA_4 0 1.3006422094145318e-02
GD_2_5 b_2 NI_2 NA_5 0 2.4205671071134452e-06
GD_2_6 b_2 NI_2 NA_6 0 5.3912438201754411e-06
GD_2_7 b_2 NI_2 NA_7 0 1.0048976273157701e-05
GD_2_8 b_2 NI_2 NA_8 0 -3.6529881331212626e-06
GD_2_9 b_2 NI_2 NA_9 0 5.6280381305120562e-06
GD_2_10 b_2 NI_2 NA_10 0 -1.8797279982086190e-06
GD_2_11 b_2 NI_2 NA_11 0 3.5860932349416339e-06
GD_2_12 b_2 NI_2 NA_12 0 -6.4862658017734116e-07
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 7.7517769892382401e-03
GC_3_2 b_3 NI_3 NS_2 0 -1.6012310598296370e-03
GC_3_3 b_3 NI_3 NS_3 0 -1.2107575693459177e-08
GC_3_4 b_3 NI_3 NS_4 0 -8.8419586339645469e-07
GC_3_5 b_3 NI_3 NS_5 0 1.0389377264044360e-04
GC_3_6 b_3 NI_3 NS_6 0 -5.1165589956097721e-04
GC_3_7 b_3 NI_3 NS_7 0 -1.9366724998170015e-03
GC_3_8 b_3 NI_3 NS_8 0 -5.9740804279262969e-04
GC_3_9 b_3 NI_3 NS_9 0 2.9415452639035252e-03
GC_3_10 b_3 NI_3 NS_10 0 2.2646130437489280e-03
GC_3_11 b_3 NI_3 NS_11 0 -3.5699577116624264e-03
GC_3_12 b_3 NI_3 NS_12 0 -3.0486836651261811e-03
GC_3_13 b_3 NI_3 NS_13 0 -1.7071501711693527e-03
GC_3_14 b_3 NI_3 NS_14 0 5.8436838894655244e-03
GC_3_15 b_3 NI_3 NS_15 0 4.3687530758664958e-03
GC_3_16 b_3 NI_3 NS_16 0 -2.4745966449742120e-03
GC_3_17 b_3 NI_3 NS_17 0 -1.1051197747859390e-04
GC_3_18 b_3 NI_3 NS_18 0 -1.0369086818087733e-04
GC_3_19 b_3 NI_3 NS_19 0 -4.4520053003454458e-03
GC_3_20 b_3 NI_3 NS_20 0 -9.2458240435421392e-04
GC_3_21 b_3 NI_3 NS_21 0 9.1257594130266829e-03
GC_3_22 b_3 NI_3 NS_22 0 1.7785327738560678e-02
GC_3_23 b_3 NI_3 NS_23 0 -4.0274380167704647e-03
GC_3_24 b_3 NI_3 NS_24 0 -1.7847943525223019e-02
GC_3_25 b_3 NI_3 NS_25 0 -8.2175435742190151e-03
GC_3_26 b_3 NI_3 NS_26 0 4.1736391870915114e-03
GC_3_27 b_3 NI_3 NS_27 0 1.7064439478491979e-02
GC_3_28 b_3 NI_3 NS_28 0 -4.4005704986626150e-04
GC_3_29 b_3 NI_3 NS_29 0 -9.2787949549096443e-03
GC_3_30 b_3 NI_3 NS_30 0 -3.2071945491397255e-03
GC_3_31 b_3 NI_3 NS_31 0 -1.3712651080767781e-02
GC_3_32 b_3 NI_3 NS_32 0 2.2836662084688212e-02
GC_3_33 b_3 NI_3 NS_33 0 2.2839357207909895e-02
GC_3_34 b_3 NI_3 NS_34 0 -2.2670702950854743e-02
GC_3_35 b_3 NI_3 NS_35 0 -9.2392572608969731e-03
GC_3_36 b_3 NI_3 NS_36 0 9.0801439911172225e-04
GC_3_37 b_3 NI_3 NS_37 0 1.8480442582964073e-02
GC_3_38 b_3 NI_3 NS_38 0 6.2433937654513055e-03
GC_3_39 b_3 NI_3 NS_39 0 -9.1763268351323351e-03
GC_3_40 b_3 NI_3 NS_40 0 -9.4611046290123246e-03
GC_3_41 b_3 NI_3 NS_41 0 -9.9741852567373432e-03
GC_3_42 b_3 NI_3 NS_42 0 6.3961382742325013e-03
GC_3_43 b_3 NI_3 NS_43 0 1.6838377600001394e-02
GC_3_44 b_3 NI_3 NS_44 0 -4.8507523893213311e-03
GC_3_45 b_3 NI_3 NS_45 0 -7.2149762194087903e-03
GC_3_46 b_3 NI_3 NS_46 0 -3.4093174659699374e-03
GC_3_47 b_3 NI_3 NS_47 0 6.8284576766921672e-03
GC_3_48 b_3 NI_3 NS_48 0 1.3296720246113598e-02
GC_3_49 b_3 NI_3 NS_49 0 -1.8198397302064510e-03
GC_3_50 b_3 NI_3 NS_50 0 -1.4401884745089921e-02
GC_3_51 b_3 NI_3 NS_51 0 -4.9859625636908614e-03
GC_3_52 b_3 NI_3 NS_52 0 1.0394190580275270e-03
GC_3_53 b_3 NI_3 NS_53 0 6.0026878822323892e-03
GC_3_54 b_3 NI_3 NS_54 0 -1.1033368521321026e-03
GC_3_55 b_3 NI_3 NS_55 0 -3.4642734690642769e-03
GC_3_56 b_3 NI_3 NS_56 0 -1.0877136339809536e-03
GC_3_57 b_3 NI_3 NS_57 0 2.7180843308076442e-03
GC_3_58 b_3 NI_3 NS_58 0 -5.0793037662505045e-04
GC_3_59 b_3 NI_3 NS_59 0 -3.2964042584180250e-03
GC_3_60 b_3 NI_3 NS_60 0 -2.8952144389030421e-03
GC_3_61 b_3 NI_3 NS_61 0 2.0160578413310911e-03
GC_3_62 b_3 NI_3 NS_62 0 7.7561498585427267e-04
GC_3_63 b_3 NI_3 NS_63 0 -2.0162392207238701e-03
GC_3_64 b_3 NI_3 NS_64 0 -9.6653809099726470e-04
GC_3_65 b_3 NI_3 NS_65 0 2.1216790656726813e-03
GC_3_66 b_3 NI_3 NS_66 0 -1.4710183178582874e-03
GC_3_67 b_3 NI_3 NS_67 0 -4.1846675847278135e-03
GC_3_68 b_3 NI_3 NS_68 0 -1.8129776189995989e-03
GC_3_69 b_3 NI_3 NS_69 0 2.3699535088033278e-03
GC_3_70 b_3 NI_3 NS_70 0 -3.7091488689194684e-04
GC_3_71 b_3 NI_3 NS_71 0 -3.0171270802953872e-03
GC_3_72 b_3 NI_3 NS_72 0 4.6227948182475231e-04
GC_3_73 b_3 NI_3 NS_73 0 2.7066174872838588e-03
GC_3_74 b_3 NI_3 NS_74 0 -2.7283517220472613e-03
GC_3_75 b_3 NI_3 NS_75 0 -5.0391208837133163e-03
GC_3_76 b_3 NI_3 NS_76 0 -1.2777727075539164e-04
GC_3_77 b_3 NI_3 NS_77 0 2.4350414796758925e-03
GC_3_78 b_3 NI_3 NS_78 0 -2.1722387246576194e-03
GC_3_79 b_3 NI_3 NS_79 0 -3.2447311778377049e-03
GC_3_80 b_3 NI_3 NS_80 0 2.6004814309470046e-03
GC_3_81 b_3 NI_3 NS_81 0 1.7440027553753746e-03
GC_3_82 b_3 NI_3 NS_82 0 -4.7506655304887643e-03
GC_3_83 b_3 NI_3 NS_83 0 -3.6334488805848104e-03
GC_3_84 b_3 NI_3 NS_84 0 2.5968948699984350e-03
GC_3_85 b_3 NI_3 NS_85 0 -2.8337756435550185e-03
GC_3_86 b_3 NI_3 NS_86 0 3.9869978363562290e-03
GC_3_87 b_3 NI_3 NS_87 0 -2.2097304216610415e-04
GC_3_88 b_3 NI_3 NS_88 0 -4.2143932075885916e-03
GC_3_89 b_3 NI_3 NS_89 0 -9.9004949439867979e-06
GC_3_90 b_3 NI_3 NS_90 0 7.5068447616220956e-06
GC_3_91 b_3 NI_3 NS_91 0 -1.3536752743014851e-03
GC_3_92 b_3 NI_3 NS_92 0 3.3750369237701989e-03
GC_3_93 b_3 NI_3 NS_93 0 -9.6981086333022349e-04
GC_3_94 b_3 NI_3 NS_94 0 -4.3483886235214436e-03
GC_3_95 b_3 NI_3 NS_95 0 -1.0004295435909370e-03
GC_3_96 b_3 NI_3 NS_96 0 2.2215355649961854e-03
GC_3_97 b_3 NI_3 NS_97 0 -1.6509350054067929e-03
GC_3_98 b_3 NI_3 NS_98 0 -4.4091720645970207e-03
GC_3_99 b_3 NI_3 NS_99 0 -1.4483889277918862e-03
GC_3_100 b_3 NI_3 NS_100 0 -2.4971171243885299e-03
GC_3_101 b_3 NI_3 NS_101 0 7.8206441137250839e-04
GC_3_102 b_3 NI_3 NS_102 0 2.5934686440194435e-03
GC_3_103 b_3 NI_3 NS_103 0 -6.9629932708796950e-04
GC_3_104 b_3 NI_3 NS_104 0 2.8791308473661288e-03
GC_3_105 b_3 NI_3 NS_105 0 -1.4354331588806500e-03
GC_3_106 b_3 NI_3 NS_106 0 -2.7718926022085749e-03
GC_3_107 b_3 NI_3 NS_107 0 -1.1678459039075461e-03
GC_3_108 b_3 NI_3 NS_108 0 2.6661739433018637e-03
GC_3_109 b_3 NI_3 NS_109 0 7.8077002198028551e-04
GC_3_110 b_3 NI_3 NS_110 0 -1.8746307422856296e-03
GC_3_111 b_3 NI_3 NS_111 0 2.3791410540050171e-08
GC_3_112 b_3 NI_3 NS_112 0 -6.0255378893479960e-08
GC_3_113 b_3 NI_3 NS_113 0 -9.0379195267616550e-07
GC_3_114 b_3 NI_3 NS_114 0 3.2032331566090646e-06
GC_3_115 b_3 NI_3 NS_115 0 2.9495780771876161e-03
GC_3_116 b_3 NI_3 NS_116 0 -6.1234120038294231e-04
GC_3_117 b_3 NI_3 NS_117 0 2.7949880405130853e-08
GC_3_118 b_3 NI_3 NS_118 0 -3.1702428509748000e-08
GC_3_119 b_3 NI_3 NS_119 0 2.0347277955968312e-04
GC_3_120 b_3 NI_3 NS_120 0 1.3799474012533288e-04
GC_3_121 b_3 NI_3 NS_121 0 5.6259278157525829e-04
GC_3_122 b_3 NI_3 NS_122 0 2.6570818081323577e-04
GC_3_123 b_3 NI_3 NS_123 0 3.1064667490479213e-03
GC_3_124 b_3 NI_3 NS_124 0 -2.2048923669259839e-03
GC_3_125 b_3 NI_3 NS_125 0 -1.5822543587228545e-03
GC_3_126 b_3 NI_3 NS_126 0 -2.6870784628982231e-03
GC_3_127 b_3 NI_3 NS_127 0 -2.0496561789789657e-03
GC_3_128 b_3 NI_3 NS_128 0 -3.7885102939486178e-03
GC_3_129 b_3 NI_3 NS_129 0 -4.9745615281467630e-03
GC_3_130 b_3 NI_3 NS_130 0 -1.5415296228933743e-03
GC_3_131 b_3 NI_3 NS_131 0 2.9290597692236916e-04
GC_3_132 b_3 NI_3 NS_132 0 1.9565110676163995e-04
GC_3_133 b_3 NI_3 NS_133 0 -2.8663287023517753e-03
GC_3_134 b_3 NI_3 NS_134 0 -9.5746369995463492e-04
GC_3_135 b_3 NI_3 NS_135 0 -2.2151869997411762e-02
GC_3_136 b_3 NI_3 NS_136 0 -1.0226316081185899e-02
GC_3_137 b_3 NI_3 NS_137 0 1.1324964603897703e-03
GC_3_138 b_3 NI_3 NS_138 0 2.0395319725874377e-02
GC_3_139 b_3 NI_3 NS_139 0 -5.8416210211683205e-03
GC_3_140 b_3 NI_3 NS_140 0 4.6116288203687465e-03
GC_3_141 b_3 NI_3 NS_141 0 5.7171497801127577e-03
GC_3_142 b_3 NI_3 NS_142 0 3.4516070767437630e-02
GC_3_143 b_3 NI_3 NS_143 0 8.0342761942350412e-03
GC_3_144 b_3 NI_3 NS_144 0 2.7930240341847603e-03
GC_3_145 b_3 NI_3 NS_145 0 -7.7724215056918745e-03
GC_3_146 b_3 NI_3 NS_146 0 2.9556754316452234e-02
GC_3_147 b_3 NI_3 NS_147 0 5.0768430140120953e-02
GC_3_148 b_3 NI_3 NS_148 0 -2.0072961081372680e-02
GC_3_149 b_3 NI_3 NS_149 0 7.9195785247055343e-03
GC_3_150 b_3 NI_3 NS_150 0 -1.6364409960749717e-03
GC_3_151 b_3 NI_3 NS_151 0 2.9084859999523156e-02
GC_3_152 b_3 NI_3 NS_152 0 -2.6464736579857914e-02
GC_3_153 b_3 NI_3 NS_153 0 -6.7250676971983159e-03
GC_3_154 b_3 NI_3 NS_154 0 -9.8822057161725898e-03
GC_3_155 b_3 NI_3 NS_155 0 8.4630826858443364e-03
GC_3_156 b_3 NI_3 NS_156 0 -8.0277980819230942e-03
GC_3_157 b_3 NI_3 NS_157 0 -1.8994952659545723e-02
GC_3_158 b_3 NI_3 NS_158 0 -2.5238422114712968e-02
GC_3_159 b_3 NI_3 NS_159 0 -5.4717850907585602e-03
GC_3_160 b_3 NI_3 NS_160 0 -2.8547841777828140e-03
GC_3_161 b_3 NI_3 NS_161 0 -1.7741074128875482e-02
GC_3_162 b_3 NI_3 NS_162 0 -1.3132230468874805e-02
GC_3_163 b_3 NI_3 NS_163 0 -4.8178007864756759e-03
GC_3_164 b_3 NI_3 NS_164 0 1.2541404248319052e-02
GC_3_165 b_3 NI_3 NS_165 0 -3.4590901695808660e-03
GC_3_166 b_3 NI_3 NS_166 0 1.5412380182272221e-03
GC_3_167 b_3 NI_3 NS_167 0 -7.1865217804843783e-04
GC_3_168 b_3 NI_3 NS_168 0 7.0058606362865114e-03
GC_3_169 b_3 NI_3 NS_169 0 1.8820411282429721e-03
GC_3_170 b_3 NI_3 NS_170 0 8.5748801406228427e-05
GC_3_171 b_3 NI_3 NS_171 0 3.1400256708056102e-04
GC_3_172 b_3 NI_3 NS_172 0 -1.9467011502516422e-03
GC_3_173 b_3 NI_3 NS_173 0 -1.8563356146475041e-03
GC_3_174 b_3 NI_3 NS_174 0 -1.6182086466213538e-03
GC_3_175 b_3 NI_3 NS_175 0 -2.1290963626111343e-03
GC_3_176 b_3 NI_3 NS_176 0 1.6850438900593251e-03
GC_3_177 b_3 NI_3 NS_177 0 7.6361034735872334e-04
GC_3_178 b_3 NI_3 NS_178 0 1.8527544698305616e-04
GC_3_179 b_3 NI_3 NS_179 0 -6.9730352416525398e-04
GC_3_180 b_3 NI_3 NS_180 0 -1.6780698218557763e-03
GC_3_181 b_3 NI_3 NS_181 0 -2.6815283765594714e-03
GC_3_182 b_3 NI_3 NS_182 0 -8.2749104602475028e-04
GC_3_183 b_3 NI_3 NS_183 0 -4.9989643487842689e-04
GC_3_184 b_3 NI_3 NS_184 0 2.9288646763956845e-03
GC_3_185 b_3 NI_3 NS_185 0 1.3533577793804590e-03
GC_3_186 b_3 NI_3 NS_186 0 -8.5805557058709974e-04
GC_3_187 b_3 NI_3 NS_187 0 -2.4189241797636847e-03
GC_3_188 b_3 NI_3 NS_188 0 -2.2676207872960748e-03
GC_3_189 b_3 NI_3 NS_189 0 -3.5540452695985770e-03
GC_3_190 b_3 NI_3 NS_190 0 7.4852702289969258e-04
GC_3_191 b_3 NI_3 NS_191 0 2.4633835860143798e-03
GC_3_192 b_3 NI_3 NS_192 0 3.0182798446697673e-03
GC_3_193 b_3 NI_3 NS_193 0 9.8455419001531003e-04
GC_3_194 b_3 NI_3 NS_194 0 -2.9418100597726846e-03
GC_3_195 b_3 NI_3 NS_195 0 -4.7678000282342231e-03
GC_3_196 b_3 NI_3 NS_196 0 5.4340226341034482e-05
GC_3_197 b_3 NI_3 NS_197 0 -1.7083703559314400e-03
GC_3_198 b_3 NI_3 NS_198 0 3.7124270186457320e-03
GC_3_199 b_3 NI_3 NS_199 0 -7.6587642478235444e-04
GC_3_200 b_3 NI_3 NS_200 0 1.5006814281130426e-03
GC_3_201 b_3 NI_3 NS_201 0 3.2213016762664623e-03
GC_3_202 b_3 NI_3 NS_202 0 -1.3508683618631398e-03
GC_3_203 b_3 NI_3 NS_203 0 -2.9326073204834440e-06
GC_3_204 b_3 NI_3 NS_204 0 8.7469700940414424e-06
GC_3_205 b_3 NI_3 NS_205 0 -1.8200418589312810e-03
GC_3_206 b_3 NI_3 NS_206 0 -2.5277363330337846e-03
GC_3_207 b_3 NI_3 NS_207 0 -2.4072534022134932e-03
GC_3_208 b_3 NI_3 NS_208 0 2.4886635219990255e-03
GC_3_209 b_3 NI_3 NS_209 0 1.0142619058303764e-03
GC_3_210 b_3 NI_3 NS_210 0 2.4256812106000798e-03
GC_3_211 b_3 NI_3 NS_211 0 8.5775930731191098e-04
GC_3_212 b_3 NI_3 NS_212 0 -2.6994852838280107e-03
GC_3_213 b_3 NI_3 NS_213 0 -3.0644787427663042e-04
GC_3_214 b_3 NI_3 NS_214 0 1.6741356684409332e-03
GC_3_215 b_3 NI_3 NS_215 0 -1.7840540721603864e-03
GC_3_216 b_3 NI_3 NS_216 0 -3.1181081265208580e-04
GC_3_217 b_3 NI_3 NS_217 0 1.4004539639447993e-03
GC_3_218 b_3 NI_3 NS_218 0 1.9709615764259185e-03
GC_3_219 b_3 NI_3 NS_219 0 1.0449287327084374e-03
GC_3_220 b_3 NI_3 NS_220 0 -2.2998045694717106e-03
GC_3_221 b_3 NI_3 NS_221 0 -6.9799494695637059e-04
GC_3_222 b_3 NI_3 NS_222 0 -1.4668898807674452e-03
GC_3_223 b_3 NI_3 NS_223 0 -1.3735491340989556e-03
GC_3_224 b_3 NI_3 NS_224 0 -3.1252861594881979e-04
GC_3_225 b_3 NI_3 NS_225 0 7.1030059129532425e-09
GC_3_226 b_3 NI_3 NS_226 0 -2.4710001567883010e-08
GC_3_227 b_3 NI_3 NS_227 0 -4.5275408315141393e-07
GC_3_228 b_3 NI_3 NS_228 0 1.6341838969925549e-06
GC_3_229 b_3 NI_3 NS_229 0 -1.4190097407435300e-02
GC_3_230 b_3 NI_3 NS_230 0 1.3879298607381572e-03
GC_3_231 b_3 NI_3 NS_231 0 -2.6214589268038936e-07
GC_3_232 b_3 NI_3 NS_232 0 -3.7469053601664712e-06
GC_3_233 b_3 NI_3 NS_233 0 -2.9950712352343694e-04
GC_3_234 b_3 NI_3 NS_234 0 4.7112868964960524e-04
GC_3_235 b_3 NI_3 NS_235 0 1.2936041298229283e-03
GC_3_236 b_3 NI_3 NS_236 0 5.6342135820495369e-04
GC_3_237 b_3 NI_3 NS_237 0 -2.7928189552435317e-03
GC_3_238 b_3 NI_3 NS_238 0 -7.1086086409688195e-04
GC_3_239 b_3 NI_3 NS_239 0 3.5977247957131326e-03
GC_3_240 b_3 NI_3 NS_240 0 2.5454554772647471e-03
GC_3_241 b_3 NI_3 NS_241 0 1.1770627409826854e-03
GC_3_242 b_3 NI_3 NS_242 0 -4.1367871145994196e-03
GC_3_243 b_3 NI_3 NS_243 0 -1.5548935818197106e-03
GC_3_244 b_3 NI_3 NS_244 0 2.7530038112826439e-03
GC_3_245 b_3 NI_3 NS_245 0 -3.5992609246651252e-04
GC_3_246 b_3 NI_3 NS_246 0 -2.1737785181827045e-04
GC_3_247 b_3 NI_3 NS_247 0 4.0014076268810655e-03
GC_3_248 b_3 NI_3 NS_248 0 2.5737083876034187e-04
GC_3_249 b_3 NI_3 NS_249 0 -7.3983785450492633e-03
GC_3_250 b_3 NI_3 NS_250 0 -1.3542083605378757e-02
GC_3_251 b_3 NI_3 NS_251 0 4.4843084901327480e-03
GC_3_252 b_3 NI_3 NS_252 0 1.3402111987595930e-02
GC_3_253 b_3 NI_3 NS_253 0 6.7170381911766195e-03
GC_3_254 b_3 NI_3 NS_254 0 -4.0292251491291665e-03
GC_3_255 b_3 NI_3 NS_255 0 -1.3321384901694924e-02
GC_3_256 b_3 NI_3 NS_256 0 6.8614002187367097e-04
GC_3_257 b_3 NI_3 NS_257 0 7.8581343523568201e-03
GC_3_258 b_3 NI_3 NS_258 0 1.8345313325804735e-03
GC_3_259 b_3 NI_3 NS_259 0 1.0514025121400934e-02
GC_3_260 b_3 NI_3 NS_260 0 -1.9642822930251404e-02
GC_3_261 b_3 NI_3 NS_261 0 -1.7746432280186474e-02
GC_3_262 b_3 NI_3 NS_262 0 1.9129827664865109e-02
GC_3_263 b_3 NI_3 NS_263 0 7.6846954657520698e-03
GC_3_264 b_3 NI_3 NS_264 0 -1.4647961155202314e-03
GC_3_265 b_3 NI_3 NS_265 0 -1.5663694621543784e-02
GC_3_266 b_3 NI_3 NS_266 0 -4.7646805759046984e-03
GC_3_267 b_3 NI_3 NS_267 0 8.0859900445670249e-03
GC_3_268 b_3 NI_3 NS_268 0 7.2458421625027671e-03
GC_3_269 b_3 NI_3 NS_269 0 8.1137552717649320e-03
GC_3_270 b_3 NI_3 NS_270 0 -6.0473597232078811e-03
GC_3_271 b_3 NI_3 NS_271 0 -1.3987021078502184e-02
GC_3_272 b_3 NI_3 NS_272 0 4.5766954769181798e-03
GC_3_273 b_3 NI_3 NS_273 0 6.2436852783541840e-03
GC_3_274 b_3 NI_3 NS_274 0 2.3779905771676609e-03
GC_3_275 b_3 NI_3 NS_275 0 -6.3098278837882514e-03
GC_3_276 b_3 NI_3 NS_276 0 -1.1127822870543303e-02
GC_3_277 b_3 NI_3 NS_277 0 2.1503423919028179e-03
GC_3_278 b_3 NI_3 NS_278 0 1.1938071371307748e-02
GC_3_279 b_3 NI_3 NS_279 0 4.2146499023713591e-03
GC_3_280 b_3 NI_3 NS_280 0 -1.1800102681177004e-03
GC_3_281 b_3 NI_3 NS_281 0 -4.9267499346084447e-03
GC_3_282 b_3 NI_3 NS_282 0 1.0434774616390379e-03
GC_3_283 b_3 NI_3 NS_283 0 3.0295902964153701e-03
GC_3_284 b_3 NI_3 NS_284 0 6.8509536985503065e-04
GC_3_285 b_3 NI_3 NS_285 0 -2.2185452352903035e-03
GC_3_286 b_3 NI_3 NS_286 0 4.8987912710520085e-04
GC_3_287 b_3 NI_3 NS_287 0 3.0814361201426670e-03
GC_3_288 b_3 NI_3 NS_288 0 2.2937716711490682e-03
GC_3_289 b_3 NI_3 NS_289 0 -1.5261901203590758e-03
GC_3_290 b_3 NI_3 NS_290 0 -6.8311371182555743e-04
GC_3_291 b_3 NI_3 NS_291 0 1.8943361597397530e-03
GC_3_292 b_3 NI_3 NS_292 0 6.7631458979500419e-04
GC_3_293 b_3 NI_3 NS_293 0 -1.5560152057580235e-03
GC_3_294 b_3 NI_3 NS_294 0 1.2187733574392601e-03
GC_3_295 b_3 NI_3 NS_295 0 3.9927794716663675e-03
GC_3_296 b_3 NI_3 NS_296 0 1.4034783070292723e-03
GC_3_297 b_3 NI_3 NS_297 0 -1.5356610430749700e-03
GC_3_298 b_3 NI_3 NS_298 0 5.9545100615131318e-05
GC_3_299 b_3 NI_3 NS_299 0 2.8410904467837195e-03
GC_3_300 b_3 NI_3 NS_300 0 -6.9178188501826401e-04
GC_3_301 b_3 NI_3 NS_301 0 -1.8626355231402562e-03
GC_3_302 b_3 NI_3 NS_302 0 1.9986033064253060e-03
GC_3_303 b_3 NI_3 NS_303 0 4.9308303887853518e-03
GC_3_304 b_3 NI_3 NS_304 0 -1.7294499576135680e-04
GC_3_305 b_3 NI_3 NS_305 0 -1.6210986159472445e-03
GC_3_306 b_3 NI_3 NS_306 0 9.0628943582777308e-04
GC_3_307 b_3 NI_3 NS_307 0 3.0921495452636998e-03
GC_3_308 b_3 NI_3 NS_308 0 -2.8475032012458220e-03
GC_3_309 b_3 NI_3 NS_309 0 -1.4246752536775250e-03
GC_3_310 b_3 NI_3 NS_310 0 3.1958050728670873e-03
GC_3_311 b_3 NI_3 NS_311 0 3.8550118525597847e-03
GC_3_312 b_3 NI_3 NS_312 0 -2.9522342675832557e-03
GC_3_313 b_3 NI_3 NS_313 0 -2.0071644383908970e-03
GC_3_314 b_3 NI_3 NS_314 0 -4.1861153497111765e-03
GC_3_315 b_3 NI_3 NS_315 0 -3.5104564331051198e-04
GC_3_316 b_3 NI_3 NS_316 0 2.2864791444868111e-03
GC_3_317 b_3 NI_3 NS_317 0 -1.0763134239394421e-05
GC_3_318 b_3 NI_3 NS_318 0 -2.3358060973476260e-05
GC_3_319 b_3 NI_3 NS_319 0 8.7769866723416494e-04
GC_3_320 b_3 NI_3 NS_320 0 -3.8352026116396528e-03
GC_3_321 b_3 NI_3 NS_321 0 3.5234563946015437e-04
GC_3_322 b_3 NI_3 NS_322 0 3.3067902032369221e-03
GC_3_323 b_3 NI_3 NS_323 0 1.3988544772359651e-03
GC_3_324 b_3 NI_3 NS_324 0 -2.3422177471358872e-03
GC_3_325 b_3 NI_3 NS_325 0 2.2595445985145873e-03
GC_3_326 b_3 NI_3 NS_326 0 3.3689528580504711e-03
GC_3_327 b_3 NI_3 NS_327 0 1.1614257540535577e-03
GC_3_328 b_3 NI_3 NS_328 0 2.4048218341710145e-03
GC_3_329 b_3 NI_3 NS_329 0 -8.2758873323753349e-04
GC_3_330 b_3 NI_3 NS_330 0 -1.9684501755091719e-03
GC_3_331 b_3 NI_3 NS_331 0 3.9844979260028602e-04
GC_3_332 b_3 NI_3 NS_332 0 -2.6910253245430076e-03
GC_3_333 b_3 NI_3 NS_333 0 9.7822596634247641e-04
GC_3_334 b_3 NI_3 NS_334 0 2.7413579780172590e-03
GC_3_335 b_3 NI_3 NS_335 0 1.0427092325713877e-03
GC_3_336 b_3 NI_3 NS_336 0 -2.4233094973752515e-03
GC_3_337 b_3 NI_3 NS_337 0 -1.0796403751135034e-03
GC_3_338 b_3 NI_3 NS_338 0 1.5897875189545480e-03
GC_3_339 b_3 NI_3 NS_339 0 -1.0824816241029396e-08
GC_3_340 b_3 NI_3 NS_340 0 -2.6618453096243945e-09
GC_3_341 b_3 NI_3 NS_341 0 2.3026497631555775e-06
GC_3_342 b_3 NI_3 NS_342 0 5.5056417255638653e-07
GC_3_343 b_3 NI_3 NS_343 0 1.8439732050886663e-02
GC_3_344 b_3 NI_3 NS_344 0 6.7473516467850912e-03
GC_3_345 b_3 NI_3 NS_345 0 4.6777094553014474e-07
GC_3_346 b_3 NI_3 NS_346 0 1.4628681236597617e-06
GC_3_347 b_3 NI_3 NS_347 0 6.0883416002558664e-03
GC_3_348 b_3 NI_3 NS_348 0 1.8079590327079135e-03
GC_3_349 b_3 NI_3 NS_349 0 -6.0693295988834273e-03
GC_3_350 b_3 NI_3 NS_350 0 -6.1755942167906021e-04
GC_3_351 b_3 NI_3 NS_351 0 7.3051642846782309e-03
GC_3_352 b_3 NI_3 NS_352 0 -1.2868565260674505e-02
GC_3_353 b_3 NI_3 NS_353 0 8.4478581794454333e-03
GC_3_354 b_3 NI_3 NS_354 0 -2.4311026053824210e-04
GC_3_355 b_3 NI_3 NS_355 0 -9.6438123284267145e-03
GC_3_356 b_3 NI_3 NS_356 0 2.6146474934407994e-03
GC_3_357 b_3 NI_3 NS_357 0 -8.8620363499959786e-03
GC_3_358 b_3 NI_3 NS_358 0 -2.4394077892382376e-02
GC_3_359 b_3 NI_3 NS_359 0 -8.6181026448399771e-04
GC_3_360 b_3 NI_3 NS_360 0 4.1810317531879209e-03
GC_3_361 b_3 NI_3 NS_361 0 7.1874271616436912e-03
GC_3_362 b_3 NI_3 NS_362 0 -1.0295512874949240e-03
GC_3_363 b_3 NI_3 NS_363 0 -2.5160943084511167e-02
GC_3_364 b_3 NI_3 NS_364 0 4.8305095271545823e-03
GC_3_365 b_3 NI_3 NS_365 0 -1.9677178361332145e-02
GC_3_366 b_3 NI_3 NS_366 0 8.9681213462700310e-04
GC_3_367 b_3 NI_3 NS_367 0 1.0760395267912655e-02
GC_3_368 b_3 NI_3 NS_368 0 -2.7835058051904320e-03
GC_3_369 b_3 NI_3 NS_369 0 -4.7876583750650009e-03
GC_3_370 b_3 NI_3 NS_370 0 4.5022298525782094e-02
GC_3_371 b_3 NI_3 NS_371 0 -1.2656498028025860e-02
GC_3_372 b_3 NI_3 NS_372 0 -2.7342535053084116e-04
GC_3_373 b_3 NI_3 NS_373 0 1.5916844056148061e-02
GC_3_374 b_3 NI_3 NS_374 0 -4.0521908129402288e-03
GC_3_375 b_3 NI_3 NS_375 0 3.2200863646357887e-02
GC_3_376 b_3 NI_3 NS_376 0 1.8584663883318416e-02
GC_3_377 b_3 NI_3 NS_377 0 -1.2597877463723353e-02
GC_3_378 b_3 NI_3 NS_378 0 1.6054731149283208e-04
GC_3_379 b_3 NI_3 NS_379 0 1.7204374242405764e-02
GC_3_380 b_3 NI_3 NS_380 0 -3.5163088457902440e-02
GC_3_381 b_3 NI_3 NS_381 0 1.4015863108230497e-02
GC_3_382 b_3 NI_3 NS_382 0 4.7859367525480189e-03
GC_3_383 b_3 NI_3 NS_383 0 -1.4402596582444907e-02
GC_3_384 b_3 NI_3 NS_384 0 2.3855243174216744e-04
GC_3_385 b_3 NI_3 NS_385 0 -2.0144415228540553e-02
GC_3_386 b_3 NI_3 NS_386 0 -3.0186763265967857e-02
GC_3_387 b_3 NI_3 NS_387 0 1.0530804791871609e-02
GC_3_388 b_3 NI_3 NS_388 0 3.5935490856946290e-03
GC_3_389 b_3 NI_3 NS_389 0 -2.6797826099077049e-02
GC_3_390 b_3 NI_3 NS_390 0 1.1150421168090745e-02
GC_3_391 b_3 NI_3 NS_391 0 -1.4133899634061442e-02
GC_3_392 b_3 NI_3 NS_392 0 -2.5194465683331915e-03
GC_3_393 b_3 NI_3 NS_393 0 7.5552516111377912e-03
GC_3_394 b_3 NI_3 NS_394 0 1.5923641786957760e-03
GC_3_395 b_3 NI_3 NS_395 0 -8.5561070558516346e-04
GC_3_396 b_3 NI_3 NS_396 0 2.4403099822878860e-02
GC_3_397 b_3 NI_3 NS_397 0 -7.6201959656694027e-03
GC_3_398 b_3 NI_3 NS_398 0 2.8212556097770064e-04
GC_3_399 b_3 NI_3 NS_399 0 -5.5980892342308514e-04
GC_3_400 b_3 NI_3 NS_400 0 -5.5368739005439670e-03
GC_3_401 b_3 NI_3 NS_401 0 8.2659996006846370e-03
GC_3_402 b_3 NI_3 NS_402 0 7.0201265002174419e-03
GC_3_403 b_3 NI_3 NS_403 0 -7.1918032335592974e-04
GC_3_404 b_3 NI_3 NS_404 0 1.2092493381636669e-02
GC_3_405 b_3 NI_3 NS_405 0 -5.1474392801595346e-03
GC_3_406 b_3 NI_3 NS_406 0 -1.3699545860260928e-04
GC_3_407 b_3 NI_3 NS_407 0 -1.8303992654257152e-03
GC_3_408 b_3 NI_3 NS_408 0 -5.1700675470025140e-03
GC_3_409 b_3 NI_3 NS_409 0 9.2878958000223895e-03
GC_3_410 b_3 NI_3 NS_410 0 5.4154508517489887e-03
GC_3_411 b_3 NI_3 NS_411 0 3.5152715797918638e-03
GC_3_412 b_3 NI_3 NS_412 0 1.1689821183028292e-02
GC_3_413 b_3 NI_3 NS_413 0 -6.1370084907515603e-03
GC_3_414 b_3 NI_3 NS_414 0 1.4286475674857805e-03
GC_3_415 b_3 NI_3 NS_415 0 -2.8171558770673970e-03
GC_3_416 b_3 NI_3 NS_416 0 -7.3462416947635244e-03
GC_3_417 b_3 NI_3 NS_417 0 9.9561294098873994e-03
GC_3_418 b_3 NI_3 NS_418 0 3.3689204907705575e-03
GC_3_419 b_3 NI_3 NS_419 0 8.1686018875512766e-03
GC_3_420 b_3 NI_3 NS_420 0 1.0244021308385393e-02
GC_3_421 b_3 NI_3 NS_421 0 -6.9844576983856023e-03
GC_3_422 b_3 NI_3 NS_422 0 2.9355127668043266e-03
GC_3_423 b_3 NI_3 NS_423 0 -5.6336298361881467e-03
GC_3_424 b_3 NI_3 NS_424 0 -8.0966182198784174e-03
GC_3_425 b_3 NI_3 NS_425 0 9.8584915540587160e-03
GC_3_426 b_3 NI_3 NS_426 0 5.4631017419306410e-04
GC_3_427 b_3 NI_3 NS_427 0 -1.0941995599537969e-02
GC_3_428 b_3 NI_3 NS_428 0 1.2300363994202089e-02
GC_3_429 b_3 NI_3 NS_429 0 9.6442553828806222e-03
GC_3_430 b_3 NI_3 NS_430 0 5.0348588902566572e-03
GC_3_431 b_3 NI_3 NS_431 0 -1.9883985200320440e-05
GC_3_432 b_3 NI_3 NS_432 0 3.1661966432011716e-05
GC_3_433 b_3 NI_3 NS_433 0 -7.1319613163818027e-03
GC_3_434 b_3 NI_3 NS_434 0 4.4777052052050416e-03
GC_3_435 b_3 NI_3 NS_435 0 -7.6765708540058762e-03
GC_3_436 b_3 NI_3 NS_436 0 -5.3213603664122051e-03
GC_3_437 b_3 NI_3 NS_437 0 9.5165623812701033e-03
GC_3_438 b_3 NI_3 NS_438 0 -1.7362126108751968e-03
GC_3_439 b_3 NI_3 NS_439 0 1.2475059192430610e-02
GC_3_440 b_3 NI_3 NS_440 0 -1.4048329693611642e-03
GC_3_441 b_3 NI_3 NS_441 0 -5.0716635897051854e-03
GC_3_442 b_3 NI_3 NS_442 0 -2.7496733966124337e-03
GC_3_443 b_3 NI_3 NS_443 0 -2.2243978909363073e-03
GC_3_444 b_3 NI_3 NS_444 0 6.6017968403823046e-03
GC_3_445 b_3 NI_3 NS_445 0 8.9571109105278639e-03
GC_3_446 b_3 NI_3 NS_446 0 1.3095527017938465e-04
GC_3_447 b_3 NI_3 NS_447 0 1.2487335323276505e-02
GC_3_448 b_3 NI_3 NS_448 0 1.7801045114246357e-03
GC_3_449 b_3 NI_3 NS_449 0 -5.3781336503785663e-03
GC_3_450 b_3 NI_3 NS_450 0 4.1549302308158936e-03
GC_3_451 b_3 NI_3 NS_451 0 -1.8500372706359753e-03
GC_3_452 b_3 NI_3 NS_452 0 -5.6869514769111260e-03
GC_3_453 b_3 NI_3 NS_453 0 2.0790311028928447e-07
GC_3_454 b_3 NI_3 NS_454 0 -2.4564428159685921e-07
GC_3_455 b_3 NI_3 NS_455 0 -1.1505423429803206e-05
GC_3_456 b_3 NI_3 NS_456 0 1.8244723149695260e-05
GC_3_457 b_3 NI_3 NS_457 0 3.0649014469929744e-04
GC_3_458 b_3 NI_3 NS_458 0 -1.4375818013946109e-05
GC_3_459 b_3 NI_3 NS_459 0 -1.2385100371115240e-09
GC_3_460 b_3 NI_3 NS_460 0 -1.9194463731832676e-08
GC_3_461 b_3 NI_3 NS_461 0 3.1995090956094945e-06
GC_3_462 b_3 NI_3 NS_462 0 -3.9682765051531092e-06
GC_3_463 b_3 NI_3 NS_463 0 -1.2574826182039560e-05
GC_3_464 b_3 NI_3 NS_464 0 -1.0246050136219216e-06
GC_3_465 b_3 NI_3 NS_465 0 3.9886438467524113e-05
GC_3_466 b_3 NI_3 NS_466 0 8.6693182335041387e-07
GC_3_467 b_3 NI_3 NS_467 0 -4.2799424677546528e-05
GC_3_468 b_3 NI_3 NS_468 0 -2.4449725198996702e-05
GC_3_469 b_3 NI_3 NS_469 0 1.1879750984604558e-06
GC_3_470 b_3 NI_3 NS_470 0 4.3287498697819369e-05
GC_3_471 b_3 NI_3 NS_471 0 1.0659389702693420e-05
GC_3_472 b_3 NI_3 NS_472 0 -4.8918960812767755e-05
GC_3_473 b_3 NI_3 NS_473 0 2.9240464284899215e-06
GC_3_474 b_3 NI_3 NS_474 0 6.2438628283825488e-06
GC_3_475 b_3 NI_3 NS_475 0 -4.5617839029301345e-05
GC_3_476 b_3 NI_3 NS_476 0 1.8881729453428681e-06
GC_3_477 b_3 NI_3 NS_477 0 1.0003674656241523e-04
GC_3_478 b_3 NI_3 NS_478 0 1.2285988350050608e-04
GC_3_479 b_3 NI_3 NS_479 0 -7.5037904375757462e-05
GC_3_480 b_3 NI_3 NS_480 0 -1.3519685186528699e-04
GC_3_481 b_3 NI_3 NS_481 0 -6.7762987393431699e-05
GC_3_482 b_3 NI_3 NS_482 0 4.9170696667270291e-05
GC_3_483 b_3 NI_3 NS_483 0 1.3378660924829309e-04
GC_3_484 b_3 NI_3 NS_484 0 -2.6377115157295681e-05
GC_3_485 b_3 NI_3 NS_485 0 -8.7279468040578437e-05
GC_3_486 b_3 NI_3 NS_486 0 -1.1629395884490385e-05
GC_3_487 b_3 NI_3 NS_487 0 -9.6761214371615420e-05
GC_3_488 b_3 NI_3 NS_488 0 2.1083875757578940e-04
GC_3_489 b_3 NI_3 NS_489 0 1.6568017167332939e-04
GC_3_490 b_3 NI_3 NS_490 0 -2.1189014283367016e-04
GC_3_491 b_3 NI_3 NS_491 0 -8.1910387861866926e-05
GC_3_492 b_3 NI_3 NS_492 0 1.9157070171098780e-05
GC_3_493 b_3 NI_3 NS_493 0 1.6054550553048152e-04
GC_3_494 b_3 NI_3 NS_494 0 4.4267034224804477e-05
GC_3_495 b_3 NI_3 NS_495 0 -8.8293784339272841e-05
GC_3_496 b_3 NI_3 NS_496 0 -7.2083231838471063e-05
GC_3_497 b_3 NI_3 NS_497 0 -8.5464792256415725e-05
GC_3_498 b_3 NI_3 NS_498 0 6.3490319919371421e-05
GC_3_499 b_3 NI_3 NS_499 0 1.4126734934239370e-04
GC_3_500 b_3 NI_3 NS_500 0 -4.6884427744525991e-05
GC_3_501 b_3 NI_3 NS_501 0 -6.6094061791706688e-05
GC_3_502 b_3 NI_3 NS_502 0 -2.4355974473400084e-05
GC_3_503 b_3 NI_3 NS_503 0 6.0403144611207921e-05
GC_3_504 b_3 NI_3 NS_504 0 1.1474521609425703e-04
GC_3_505 b_3 NI_3 NS_505 0 -2.2018823439197774e-05
GC_3_506 b_3 NI_3 NS_506 0 -1.2143064039939254e-04
GC_3_507 b_3 NI_3 NS_507 0 -4.4471467126523004e-05
GC_3_508 b_3 NI_3 NS_508 0 1.0923645233293983e-05
GC_3_509 b_3 NI_3 NS_509 0 4.7465213081754004e-05
GC_3_510 b_3 NI_3 NS_510 0 -9.9250319555159098e-06
GC_3_511 b_3 NI_3 NS_511 0 -3.2079696520982190e-05
GC_3_512 b_3 NI_3 NS_512 0 -7.5861025176683511e-06
GC_3_513 b_3 NI_3 NS_513 0 2.1298742125805790e-05
GC_3_514 b_3 NI_3 NS_514 0 -4.6124679563248106e-06
GC_3_515 b_3 NI_3 NS_515 0 -3.2316439369767654e-05
GC_3_516 b_3 NI_3 NS_516 0 -2.5188454948368593e-05
GC_3_517 b_3 NI_3 NS_517 0 1.2511646345921906e-05
GC_3_518 b_3 NI_3 NS_518 0 6.5127524800000128e-06
GC_3_519 b_3 NI_3 NS_519 0 -2.0423934957688914e-05
GC_3_520 b_3 NI_3 NS_520 0 -7.6317420445111308e-06
GC_3_521 b_3 NI_3 NS_521 0 1.3991873368839516e-05
GC_3_522 b_3 NI_3 NS_522 0 -1.2277807416821980e-05
GC_3_523 b_3 NI_3 NS_523 0 -4.1514156812882472e-05
GC_3_524 b_3 NI_3 NS_524 0 -1.6952622022818808e-05
GC_3_525 b_3 NI_3 NS_525 0 1.1564886106937286e-05
GC_3_526 b_3 NI_3 NS_526 0 -1.4317484316671382e-06
GC_3_527 b_3 NI_3 NS_527 0 -3.0400739246435405e-05
GC_3_528 b_3 NI_3 NS_528 0 5.6250432972654645e-06
GC_3_529 b_3 NI_3 NS_529 0 1.6017175717592890e-05
GC_3_530 b_3 NI_3 NS_530 0 -2.0571749040691448e-05
GC_3_531 b_3 NI_3 NS_531 0 -5.0238949094566849e-05
GC_3_532 b_3 NI_3 NS_532 0 -1.7712123434383629e-06
GC_3_533 b_3 NI_3 NS_533 0 1.1586538840626309e-05
GC_3_534 b_3 NI_3 NS_534 0 -1.1192321951074001e-05
GC_3_535 b_3 NI_3 NS_535 0 -3.2362723135694858e-05
GC_3_536 b_3 NI_3 NS_536 0 2.5180884348485988e-05
GC_3_537 b_3 NI_3 NS_537 0 1.0238935366203533e-05
GC_3_538 b_3 NI_3 NS_538 0 -3.5897419939861997e-05
GC_3_539 b_3 NI_3 NS_539 0 -3.4867048802824876e-05
GC_3_540 b_3 NI_3 NS_540 0 1.8379095255693627e-05
GC_3_541 b_3 NI_3 NS_541 0 -5.6371123367503143e-05
GC_3_542 b_3 NI_3 NS_542 0 1.3313686501379785e-04
GC_3_543 b_3 NI_3 NS_543 0 -1.5277017031428080e-05
GC_3_544 b_3 NI_3 NS_544 0 -3.1721916803075226e-05
GC_3_545 b_3 NI_3 NS_545 0 -3.7761113317399649e-07
GC_3_546 b_3 NI_3 NS_546 0 3.9607644817420515e-07
GC_3_547 b_3 NI_3 NS_547 0 -2.0156821510969414e-05
GC_3_548 b_3 NI_3 NS_548 0 3.2120813892119232e-05
GC_3_549 b_3 NI_3 NS_549 0 -1.4301601693077072e-05
GC_3_550 b_3 NI_3 NS_550 0 -3.3397592519392633e-05
GC_3_551 b_3 NI_3 NS_551 0 -6.1607147560229697e-06
GC_3_552 b_3 NI_3 NS_552 0 5.1177418527893296e-06
GC_3_553 b_3 NI_3 NS_553 0 -2.1208244191657411e-05
GC_3_554 b_3 NI_3 NS_554 0 -6.5712469316889046e-05
GC_3_555 b_3 NI_3 NS_555 0 -9.1589652472161583e-06
GC_3_556 b_3 NI_3 NS_556 0 -2.0643900415547212e-05
GC_3_557 b_3 NI_3 NS_557 0 1.5019857709165147e-05
GC_3_558 b_3 NI_3 NS_558 0 2.2754441222959755e-05
GC_3_559 b_3 NI_3 NS_559 0 -6.7861489750651491e-06
GC_3_560 b_3 NI_3 NS_560 0 2.7711939325075522e-05
GC_3_561 b_3 NI_3 NS_561 0 -1.1040735791539848e-05
GC_3_562 b_3 NI_3 NS_562 0 -2.1529802259453545e-05
GC_3_563 b_3 NI_3 NS_563 0 -1.1040032893846277e-05
GC_3_564 b_3 NI_3 NS_564 0 2.3841805447653507e-05
GC_3_565 b_3 NI_3 NS_565 0 5.1225288501658066e-06
GC_3_566 b_3 NI_3 NS_566 0 -1.5323283050338317e-05
GC_3_567 b_3 NI_3 NS_567 0 -4.7531527920949216e-10
GC_3_568 b_3 NI_3 NS_568 0 -9.1476844985451802e-10
GC_3_569 b_3 NI_3 NS_569 0 -5.5313689436814466e-08
GC_3_570 b_3 NI_3 NS_570 0 7.4255347324336934e-09
GC_3_571 b_3 NI_3 NS_571 0 -2.0465924711883491e-04
GC_3_572 b_3 NI_3 NS_572 0 -3.3255116830617994e-06
GC_3_573 b_3 NI_3 NS_573 0 1.2945489070889762e-09
GC_3_574 b_3 NI_3 NS_574 0 9.6766135775247091e-09
GC_3_575 b_3 NI_3 NS_575 0 -4.2560823378567742e-06
GC_3_576 b_3 NI_3 NS_576 0 6.2139744073949615e-06
GC_3_577 b_3 NI_3 NS_577 0 3.7169291381139890e-06
GC_3_578 b_3 NI_3 NS_578 0 -8.0226842979537442e-06
GC_3_579 b_3 NI_3 NS_579 0 2.1711139613155058e-05
GC_3_580 b_3 NI_3 NS_580 0 -8.4068393612986719e-06
GC_3_581 b_3 NI_3 NS_581 0 -2.1213735891461894e-05
GC_3_582 b_3 NI_3 NS_582 0 -1.2028684245006803e-06
GC_3_583 b_3 NI_3 NS_583 0 -2.9295838686155297e-05
GC_3_584 b_3 NI_3 NS_584 0 -2.8036655938407405e-05
GC_3_585 b_3 NI_3 NS_585 0 -4.8461134704412288e-06
GC_3_586 b_3 NI_3 NS_586 0 1.6200691785524323e-05
GC_3_587 b_3 NI_3 NS_587 0 -2.6737682723069671e-06
GC_3_588 b_3 NI_3 NS_588 0 -7.1113069843625868e-06
GC_3_589 b_3 NI_3 NS_589 0 -2.2547101883084176e-05
GC_3_590 b_3 NI_3 NS_590 0 5.7325226522067262e-06
GC_3_591 b_3 NI_3 NS_591 0 -1.8497083567226076e-04
GC_3_592 b_3 NI_3 NS_592 0 -4.4589107999867990e-05
GC_3_593 b_3 NI_3 NS_593 0 6.1993812843676808e-05
GC_3_594 b_3 NI_3 NS_594 0 1.3751678866234945e-04
GC_3_595 b_3 NI_3 NS_595 0 -3.7420883115908971e-05
GC_3_596 b_3 NI_3 NS_596 0 5.6316425443601031e-05
GC_3_597 b_3 NI_3 NS_597 0 9.5006449750773385e-05
GC_3_598 b_3 NI_3 NS_598 0 2.4592086909545999e-04
GC_3_599 b_3 NI_3 NS_599 0 7.3727691183909716e-05
GC_3_600 b_3 NI_3 NS_600 0 8.1340869169519900e-07
GC_3_601 b_3 NI_3 NS_601 0 -1.6013488611784134e-05
GC_3_602 b_3 NI_3 NS_602 0 2.6083742161305538e-04
GC_3_603 b_3 NI_3 NS_603 0 3.6487195440239041e-04
GC_3_604 b_3 NI_3 NS_604 0 -2.4275812290787003e-04
GC_3_605 b_3 NI_3 NS_605 0 6.5712947292076849e-05
GC_3_606 b_3 NI_3 NS_606 0 -2.8184590609336607e-05
GC_3_607 b_3 NI_3 NS_607 0 2.0799642788529849e-04
GC_3_608 b_3 NI_3 NS_608 0 -2.4122513636738399e-04
GC_3_609 b_3 NI_3 NS_609 0 -7.1069705111480292e-05
GC_3_610 b_3 NI_3 NS_610 0 -7.1882656785808710e-05
GC_3_611 b_3 NI_3 NS_611 0 6.4720731034706474e-05
GC_3_612 b_3 NI_3 NS_612 0 -7.5166912716703423e-05
GC_3_613 b_3 NI_3 NS_613 0 -1.7062494745988651e-04
GC_3_614 b_3 NI_3 NS_614 0 -1.8331083913722483e-04
GC_3_615 b_3 NI_3 NS_615 0 -4.8753415333357332e-05
GC_3_616 b_3 NI_3 NS_616 0 -1.9422271967077200e-05
GC_3_617 b_3 NI_3 NS_617 0 -1.4456137574137560e-04
GC_3_618 b_3 NI_3 NS_618 0 -9.5399247564629955e-05
GC_3_619 b_3 NI_3 NS_619 0 -2.7694032879901671e-05
GC_3_620 b_3 NI_3 NS_620 0 1.0380547924474076e-04
GC_3_621 b_3 NI_3 NS_621 0 -2.7258367655581769e-05
GC_3_622 b_3 NI_3 NS_622 0 1.3718071693849103e-05
GC_3_623 b_3 NI_3 NS_623 0 2.3543137291152653e-06
GC_3_624 b_3 NI_3 NS_624 0 5.0802587989043759e-05
GC_3_625 b_3 NI_3 NS_625 0 1.6821899088470406e-05
GC_3_626 b_3 NI_3 NS_626 0 -4.6940276499444392e-07
GC_3_627 b_3 NI_3 NS_627 0 1.7925283712577277e-06
GC_3_628 b_3 NI_3 NS_628 0 -1.5480347570582047e-05
GC_3_629 b_3 NI_3 NS_629 0 -1.4962445078380682e-05
GC_3_630 b_3 NI_3 NS_630 0 -1.3719795215391290e-05
GC_3_631 b_3 NI_3 NS_631 0 -1.2980299454703587e-05
GC_3_632 b_3 NI_3 NS_632 0 1.2291504010766836e-05
GC_3_633 b_3 NI_3 NS_633 0 7.7935024248751446e-06
GC_3_634 b_3 NI_3 NS_634 0 1.2794176646672751e-06
GC_3_635 b_3 NI_3 NS_635 0 -5.1334665923570329e-06
GC_3_636 b_3 NI_3 NS_636 0 -1.2739690861806197e-05
GC_3_637 b_3 NI_3 NS_637 0 -2.0684368992677153e-05
GC_3_638 b_3 NI_3 NS_638 0 -5.9679191800773483e-06
GC_3_639 b_3 NI_3 NS_639 0 1.1830383722591569e-06
GC_3_640 b_3 NI_3 NS_640 0 2.1729586076454957e-05
GC_3_641 b_3 NI_3 NS_641 0 1.2901795489733608e-05
GC_3_642 b_3 NI_3 NS_642 0 -6.8764804997816952e-06
GC_3_643 b_3 NI_3 NS_643 0 -1.7239594347304546e-05
GC_3_644 b_3 NI_3 NS_644 0 -1.6087364554722395e-05
GC_3_645 b_3 NI_3 NS_645 0 -2.7000607259752654e-05
GC_3_646 b_3 NI_3 NS_646 0 8.7818313629167679e-06
GC_3_647 b_3 NI_3 NS_647 0 2.7184785548216861e-05
GC_3_648 b_3 NI_3 NS_648 0 2.2283570225192131e-05
GC_3_649 b_3 NI_3 NS_649 0 1.1017161633763587e-05
GC_3_650 b_3 NI_3 NS_650 0 -2.1371412190780910e-05
GC_3_651 b_3 NI_3 NS_651 0 -3.0546769742005021e-05
GC_3_652 b_3 NI_3 NS_652 0 3.7146577009725459e-06
GC_3_653 b_3 NI_3 NS_653 0 -9.5336410837867883e-06
GC_3_654 b_3 NI_3 NS_654 0 3.9207837066975832e-05
GC_3_655 b_3 NI_3 NS_655 0 1.8462470006090607e-05
GC_3_656 b_3 NI_3 NS_656 0 -6.8326581635949943e-05
GC_3_657 b_3 NI_3 NS_657 0 4.3338394090484927e-05
GC_3_658 b_3 NI_3 NS_658 0 -1.7306953940697546e-05
GC_3_659 b_3 NI_3 NS_659 0 1.9831835268566361e-07
GC_3_660 b_3 NI_3 NS_660 0 -2.4930649680851481e-07
GC_3_661 b_3 NI_3 NS_661 0 -3.6889333819601574e-06
GC_3_662 b_3 NI_3 NS_662 0 -2.1088368866046044e-05
GC_3_663 b_3 NI_3 NS_663 0 -1.0619647434233235e-05
GC_3_664 b_3 NI_3 NS_664 0 1.6523072874606205e-05
GC_3_665 b_3 NI_3 NS_665 0 9.4073706782430947e-06
GC_3_666 b_3 NI_3 NS_666 0 3.1757011385023296e-05
GC_3_667 b_3 NI_3 NS_667 0 1.4489703787008575e-05
GC_3_668 b_3 NI_3 NS_668 0 -3.2770643984440729e-06
GC_3_669 b_3 NI_3 NS_669 0 -3.8741493362292013e-06
GC_3_670 b_3 NI_3 NS_670 0 1.2514850254492605e-05
GC_3_671 b_3 NI_3 NS_671 0 -1.8542555312356906e-05
GC_3_672 b_3 NI_3 NS_672 0 -3.5697553510284904e-06
GC_3_673 b_3 NI_3 NS_673 0 1.3189260563169996e-05
GC_3_674 b_3 NI_3 NS_674 0 1.3199110180773637e-05
GC_3_675 b_3 NI_3 NS_675 0 7.6293358802796637e-06
GC_3_676 b_3 NI_3 NS_676 0 -2.3004658301504690e-05
GC_3_677 b_3 NI_3 NS_677 0 -3.8543187146119047e-06
GC_3_678 b_3 NI_3 NS_678 0 -1.1714815665584061e-05
GC_3_679 b_3 NI_3 NS_679 0 -8.7383824714374016e-06
GC_3_680 b_3 NI_3 NS_680 0 -2.6220831285732038e-06
GC_3_681 b_3 NI_3 NS_681 0 5.5128498742437658e-10
GC_3_682 b_3 NI_3 NS_682 0 2.9325602419775103e-10
GC_3_683 b_3 NI_3 NS_683 0 4.2108235304711091e-08
GC_3_684 b_3 NI_3 NS_684 0 3.6979686990901636e-08
GC_3_685 b_3 NI_3 NS_685 0 -1.0995071658319755e-04
GC_3_686 b_3 NI_3 NS_686 0 -2.1492391553394247e-06
GC_3_687 b_3 NI_3 NS_687 0 -2.5033371285226215e-10
GC_3_688 b_3 NI_3 NS_688 0 2.6123672988752566e-09
GC_3_689 b_3 NI_3 NS_689 0 1.8909815545965308e-06
GC_3_690 b_3 NI_3 NS_690 0 -1.6338261398097897e-06
GC_3_691 b_3 NI_3 NS_691 0 3.4328438770107056e-07
GC_3_692 b_3 NI_3 NS_692 0 -6.5685023897939638e-06
GC_3_693 b_3 NI_3 NS_693 0 -7.5232094597130009e-06
GC_3_694 b_3 NI_3 NS_694 0 -5.2405427509015949e-07
GC_3_695 b_3 NI_3 NS_695 0 -1.5644387221847511e-06
GC_3_696 b_3 NI_3 NS_696 0 -4.8503531791645673e-06
GC_3_697 b_3 NI_3 NS_697 0 -1.6089131276921545e-05
GC_3_698 b_3 NI_3 NS_698 0 -2.1861625286453285e-06
GC_3_699 b_3 NI_3 NS_699 0 -7.5367534063675820e-06
GC_3_700 b_3 NI_3 NS_700 0 1.8919009302429557e-05
GC_3_701 b_3 NI_3 NS_701 0 5.0282700012095641e-06
GC_3_702 b_3 NI_3 NS_702 0 -2.8006235176684077e-06
GC_3_703 b_3 NI_3 NS_703 0 -2.3106472534723684e-07
GC_3_704 b_3 NI_3 NS_704 0 -2.4616851259300322e-06
GC_3_705 b_3 NI_3 NS_705 0 -2.6994515037914213e-05
GC_3_706 b_3 NI_3 NS_706 0 2.8300303426634692e-05
GC_3_707 b_3 NI_3 NS_707 0 2.8448288981549877e-05
GC_3_708 b_3 NI_3 NS_708 0 -7.8440793707640571e-06
GC_3_709 b_3 NI_3 NS_709 0 -8.2731830366799393e-06
GC_3_710 b_3 NI_3 NS_710 0 -4.3391056033875800e-06
GC_3_711 b_3 NI_3 NS_711 0 1.2150359263408708e-05
GC_3_712 b_3 NI_3 NS_712 0 2.7749141914301770e-05
GC_3_713 b_3 NI_3 NS_713 0 1.4969706447569881e-06
GC_3_714 b_3 NI_3 NS_714 0 -8.9353110944226631e-06
GC_3_715 b_3 NI_3 NS_715 0 -2.9031332100972794e-05
GC_3_716 b_3 NI_3 NS_716 0 4.5480859297515018e-06
GC_3_717 b_3 NI_3 NS_717 0 4.1816724942698727e-05
GC_3_718 b_3 NI_3 NS_718 0 1.1681511468032412e-05
GC_3_719 b_3 NI_3 NS_719 0 -3.0448947307726491e-06
GC_3_720 b_3 NI_3 NS_720 0 -4.4842326053635404e-06
GC_3_721 b_3 NI_3 NS_721 0 1.2838682369610030e-05
GC_3_722 b_3 NI_3 NS_722 0 1.9718563319314308e-05
GC_3_723 b_3 NI_3 NS_723 0 3.9956459581740945e-06
GC_3_724 b_3 NI_3 NS_724 0 -1.0979149548758579e-05
GC_3_725 b_3 NI_3 NS_725 0 -6.6146714106323802e-06
GC_3_726 b_3 NI_3 NS_726 0 8.3775266086306512e-07
GC_3_727 b_3 NI_3 NS_727 0 1.9105219145631208e-05
GC_3_728 b_3 NI_3 NS_728 0 5.9545117395987191e-06
GC_3_729 b_3 NI_3 NS_729 0 -4.3481125736982748e-08
GC_3_730 b_3 NI_3 NS_730 0 -4.2143336895628874e-06
GC_3_731 b_3 NI_3 NS_731 0 4.6805666915879934e-06
GC_3_732 b_3 NI_3 NS_732 0 1.4625900227545052e-05
GC_3_733 b_3 NI_3 NS_733 0 8.1127082587652768e-06
GC_3_734 b_3 NI_3 NS_734 0 -1.1159021727283026e-05
GC_3_735 b_3 NI_3 NS_735 0 -1.4428375333318430e-06
GC_3_736 b_3 NI_3 NS_736 0 9.3170776315321842e-07
GC_3_737 b_3 NI_3 NS_737 0 1.0891210600660229e-05
GC_3_738 b_3 NI_3 NS_738 0 4.3456003269171648e-06
GC_3_739 b_3 NI_3 NS_739 0 1.7188897527880696e-06
GC_3_740 b_3 NI_3 NS_740 0 -6.0609921075008600e-07
GC_3_741 b_3 NI_3 NS_741 0 5.6777116782324429e-06
GC_3_742 b_3 NI_3 NS_742 0 1.7899370625629643e-06
GC_3_743 b_3 NI_3 NS_743 0 3.3742923173757845e-06
GC_3_744 b_3 NI_3 NS_744 0 2.0720323034137567e-06
GC_3_745 b_3 NI_3 NS_745 0 1.0916608323005554e-05
GC_3_746 b_3 NI_3 NS_746 0 3.9123303080877349e-06
GC_3_747 b_3 NI_3 NS_747 0 4.8432409496433256e-06
GC_3_748 b_3 NI_3 NS_748 0 -4.2628894688401573e-08
GC_3_749 b_3 NI_3 NS_749 0 9.9680749825861481e-06
GC_3_750 b_3 NI_3 NS_750 0 -9.9862875253092699e-07
GC_3_751 b_3 NI_3 NS_751 0 8.1884655851505216e-06
GC_3_752 b_3 NI_3 NS_752 0 2.9679944661648354e-06
GC_3_753 b_3 NI_3 NS_753 0 1.8986720063351001e-05
GC_3_754 b_3 NI_3 NS_754 0 -5.4365283869611755e-06
GC_3_755 b_3 NI_3 NS_755 0 7.1694241924664644e-06
GC_3_756 b_3 NI_3 NS_756 0 -3.9853757566060747e-06
GC_3_757 b_3 NI_3 NS_757 0 1.3685887051375825e-05
GC_3_758 b_3 NI_3 NS_758 0 -1.1804061813241060e-05
GC_3_759 b_3 NI_3 NS_759 0 1.2305622388236030e-05
GC_3_760 b_3 NI_3 NS_760 0 -3.9592531259690731e-06
GC_3_761 b_3 NI_3 NS_761 0 9.0879427022406556e-06
GC_3_762 b_3 NI_3 NS_762 0 -2.6621762459780410e-05
GC_3_763 b_3 NI_3 NS_763 0 2.2848314601902371e-06
GC_3_764 b_3 NI_3 NS_764 0 -1.2337140459447173e-05
GC_3_765 b_3 NI_3 NS_765 0 -8.3397817167145319e-06
GC_3_766 b_3 NI_3 NS_766 0 -1.8510652616959135e-05
GC_3_767 b_3 NI_3 NS_767 0 -5.0670740911096453e-06
GC_3_768 b_3 NI_3 NS_768 0 -1.2091739050035339e-05
GC_3_769 b_3 NI_3 NS_769 0 5.5654557616292001e-05
GC_3_770 b_3 NI_3 NS_770 0 -8.7608662941574797e-05
GC_3_771 b_3 NI_3 NS_771 0 -1.0050338247931526e-05
GC_3_772 b_3 NI_3 NS_772 0 1.5956335333789003e-06
GC_3_773 b_3 NI_3 NS_773 0 3.9373702446578515e-07
GC_3_774 b_3 NI_3 NS_774 0 -1.2103088307101328e-07
GC_3_775 b_3 NI_3 NS_775 0 -2.7541894813640104e-06
GC_3_776 b_3 NI_3 NS_776 0 -1.8116236091766328e-06
GC_3_777 b_3 NI_3 NS_777 0 -4.3434368544254476e-06
GC_3_778 b_3 NI_3 NS_778 0 6.8569496277354945e-07
GC_3_779 b_3 NI_3 NS_779 0 -1.7627011910660767e-05
GC_3_780 b_3 NI_3 NS_780 0 9.5650470227720803e-06
GC_3_781 b_3 NI_3 NS_781 0 -9.4006794355537305e-06
GC_3_782 b_3 NI_3 NS_782 0 3.7414743909207805e-05
GC_3_783 b_3 NI_3 NS_783 0 -7.2091677047789418e-06
GC_3_784 b_3 NI_3 NS_784 0 3.1130503356622155e-07
GC_3_785 b_3 NI_3 NS_785 0 -1.3385611476398891e-05
GC_3_786 b_3 NI_3 NS_786 0 1.8110377163175244e-06
GC_3_787 b_3 NI_3 NS_787 0 -4.6173104119446268e-06
GC_3_788 b_3 NI_3 NS_788 0 -3.3928411351718128e-06
GC_3_789 b_3 NI_3 NS_789 0 -6.3738661871990090e-06
GC_3_790 b_3 NI_3 NS_790 0 1.0329455367702135e-06
GC_3_791 b_3 NI_3 NS_791 0 -3.0262566137034831e-06
GC_3_792 b_3 NI_3 NS_792 0 8.9218041036595846e-07
GC_3_793 b_3 NI_3 NS_793 0 -1.7748343322979847e-06
GC_3_794 b_3 NI_3 NS_794 0 -9.4793263917008579e-07
GC_3_795 b_3 NI_3 NS_795 0 -2.6182138817604382e-10
GC_3_796 b_3 NI_3 NS_796 0 4.2365478344801116e-10
GC_3_797 b_3 NI_3 NS_797 0 2.2745899873363352e-09
GC_3_798 b_3 NI_3 NS_798 0 -2.6878269256795161e-08
GC_3_799 b_3 NI_3 NS_799 0 -3.2372655403145934e-05
GC_3_800 b_3 NI_3 NS_800 0 2.2170618685418072e-06
GC_3_801 b_3 NI_3 NS_801 0 6.8027667763796748e-11
GC_3_802 b_3 NI_3 NS_802 0 3.0563865772536732e-09
GC_3_803 b_3 NI_3 NS_803 0 -1.7154486229367010e-06
GC_3_804 b_3 NI_3 NS_804 0 -1.8282392082159797e-06
GC_3_805 b_3 NI_3 NS_805 0 -5.3489861316351448e-06
GC_3_806 b_3 NI_3 NS_806 0 2.8545579865546766e-06
GC_3_807 b_3 NI_3 NS_807 0 -1.6536858483337460e-05
GC_3_808 b_3 NI_3 NS_808 0 1.8376536162785947e-05
GC_3_809 b_3 NI_3 NS_809 0 1.5065514918522059e-05
GC_3_810 b_3 NI_3 NS_810 0 9.7699993143859924e-06
GC_3_811 b_3 NI_3 NS_811 0 1.7310070878716194e-05
GC_3_812 b_3 NI_3 NS_812 0 2.2719510770004336e-05
GC_3_813 b_3 NI_3 NS_813 0 2.9106417144399645e-05
GC_3_814 b_3 NI_3 NS_814 0 4.9740901250459558e-06
GC_3_815 b_3 NI_3 NS_815 0 -2.9664972750972257e-06
GC_3_816 b_3 NI_3 NS_816 0 -1.8803100698606446e-06
GC_3_817 b_3 NI_3 NS_817 0 1.6935351026235019e-05
GC_3_818 b_3 NI_3 NS_818 0 -2.2272197858420127e-06
GC_3_819 b_3 NI_3 NS_819 0 1.2887338340415521e-04
GC_3_820 b_3 NI_3 NS_820 0 3.4716980738199139e-05
GC_3_821 b_3 NI_3 NS_821 0 -2.8880068552649602e-05
GC_3_822 b_3 NI_3 NS_822 0 -9.8668878154862383e-05
GC_3_823 b_3 NI_3 NS_823 0 2.4897332358078696e-05
GC_3_824 b_3 NI_3 NS_824 0 -3.1464745687811739e-05
GC_3_825 b_3 NI_3 NS_825 0 -4.1613532180863162e-05
GC_3_826 b_3 NI_3 NS_826 0 -1.6650660315292002e-04
GC_3_827 b_3 NI_3 NS_827 0 -4.1829247141262047e-05
GC_3_828 b_3 NI_3 NS_828 0 -4.8975538791137747e-06
GC_3_829 b_3 NI_3 NS_829 0 2.1413279428411633e-05
GC_3_830 b_3 NI_3 NS_830 0 -1.5190691064318927e-04
GC_3_831 b_3 NI_3 NS_831 0 -2.3047172936127621e-04
GC_3_832 b_3 NI_3 NS_832 0 1.1445428517724246e-04
GC_3_833 b_3 NI_3 NS_833 0 -3.7402323983897543e-05
GC_3_834 b_3 NI_3 NS_834 0 1.4353147932653330e-05
GC_3_835 b_3 NI_3 NS_835 0 -1.3776506428070929e-04
GC_3_836 b_3 NI_3 NS_836 0 1.3054866548982562e-04
GC_3_837 b_3 NI_3 NS_837 0 3.6495595296496094e-05
GC_3_838 b_3 NI_3 NS_838 0 4.1231366661423160e-05
GC_3_839 b_3 NI_3 NS_839 0 -3.8131820905035908e-05
GC_3_840 b_3 NI_3 NS_840 0 4.3361763755321303e-05
GC_3_841 b_3 NI_3 NS_841 0 8.7557356471313705e-05
GC_3_842 b_3 NI_3 NS_842 0 1.1842875785047131e-04
GC_3_843 b_3 NI_3 NS_843 0 2.7361987208821612e-05
GC_3_844 b_3 NI_3 NS_844 0 1.0121129557525837e-05
GC_3_845 b_3 NI_3 NS_845 0 8.7345259116927416e-05
GC_3_846 b_3 NI_3 NS_846 0 6.5655783842958430e-05
GC_3_847 b_3 NI_3 NS_847 0 2.0320867692998427e-05
GC_3_848 b_3 NI_3 NS_848 0 -5.7039455048417195e-05
GC_3_849 b_3 NI_3 NS_849 0 1.6979052262970581e-05
GC_3_850 b_3 NI_3 NS_850 0 -8.9186494634914333e-06
GC_3_851 b_3 NI_3 NS_851 0 8.5888397724407999e-06
GC_3_852 b_3 NI_3 NS_852 0 -3.2921175971523586e-05
GC_3_853 b_3 NI_3 NS_853 0 -8.8489279238482119e-06
GC_3_854 b_3 NI_3 NS_854 0 5.5973408174814575e-07
GC_3_855 b_3 NI_3 NS_855 0 -2.4313525796701676e-06
GC_3_856 b_3 NI_3 NS_856 0 8.5078738942685965e-06
GC_3_857 b_3 NI_3 NS_857 0 1.0241025438727897e-05
GC_3_858 b_3 NI_3 NS_858 0 6.0555287800386642e-06
GC_3_859 b_3 NI_3 NS_859 0 1.2188367760176635e-05
GC_3_860 b_3 NI_3 NS_860 0 -7.8214178877504860e-06
GC_3_861 b_3 NI_3 NS_861 0 -3.4896526587819412e-06
GC_3_862 b_3 NI_3 NS_862 0 -4.3242939995868031e-07
GC_3_863 b_3 NI_3 NS_863 0 2.4744423179454227e-06
GC_3_864 b_3 NI_3 NS_864 0 7.4084005970259214e-06
GC_3_865 b_3 NI_3 NS_865 0 1.3659439484128667e-05
GC_3_866 b_3 NI_3 NS_866 0 2.6169974730069272e-06
GC_3_867 b_3 NI_3 NS_867 0 4.5330335034080087e-06
GC_3_868 b_3 NI_3 NS_868 0 -1.4186448992106106e-05
GC_3_869 b_3 NI_3 NS_869 0 -5.9288408075792013e-06
GC_3_870 b_3 NI_3 NS_870 0 4.2661993909303840e-06
GC_3_871 b_3 NI_3 NS_871 0 1.0298080426193288e-05
GC_3_872 b_3 NI_3 NS_872 0 9.9363539433707410e-06
GC_3_873 b_3 NI_3 NS_873 0 1.7307569443219373e-05
GC_3_874 b_3 NI_3 NS_874 0 -4.2766756757517985e-06
GC_3_875 b_3 NI_3 NS_875 0 -9.2960026011259953e-06
GC_3_876 b_3 NI_3 NS_876 0 -1.5305295657661056e-05
GC_3_877 b_3 NI_3 NS_877 0 -4.0930044328704479e-06
GC_3_878 b_3 NI_3 NS_878 0 1.3520441879926605e-05
GC_3_879 b_3 NI_3 NS_879 0 2.0923707008858084e-05
GC_3_880 b_3 NI_3 NS_880 0 -5.4861471625659523e-07
GC_3_881 b_3 NI_3 NS_881 0 8.8628354075700043e-06
GC_3_882 b_3 NI_3 NS_882 0 -1.7438302579169407e-05
GC_3_883 b_3 NI_3 NS_883 0 2.5769314431633821e-06
GC_3_884 b_3 NI_3 NS_884 0 -1.3773136071740682e-05
GC_3_885 b_3 NI_3 NS_885 0 -1.3801285799065907e-05
GC_3_886 b_3 NI_3 NS_886 0 4.4172114799754868e-06
GC_3_887 b_3 NI_3 NS_887 0 1.6026718765365698e-08
GC_3_888 b_3 NI_3 NS_888 0 -4.1748051403027869e-08
GC_3_889 b_3 NI_3 NS_889 0 8.6200526743100843e-06
GC_3_890 b_3 NI_3 NS_890 0 1.1611777456489526e-05
GC_3_891 b_3 NI_3 NS_891 0 1.0921474389740512e-05
GC_3_892 b_3 NI_3 NS_892 0 -1.1277713964077684e-05
GC_3_893 b_3 NI_3 NS_893 0 -3.7556061023648539e-06
GC_3_894 b_3 NI_3 NS_894 0 -1.0184122378552973e-05
GC_3_895 b_3 NI_3 NS_895 0 -2.3203085548080181e-06
GC_3_896 b_3 NI_3 NS_896 0 1.2932004457856330e-05
GC_3_897 b_3 NI_3 NS_897 0 9.7592890217573124e-07
GC_3_898 b_3 NI_3 NS_898 0 -7.2834869278424407e-06
GC_3_899 b_3 NI_3 NS_899 0 7.5033949889472675e-06
GC_3_900 b_3 NI_3 NS_900 0 1.6764895569629028e-06
GC_3_901 b_3 NI_3 NS_901 0 -6.0990787888875172e-06
GC_3_902 b_3 NI_3 NS_902 0 -8.8899505038446546e-06
GC_3_903 b_3 NI_3 NS_903 0 -4.1231984090056245e-06
GC_3_904 b_3 NI_3 NS_904 0 9.6572580478477900e-06
GC_3_905 b_3 NI_3 NS_905 0 3.3299265004533529e-06
GC_3_906 b_3 NI_3 NS_906 0 6.0429567321399008e-06
GC_3_907 b_3 NI_3 NS_907 0 5.6621067730978258e-06
GC_3_908 b_3 NI_3 NS_908 0 5.1491141523601244e-07
GC_3_909 b_3 NI_3 NS_909 0 6.1217210890633393e-11
GC_3_910 b_3 NI_3 NS_910 0 1.4945703099566448e-10
GC_3_911 b_3 NI_3 NS_911 0 5.9799816901013211e-09
GC_3_912 b_3 NI_3 NS_912 0 -8.3554729968812590e-09
GC_3_913 b_3 NI_3 NS_913 0 4.4177060865611725e-05
GC_3_914 b_3 NI_3 NS_914 0 -2.5097186638868947e-07
GC_3_915 b_3 NI_3 NS_915 0 -1.3616152683812551e-11
GC_3_916 b_3 NI_3 NS_916 0 3.6730829590821991e-10
GC_3_917 b_3 NI_3 NS_917 0 9.4985818741056539e-07
GC_3_918 b_3 NI_3 NS_918 0 -2.0373723275503674e-07
GC_3_919 b_3 NI_3 NS_919 0 1.1052050607945503e-06
GC_3_920 b_3 NI_3 NS_920 0 -6.5605003538830031e-07
GC_3_921 b_3 NI_3 NS_921 0 1.6285499628442734e-06
GC_3_922 b_3 NI_3 NS_922 0 -3.6724997221192830e-06
GC_3_923 b_3 NI_3 NS_923 0 -2.3667652651887931e-06
GC_3_924 b_3 NI_3 NS_924 0 -1.3304689318962937e-06
GC_3_925 b_3 NI_3 NS_925 0 -2.0333779839636171e-07
GC_3_926 b_3 NI_3 NS_926 0 -2.4445406920546318e-06
GC_3_927 b_3 NI_3 NS_927 0 -7.1157299120281041e-06
GC_3_928 b_3 NI_3 NS_928 0 -2.8107547510678335e-06
GC_3_929 b_3 NI_3 NS_929 0 1.7244824603418727e-06
GC_3_930 b_3 NI_3 NS_930 0 1.3116575558375586e-06
GC_3_931 b_3 NI_3 NS_931 0 -1.6513152052959692e-06
GC_3_932 b_3 NI_3 NS_932 0 9.9666912661412106e-07
GC_3_933 b_3 NI_3 NS_933 0 -2.8707134907200220e-06
GC_3_934 b_3 NI_3 NS_934 0 -1.6218900706569080e-06
GC_3_935 b_3 NI_3 NS_935 0 -2.0401142360180258e-06
GC_3_936 b_3 NI_3 NS_936 0 2.9683224547563123e-06
GC_3_937 b_3 NI_3 NS_937 0 -1.1731161052972225e-06
GC_3_938 b_3 NI_3 NS_938 0 1.1051280936939885e-06
GC_3_939 b_3 NI_3 NS_939 0 -2.0978467059781227e-06
GC_3_940 b_3 NI_3 NS_940 0 1.5286386186653615e-06
GC_3_941 b_3 NI_3 NS_941 0 -9.4302697387863662e-07
GC_3_942 b_3 NI_3 NS_942 0 1.4307778991596463e-06
GC_3_943 b_3 NI_3 NS_943 0 -1.4824681294939226e-06
GC_3_944 b_3 NI_3 NS_944 0 1.7943987626761130e-06
GC_3_945 b_3 NI_3 NS_945 0 2.5484730974979390e-07
GC_3_946 b_3 NI_3 NS_946 0 1.3612752466576283e-06
GC_3_947 b_3 NI_3 NS_947 0 -8.4240911635689353e-07
GC_3_948 b_3 NI_3 NS_948 0 1.3600820798292787e-06
GC_3_949 b_3 NI_3 NS_949 0 9.0836753353544682e-07
GC_3_950 b_3 NI_3 NS_950 0 1.8504787199215935e-06
GC_3_951 b_3 NI_3 NS_951 0 -7.6710521753919026e-07
GC_3_952 b_3 NI_3 NS_952 0 5.7087098527675457e-07
GC_3_953 b_3 NI_3 NS_953 0 -8.0356113212018927e-07
GC_3_954 b_3 NI_3 NS_954 0 1.5919271308684389e-06
GC_3_955 b_3 NI_3 NS_955 0 1.2779890713338251e-06
GC_3_956 b_3 NI_3 NS_956 0 5.6822829760383927e-07
GC_3_957 b_3 NI_3 NS_957 0 -6.6680311365602551e-07
GC_3_958 b_3 NI_3 NS_958 0 6.5598676699021202e-07
GC_3_959 b_3 NI_3 NS_959 0 5.3996086811349707e-07
GC_3_960 b_3 NI_3 NS_960 0 1.7896995378621174e-06
GC_3_961 b_3 NI_3 NS_961 0 -2.5639123668799729e-07
GC_3_962 b_3 NI_3 NS_962 0 -3.2550611217580332e-07
GC_3_963 b_3 NI_3 NS_963 0 -4.7492380634407808e-07
GC_3_964 b_3 NI_3 NS_964 0 6.1074267645079289e-07
GC_3_965 b_3 NI_3 NS_965 0 1.1438518183421884e-07
GC_3_966 b_3 NI_3 NS_966 0 5.8913309567934370e-07
GC_3_967 b_3 NI_3 NS_967 0 -3.1820155663074346e-07
GC_3_968 b_3 NI_3 NS_968 0 4.4618015125325984e-07
GC_3_969 b_3 NI_3 NS_969 0 6.3950178039105934e-08
GC_3_970 b_3 NI_3 NS_970 0 2.2647527320377170e-07
GC_3_971 b_3 NI_3 NS_971 0 -6.7253827992132606e-07
GC_3_972 b_3 NI_3 NS_972 0 2.4744285264853228e-07
GC_3_973 b_3 NI_3 NS_973 0 -1.6416035217875502e-07
GC_3_974 b_3 NI_3 NS_974 0 5.7606106274174895e-07
GC_3_975 b_3 NI_3 NS_975 0 -3.0458069507785400e-07
GC_3_976 b_3 NI_3 NS_976 0 2.5969235005585639e-07
GC_3_977 b_3 NI_3 NS_977 0 -9.8767048196711519e-08
GC_3_978 b_3 NI_3 NS_978 0 2.0869421631215413e-07
GC_3_979 b_3 NI_3 NS_979 0 -7.6623277193570601e-07
GC_3_980 b_3 NI_3 NS_980 0 5.3639653787766106e-08
GC_3_981 b_3 NI_3 NS_981 0 -4.8039118803191450e-07
GC_3_982 b_3 NI_3 NS_982 0 4.3217421540659633e-07
GC_3_983 b_3 NI_3 NS_983 0 -5.3152819138060208e-07
GC_3_984 b_3 NI_3 NS_984 0 2.1427235146615236e-07
GC_3_985 b_3 NI_3 NS_985 0 -5.2278848993715626e-07
GC_3_986 b_3 NI_3 NS_986 0 1.4454166133218744e-07
GC_3_987 b_3 NI_3 NS_987 0 -1.0033849855108283e-06
GC_3_988 b_3 NI_3 NS_988 0 -3.4734940094131252e-07
GC_3_989 b_3 NI_3 NS_989 0 -1.4397698721732006e-06
GC_3_990 b_3 NI_3 NS_990 0 5.4836666380478718e-07
GC_3_991 b_3 NI_3 NS_991 0 -1.1943884880207086e-06
GC_3_992 b_3 NI_3 NS_992 0 1.3609839795645726e-07
GC_3_993 b_3 NI_3 NS_993 0 -1.4806568520943862e-06
GC_3_994 b_3 NI_3 NS_994 0 7.7902411555177812e-07
GC_3_995 b_3 NI_3 NS_995 0 -2.2609435353423528e-06
GC_3_996 b_3 NI_3 NS_996 0 -8.4608337541737472e-07
GC_3_997 b_3 NI_3 NS_997 0 5.6638039775549932e-06
GC_3_998 b_3 NI_3 NS_998 0 1.1197138908282034e-05
GC_3_999 b_3 NI_3 NS_999 0 -2.2219658670416656e-06
GC_3_1000 b_3 NI_3 NS_1000 0 3.0963833595659916e-06
GC_3_1001 b_3 NI_3 NS_1001 0 1.1649812711249133e-08
GC_3_1002 b_3 NI_3 NS_1002 0 7.3477932810202773e-08
GC_3_1003 b_3 NI_3 NS_1003 0 -1.2473679226794471e-06
GC_3_1004 b_3 NI_3 NS_1004 0 1.6458031996802141e-06
GC_3_1005 b_3 NI_3 NS_1005 0 -6.3373480320561619e-07
GC_3_1006 b_3 NI_3 NS_1006 0 1.4520521693953957e-06
GC_3_1007 b_3 NI_3 NS_1007 0 -1.6479512760434973e-06
GC_3_1008 b_3 NI_3 NS_1008 0 -1.2214123858808082e-06
GC_3_1009 b_3 NI_3 NS_1009 0 -3.3894900201242256e-06
GC_3_1010 b_3 NI_3 NS_1010 0 -1.1083936800717308e-06
GC_3_1011 b_3 NI_3 NS_1011 0 7.1945204939936739e-09
GC_3_1012 b_3 NI_3 NS_1012 0 -1.2021669254395325e-07
GC_3_1013 b_3 NI_3 NS_1013 0 6.2008602208056386e-07
GC_3_1014 b_3 NI_3 NS_1014 0 -3.6780548142135339e-07
GC_3_1015 b_3 NI_3 NS_1015 0 -4.6880507985864784e-08
GC_3_1016 b_3 NI_3 NS_1016 0 3.9700351944666724e-07
GC_3_1017 b_3 NI_3 NS_1017 0 -5.1636680025940568e-08
GC_3_1018 b_3 NI_3 NS_1018 0 2.9619692294955124e-08
GC_3_1019 b_3 NI_3 NS_1019 0 -2.7362373296513165e-07
GC_3_1020 b_3 NI_3 NS_1020 0 1.7742433675872382e-07
GC_3_1021 b_3 NI_3 NS_1021 0 -2.2775884838723959e-07
GC_3_1022 b_3 NI_3 NS_1022 0 -6.5495297870191421e-09
GC_3_1023 b_3 NI_3 NS_1023 0 -8.0167911197669566e-12
GC_3_1024 b_3 NI_3 NS_1024 0 -8.1401124711970268e-13
GC_3_1025 b_3 NI_3 NS_1025 0 -1.1403329678457205e-09
GC_3_1026 b_3 NI_3 NS_1026 0 -2.4259802141212357e-09
GC_3_1027 b_3 NI_3 NS_1027 0 -2.1854833916839877e-05
GC_3_1028 b_3 NI_3 NS_1028 0 2.4289006161172072e-07
GC_3_1029 b_3 NI_3 NS_1029 0 1.6216376315217918e-11
GC_3_1030 b_3 NI_3 NS_1030 0 -4.8482427783474362e-10
GC_3_1031 b_3 NI_3 NS_1031 0 3.7396450755763121e-07
GC_3_1032 b_3 NI_3 NS_1032 0 -1.3861159034772247e-06
GC_3_1033 b_3 NI_3 NS_1033 0 -1.4309718016943832e-07
GC_3_1034 b_3 NI_3 NS_1034 0 1.1186853835911725e-06
GC_3_1035 b_3 NI_3 NS_1035 0 -3.5071031713927747e-06
GC_3_1036 b_3 NI_3 NS_1036 0 -2.2368614843726807e-06
GC_3_1037 b_3 NI_3 NS_1037 0 -7.4899853345431133e-07
GC_3_1038 b_3 NI_3 NS_1038 0 -1.1228926603116274e-06
GC_3_1039 b_3 NI_3 NS_1039 0 -6.8318113371680019e-07
GC_3_1040 b_3 NI_3 NS_1040 0 2.6597400275025363e-06
GC_3_1041 b_3 NI_3 NS_1041 0 -5.0808607070636255e-06
GC_3_1042 b_3 NI_3 NS_1042 0 3.8731854316074817e-06
GC_3_1043 b_3 NI_3 NS_1043 0 9.5027454279433163e-07
GC_3_1044 b_3 NI_3 NS_1044 0 -1.5539572419579908e-07
GC_3_1045 b_3 NI_3 NS_1045 0 -2.6330818123314943e-07
GC_3_1046 b_3 NI_3 NS_1046 0 -5.2973881055152311e-07
GC_3_1047 b_3 NI_3 NS_1047 0 -1.4734433088954404e-06
GC_3_1048 b_3 NI_3 NS_1048 0 1.1165094942074517e-05
GC_3_1049 b_3 NI_3 NS_1049 0 5.7514554652619234e-06
GC_3_1050 b_3 NI_3 NS_1050 0 2.9696775351562493e-06
GC_3_1051 b_3 NI_3 NS_1051 0 7.6119473594551712e-07
GC_3_1052 b_3 NI_3 NS_1052 0 -4.0129821364163212e-07
GC_3_1053 b_3 NI_3 NS_1053 0 1.7102516135620666e-05
GC_3_1054 b_3 NI_3 NS_1054 0 -2.9720072801065402e-07
GC_3_1055 b_3 NI_3 NS_1055 0 6.9918325192707569e-07
GC_3_1056 b_3 NI_3 NS_1056 0 1.7755160349321875e-07
GC_3_1057 b_3 NI_3 NS_1057 0 6.4112195712857293e-06
GC_3_1058 b_3 NI_3 NS_1058 0 -4.4581809915092639e-07
GC_3_1059 b_3 NI_3 NS_1059 0 -8.2284108182883289e-07
GC_3_1060 b_3 NI_3 NS_1060 0 -1.7742554150705101e-05
GC_3_1061 b_3 NI_3 NS_1061 0 -2.8403935440038478e-07
GC_3_1062 b_3 NI_3 NS_1062 0 2.3076377879487017e-07
GC_3_1063 b_3 NI_3 NS_1063 0 -1.0767530077562390e-05
GC_3_1064 b_3 NI_3 NS_1064 0 -9.4785309496369869e-06
GC_3_1065 b_3 NI_3 NS_1065 0 -1.3407996095751213e-06
GC_3_1066 b_3 NI_3 NS_1066 0 -8.1236735986811678e-07
GC_3_1067 b_3 NI_3 NS_1067 0 -1.6041529567043698e-06
GC_3_1068 b_3 NI_3 NS_1068 0 4.5798552753772628e-07
GC_3_1069 b_3 NI_3 NS_1069 0 -9.3315609161291004e-06
GC_3_1070 b_3 NI_3 NS_1070 0 6.4364178034936087e-06
GC_3_1071 b_3 NI_3 NS_1071 0 6.8137844921972216e-08
GC_3_1072 b_3 NI_3 NS_1072 0 -4.0002759668406791e-07
GC_3_1073 b_3 NI_3 NS_1073 0 -7.1694041684007398e-07
GC_3_1074 b_3 NI_3 NS_1074 0 7.2315333590394443e-06
GC_3_1075 b_3 NI_3 NS_1075 0 2.0724130263129315e-06
GC_3_1076 b_3 NI_3 NS_1076 0 2.4601621450913063e-06
GC_3_1077 b_3 NI_3 NS_1077 0 6.1987306347716987e-07
GC_3_1078 b_3 NI_3 NS_1078 0 -2.5283446981464403e-07
GC_3_1079 b_3 NI_3 NS_1079 0 4.6121006100660666e-06
GC_3_1080 b_3 NI_3 NS_1080 0 3.3416119348159197e-07
GC_3_1081 b_3 NI_3 NS_1081 0 1.7600652659148247e-07
GC_3_1082 b_3 NI_3 NS_1082 0 5.3884781661101352e-07
GC_3_1083 b_3 NI_3 NS_1083 0 -7.4062907440798735e-07
GC_3_1084 b_3 NI_3 NS_1084 0 -4.2130860863351629e-08
GC_3_1085 b_3 NI_3 NS_1085 0 7.4630668274184051e-07
GC_3_1086 b_3 NI_3 NS_1086 0 -5.2040215538456747e-07
GC_3_1087 b_3 NI_3 NS_1087 0 1.8297447412316341e-06
GC_3_1088 b_3 NI_3 NS_1088 0 4.7558514262942340e-07
GC_3_1089 b_3 NI_3 NS_1089 0 1.7694656183618092e-07
GC_3_1090 b_3 NI_3 NS_1090 0 4.5204738374169875e-07
GC_3_1091 b_3 NI_3 NS_1091 0 -4.4611196905913837e-07
GC_3_1092 b_3 NI_3 NS_1092 0 2.3590712449105618e-07
GC_3_1093 b_3 NI_3 NS_1093 0 6.5001055182241062e-07
GC_3_1094 b_3 NI_3 NS_1094 0 -3.4566770445980366e-07
GC_3_1095 b_3 NI_3 NS_1095 0 1.8731712155427387e-06
GC_3_1096 b_3 NI_3 NS_1096 0 -2.9453557855618551e-08
GC_3_1097 b_3 NI_3 NS_1097 0 2.9820909240609741e-07
GC_3_1098 b_3 NI_3 NS_1098 0 5.0989358305567060e-07
GC_3_1099 b_3 NI_3 NS_1099 0 -3.1510652258649679e-07
GC_3_1100 b_3 NI_3 NS_1100 0 4.5573818822392562e-07
GC_3_1101 b_3 NI_3 NS_1101 0 5.5362439431607750e-07
GC_3_1102 b_3 NI_3 NS_1102 0 -4.4923655012113536e-08
GC_3_1103 b_3 NI_3 NS_1103 0 1.9806774378712053e-06
GC_3_1104 b_3 NI_3 NS_1104 0 -4.0116316196502819e-07
GC_3_1105 b_3 NI_3 NS_1105 0 4.1707219294372835e-07
GC_3_1106 b_3 NI_3 NS_1106 0 7.7173675522300544e-07
GC_3_1107 b_3 NI_3 NS_1107 0 5.0608309900710873e-07
GC_3_1108 b_3 NI_3 NS_1108 0 7.2744621090448871e-07
GC_3_1109 b_3 NI_3 NS_1109 0 9.0286388904487120e-07
GC_3_1110 b_3 NI_3 NS_1110 0 9.8962342683309828e-07
GC_3_1111 b_3 NI_3 NS_1111 0 1.6379049827481174e-06
GC_3_1112 b_3 NI_3 NS_1112 0 -9.9913773058552313e-06
GC_3_1113 b_3 NI_3 NS_1113 0 2.8722296552602965e-06
GC_3_1114 b_3 NI_3 NS_1114 0 -1.2252699164075661e-06
GC_3_1115 b_3 NI_3 NS_1115 0 3.1662845927222963e-08
GC_3_1116 b_3 NI_3 NS_1116 0 -4.6442983968559331e-08
GC_3_1117 b_3 NI_3 NS_1117 0 1.4053571982135720e-06
GC_3_1118 b_3 NI_3 NS_1118 0 1.6962825771210313e-07
GC_3_1119 b_3 NI_3 NS_1119 0 9.7886501749551862e-07
GC_3_1120 b_3 NI_3 NS_1120 0 -4.9523763139335020e-07
GC_3_1121 b_3 NI_3 NS_1121 0 6.9365036086722203e-07
GC_3_1122 b_3 NI_3 NS_1122 0 1.3037895393861259e-06
GC_3_1123 b_3 NI_3 NS_1123 0 1.3369635426314440e-06
GC_3_1124 b_3 NI_3 NS_1124 0 1.9872947531758050e-06
GC_3_1125 b_3 NI_3 NS_1125 0 -9.2421497664907159e-08
GC_3_1126 b_3 NI_3 NS_1126 0 -2.7687295988050489e-08
GC_3_1127 b_3 NI_3 NS_1127 0 -5.3468419616295960e-07
GC_3_1128 b_3 NI_3 NS_1128 0 1.8254478172399365e-07
GC_3_1129 b_3 NI_3 NS_1129 0 3.1918784378970951e-07
GC_3_1130 b_3 NI_3 NS_1130 0 -3.6116449475131514e-07
GC_3_1131 b_3 NI_3 NS_1131 0 1.1497922852441639e-08
GC_3_1132 b_3 NI_3 NS_1132 0 -6.0654716672725754e-07
GC_3_1133 b_3 NI_3 NS_1133 0 5.2303159743021169e-08
GC_3_1134 b_3 NI_3 NS_1134 0 1.0683521734373943e-07
GC_3_1135 b_3 NI_3 NS_1135 0 2.9593147580000381e-07
GC_3_1136 b_3 NI_3 NS_1136 0 -1.4165766505665311e-09
GC_3_1137 b_3 NI_3 NS_1137 0 -2.9851551078523995e-12
GC_3_1138 b_3 NI_3 NS_1138 0 -1.0058610796764704e-11
GC_3_1139 b_3 NI_3 NS_1139 0 9.3171691239647071e-10
GC_3_1140 b_3 NI_3 NS_1140 0 3.3553230155536144e-09
GC_3_1141 b_3 NI_3 NS_1141 0 1.3355928779924241e-05
GC_3_1142 b_3 NI_3 NS_1142 0 -5.8997575843653977e-08
GC_3_1143 b_3 NI_3 NS_1143 0 -1.4899441856949840e-11
GC_3_1144 b_3 NI_3 NS_1144 0 1.3547829277727867e-10
GC_3_1145 b_3 NI_3 NS_1145 0 3.5636791814970023e-07
GC_3_1146 b_3 NI_3 NS_1146 0 -1.8177455202896949e-07
GC_3_1147 b_3 NI_3 NS_1147 0 2.7825888932095555e-07
GC_3_1148 b_3 NI_3 NS_1148 0 -3.4971824928940547e-07
GC_3_1149 b_3 NI_3 NS_1149 0 4.9250083158441482e-07
GC_3_1150 b_3 NI_3 NS_1150 0 -1.4213854174470790e-06
GC_3_1151 b_3 NI_3 NS_1151 0 -1.1592228389141460e-06
GC_3_1152 b_3 NI_3 NS_1152 0 -4.5897559803955047e-07
GC_3_1153 b_3 NI_3 NS_1153 0 -3.4112976087247571e-07
GC_3_1154 b_3 NI_3 NS_1154 0 -6.2118969777542360e-07
GC_3_1155 b_3 NI_3 NS_1155 0 -2.5796967972792178e-06
GC_3_1156 b_3 NI_3 NS_1156 0 -6.4054838805611215e-07
GC_3_1157 b_3 NI_3 NS_1157 0 7.1614975244652757e-07
GC_3_1158 b_3 NI_3 NS_1158 0 3.5572596464849419e-07
GC_3_1159 b_3 NI_3 NS_1159 0 -7.3376226715232976e-07
GC_3_1160 b_3 NI_3 NS_1160 0 3.7327428235125935e-07
GC_3_1161 b_3 NI_3 NS_1161 0 -9.8858906882211567e-07
GC_3_1162 b_3 NI_3 NS_1162 0 5.8562385369982251e-07
GC_3_1163 b_3 NI_3 NS_1163 0 -4.3258656989175277e-07
GC_3_1164 b_3 NI_3 NS_1164 0 2.6363656191994604e-07
GC_3_1165 b_3 NI_3 NS_1165 0 -8.4568601088799554e-07
GC_3_1166 b_3 NI_3 NS_1166 0 4.5886027767438341e-07
GC_3_1167 b_3 NI_3 NS_1167 0 1.6312891923678258e-07
GC_3_1168 b_3 NI_3 NS_1168 0 1.1048465325664357e-06
GC_3_1169 b_3 NI_3 NS_1169 0 -5.9745441796363744e-07
GC_3_1170 b_3 NI_3 NS_1170 0 1.3142479523639729e-07
GC_3_1171 b_3 NI_3 NS_1171 0 -1.8757719219047504e-06
GC_3_1172 b_3 NI_3 NS_1172 0 1.2999561359164899e-06
GC_3_1173 b_3 NI_3 NS_1173 0 2.0548080279058990e-06
GC_3_1174 b_3 NI_3 NS_1174 0 2.3036184858318379e-07
GC_3_1175 b_3 NI_3 NS_1175 0 -6.8567139074755796e-07
GC_3_1176 b_3 NI_3 NS_1176 0 2.0176516555353288e-07
GC_3_1177 b_3 NI_3 NS_1177 0 1.0020787945142575e-06
GC_3_1178 b_3 NI_3 NS_1178 0 1.6689079961481677e-06
GC_3_1179 b_3 NI_3 NS_1179 0 -2.4458558293495402e-07
GC_3_1180 b_3 NI_3 NS_1180 0 -5.7788288060943317e-07
GC_3_1181 b_3 NI_3 NS_1181 0 -9.1772841285059987e-07
GC_3_1182 b_3 NI_3 NS_1182 0 4.3231178804327360e-07
GC_3_1183 b_3 NI_3 NS_1183 0 1.4296286993438959e-06
GC_3_1184 b_3 NI_3 NS_1184 0 6.7975816412396317e-07
GC_3_1185 b_3 NI_3 NS_1185 0 -3.4205146343261994e-07
GC_3_1186 b_3 NI_3 NS_1186 0 -2.1142722236866814e-07
GC_3_1187 b_3 NI_3 NS_1187 0 -2.7750028411562343e-08
GC_3_1188 b_3 NI_3 NS_1188 0 1.4222467437740106e-06
GC_3_1189 b_3 NI_3 NS_1189 0 4.6031318011848701e-07
GC_3_1190 b_3 NI_3 NS_1190 0 -7.6889132001462161e-07
GC_3_1191 b_3 NI_3 NS_1191 0 -3.5271748362096316e-07
GC_3_1192 b_3 NI_3 NS_1192 0 4.9305938884831837e-08
GC_3_1193 b_3 NI_3 NS_1193 0 3.2510584976581727e-07
GC_3_1194 b_3 NI_3 NS_1194 0 3.7853226377604676e-07
GC_3_1195 b_3 NI_3 NS_1195 0 -1.4616429277788368e-07
GC_3_1196 b_3 NI_3 NS_1196 0 -8.4907404384046290e-09
GC_3_1197 b_3 NI_3 NS_1197 0 1.4143255035027092e-07
GC_3_1198 b_3 NI_3 NS_1198 0 1.2099134828375291e-07
GC_3_1199 b_3 NI_3 NS_1199 0 -1.9313702359837866e-07
GC_3_1200 b_3 NI_3 NS_1200 0 -6.8313867170881862e-08
GC_3_1201 b_3 NI_3 NS_1201 0 4.1149209533247286e-08
GC_3_1202 b_3 NI_3 NS_1202 0 1.9490945962711809e-07
GC_3_1203 b_3 NI_3 NS_1203 0 -1.1272486331833694e-07
GC_3_1204 b_3 NI_3 NS_1204 0 1.0158074531120513e-08
GC_3_1205 b_3 NI_3 NS_1205 0 4.5539164385144883e-08
GC_3_1206 b_3 NI_3 NS_1206 0 4.4122148194239485e-09
GC_3_1207 b_3 NI_3 NS_1207 0 -2.9983399061206948e-07
GC_3_1208 b_3 NI_3 NS_1208 0 -5.1244868827055448e-08
GC_3_1209 b_3 NI_3 NS_1209 0 -9.0042054298672344e-08
GC_3_1210 b_3 NI_3 NS_1210 0 6.0468737797561971e-08
GC_3_1211 b_3 NI_3 NS_1211 0 -2.3102780706098720e-07
GC_3_1212 b_3 NI_3 NS_1212 0 8.0940910035913113e-08
GC_3_1213 b_3 NI_3 NS_1213 0 -1.3243196578118853e-07
GC_3_1214 b_3 NI_3 NS_1214 0 -7.1040466929569825e-08
GC_3_1215 b_3 NI_3 NS_1215 0 -4.3092867016865744e-07
GC_3_1216 b_3 NI_3 NS_1216 0 -5.3209705755778633e-08
GC_3_1217 b_3 NI_3 NS_1217 0 -4.1895467943399529e-07
GC_3_1218 b_3 NI_3 NS_1218 0 6.1480670897006409e-08
GC_3_1219 b_3 NI_3 NS_1219 0 -4.4023004427610444e-07
GC_3_1220 b_3 NI_3 NS_1220 0 1.4721721019710926e-07
GC_3_1221 b_3 NI_3 NS_1221 0 -5.1067934735299270e-07
GC_3_1222 b_3 NI_3 NS_1222 0 9.9880054546952523e-08
GC_3_1223 b_3 NI_3 NS_1223 0 -9.6150363769223957e-07
GC_3_1224 b_3 NI_3 NS_1224 0 -9.5716339347894795e-08
GC_3_1225 b_3 NI_3 NS_1225 0 2.6176288262825442e-06
GC_3_1226 b_3 NI_3 NS_1226 0 2.9785672045804833e-06
GC_3_1227 b_3 NI_3 NS_1227 0 -6.1418730955583245e-07
GC_3_1228 b_3 NI_3 NS_1228 0 1.0336821957393965e-06
GC_3_1229 b_3 NI_3 NS_1229 0 9.1644536949046858e-09
GC_3_1230 b_3 NI_3 NS_1230 0 2.5329123382461496e-08
GC_3_1231 b_3 NI_3 NS_1231 0 -4.6836661294466355e-07
GC_3_1232 b_3 NI_3 NS_1232 0 8.2780362337887810e-07
GC_3_1233 b_3 NI_3 NS_1233 0 8.8696459981831150e-09
GC_3_1234 b_3 NI_3 NS_1234 0 3.8273363163960832e-07
GC_3_1235 b_3 NI_3 NS_1235 0 -8.6693344593613361e-07
GC_3_1236 b_3 NI_3 NS_1236 0 -7.0542492973445490e-08
GC_3_1237 b_3 NI_3 NS_1237 0 -9.7666778363759561e-07
GC_3_1238 b_3 NI_3 NS_1238 0 -1.7992953708276506e-07
GC_3_1239 b_3 NI_3 NS_1239 0 1.0735188325266170e-07
GC_3_1240 b_3 NI_3 NS_1240 0 -1.4754516656861407e-07
GC_3_1241 b_3 NI_3 NS_1241 0 6.6793592072872095e-08
GC_3_1242 b_3 NI_3 NS_1242 0 1.4683466627919087e-08
GC_3_1243 b_3 NI_3 NS_1243 0 -6.9788036865501535e-08
GC_3_1244 b_3 NI_3 NS_1244 0 1.6094615098681515e-07
GC_3_1245 b_3 NI_3 NS_1245 0 2.7671234455170610e-08
GC_3_1246 b_3 NI_3 NS_1246 0 -4.0810114302600088e-08
GC_3_1247 b_3 NI_3 NS_1247 0 -8.1264117299518983e-08
GC_3_1248 b_3 NI_3 NS_1248 0 1.6048702555422177e-07
GC_3_1249 b_3 NI_3 NS_1249 0 5.6542114187423213e-08
GC_3_1250 b_3 NI_3 NS_1250 0 -1.6756790926251196e-08
GC_3_1251 b_3 NI_3 NS_1251 0 -1.1794878453629393e-11
GC_3_1252 b_3 NI_3 NS_1252 0 5.2725089488218524e-12
GC_3_1253 b_3 NI_3 NS_1253 0 -3.4161779494748779e-10
GC_3_1254 b_3 NI_3 NS_1254 0 -9.7247739979151361e-10
GC_3_1255 b_3 NI_3 NS_1255 0 -2.7457099510083907e-05
GC_3_1256 b_3 NI_3 NS_1256 0 -1.0861478791027058e-08
GC_3_1257 b_3 NI_3 NS_1257 0 1.0271907587114943e-11
GC_3_1258 b_3 NI_3 NS_1258 0 -5.9963266062516298e-11
GC_3_1259 b_3 NI_3 NS_1259 0 -6.3441211531843190e-07
GC_3_1260 b_3 NI_3 NS_1260 0 -1.0701452793679695e-06
GC_3_1261 b_3 NI_3 NS_1261 0 -1.4351350423279812e-06
GC_3_1262 b_3 NI_3 NS_1262 0 2.3180834773562908e-06
GC_3_1263 b_3 NI_3 NS_1263 0 -3.8038650900736769e-06
GC_3_1264 b_3 NI_3 NS_1264 0 2.1755692185514793e-06
GC_3_1265 b_3 NI_3 NS_1265 0 1.9264441242360036e-06
GC_3_1266 b_3 NI_3 NS_1266 0 -2.2569410511151593e-07
GC_3_1267 b_3 NI_3 NS_1267 0 1.3997827429552893e-06
GC_3_1268 b_3 NI_3 NS_1268 0 5.7146480618049405e-06
GC_3_1269 b_3 NI_3 NS_1269 0 3.7149719486471843e-06
GC_3_1270 b_3 NI_3 NS_1270 0 3.2450720541167335e-06
GC_3_1271 b_3 NI_3 NS_1271 0 -1.4756029610803270e-06
GC_3_1272 b_3 NI_3 NS_1272 0 -9.4893618966407163e-07
GC_3_1273 b_3 NI_3 NS_1273 0 9.7598934374769382e-07
GC_3_1274 b_3 NI_3 NS_1274 0 -2.1769782531005905e-06
GC_3_1275 b_3 NI_3 NS_1275 0 6.4144581749583732e-06
GC_3_1276 b_3 NI_3 NS_1276 0 8.5314135250929441e-06
GC_3_1277 b_3 NI_3 NS_1277 0 1.3418228821299207e-06
GC_3_1278 b_3 NI_3 NS_1278 0 -9.5630748516469349e-07
GC_3_1279 b_3 NI_3 NS_1279 0 1.0785520168783401e-06
GC_3_1280 b_3 NI_3 NS_1280 0 -1.8906356486533086e-06
GC_3_1281 b_3 NI_3 NS_1281 0 1.4514945754946443e-05
GC_3_1282 b_3 NI_3 NS_1282 0 -4.1896499976164626e-06
GC_3_1283 b_3 NI_3 NS_1283 0 -2.0072732425756435e-07
GC_3_1284 b_3 NI_3 NS_1284 0 6.6359849088599658e-07
GC_3_1285 b_3 NI_3 NS_1285 0 4.9434709644091452e-06
GC_3_1286 b_3 NI_3 NS_1286 0 -2.1797969805400931e-06
GC_3_1287 b_3 NI_3 NS_1287 0 -7.7232717742966298e-07
GC_3_1288 b_3 NI_3 NS_1288 0 -1.5002602308229277e-05
GC_3_1289 b_3 NI_3 NS_1289 0 -7.8146230778624731e-08
GC_3_1290 b_3 NI_3 NS_1290 0 9.5809245687976838e-07
GC_3_1291 b_3 NI_3 NS_1291 0 -7.9221105587554165e-06
GC_3_1292 b_3 NI_3 NS_1292 0 -8.5842983504962023e-06
GC_3_1293 b_3 NI_3 NS_1293 0 -6.3256724637475604e-07
GC_3_1294 b_3 NI_3 NS_1294 0 -2.1422062831179413e-06
GC_3_1295 b_3 NI_3 NS_1295 0 -1.4556512303338171e-08
GC_3_1296 b_3 NI_3 NS_1296 0 1.1898573444286794e-06
GC_3_1297 b_3 NI_3 NS_1297 0 -7.7141138085066465e-06
GC_3_1298 b_3 NI_3 NS_1298 0 1.9653040851883898e-06
GC_3_1299 b_3 NI_3 NS_1299 0 2.3902170250166915e-07
GC_3_1300 b_3 NI_3 NS_1300 0 -1.6696989031789351e-06
GC_3_1301 b_3 NI_3 NS_1301 0 1.1429316660081859e-06
GC_3_1302 b_3 NI_3 NS_1302 0 3.0633318614611127e-06
GC_3_1303 b_3 NI_3 NS_1303 0 -9.6195302680345090e-07
GC_3_1304 b_3 NI_3 NS_1304 0 2.0271908840629301e-06
GC_3_1305 b_3 NI_3 NS_1305 0 4.5489752459104979e-07
GC_3_1306 b_3 NI_3 NS_1306 0 -1.2226879406804894e-06
GC_3_1307 b_3 NI_3 NS_1307 0 3.2356557403414747e-06
GC_3_1308 b_3 NI_3 NS_1308 0 -8.8238422670244767e-07
GC_3_1309 b_3 NI_3 NS_1309 0 -1.6005496647670098e-07
GC_3_1310 b_3 NI_3 NS_1310 0 5.0797650344394727e-07
GC_3_1311 b_3 NI_3 NS_1311 0 -8.4404626621265651e-07
GC_3_1312 b_3 NI_3 NS_1312 0 -4.1916142125100484e-07
GC_3_1313 b_3 NI_3 NS_1313 0 9.8705305615510593e-07
GC_3_1314 b_3 NI_3 NS_1314 0 -1.2634880496292523e-06
GC_3_1315 b_3 NI_3 NS_1315 0 1.4385530462802324e-06
GC_3_1316 b_3 NI_3 NS_1316 0 -5.6892575054487458e-07
GC_3_1317 b_3 NI_3 NS_1317 0 -3.3372296134157854e-08
GC_3_1318 b_3 NI_3 NS_1318 0 9.4898114912483485e-08
GC_3_1319 b_3 NI_3 NS_1319 0 -5.9608893443382612e-07
GC_3_1320 b_3 NI_3 NS_1320 0 -3.3988583218085019e-07
GC_3_1321 b_3 NI_3 NS_1321 0 9.6297769847572539e-07
GC_3_1322 b_3 NI_3 NS_1322 0 -1.0755627528279551e-06
GC_3_1323 b_3 NI_3 NS_1323 0 1.3913823101534867e-06
GC_3_1324 b_3 NI_3 NS_1324 0 -1.2415325144054453e-06
GC_3_1325 b_3 NI_3 NS_1325 0 1.6086340407201491e-07
GC_3_1326 b_3 NI_3 NS_1326 0 -4.5335282303180441e-08
GC_3_1327 b_3 NI_3 NS_1327 0 -4.8806037852542490e-07
GC_3_1328 b_3 NI_3 NS_1328 0 -5.0217567844356353e-07
GC_3_1329 b_3 NI_3 NS_1329 0 1.0601441219523552e-06
GC_3_1330 b_3 NI_3 NS_1330 0 -7.9957717039042260e-07
GC_3_1331 b_3 NI_3 NS_1331 0 1.2253761506320211e-06
GC_3_1332 b_3 NI_3 NS_1332 0 -2.1157340415443674e-06
GC_3_1333 b_3 NI_3 NS_1333 0 4.9451683030933754e-07
GC_3_1334 b_3 NI_3 NS_1334 0 -2.5501268423346859e-07
GC_3_1335 b_3 NI_3 NS_1335 0 -2.4640565269127777e-07
GC_3_1336 b_3 NI_3 NS_1336 0 -9.1750762572453581e-07
GC_3_1337 b_3 NI_3 NS_1337 0 1.9158084970491687e-06
GC_3_1338 b_3 NI_3 NS_1338 0 -9.9682757765938075e-07
GC_3_1339 b_3 NI_3 NS_1339 0 -8.0875088346273894e-06
GC_3_1340 b_3 NI_3 NS_1340 0 -9.1346814494608813e-07
GC_3_1341 b_3 NI_3 NS_1341 0 -3.1591125772568699e-07
GC_3_1342 b_3 NI_3 NS_1342 0 -3.6199105438333280e-06
GC_3_1343 b_3 NI_3 NS_1343 0 -4.8932411436626737e-08
GC_3_1344 b_3 NI_3 NS_1344 0 -3.3150758983546679e-08
GC_3_1345 b_3 NI_3 NS_1345 0 -1.0396024639549672e-07
GC_3_1346 b_3 NI_3 NS_1346 0 -1.2351431339897209e-06
GC_3_1347 b_3 NI_3 NS_1347 0 -1.0202889883578535e-06
GC_3_1348 b_3 NI_3 NS_1348 0 -6.6669642922159300e-07
GC_3_1349 b_3 NI_3 NS_1349 0 1.4550417169071718e-06
GC_3_1350 b_3 NI_3 NS_1350 0 -7.5894691255911763e-07
GC_3_1351 b_3 NI_3 NS_1351 0 1.9403522662374919e-06
GC_3_1352 b_3 NI_3 NS_1352 0 -1.8687522571719934e-06
GC_3_1353 b_3 NI_3 NS_1353 0 -2.2166647943887367e-07
GC_3_1354 b_3 NI_3 NS_1354 0 3.2466588246765102e-07
GC_3_1355 b_3 NI_3 NS_1355 0 2.1427942366090408e-07
GC_3_1356 b_3 NI_3 NS_1356 0 5.2885352493133305e-07
GC_3_1357 b_3 NI_3 NS_1357 0 -1.0742406791840054e-07
GC_3_1358 b_3 NI_3 NS_1358 0 -2.8271622058946143e-07
GC_3_1359 b_3 NI_3 NS_1359 0 7.8977422832126255e-09
GC_3_1360 b_3 NI_3 NS_1360 0 -9.5823911353544094e-08
GC_3_1361 b_3 NI_3 NS_1361 0 -8.8821567292426217e-08
GC_3_1362 b_3 NI_3 NS_1362 0 4.1483700995514124e-08
GC_3_1363 b_3 NI_3 NS_1363 0 -1.2204426605143805e-07
GC_3_1364 b_3 NI_3 NS_1364 0 -5.3450742015195159e-08
GC_3_1365 b_3 NI_3 NS_1365 0 6.1485649351581913e-12
GC_3_1366 b_3 NI_3 NS_1366 0 -1.7071122529261468e-12
GC_3_1367 b_3 NI_3 NS_1367 0 3.5216523701673846e-10
GC_3_1368 b_3 NI_3 NS_1368 0 6.9300684425809031e-10
GD_3_1 b_3 NI_3 NA_1 0 1.3006422144172181e-02
GD_3_2 b_3 NI_3 NA_2 0 5.9084066587420487e-04
GD_3_3 b_3 NI_3 NA_3 0 -8.6867583427960773e-03
GD_3_4 b_3 NI_3 NA_4 0 -4.2441749448996948e-03
GD_3_5 b_3 NI_3 NA_5 0 1.0032020473432268e-04
GD_3_6 b_3 NI_3 NA_6 0 2.7000168285998986e-05
GD_3_7 b_3 NI_3 NA_7 0 3.4014531115666674e-06
GD_3_8 b_3 NI_3 NA_8 0 1.1832415158620740e-06
GD_3_9 b_3 NI_3 NA_9 0 -5.5534209837450566e-06
GD_3_10 b_3 NI_3 NA_10 0 4.7471719663156571e-07
GD_3_11 b_3 NI_3 NA_11 0 -1.8690895286311346e-06
GD_3_12 b_3 NI_3 NA_12 0 5.6258463865609864e-06
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 2.9495792000684591e-03
GC_4_2 b_4 NI_4 NS_2 0 -6.1234121802852890e-04
GC_4_3 b_4 NI_4 NS_3 0 2.7949878545371285e-08
GC_4_4 b_4 NI_4 NS_4 0 -3.1702392990733477e-08
GC_4_5 b_4 NI_4 NS_5 0 2.0347269738621966e-04
GC_4_6 b_4 NI_4 NS_6 0 1.3799469265289848e-04
GC_4_7 b_4 NI_4 NS_7 0 5.6259274658273855e-04
GC_4_8 b_4 NI_4 NS_8 0 2.6570823116899890e-04
GC_4_9 b_4 NI_4 NS_9 0 3.1064666446230099e-03
GC_4_10 b_4 NI_4 NS_10 0 -2.2048919836966628e-03
GC_4_11 b_4 NI_4 NS_11 0 -1.5822541471011678e-03
GC_4_12 b_4 NI_4 NS_12 0 -2.6870784037591440e-03
GC_4_13 b_4 NI_4 NS_13 0 -2.0496554919685519e-03
GC_4_14 b_4 NI_4 NS_14 0 -3.7885102461833885e-03
GC_4_15 b_4 NI_4 NS_15 0 -4.9745613813943958e-03
GC_4_16 b_4 NI_4 NS_16 0 -1.5415311515132994e-03
GC_4_17 b_4 NI_4 NS_17 0 2.9290575022278108e-04
GC_4_18 b_4 NI_4 NS_18 0 1.9565159751352873e-04
GC_4_19 b_4 NI_4 NS_19 0 -2.8663291493454743e-03
GC_4_20 b_4 NI_4 NS_20 0 -9.5746385289233443e-04
GC_4_21 b_4 NI_4 NS_21 0 -2.2151871598365583e-02
GC_4_22 b_4 NI_4 NS_22 0 -1.0226316681973850e-02
GC_4_23 b_4 NI_4 NS_23 0 1.1324969823597005e-03
GC_4_24 b_4 NI_4 NS_24 0 2.0395321152750463e-02
GC_4_25 b_4 NI_4 NS_25 0 -5.8416211655905707e-03
GC_4_26 b_4 NI_4 NS_26 0 4.6116292314381862e-03
GC_4_27 b_4 NI_4 NS_27 0 5.7171509138104959e-03
GC_4_28 b_4 NI_4 NS_28 0 3.4516071269026734e-02
GC_4_29 b_4 NI_4 NS_29 0 8.0342763895865747e-03
GC_4_30 b_4 NI_4 NS_30 0 2.7930238811015983e-03
GC_4_31 b_4 NI_4 NS_31 0 -7.7724209734374100e-03
GC_4_32 b_4 NI_4 NS_32 0 2.9556754670475062e-02
GC_4_33 b_4 NI_4 NS_33 0 5.0768429833649605e-02
GC_4_34 b_4 NI_4 NS_34 0 -2.0072962229514092e-02
GC_4_35 b_4 NI_4 NS_35 0 7.9195784236166349e-03
GC_4_36 b_4 NI_4 NS_36 0 -1.6364410927427924e-03
GC_4_37 b_4 NI_4 NS_37 0 2.9084859403911607e-02
GC_4_38 b_4 NI_4 NS_38 0 -2.6464736322709379e-02
GC_4_39 b_4 NI_4 NS_39 0 -6.7250675992636885e-03
GC_4_40 b_4 NI_4 NS_40 0 -9.8822055516598253e-03
GC_4_41 b_4 NI_4 NS_41 0 8.4630825871619113e-03
GC_4_42 b_4 NI_4 NS_42 0 -8.0277978646210672e-03
GC_4_43 b_4 NI_4 NS_43 0 -1.8994952132973579e-02
GC_4_44 b_4 NI_4 NS_44 0 -2.5238421796827698e-02
GC_4_45 b_4 NI_4 NS_45 0 -5.4717849928970601e-03
GC_4_46 b_4 NI_4 NS_46 0 -2.8547841807847474e-03
GC_4_47 b_4 NI_4 NS_47 0 -1.7741073793125079e-02
GC_4_48 b_4 NI_4 NS_48 0 -1.3132230193186241e-02
GC_4_49 b_4 NI_4 NS_49 0 -4.8178005931692192e-03
GC_4_50 b_4 NI_4 NS_50 0 1.2541404083866248e-02
GC_4_51 b_4 NI_4 NS_51 0 -3.4590900573936768e-03
GC_4_52 b_4 NI_4 NS_52 0 1.5412381717933149e-03
GC_4_53 b_4 NI_4 NS_53 0 -7.1865143851114661e-04
GC_4_54 b_4 NI_4 NS_54 0 7.0058605723982261e-03
GC_4_55 b_4 NI_4 NS_55 0 1.8820413852480909e-03
GC_4_56 b_4 NI_4 NS_56 0 8.5748616983273912e-05
GC_4_57 b_4 NI_4 NS_57 0 3.1400281668075175e-04
GC_4_58 b_4 NI_4 NS_58 0 -1.9467014138642843e-03
GC_4_59 b_4 NI_4 NS_59 0 -1.8563352620861407e-03
GC_4_60 b_4 NI_4 NS_60 0 -1.6182088780022431e-03
GC_4_61 b_4 NI_4 NS_61 0 -2.1290960678084334e-03
GC_4_62 b_4 NI_4 NS_62 0 1.6850433436621393e-03
GC_4_63 b_4 NI_4 NS_63 0 7.6361045457538641e-04
GC_4_64 b_4 NI_4 NS_64 0 1.8527512955730910e-04
GC_4_65 b_4 NI_4 NS_65 0 -6.9730354299662772e-04
GC_4_66 b_4 NI_4 NS_66 0 -1.6780703351843985e-03
GC_4_67 b_4 NI_4 NS_67 0 -2.6815282153668154e-03
GC_4_68 b_4 NI_4 NS_68 0 -8.2749160389724663e-04
GC_4_69 b_4 NI_4 NS_69 0 -4.9989688347921264e-04
GC_4_70 b_4 NI_4 NS_70 0 2.9288639052344376e-03
GC_4_71 b_4 NI_4 NS_71 0 1.3533574681095025e-03
GC_4_72 b_4 NI_4 NS_72 0 -8.5805587491199098e-04
GC_4_73 b_4 NI_4 NS_73 0 -2.4189247490921167e-03
GC_4_74 b_4 NI_4 NS_74 0 -2.2676209715785317e-03
GC_4_75 b_4 NI_4 NS_75 0 -3.5540455350823725e-03
GC_4_76 b_4 NI_4 NS_76 0 7.4852673594070259e-04
GC_4_77 b_4 NI_4 NS_77 0 2.4633829809719010e-03
GC_4_78 b_4 NI_4 NS_78 0 3.0182799545515294e-03
GC_4_79 b_4 NI_4 NS_79 0 9.8455399573227722e-04
GC_4_80 b_4 NI_4 NS_80 0 -2.9418100013680337e-03
GC_4_81 b_4 NI_4 NS_81 0 -4.7678001553018729e-03
GC_4_82 b_4 NI_4 NS_82 0 5.4340315943759746e-05
GC_4_83 b_4 NI_4 NS_83 0 -1.7083702904996689e-03
GC_4_84 b_4 NI_4 NS_84 0 3.7124268883669651e-03
GC_4_85 b_4 NI_4 NS_85 0 -7.6587733078630046e-04
GC_4_86 b_4 NI_4 NS_86 0 1.5006835018716784e-03
GC_4_87 b_4 NI_4 NS_87 0 3.2213013519404440e-03
GC_4_88 b_4 NI_4 NS_88 0 -1.3508686604321795e-03
GC_4_89 b_4 NI_4 NS_89 0 -2.9326239323711017e-06
GC_4_90 b_4 NI_4 NS_90 0 8.7469590733944450e-06
GC_4_91 b_4 NI_4 NS_91 0 -1.8200422811098234e-03
GC_4_92 b_4 NI_4 NS_92 0 -2.5277365471798839e-03
GC_4_93 b_4 NI_4 NS_93 0 -2.4072537620752968e-03
GC_4_94 b_4 NI_4 NS_94 0 2.4886636542996187e-03
GC_4_95 b_4 NI_4 NS_95 0 1.0142618786233573e-03
GC_4_96 b_4 NI_4 NS_96 0 2.4256808564866224e-03
GC_4_97 b_4 NI_4 NS_97 0 8.5775914850749670e-04
GC_4_98 b_4 NI_4 NS_98 0 -2.6994858278521056e-03
GC_4_99 b_4 NI_4 NS_99 0 -3.0644780784384336e-04
GC_4_100 b_4 NI_4 NS_100 0 1.6741356971131619e-03
GC_4_101 b_4 NI_4 NS_101 0 -1.7840539173598236e-03
GC_4_102 b_4 NI_4 NS_102 0 -3.1181076983861195e-04
GC_4_103 b_4 NI_4 NS_103 0 1.4004539394093650e-03
GC_4_104 b_4 NI_4 NS_104 0 1.9709616314733010e-03
GC_4_105 b_4 NI_4 NS_105 0 1.0449287584058720e-03
GC_4_106 b_4 NI_4 NS_106 0 -2.2998045206167159e-03
GC_4_107 b_4 NI_4 NS_107 0 -6.9799496549654389e-04
GC_4_108 b_4 NI_4 NS_108 0 -1.4668898646361325e-03
GC_4_109 b_4 NI_4 NS_109 0 -1.3735491569299017e-03
GC_4_110 b_4 NI_4 NS_110 0 -3.1252860486514025e-04
GC_4_111 b_4 NI_4 NS_111 0 7.1030031780261722e-09
GC_4_112 b_4 NI_4 NS_112 0 -2.4709996914266187e-08
GC_4_113 b_4 NI_4 NS_113 0 -4.5275395999440338e-07
GC_4_114 b_4 NI_4 NS_114 0 1.6341836862293618e-06
GC_4_115 b_4 NI_4 NS_115 0 7.7623631688561491e-03
GC_4_116 b_4 NI_4 NS_116 0 -1.6012429819176404e-03
GC_4_117 b_4 NI_4 NS_117 0 -1.2109163074591947e-08
GC_4_118 b_4 NI_4 NS_118 0 -8.8417590504104604e-07
GC_4_119 b_4 NI_4 NS_119 0 1.0417924325171096e-04
GC_4_120 b_4 NI_4 NS_120 0 -5.1170037849583583e-04
GC_4_121 b_4 NI_4 NS_121 0 -1.9362887985216318e-03
GC_4_122 b_4 NI_4 NS_122 0 -5.9765172108031453e-04
GC_4_123 b_4 NI_4 NS_123 0 2.9418128645987730e-03
GC_4_124 b_4 NI_4 NS_124 0 2.2635993047106233e-03
GC_4_125 b_4 NI_4 NS_125 0 -3.5704327589433219e-03
GC_4_126 b_4 NI_4 NS_126 0 -3.0490673763529279e-03
GC_4_127 b_4 NI_4 NS_127 0 -1.7073725775676538e-03
GC_4_128 b_4 NI_4 NS_128 0 5.8427846668897346e-03
GC_4_129 b_4 NI_4 NS_129 0 4.3666970100515942e-03
GC_4_130 b_4 NI_4 NS_130 0 -2.4750965250182272e-03
GC_4_131 b_4 NI_4 NS_131 0 -1.1000888431063059e-04
GC_4_132 b_4 NI_4 NS_132 0 -1.0334512900322201e-04
GC_4_133 b_4 NI_4 NS_133 0 -4.4523052985084429e-03
GC_4_134 b_4 NI_4 NS_134 0 -9.2440307397423024e-04
GC_4_135 b_4 NI_4 NS_135 0 9.1241543833593206e-03
GC_4_136 b_4 NI_4 NS_136 0 1.7784746375376241e-02
GC_4_137 b_4 NI_4 NS_137 0 -4.0272971001971162e-03
GC_4_138 b_4 NI_4 NS_138 0 -1.7846771806133508e-02
GC_4_139 b_4 NI_4 NS_139 0 -8.2177715191633569e-03
GC_4_140 b_4 NI_4 NS_140 0 4.1736008749428703e-03
GC_4_141 b_4 NI_4 NS_141 0 1.7063484686914848e-02
GC_4_142 b_4 NI_4 NS_142 0 -4.3909977323247477e-04
GC_4_143 b_4 NI_4 NS_143 0 -9.2787160081969702e-03
GC_4_144 b_4 NI_4 NS_144 0 -3.2069945516611481e-03
GC_4_145 b_4 NI_4 NS_145 0 -1.3713361965252649e-02
GC_4_146 b_4 NI_4 NS_146 0 2.2836239953912263e-02
GC_4_147 b_4 NI_4 NS_147 0 2.2839552393873409e-02
GC_4_148 b_4 NI_4 NS_148 0 -2.2669171312837626e-02
GC_4_149 b_4 NI_4 NS_149 0 -9.2392853314965575e-03
GC_4_150 b_4 NI_4 NS_150 0 9.0811376156037162e-04
GC_4_151 b_4 NI_4 NS_151 0 1.8480132532700803e-02
GC_4_152 b_4 NI_4 NS_152 0 6.2442241031404194e-03
GC_4_153 b_4 NI_4 NS_153 0 -9.1760808824884622e-03
GC_4_154 b_4 NI_4 NS_154 0 -9.4609794904917510e-03
GC_4_155 b_4 NI_4 NS_155 0 -9.9743264482778839e-03
GC_4_156 b_4 NI_4 NS_156 0 6.3961885386921791e-03
GC_4_157 b_4 NI_4 NS_157 0 1.6838481102828842e-02
GC_4_158 b_4 NI_4 NS_158 0 -4.8501205082519955e-03
GC_4_159 b_4 NI_4 NS_159 0 -7.2149225369588328e-03
GC_4_160 b_4 NI_4 NS_160 0 -3.4092354578831243e-03
GC_4_161 b_4 NI_4 NS_161 0 6.8281954720174716e-03
GC_4_162 b_4 NI_4 NS_162 0 1.3297053324887518e-02
GC_4_163 b_4 NI_4 NS_163 0 -1.8195824533954650e-03
GC_4_164 b_4 NI_4 NS_164 0 -1.4401720113427167e-02
GC_4_165 b_4 NI_4 NS_165 0 -4.9860069971144885e-03
GC_4_166 b_4 NI_4 NS_166 0 1.0394629019383924e-03
GC_4_167 b_4 NI_4 NS_167 0 6.0026097697613769e-03
GC_4_168 b_4 NI_4 NS_168 0 -1.1030574878134907e-03
GC_4_169 b_4 NI_4 NS_169 0 -3.4642734364297044e-03
GC_4_170 b_4 NI_4 NS_170 0 -1.0876297929216018e-03
GC_4_171 b_4 NI_4 NS_171 0 2.7180517521858422e-03
GC_4_172 b_4 NI_4 NS_172 0 -5.0782105589794707e-04
GC_4_173 b_4 NI_4 NS_173 0 -3.2964856509058501e-03
GC_4_174 b_4 NI_4 NS_174 0 -2.8951315922029681e-03
GC_4_175 b_4 NI_4 NS_175 0 2.0159621881415679e-03
GC_4_176 b_4 NI_4 NS_176 0 7.7577849499975698e-04
GC_4_177 b_4 NI_4 NS_177 0 -2.0162760629968343e-03
GC_4_178 b_4 NI_4 NS_178 0 -9.6646512748903843e-04
GC_4_179 b_4 NI_4 NS_179 0 2.1216220343240077e-03
GC_4_180 b_4 NI_4 NS_180 0 -1.4709118335064430e-03
GC_4_181 b_4 NI_4 NS_181 0 -4.1847944562860223e-03
GC_4_182 b_4 NI_4 NS_182 0 -1.8129441562800082e-03
GC_4_183 b_4 NI_4 NS_183 0 2.3697817652706642e-03
GC_4_184 b_4 NI_4 NS_184 0 -3.7075719351620272e-04
GC_4_185 b_4 NI_4 NS_185 0 -3.0172215283794366e-03
GC_4_186 b_4 NI_4 NS_186 0 4.6233692494282083e-04
GC_4_187 b_4 NI_4 NS_187 0 2.7064446320437131e-03
GC_4_188 b_4 NI_4 NS_188 0 -2.7282256796781223e-03
GC_4_189 b_4 NI_4 NS_189 0 -5.0393282341870465e-03
GC_4_190 b_4 NI_4 NS_190 0 -1.2783040350739932e-04
GC_4_191 b_4 NI_4 NS_191 0 2.4346778108655033e-03
GC_4_192 b_4 NI_4 NS_192 0 -2.1719821015915575e-03
GC_4_193 b_4 NI_4 NS_193 0 -3.2449804044218924e-03
GC_4_194 b_4 NI_4 NS_194 0 2.6005310513343934e-03
GC_4_195 b_4 NI_4 NS_195 0 1.7436680446392184e-03
GC_4_196 b_4 NI_4 NS_196 0 -4.7503555602724798e-03
GC_4_197 b_4 NI_4 NS_197 0 -3.6339959509179673e-03
GC_4_198 b_4 NI_4 NS_198 0 2.5967283187582329e-03
GC_4_199 b_4 NI_4 NS_199 0 -2.8319057300752160e-03
GC_4_200 b_4 NI_4 NS_200 0 3.9895611144148083e-03
GC_4_201 b_4 NI_4 NS_201 0 -2.2141465850228584e-04
GC_4_202 b_4 NI_4 NS_202 0 -4.2135156478536285e-03
GC_4_203 b_4 NI_4 NS_203 0 -9.8958396329086554e-06
GC_4_204 b_4 NI_4 NS_204 0 7.5257580403191724e-06
GC_4_205 b_4 NI_4 NS_205 0 -1.3539532717195106e-03
GC_4_206 b_4 NI_4 NS_206 0 3.3754867364945342e-03
GC_4_207 b_4 NI_4 NS_207 0 -9.6985114954640226e-04
GC_4_208 b_4 NI_4 NS_208 0 -4.3479519129108633e-03
GC_4_209 b_4 NI_4 NS_209 0 -1.0009104611071349e-03
GC_4_210 b_4 NI_4 NS_210 0 2.2213067654426079e-03
GC_4_211 b_4 NI_4 NS_211 0 -1.6517261451241970e-03
GC_4_212 b_4 NI_4 NS_212 0 -4.4093120919240260e-03
GC_4_213 b_4 NI_4 NS_213 0 -1.4483164113464715e-03
GC_4_214 b_4 NI_4 NS_214 0 -2.4971461095295100e-03
GC_4_215 b_4 NI_4 NS_215 0 7.8219531513637388e-04
GC_4_216 b_4 NI_4 NS_216 0 2.5933467042086496e-03
GC_4_217 b_4 NI_4 NS_217 0 -6.9628504516106742e-04
GC_4_218 b_4 NI_4 NS_218 0 2.8792034901524276e-03
GC_4_219 b_4 NI_4 NS_219 0 -1.4353710703652587e-03
GC_4_220 b_4 NI_4 NS_220 0 -2.7718619392436326e-03
GC_4_221 b_4 NI_4 NS_221 0 -1.1678495857963560e-03
GC_4_222 b_4 NI_4 NS_222 0 2.6661993124948834e-03
GC_4_223 b_4 NI_4 NS_223 0 7.8075943466382914e-04
GC_4_224 b_4 NI_4 NS_224 0 -1.8746156136013046e-03
GC_4_225 b_4 NI_4 NS_225 0 2.3789690379723077e-08
GC_4_226 b_4 NI_4 NS_226 0 -6.0253482765116211e-08
GC_4_227 b_4 NI_4 NS_227 0 -9.0373275434108698e-07
GC_4_228 b_4 NI_4 NS_228 0 3.2031385932389857e-06
GC_4_229 b_4 NI_4 NS_229 0 1.8439409624874996e-02
GC_4_230 b_4 NI_4 NS_230 0 6.7473522172684002e-03
GC_4_231 b_4 NI_4 NS_231 0 4.6777105134428026e-07
GC_4_232 b_4 NI_4 NS_232 0 1.4628662474477701e-06
GC_4_233 b_4 NI_4 NS_233 0 6.0883192874167024e-03
GC_4_234 b_4 NI_4 NS_234 0 1.8079505775020098e-03
GC_4_235 b_4 NI_4 NS_235 0 -6.0692963087718961e-03
GC_4_236 b_4 NI_4 NS_236 0 -6.1756069281944891e-04
GC_4_237 b_4 NI_4 NS_237 0 7.3051306825333050e-03
GC_4_238 b_4 NI_4 NS_238 0 -1.2868558987382010e-02
GC_4_239 b_4 NI_4 NS_239 0 8.4477910503870553e-03
GC_4_240 b_4 NI_4 NS_240 0 -2.4311197144477102e-04
GC_4_241 b_4 NI_4 NS_241 0 -9.6438190479626040e-03
GC_4_242 b_4 NI_4 NS_242 0 2.6146352919277104e-03
GC_4_243 b_4 NI_4 NS_243 0 -8.8620581363026835e-03
GC_4_244 b_4 NI_4 NS_244 0 -2.4393956645971427e-02
GC_4_245 b_4 NI_4 NS_245 0 -8.6179941024843842e-04
GC_4_246 b_4 NI_4 NS_246 0 4.1810183765506603e-03
GC_4_247 b_4 NI_4 NS_247 0 7.1873813893271162e-03
GC_4_248 b_4 NI_4 NS_248 0 -1.0295269902994800e-03
GC_4_249 b_4 NI_4 NS_249 0 -2.5161037733684031e-02
GC_4_250 b_4 NI_4 NS_250 0 4.8306268573339852e-03
GC_4_251 b_4 NI_4 NS_251 0 -1.9676958705501062e-02
GC_4_252 b_4 NI_4 NS_252 0 8.9689435040783715e-04
GC_4_253 b_4 NI_4 NS_253 0 1.0760365757916583e-02
GC_4_254 b_4 NI_4 NS_254 0 -2.7834372363887113e-03
GC_4_255 b_4 NI_4 NS_255 0 -4.7873570543613495e-03
GC_4_256 b_4 NI_4 NS_256 0 4.5022305268941458e-02
GC_4_257 b_4 NI_4 NS_257 0 -1.2656403541193396e-02
GC_4_258 b_4 NI_4 NS_258 0 -2.7346933271607386e-04
GC_4_259 b_4 NI_4 NS_259 0 1.5916984819721369e-02
GC_4_260 b_4 NI_4 NS_260 0 -4.0520132544199739e-03
GC_4_261 b_4 NI_4 NS_261 0 3.2200849067182943e-02
GC_4_262 b_4 NI_4 NS_262 0 1.8584186257918040e-02
GC_4_263 b_4 NI_4 NS_263 0 -1.2597834021689298e-02
GC_4_264 b_4 NI_4 NS_264 0 1.6049566381409928e-04
GC_4_265 b_4 NI_4 NS_265 0 1.7204281161243330e-02
GC_4_266 b_4 NI_4 NS_266 0 -3.5163275043345134e-02
GC_4_267 b_4 NI_4 NS_267 0 1.4015762398782293e-02
GC_4_268 b_4 NI_4 NS_268 0 4.7859300813441943e-03
GC_4_269 b_4 NI_4 NS_269 0 -1.4402586569019035e-02
GC_4_270 b_4 NI_4 NS_270 0 2.3849088542255193e-04
GC_4_271 b_4 NI_4 NS_271 0 -2.0144561931922683e-02
GC_4_272 b_4 NI_4 NS_272 0 -3.0186695167525677e-02
GC_4_273 b_4 NI_4 NS_273 0 1.0530763157968616e-02
GC_4_274 b_4 NI_4 NS_274 0 3.5935602272290984e-03
GC_4_275 b_4 NI_4 NS_275 0 -2.6797879283576832e-02
GC_4_276 b_4 NI_4 NS_276 0 1.1150463481418066e-02
GC_4_277 b_4 NI_4 NS_277 0 -1.4133838396323400e-02
GC_4_278 b_4 NI_4 NS_278 0 -2.5194000435845095e-03
GC_4_279 b_4 NI_4 NS_279 0 7.5552452397437825e-03
GC_4_280 b_4 NI_4 NS_280 0 1.5923785527835652e-03
GC_4_281 b_4 NI_4 NS_281 0 -8.5556981780459849e-04
GC_4_282 b_4 NI_4 NS_282 0 2.4403095578915977e-02
GC_4_283 b_4 NI_4 NS_283 0 -7.6201794021305965e-03
GC_4_284 b_4 NI_4 NS_284 0 2.8212088392895511e-04
GC_4_285 b_4 NI_4 NS_285 0 -5.5980342287930264e-04
GC_4_286 b_4 NI_4 NS_286 0 -5.5368776786066803e-03
GC_4_287 b_4 NI_4 NS_287 0 8.2660041907530839e-03
GC_4_288 b_4 NI_4 NS_288 0 7.0201199312176039e-03
GC_4_289 b_4 NI_4 NS_289 0 -7.1916634664827902e-04
GC_4_290 b_4 NI_4 NS_290 0 1.2092481870869795e-02
GC_4_291 b_4 NI_4 NS_291 0 -5.1474318566086209e-03
GC_4_292 b_4 NI_4 NS_292 0 -1.3699948903729829e-04
GC_4_293 b_4 NI_4 NS_293 0 -1.8303920056844494e-03
GC_4_294 b_4 NI_4 NS_294 0 -5.1700766224467226e-03
GC_4_295 b_4 NI_4 NS_295 0 9.2879112937599186e-03
GC_4_296 b_4 NI_4 NS_296 0 5.4154418169098670e-03
GC_4_297 b_4 NI_4 NS_297 0 3.5152834491960303e-03
GC_4_298 b_4 NI_4 NS_298 0 1.1689789824763288e-02
GC_4_299 b_4 NI_4 NS_299 0 -6.1370069651302869e-03
GC_4_300 b_4 NI_4 NS_300 0 1.4286277741343476e-03
GC_4_301 b_4 NI_4 NS_301 0 -2.8171746200841273e-03
GC_4_302 b_4 NI_4 NS_302 0 -7.3462681257854077e-03
GC_4_303 b_4 NI_4 NS_303 0 9.9561207557705977e-03
GC_4_304 b_4 NI_4 NS_304 0 3.3689015303838168e-03
GC_4_305 b_4 NI_4 NS_305 0 8.1685764162415467e-03
GC_4_306 b_4 NI_4 NS_306 0 1.0244024154684108e-02
GC_4_307 b_4 NI_4 NS_307 0 -6.9844654808815243e-03
GC_4_308 b_4 NI_4 NS_308 0 2.9355138333100263e-03
GC_4_309 b_4 NI_4 NS_309 0 -5.6336390414053750e-03
GC_4_310 b_4 NI_4 NS_310 0 -8.0966143239036472e-03
GC_4_311 b_4 NI_4 NS_311 0 9.8584761748458111e-03
GC_4_312 b_4 NI_4 NS_312 0 5.4631783153492636e-04
GC_4_313 b_4 NI_4 NS_313 0 -1.0941980381302022e-02
GC_4_314 b_4 NI_4 NS_314 0 1.2300248078408047e-02
GC_4_315 b_4 NI_4 NS_315 0 9.6442776560288282e-03
GC_4_316 b_4 NI_4 NS_316 0 5.0348793921206432e-03
GC_4_317 b_4 NI_4 NS_317 0 -1.9883257539694807e-05
GC_4_318 b_4 NI_4 NS_318 0 3.1661380921318448e-05
GC_4_319 b_4 NI_4 NS_319 0 -7.1319479659557134e-03
GC_4_320 b_4 NI_4 NS_320 0 4.4777063058622051e-03
GC_4_321 b_4 NI_4 NS_321 0 -7.6765613911509035e-03
GC_4_322 b_4 NI_4 NS_322 0 -5.3213649992725461e-03
GC_4_323 b_4 NI_4 NS_323 0 9.5165634682715800e-03
GC_4_324 b_4 NI_4 NS_324 0 -1.7361931039336824e-03
GC_4_325 b_4 NI_4 NS_325 0 1.2475075402011489e-02
GC_4_326 b_4 NI_4 NS_326 0 -1.4048039409351501e-03
GC_4_327 b_4 NI_4 NS_327 0 -5.0716681954236387e-03
GC_4_328 b_4 NI_4 NS_328 0 -2.7496731600631782e-03
GC_4_329 b_4 NI_4 NS_329 0 -2.2244068800202697e-03
GC_4_330 b_4 NI_4 NS_330 0 6.6017975307154702e-03
GC_4_331 b_4 NI_4 NS_331 0 8.9571101847764432e-03
GC_4_332 b_4 NI_4 NS_332 0 1.3095225880173375e-04
GC_4_333 b_4 NI_4 NS_333 0 1.2487333296179350e-02
GC_4_334 b_4 NI_4 NS_334 0 1.7801034493617896e-03
GC_4_335 b_4 NI_4 NS_335 0 -5.3781333782729002e-03
GC_4_336 b_4 NI_4 NS_336 0 4.1549292859347957e-03
GC_4_337 b_4 NI_4 NS_337 0 -1.8500367292116242e-03
GC_4_338 b_4 NI_4 NS_338 0 -5.6869519876894658e-03
GC_4_339 b_4 NI_4 NS_339 0 2.0790328499661129e-07
GC_4_340 b_4 NI_4 NS_340 0 -2.4564439341175698e-07
GC_4_341 b_4 NI_4 NS_341 0 -1.1505429974016690e-05
GC_4_342 b_4 NI_4 NS_342 0 1.8244729530072067e-05
GC_4_343 b_4 NI_4 NS_343 0 -1.4190097407436177e-02
GC_4_344 b_4 NI_4 NS_344 0 1.3879298607381090e-03
GC_4_345 b_4 NI_4 NS_345 0 -2.6214589268034229e-07
GC_4_346 b_4 NI_4 NS_346 0 -3.7469053601666173e-06
GC_4_347 b_4 NI_4 NS_347 0 -2.9950712352338170e-04
GC_4_348 b_4 NI_4 NS_348 0 4.7112868964953406e-04
GC_4_349 b_4 NI_4 NS_349 0 1.2936041298229365e-03
GC_4_350 b_4 NI_4 NS_350 0 5.6342135820482663e-04
GC_4_351 b_4 NI_4 NS_351 0 -2.7928189552436206e-03
GC_4_352 b_4 NI_4 NS_352 0 -7.1086086409722119e-04
GC_4_353 b_4 NI_4 NS_353 0 3.5977247957128668e-03
GC_4_354 b_4 NI_4 NS_354 0 2.5454554772646994e-03
GC_4_355 b_4 NI_4 NS_355 0 1.1770627409822794e-03
GC_4_356 b_4 NI_4 NS_356 0 -4.1367871145997943e-03
GC_4_357 b_4 NI_4 NS_357 0 -1.5548935818210012e-03
GC_4_358 b_4 NI_4 NS_358 0 2.7530038112833473e-03
GC_4_359 b_4 NI_4 NS_359 0 -3.5992609246607939e-04
GC_4_360 b_4 NI_4 NS_360 0 -2.1737785181832333e-04
GC_4_361 b_4 NI_4 NS_361 0 4.0014076268810213e-03
GC_4_362 b_4 NI_4 NS_362 0 2.5737083876065461e-04
GC_4_363 b_4 NI_4 NS_363 0 -7.3983785450501185e-03
GC_4_364 b_4 NI_4 NS_364 0 -1.3542083605377961e-02
GC_4_365 b_4 NI_4 NS_365 0 4.4843084901334661e-03
GC_4_366 b_4 NI_4 NS_366 0 1.3402111987596320e-02
GC_4_367 b_4 NI_4 NS_367 0 6.7170381911765354e-03
GC_4_368 b_4 NI_4 NS_368 0 -4.0292251491289488e-03
GC_4_369 b_4 NI_4 NS_369 0 -1.3321384901694423e-02
GC_4_370 b_4 NI_4 NS_370 0 6.8614002187479951e-04
GC_4_371 b_4 NI_4 NS_371 0 7.8581343523570855e-03
GC_4_372 b_4 NI_4 NS_372 0 1.8345313325805557e-03
GC_4_373 b_4 NI_4 NS_373 0 1.0514025121400426e-02
GC_4_374 b_4 NI_4 NS_374 0 -1.9642822930250468e-02
GC_4_375 b_4 NI_4 NS_375 0 -1.7746432280184517e-02
GC_4_376 b_4 NI_4 NS_376 0 1.9129827664864821e-02
GC_4_377 b_4 NI_4 NS_377 0 7.6846954657522806e-03
GC_4_378 b_4 NI_4 NS_378 0 -1.4647961155201780e-03
GC_4_379 b_4 NI_4 NS_379 0 -1.5663694621542504e-02
GC_4_380 b_4 NI_4 NS_380 0 -4.7646805759049430e-03
GC_4_381 b_4 NI_4 NS_381 0 8.0859900445670058e-03
GC_4_382 b_4 NI_4 NS_382 0 7.2458421625024184e-03
GC_4_383 b_4 NI_4 NS_383 0 8.1137552717652148e-03
GC_4_384 b_4 NI_4 NS_384 0 -6.0473597232078560e-03
GC_4_385 b_4 NI_4 NS_385 0 -1.3987021078501909e-02
GC_4_386 b_4 NI_4 NS_386 0 4.5766954769174617e-03
GC_4_387 b_4 NI_4 NS_387 0 6.2436852783542265e-03
GC_4_388 b_4 NI_4 NS_388 0 2.3779905771675394e-03
GC_4_389 b_4 NI_4 NS_389 0 -6.3098278837879149e-03
GC_4_390 b_4 NI_4 NS_390 0 -1.1127822870543652e-02
GC_4_391 b_4 NI_4 NS_391 0 2.1503423919025898e-03
GC_4_392 b_4 NI_4 NS_392 0 1.1938071371307571e-02
GC_4_393 b_4 NI_4 NS_393 0 4.2146499023713755e-03
GC_4_394 b_4 NI_4 NS_394 0 -1.1800102681177715e-03
GC_4_395 b_4 NI_4 NS_395 0 -4.9267499346085097e-03
GC_4_396 b_4 NI_4 NS_396 0 1.0434774616388919e-03
GC_4_397 b_4 NI_4 NS_397 0 3.0295902964153159e-03
GC_4_398 b_4 NI_4 NS_398 0 6.8509536985502414e-04
GC_4_399 b_4 NI_4 NS_399 0 -2.2185452352903594e-03
GC_4_400 b_4 NI_4 NS_400 0 4.8987912710523620e-04
GC_4_401 b_4 NI_4 NS_401 0 3.0814361201425664e-03
GC_4_402 b_4 NI_4 NS_402 0 2.2937716711491510e-03
GC_4_403 b_4 NI_4 NS_403 0 -1.5261901203591345e-03
GC_4_404 b_4 NI_4 NS_404 0 -6.8311371182526437e-04
GC_4_405 b_4 NI_4 NS_405 0 1.8943361597397752e-03
GC_4_406 b_4 NI_4 NS_406 0 6.7631458979521409e-04
GC_4_407 b_4 NI_4 NS_407 0 -1.5560152057578775e-03
GC_4_408 b_4 NI_4 NS_408 0 1.2187733574395966e-03
GC_4_409 b_4 NI_4 NS_409 0 3.9927794716663762e-03
GC_4_410 b_4 NI_4 NS_410 0 1.4034783070298270e-03
GC_4_411 b_4 NI_4 NS_411 0 -1.5356610430742232e-03
GC_4_412 b_4 NI_4 NS_412 0 5.9545100615878097e-05
GC_4_413 b_4 NI_4 NS_413 0 2.8410904467841666e-03
GC_4_414 b_4 NI_4 NS_414 0 -6.9178188501784908e-04
GC_4_415 b_4 NI_4 NS_415 0 -1.8626355231391152e-03
GC_4_416 b_4 NI_4 NS_416 0 1.9986033064257791e-03
GC_4_417 b_4 NI_4 NS_417 0 4.9308303887860908e-03
GC_4_418 b_4 NI_4 NS_418 0 -1.7294499576014309e-04
GC_4_419 b_4 NI_4 NS_419 0 -1.6210986159441478e-03
GC_4_420 b_4 NI_4 NS_420 0 9.0628943582759397e-04
GC_4_421 b_4 NI_4 NS_421 0 3.0921495452657542e-03
GC_4_422 b_4 NI_4 NS_422 0 -2.8475032012455596e-03
GC_4_423 b_4 NI_4 NS_423 0 -1.4246752536744083e-03
GC_4_424 b_4 NI_4 NS_424 0 3.1958050728646652e-03
GC_4_425 b_4 NI_4 NS_425 0 3.8550118525656693e-03
GC_4_426 b_4 NI_4 NS_426 0 -2.9522342675832067e-03
GC_4_427 b_4 NI_4 NS_427 0 -2.0071644384038081e-03
GC_4_428 b_4 NI_4 NS_428 0 -4.1861153496894803e-03
GC_4_429 b_4 NI_4 NS_429 0 -3.5104564331089996e-04
GC_4_430 b_4 NI_4 NS_430 0 2.2864791444765081e-03
GC_4_431 b_4 NI_4 NS_431 0 -1.0763134239618780e-05
GC_4_432 b_4 NI_4 NS_432 0 -2.3358060973643380e-05
GC_4_433 b_4 NI_4 NS_433 0 8.7769866723201042e-04
GC_4_434 b_4 NI_4 NS_434 0 -3.8352026116451349e-03
GC_4_435 b_4 NI_4 NS_435 0 3.5234563945573522e-04
GC_4_436 b_4 NI_4 NS_436 0 3.3067902032346917e-03
GC_4_437 b_4 NI_4 NS_437 0 1.3988544772376155e-03
GC_4_438 b_4 NI_4 NS_438 0 -2.3422177471417826e-03
GC_4_439 b_4 NI_4 NS_439 0 2.2595445985122181e-03
GC_4_440 b_4 NI_4 NS_440 0 3.3689528580423912e-03
GC_4_441 b_4 NI_4 NS_441 0 1.1614257540540143e-03
GC_4_442 b_4 NI_4 NS_442 0 2.4048218341710327e-03
GC_4_443 b_4 NI_4 NS_443 0 -8.2758873323613466e-04
GC_4_444 b_4 NI_4 NS_444 0 -1.9684501755093463e-03
GC_4_445 b_4 NI_4 NS_445 0 3.9844979260024628e-04
GC_4_446 b_4 NI_4 NS_446 0 -2.6910253245426997e-03
GC_4_447 b_4 NI_4 NS_447 0 9.7822596634266896e-04
GC_4_448 b_4 NI_4 NS_448 0 2.7413579780174403e-03
GC_4_449 b_4 NI_4 NS_449 0 1.0427092325713525e-03
GC_4_450 b_4 NI_4 NS_450 0 -2.4233094973751769e-03
GC_4_451 b_4 NI_4 NS_451 0 -1.0796403751135587e-03
GC_4_452 b_4 NI_4 NS_452 0 1.5897875189545907e-03
GC_4_453 b_4 NI_4 NS_453 0 -1.0824816241032422e-08
GC_4_454 b_4 NI_4 NS_454 0 -2.6618453096153849e-09
GC_4_455 b_4 NI_4 NS_455 0 2.3026497631558820e-06
GC_4_456 b_4 NI_4 NS_456 0 5.5056417255584358e-07
GC_4_457 b_4 NI_4 NS_457 0 -2.0458591472770791e-04
GC_4_458 b_4 NI_4 NS_458 0 -3.3255723314227729e-06
GC_4_459 b_4 NI_4 NS_459 0 1.2945373296333518e-09
GC_4_460 b_4 NI_4 NS_460 0 9.6769651223358899e-09
GC_4_461 b_4 NI_4 NS_461 0 -4.2458955218704479e-06
GC_4_462 b_4 NI_4 NS_462 0 6.2176604615697366e-06
GC_4_463 b_4 NI_4 NS_463 0 3.7003830119254581e-06
GC_4_464 b_4 NI_4 NS_464 0 -8.0289206456372794e-06
GC_4_465 b_4 NI_4 NS_465 0 2.1715338386104325e-05
GC_4_466 b_4 NI_4 NS_466 0 -8.4141862167397950e-06
GC_4_467 b_4 NI_4 NS_467 0 -2.1191980992048462e-05
GC_4_468 b_4 NI_4 NS_468 0 -1.1902108641894125e-06
GC_4_469 b_4 NI_4 NS_469 0 -2.9306370753850560e-05
GC_4_470 b_4 NI_4 NS_470 0 -2.8028717298386971e-05
GC_4_471 b_4 NI_4 NS_471 0 -4.8383588282610380e-06
GC_4_472 b_4 NI_4 NS_472 0 1.6178947812564982e-05
GC_4_473 b_4 NI_4 NS_473 0 -2.6738470529676730e-06
GC_4_474 b_4 NI_4 NS_474 0 -7.1112454190006839e-06
GC_4_475 b_4 NI_4 NS_475 0 -2.2526886440091852e-05
GC_4_476 b_4 NI_4 NS_476 0 5.7341866404320799e-06
GC_4_477 b_4 NI_4 NS_477 0 -1.8493943438930389e-04
GC_4_478 b_4 NI_4 NS_478 0 -4.4593170405377930e-05
GC_4_479 b_4 NI_4 NS_479 0 6.1949175997233754e-05
GC_4_480 b_4 NI_4 NS_480 0 1.3746856892815675e-04
GC_4_481 b_4 NI_4 NS_481 0 -3.7405897393990076e-05
GC_4_482 b_4 NI_4 NS_482 0 5.6303428532306340e-05
GC_4_483 b_4 NI_4 NS_483 0 9.4942303176110126e-05
GC_4_484 b_4 NI_4 NS_484 0 2.4590671208778105e-04
GC_4_485 b_4 NI_4 NS_485 0 7.3705223314888066e-05
GC_4_486 b_4 NI_4 NS_486 0 8.1377042767024259e-07
GC_4_487 b_4 NI_4 NS_487 0 -1.6021257958682763e-05
GC_4_488 b_4 NI_4 NS_488 0 2.6079714620377202e-04
GC_4_489 b_4 NI_4 NS_489 0 3.6483924718044765e-04
GC_4_490 b_4 NI_4 NS_490 0 -2.4267031858268769e-04
GC_4_491 b_4 NI_4 NS_491 0 6.5700690230414895e-05
GC_4_492 b_4 NI_4 NS_492 0 -2.8179948767616658e-05
GC_4_493 b_4 NI_4 NS_493 0 2.0799814204179926e-04
GC_4_494 b_4 NI_4 NS_494 0 -2.4118642815367818e-04
GC_4_495 b_4 NI_4 NS_495 0 -7.1054869040351564e-05
GC_4_496 b_4 NI_4 NS_496 0 -7.1872563714538623e-05
GC_4_497 b_4 NI_4 NS_497 0 6.4713639143108395e-05
GC_4_498 b_4 NI_4 NS_498 0 -7.5159632896137926e-05
GC_4_499 b_4 NI_4 NS_499 0 -1.7059832057214085e-04
GC_4_500 b_4 NI_4 NS_500 0 -1.8330408511182521e-04
GC_4_501 b_4 NI_4 NS_501 0 -4.8748184601824110e-05
GC_4_502 b_4 NI_4 NS_502 0 -1.9418952075242445e-05
GC_4_503 b_4 NI_4 NS_503 0 -1.4455356405647531e-04
GC_4_504 b_4 NI_4 NS_504 0 -9.5394431315477232e-05
GC_4_505 b_4 NI_4 NS_505 0 -2.7691635115826379e-05
GC_4_506 b_4 NI_4 NS_506 0 1.0379604806462821e-04
GC_4_507 b_4 NI_4 NS_507 0 -2.7256719549130272e-05
GC_4_508 b_4 NI_4 NS_508 0 1.3718670227618913e-05
GC_4_509 b_4 NI_4 NS_509 0 2.3523443899503738e-06
GC_4_510 b_4 NI_4 NS_510 0 5.0801561014577740e-05
GC_4_511 b_4 NI_4 NS_511 0 1.6821088061256221e-05
GC_4_512 b_4 NI_4 NS_512 0 -4.6980982300756002e-07
GC_4_513 b_4 NI_4 NS_513 0 1.7928537740529239e-06
GC_4_514 b_4 NI_4 NS_514 0 -1.5479233413909978e-05
GC_4_515 b_4 NI_4 NS_515 0 -1.4962773486692858e-05
GC_4_516 b_4 NI_4 NS_516 0 -1.3717819588692884e-05
GC_4_517 b_4 NI_4 NS_517 0 -1.2980733344442180e-05
GC_4_518 b_4 NI_4 NS_518 0 1.2292196880129233e-05
GC_4_519 b_4 NI_4 NS_519 0 7.7931177221999960e-06
GC_4_520 b_4 NI_4 NS_520 0 1.2794667955248025e-06
GC_4_521 b_4 NI_4 NS_521 0 -5.1332449398262119e-06
GC_4_522 b_4 NI_4 NS_522 0 -1.2738562034702455e-05
GC_4_523 b_4 NI_4 NS_523 0 -2.0684794265683525e-05
GC_4_524 b_4 NI_4 NS_524 0 -5.9665478141428838e-06
GC_4_525 b_4 NI_4 NS_525 0 1.1819038400906785e-06
GC_4_526 b_4 NI_4 NS_526 0 2.1730412818427216e-05
GC_4_527 b_4 NI_4 NS_527 0 1.2900857903941631e-05
GC_4_528 b_4 NI_4 NS_528 0 -6.8760465744730091e-06
GC_4_529 b_4 NI_4 NS_529 0 -1.7239530201706113e-05
GC_4_530 b_4 NI_4 NS_530 0 -1.6085702646261059e-05
GC_4_531 b_4 NI_4 NS_531 0 -2.7001165648797455e-05
GC_4_532 b_4 NI_4 NS_532 0 8.7823009689225932e-06
GC_4_533 b_4 NI_4 NS_533 0 2.7182345307095416e-05
GC_4_534 b_4 NI_4 NS_534 0 2.2285116165813935e-05
GC_4_535 b_4 NI_4 NS_535 0 1.1015442660457540e-05
GC_4_536 b_4 NI_4 NS_536 0 -2.1370446555678229e-05
GC_4_537 b_4 NI_4 NS_537 0 -3.0546877213807299e-05
GC_4_538 b_4 NI_4 NS_538 0 3.7167562835979045e-06
GC_4_539 b_4 NI_4 NS_539 0 -9.5362932298721817e-06
GC_4_540 b_4 NI_4 NS_540 0 3.9206795080321890e-05
GC_4_541 b_4 NI_4 NS_541 0 1.8475825447962795e-05
GC_4_542 b_4 NI_4 NS_542 0 -6.8312009718671512e-05
GC_4_543 b_4 NI_4 NS_543 0 4.3335432598292838e-05
GC_4_544 b_4 NI_4 NS_544 0 -1.7301395953052625e-05
GC_4_545 b_4 NI_4 NS_545 0 1.9835697107719915e-07
GC_4_546 b_4 NI_4 NS_546 0 -2.4920222585533091e-07
GC_4_547 b_4 NI_4 NS_547 0 -3.6902239891230522e-06
GC_4_548 b_4 NI_4 NS_548 0 -2.1085270829642796e-05
GC_4_549 b_4 NI_4 NS_549 0 -1.0619039182367857e-05
GC_4_550 b_4 NI_4 NS_550 0 1.6525264320765516e-05
GC_4_551 b_4 NI_4 NS_551 0 9.4041844202546125e-06
GC_4_552 b_4 NI_4 NS_552 0 3.1755349127666627e-05
GC_4_553 b_4 NI_4 NS_553 0 1.4484110242664668e-05
GC_4_554 b_4 NI_4 NS_554 0 -3.2769563664554577e-06
GC_4_555 b_4 NI_4 NS_555 0 -3.8735040775907662e-06
GC_4_556 b_4 NI_4 NS_556 0 1.2514302651492976e-05
GC_4_557 b_4 NI_4 NS_557 0 -1.8541635299062740e-05
GC_4_558 b_4 NI_4 NS_558 0 -3.5705365107980846e-06
GC_4_559 b_4 NI_4 NS_559 0 1.3189367709763700e-05
GC_4_560 b_4 NI_4 NS_560 0 1.3199058488625522e-05
GC_4_561 b_4 NI_4 NS_561 0 7.6290957831478631e-06
GC_4_562 b_4 NI_4 NS_562 0 -2.3004369783225720e-05
GC_4_563 b_4 NI_4 NS_563 0 -3.8544196941285046e-06
GC_4_564 b_4 NI_4 NS_564 0 -1.1714514662797809e-05
GC_4_565 b_4 NI_4 NS_565 0 -8.7383924802803534e-06
GC_4_566 b_4 NI_4 NS_566 0 -2.6219006088798647e-06
GC_4_567 b_4 NI_4 NS_567 0 5.5124513433705473e-10
GC_4_568 b_4 NI_4 NS_568 0 2.9329261987675558e-10
GC_4_569 b_4 NI_4 NS_569 0 4.2110172793532950e-08
GC_4_570 b_4 NI_4 NS_570 0 3.6978460729324487e-08
GC_4_571 b_4 NI_4 NS_571 0 3.0652005968073796e-04
GC_4_572 b_4 NI_4 NS_572 0 -1.4375835996879613e-05
GC_4_573 b_4 NI_4 NS_573 0 -1.2385117507972032e-09
GC_4_574 b_4 NI_4 NS_574 0 -1.9194439934894216e-08
GC_4_575 b_4 NI_4 NS_575 0 3.2004163046321959e-06
GC_4_576 b_4 NI_4 NS_576 0 -3.9681502933824248e-06
GC_4_577 b_4 NI_4 NS_577 0 -1.2573342362072997e-05
GC_4_578 b_4 NI_4 NS_578 0 -1.0250929510825968e-06
GC_4_579 b_4 NI_4 NS_579 0 3.9887653692699220e-05
GC_4_580 b_4 NI_4 NS_580 0 8.6396725134424087e-07
GC_4_581 b_4 NI_4 NS_581 0 -4.2800323124942070e-05
GC_4_582 b_4 NI_4 NS_582 0 -2.4451092134913065e-05
GC_4_583 b_4 NI_4 NS_583 0 1.1877311794386201e-06
GC_4_584 b_4 NI_4 NS_584 0 4.3284248250230208e-05
GC_4_585 b_4 NI_4 NS_585 0 1.0653264399137476e-05
GC_4_586 b_4 NI_4 NS_586 0 -4.8921231973351526e-05
GC_4_587 b_4 NI_4 NS_587 0 2.9254040339454532e-06
GC_4_588 b_4 NI_4 NS_588 0 6.2451616114829999e-06
GC_4_589 b_4 NI_4 NS_589 0 -4.5618512623781188e-05
GC_4_590 b_4 NI_4 NS_590 0 1.8884926620931633e-06
GC_4_591 b_4 NI_4 NS_591 0 1.0003124049204488e-04
GC_4_592 b_4 NI_4 NS_592 0 1.2285660350199053e-04
GC_4_593 b_4 NI_4 NS_593 0 -7.5037289268233126e-05
GC_4_594 b_4 NI_4 NS_594 0 -1.3519238328707199e-04
GC_4_595 b_4 NI_4 NS_595 0 -6.7763285050347741e-05
GC_4_596 b_4 NI_4 NS_596 0 4.9170014005457627e-05
GC_4_597 b_4 NI_4 NS_597 0 1.3378245709167534e-04
GC_4_598 b_4 NI_4 NS_598 0 -2.6374213657412372e-05
GC_4_599 b_4 NI_4 NS_599 0 -8.7278703315866836e-05
GC_4_600 b_4 NI_4 NS_600 0 -1.1628849221655160e-05
GC_4_601 b_4 NI_4 NS_601 0 -9.6762933255369502e-05
GC_4_602 b_4 NI_4 NS_602 0 2.1083572352645507e-04
GC_4_603 b_4 NI_4 NS_603 0 1.6567950462949215e-04
GC_4_604 b_4 NI_4 NS_604 0 -2.1188394296487830e-04
GC_4_605 b_4 NI_4 NS_605 0 -8.1910068534622157e-05
GC_4_606 b_4 NI_4 NS_606 0 1.9157059459026976e-05
GC_4_607 b_4 NI_4 NS_607 0 1.6054321642056043e-04
GC_4_608 b_4 NI_4 NS_608 0 4.4269398809320392e-05
GC_4_609 b_4 NI_4 NS_609 0 -8.8292490995040918e-05
GC_4_610 b_4 NI_4 NS_610 0 -7.2082535867593577e-05
GC_4_611 b_4 NI_4 NS_611 0 -8.5464952864777743e-05
GC_4_612 b_4 NI_4 NS_612 0 6.3489913080792048e-05
GC_4_613 b_4 NI_4 NS_613 0 1.4126679565504817e-04
GC_4_614 b_4 NI_4 NS_614 0 -4.6881954360370984e-05
GC_4_615 b_4 NI_4 NS_615 0 -6.6093588074038297e-05
GC_4_616 b_4 NI_4 NS_616 0 -2.4355716992928692e-05
GC_4_617 b_4 NI_4 NS_617 0 6.0401776679851320e-05
GC_4_618 b_4 NI_4 NS_618 0 1.1474581726381377e-04
GC_4_619 b_4 NI_4 NS_619 0 -2.2017764934415190e-05
GC_4_620 b_4 NI_4 NS_620 0 -1.2142962486917464e-04
GC_4_621 b_4 NI_4 NS_621 0 -4.4471483489060347e-05
GC_4_622 b_4 NI_4 NS_622 0 1.0923655296590391e-05
GC_4_623 b_4 NI_4 NS_623 0 4.7464787844469769e-05
GC_4_624 b_4 NI_4 NS_624 0 -9.9240657347725398e-06
GC_4_625 b_4 NI_4 NS_625 0 -3.2079591982500687e-05
GC_4_626 b_4 NI_4 NS_626 0 -7.5858717092966126e-06
GC_4_627 b_4 NI_4 NS_627 0 2.1298598177296238e-05
GC_4_628 b_4 NI_4 NS_628 0 -4.6121028733237817e-06
GC_4_629 b_4 NI_4 NS_629 0 -3.2316568226321736e-05
GC_4_630 b_4 NI_4 NS_630 0 -2.5188213132706413e-05
GC_4_631 b_4 NI_4 NS_631 0 1.2511323264674511e-05
GC_4_632 b_4 NI_4 NS_632 0 6.5132089106103619e-06
GC_4_633 b_4 NI_4 NS_633 0 -2.0424006424318454e-05
GC_4_634 b_4 NI_4 NS_634 0 -7.6315541499494252e-06
GC_4_635 b_4 NI_4 NS_635 0 1.3991693687400267e-05
GC_4_636 b_4 NI_4 NS_636 0 -1.2277477142741707e-05
GC_4_637 b_4 NI_4 NS_637 0 -4.1514445816092440e-05
GC_4_638 b_4 NI_4 NS_638 0 -1.6952575625048105e-05
GC_4_639 b_4 NI_4 NS_639 0 1.1564369764115243e-05
GC_4_640 b_4 NI_4 NS_640 0 -1.4313411166816337e-06
GC_4_641 b_4 NI_4 NS_641 0 -3.0401004496988376e-05
GC_4_642 b_4 NI_4 NS_642 0 5.6251339487485658e-06
GC_4_643 b_4 NI_4 NS_643 0 1.6016639714145846e-05
GC_4_644 b_4 NI_4 NS_644 0 -2.0571426603865386e-05
GC_4_645 b_4 NI_4 NS_645 0 -5.0239545634890681e-05
GC_4_646 b_4 NI_4 NS_646 0 -1.7714961354527389e-06
GC_4_647 b_4 NI_4 NS_647 0 1.1585346158436572e-05
GC_4_648 b_4 NI_4 NS_648 0 -1.1191608954306456e-05
GC_4_649 b_4 NI_4 NS_649 0 -3.2363535781851795e-05
GC_4_650 b_4 NI_4 NS_650 0 2.5180975813592517e-05
GC_4_651 b_4 NI_4 NS_651 0 1.0237908604543423e-05
GC_4_652 b_4 NI_4 NS_652 0 -3.5896464134055587e-05
GC_4_653 b_4 NI_4 NS_653 0 -3.4868718439033050e-05
GC_4_654 b_4 NI_4 NS_654 0 1.8378562044000126e-05
GC_4_655 b_4 NI_4 NS_655 0 -5.6366148448355959e-05
GC_4_656 b_4 NI_4 NS_656 0 1.3314460596880584e-04
GC_4_657 b_4 NI_4 NS_657 0 -1.5278315911544369e-05
GC_4_658 b_4 NI_4 NS_658 0 -3.1719297796623738e-05
GC_4_659 b_4 NI_4 NS_659 0 -3.7759711785279231e-07
GC_4_660 b_4 NI_4 NS_660 0 3.9613378469568161e-07
GC_4_661 b_4 NI_4 NS_661 0 -2.0157654431045217e-05
GC_4_662 b_4 NI_4 NS_662 0 3.2122139616021145e-05
GC_4_663 b_4 NI_4 NS_663 0 -1.4301666089613292e-05
GC_4_664 b_4 NI_4 NS_664 0 -3.3396350366747805e-05
GC_4_665 b_4 NI_4 NS_665 0 -6.1620326179370968e-06
GC_4_666 b_4 NI_4 NS_666 0 5.1170144575892619e-06
GC_4_667 b_4 NI_4 NS_667 0 -2.1210447289288519e-05
GC_4_668 b_4 NI_4 NS_668 0 -6.5713064797008226e-05
GC_4_669 b_4 NI_4 NS_669 0 -9.1587285651022905e-06
GC_4_670 b_4 NI_4 NS_670 0 -2.0643971571691208e-05
GC_4_671 b_4 NI_4 NS_671 0 1.5020247737296030e-05
GC_4_672 b_4 NI_4 NS_672 0 2.2754098215113454e-05
GC_4_673 b_4 NI_4 NS_673 0 -6.7861253119117845e-06
GC_4_674 b_4 NI_4 NS_674 0 2.7712147630292009e-05
GC_4_675 b_4 NI_4 NS_675 0 -1.1040554557256371e-05
GC_4_676 b_4 NI_4 NS_676 0 -2.1529685281701885e-05
GC_4_677 b_4 NI_4 NS_677 0 -1.1040049265167754e-05
GC_4_678 b_4 NI_4 NS_678 0 2.3841904690487676e-05
GC_4_679 b_4 NI_4 NS_679 0 5.1225221009544806e-06
GC_4_680 b_4 NI_4 NS_680 0 -1.5323216565660304e-05
GC_4_681 b_4 NI_4 NS_681 0 -4.7531894669303598e-10
GC_4_682 b_4 NI_4 NS_682 0 -9.1476657761055976e-10
GC_4_683 b_4 NI_4 NS_683 0 -5.5313561760909804e-08
GC_4_684 b_4 NI_4 NS_684 0 7.4254783386661199e-09
GC_4_685 b_4 NI_4 NS_685 0 -3.2373991072904635e-05
GC_4_686 b_4 NI_4 NS_686 0 2.2170618837827341e-06
GC_4_687 b_4 NI_4 NS_687 0 6.8028468605847583e-11
GC_4_688 b_4 NI_4 NS_688 0 3.0563739730857087e-09
GC_4_689 b_4 NI_4 NS_689 0 -1.7156141091610478e-06
GC_4_690 b_4 NI_4 NS_690 0 -1.8282676158673455e-06
GC_4_691 b_4 NI_4 NS_691 0 -5.3488494019361470e-06
GC_4_692 b_4 NI_4 NS_692 0 2.8545835182358181e-06
GC_4_693 b_4 NI_4 NS_693 0 -1.6536985879604681e-05
GC_4_694 b_4 NI_4 NS_694 0 1.8376724210853743e-05
GC_4_695 b_4 NI_4 NS_695 0 1.5065180464389999e-05
GC_4_696 b_4 NI_4 NS_696 0 9.7699969916961614e-06
GC_4_697 b_4 NI_4 NS_697 0 1.7310034108366761e-05
GC_4_698 b_4 NI_4 NS_698 0 2.2719451594295911e-05
GC_4_699 b_4 NI_4 NS_699 0 2.9106628079298964e-05
GC_4_700 b_4 NI_4 NS_700 0 4.9748813501102743e-06
GC_4_701 b_4 NI_4 NS_701 0 -2.9665369109552615e-06
GC_4_702 b_4 NI_4 NS_702 0 -1.8804681854300972e-06
GC_4_703 b_4 NI_4 NS_703 0 1.6935041474094395e-05
GC_4_704 b_4 NI_4 NS_704 0 -2.2271407151506645e-06
GC_4_705 b_4 NI_4 NS_705 0 1.2887257497306317e-04
GC_4_706 b_4 NI_4 NS_706 0 3.4717432331558045e-05
GC_4_707 b_4 NI_4 NS_707 0 -2.8878617632791557e-05
GC_4_708 b_4 NI_4 NS_708 0 -9.8668099822513006e-05
GC_4_709 b_4 NI_4 NS_709 0 2.4897076613978208e-05
GC_4_710 b_4 NI_4 NS_710 0 -3.1464182294100864e-05
GC_4_711 b_4 NI_4 NS_711 0 -4.1611410450250955e-05
GC_4_712 b_4 NI_4 NS_712 0 -1.6650641586582501e-04
GC_4_713 b_4 NI_4 NS_713 0 -4.1828488044338781e-05
GC_4_714 b_4 NI_4 NS_714 0 -4.8978461407216551e-06
GC_4_715 b_4 NI_4 NS_715 0 2.1414126570013536e-05
GC_4_716 b_4 NI_4 NS_716 0 -1.5190516737800285e-04
GC_4_717 b_4 NI_4 NS_717 0 -2.3047123414800887e-04
GC_4_718 b_4 NI_4 NS_718 0 1.1445044644497317e-04
GC_4_719 b_4 NI_4 NS_719 0 -3.7401825085306030e-05
GC_4_720 b_4 NI_4 NS_720 0 1.4352681834188833e-05
GC_4_721 b_4 NI_4 NS_721 0 -1.3776551048068041e-04
GC_4_722 b_4 NI_4 NS_722 0 1.3054679590277933e-04
GC_4_723 b_4 NI_4 NS_723 0 3.6494591569296241e-05
GC_4_724 b_4 NI_4 NS_724 0 4.1231203617091956e-05
GC_4_725 b_4 NI_4 NS_725 0 -3.8131631695316821e-05
GC_4_726 b_4 NI_4 NS_726 0 4.3361082479102643e-05
GC_4_727 b_4 NI_4 NS_727 0 8.7555850792653137e-05
GC_4_728 b_4 NI_4 NS_728 0 1.1842919561497462e-04
GC_4_729 b_4 NI_4 NS_729 0 2.7361533079711468e-05
GC_4_730 b_4 NI_4 NS_730 0 1.0121201461649028e-05
GC_4_731 b_4 NI_4 NS_731 0 8.7344645905777346e-05
GC_4_732 b_4 NI_4 NS_732 0 6.5655938436806732e-05
GC_4_733 b_4 NI_4 NS_733 0 2.0321375862287634e-05
GC_4_734 b_4 NI_4 NS_734 0 -5.7038893388222062e-05
GC_4_735 b_4 NI_4 NS_735 0 1.6978947316654539e-05
GC_4_736 b_4 NI_4 NS_736 0 -8.9185286752462233e-06
GC_4_737 b_4 NI_4 NS_737 0 8.5891157564320330e-06
GC_4_738 b_4 NI_4 NS_738 0 -3.2921326440757718e-05
GC_4_739 b_4 NI_4 NS_739 0 -8.8488158740551567e-06
GC_4_740 b_4 NI_4 NS_740 0 5.5965307963155810e-07
GC_4_741 b_4 NI_4 NS_741 0 -2.4314152216385347e-06
GC_4_742 b_4 NI_4 NS_742 0 8.5078369591348443e-06
GC_4_743 b_4 NI_4 NS_743 0 1.0240905620659032e-05
GC_4_744 b_4 NI_4 NS_744 0 6.0554401533370572e-06
GC_4_745 b_4 NI_4 NS_745 0 1.2188371522525288e-05
GC_4_746 b_4 NI_4 NS_746 0 -7.8214835890680922e-06
GC_4_747 b_4 NI_4 NS_747 0 -3.4896278632326202e-06
GC_4_748 b_4 NI_4 NS_748 0 -4.3246306446206885e-07
GC_4_749 b_4 NI_4 NS_749 0 2.4743799971709526e-06
GC_4_750 b_4 NI_4 NS_750 0 7.4083936693578832e-06
GC_4_751 b_4 NI_4 NS_751 0 1.3659373370396462e-05
GC_4_752 b_4 NI_4 NS_752 0 2.6169670027530936e-06
GC_4_753 b_4 NI_4 NS_753 0 4.5330444492744186e-06
GC_4_754 b_4 NI_4 NS_754 0 -1.4186507802005041e-05
GC_4_755 b_4 NI_4 NS_755 0 -5.9288346134383488e-06
GC_4_756 b_4 NI_4 NS_756 0 4.2661556335968899e-06
GC_4_757 b_4 NI_4 NS_757 0 1.0298028898535143e-05
GC_4_758 b_4 NI_4 NS_758 0 9.9363442167763027e-06
GC_4_759 b_4 NI_4 NS_759 0 1.7307568644313812e-05
GC_4_760 b_4 NI_4 NS_760 0 -4.2766864441556385e-06
GC_4_761 b_4 NI_4 NS_761 0 -9.2960013542528496e-06
GC_4_762 b_4 NI_4 NS_762 0 -1.5305387657922788e-05
GC_4_763 b_4 NI_4 NS_763 0 -4.0930045535209053e-06
GC_4_764 b_4 NI_4 NS_764 0 1.3520392245305693e-05
GC_4_765 b_4 NI_4 NS_765 0 2.0923683214338846e-05
GC_4_766 b_4 NI_4 NS_766 0 -5.4865174530504664e-07
GC_4_767 b_4 NI_4 NS_767 0 8.8629121384995132e-06
GC_4_768 b_4 NI_4 NS_768 0 -1.7438354113757084e-05
GC_4_769 b_4 NI_4 NS_769 0 2.5763808082458058e-06
GC_4_770 b_4 NI_4 NS_770 0 -1.3772984227864856e-05
GC_4_771 b_4 NI_4 NS_771 0 -1.3801385743692209e-05
GC_4_772 b_4 NI_4 NS_772 0 4.4170586868531603e-06
GC_4_773 b_4 NI_4 NS_773 0 1.6023551533126320e-08
GC_4_774 b_4 NI_4 NS_774 0 -4.1749362667368751e-08
GC_4_775 b_4 NI_4 NS_775 0 8.6199990019275025e-06
GC_4_776 b_4 NI_4 NS_776 0 1.1611706761408891e-05
GC_4_777 b_4 NI_4 NS_777 0 1.0921434486643149e-05
GC_4_778 b_4 NI_4 NS_778 0 -1.1277738045090187e-05
GC_4_779 b_4 NI_4 NS_779 0 -3.7555126538404599e-06
GC_4_780 b_4 NI_4 NS_780 0 -1.0184191551466088e-05
GC_4_781 b_4 NI_4 NS_781 0 -2.3202515573592923e-06
GC_4_782 b_4 NI_4 NS_782 0 1.2931861128342023e-05
GC_4_783 b_4 NI_4 NS_783 0 9.7593896796000073e-07
GC_4_784 b_4 NI_4 NS_784 0 -7.2834607848314593e-06
GC_4_785 b_4 NI_4 NS_785 0 7.5034060421712681e-06
GC_4_786 b_4 NI_4 NS_786 0 1.6765298929582354e-06
GC_4_787 b_4 NI_4 NS_787 0 -6.0990908760681278e-06
GC_4_788 b_4 NI_4 NS_788 0 -8.8899449060904151e-06
GC_4_789 b_4 NI_4 NS_789 0 -4.1232001850333239e-06
GC_4_790 b_4 NI_4 NS_790 0 9.6572719678201984e-06
GC_4_791 b_4 NI_4 NS_791 0 3.3299194646663430e-06
GC_4_792 b_4 NI_4 NS_792 0 6.0429586326777545e-06
GC_4_793 b_4 NI_4 NS_793 0 5.6621022398168639e-06
GC_4_794 b_4 NI_4 NS_794 0 5.1491837693620433e-07
GC_4_795 b_4 NI_4 NS_795 0 6.1218318204122838e-11
GC_4_796 b_4 NI_4 NS_796 0 1.4945631472771646e-10
GC_4_797 b_4 NI_4 NS_797 0 5.9799313799019125e-09
GC_4_798 b_4 NI_4 NS_798 0 -8.3554293382255850e-09
GC_4_799 b_4 NI_4 NS_799 0 -1.1096947998863547e-04
GC_4_800 b_4 NI_4 NS_800 0 -2.1483029994741108e-06
GC_4_801 b_4 NI_4 NS_801 0 -2.5029527534383814e-10
GC_4_802 b_4 NI_4 NS_802 0 2.6115886770322468e-09
GC_4_803 b_4 NI_4 NS_803 0 1.8723153808792502e-06
GC_4_804 b_4 NI_4 NS_804 0 -1.6074371670395565e-06
GC_4_805 b_4 NI_4 NS_805 0 3.2540214238508757e-07
GC_4_806 b_4 NI_4 NS_806 0 -6.5210481624859249e-06
GC_4_807 b_4 NI_4 NS_807 0 -7.4589937765701950e-06
GC_4_808 b_4 NI_4 NS_808 0 -4.2413692587380962e-07
GC_4_809 b_4 NI_4 NS_809 0 -1.5203211923962569e-06
GC_4_810 b_4 NI_4 NS_810 0 -4.8607527944288847e-06
GC_4_811 b_4 NI_4 NS_811 0 -1.6019419641469411e-05
GC_4_812 b_4 NI_4 NS_812 0 -2.1097788755282922e-06
GC_4_813 b_4 NI_4 NS_813 0 -7.3376620143334952e-06
GC_4_814 b_4 NI_4 NS_814 0 1.8827317385039855e-05
GC_4_815 b_4 NI_4 NS_815 0 4.9694024739769324e-06
GC_4_816 b_4 NI_4 NS_816 0 -2.7979711184245424e-06
GC_4_817 b_4 NI_4 NS_817 0 -2.3130512085197727e-07
GC_4_818 b_4 NI_4 NS_818 0 -2.4916635953630641e-06
GC_4_819 b_4 NI_4 NS_819 0 -2.6811397175482002e-05
GC_4_820 b_4 NI_4 NS_820 0 2.8304979959739748e-05
GC_4_821 b_4 NI_4 NS_821 0 2.8363183182365929e-05
GC_4_822 b_4 NI_4 NS_822 0 -7.9685185135715132e-06
GC_4_823 b_4 NI_4 NS_823 0 -8.2696309608001802e-06
GC_4_824 b_4 NI_4 NS_824 0 -4.3355265098141424e-06
GC_4_825 b_4 NI_4 NS_825 0 1.2216123036083018e-05
GC_4_826 b_4 NI_4 NS_826 0 2.7630082769161013e-05
GC_4_827 b_4 NI_4 NS_827 0 1.4665317849051245e-06
GC_4_828 b_4 NI_4 NS_828 0 -8.9517362999865315e-06
GC_4_829 b_4 NI_4 NS_829 0 -2.8979852545498683e-05
GC_4_830 b_4 NI_4 NS_830 0 4.5865777820464355e-06
GC_4_831 b_4 NI_4 NS_831 0 4.1777950668706927e-05
GC_4_832 b_4 NI_4 NS_832 0 1.1538570147852567e-05
GC_4_833 b_4 NI_4 NS_833 0 -3.0566436279661411e-06
GC_4_834 b_4 NI_4 NS_834 0 -4.4930606227095941e-06
GC_4_835 b_4 NI_4 NS_835 0 1.2853449343391978e-05
GC_4_836 b_4 NI_4 NS_836 0 1.9652908147612365e-05
GC_4_837 b_4 NI_4 NS_837 0 3.9663200204319358e-06
GC_4_838 b_4 NI_4 NS_838 0 -1.0991933378985347e-05
GC_4_839 b_4 NI_4 NS_839 0 -6.6134810425530709e-06
GC_4_840 b_4 NI_4 NS_840 0 8.3132160669319155e-07
GC_4_841 b_4 NI_4 NS_841 0 1.9091620214312028e-05
GC_4_842 b_4 NI_4 NS_842 0 5.9084922482756966e-06
GC_4_843 b_4 NI_4 NS_843 0 -5.2595655330503570e-08
GC_4_844 b_4 NI_4 NS_844 0 -4.2237277357565726e-06
GC_4_845 b_4 NI_4 NS_845 0 4.6917578401714158e-06
GC_4_846 b_4 NI_4 NS_846 0 1.4599971679091221e-05
GC_4_847 b_4 NI_4 NS_847 0 8.0921060501808895e-06
GC_4_848 b_4 NI_4 NS_848 0 -1.1172243885057634e-05
GC_4_849 b_4 NI_4 NS_849 0 -1.4419298979978210e-06
GC_4_850 b_4 NI_4 NS_850 0 9.2581090795056490e-07
GC_4_851 b_4 NI_4 NS_851 0 1.0893573879527675e-05
GC_4_852 b_4 NI_4 NS_852 0 4.3229017808078838e-06
GC_4_853 b_4 NI_4 NS_853 0 1.7169272581788999e-06
GC_4_854 b_4 NI_4 NS_854 0 -6.1401544344739865e-07
GC_4_855 b_4 NI_4 NS_855 0 5.6792608538748751e-06
GC_4_856 b_4 NI_4 NS_856 0 1.7812866317219540e-06
GC_4_857 b_4 NI_4 NS_857 0 3.3801498781542340e-06
GC_4_858 b_4 NI_4 NS_858 0 2.0631600559657637e-06
GC_4_859 b_4 NI_4 NS_859 0 1.0923423723706830e-05
GC_4_860 b_4 NI_4 NS_860 0 3.8982228899389857e-06
GC_4_861 b_4 NI_4 NS_861 0 4.8460148795581398e-06
GC_4_862 b_4 NI_4 NS_862 0 -4.9709750824881996e-08
GC_4_863 b_4 NI_4 NS_863 0 9.9733341343357675e-06
GC_4_864 b_4 NI_4 NS_864 0 -1.0087354401161255e-06
GC_4_865 b_4 NI_4 NS_865 0 8.2004986474436246e-06
GC_4_866 b_4 NI_4 NS_866 0 2.9626422883261190e-06
GC_4_867 b_4 NI_4 NS_867 0 1.9001978534868572e-05
GC_4_868 b_4 NI_4 NS_868 0 -5.4549104315747681e-06
GC_4_869 b_4 NI_4 NS_869 0 7.1770832705838115e-06
GC_4_870 b_4 NI_4 NS_870 0 -3.9934630783014532e-06
GC_4_871 b_4 NI_4 NS_871 0 1.3699651711053511e-05
GC_4_872 b_4 NI_4 NS_872 0 -1.1820624993036959e-05
GC_4_873 b_4 NI_4 NS_873 0 1.2324204826198753e-05
GC_4_874 b_4 NI_4 NS_874 0 -3.9604840079486639e-06
GC_4_875 b_4 NI_4 NS_875 0 9.1123487819147183e-06
GC_4_876 b_4 NI_4 NS_876 0 -2.6652121127434954e-05
GC_4_877 b_4 NI_4 NS_877 0 2.3022874118102274e-06
GC_4_878 b_4 NI_4 NS_878 0 -1.2345511389304781e-05
GC_4_879 b_4 NI_4 NS_879 0 -8.3181276908788775e-06
GC_4_880 b_4 NI_4 NS_880 0 -1.8540253364999637e-05
GC_4_881 b_4 NI_4 NS_881 0 -5.0234188256768768e-06
GC_4_882 b_4 NI_4 NS_882 0 -1.2083006336178865e-05
GC_4_883 b_4 NI_4 NS_883 0 5.5479940736457675e-05
GC_4_884 b_4 NI_4 NS_884 0 -8.7812851065455338e-05
GC_4_885 b_4 NI_4 NS_885 0 -1.0021971097295590e-05
GC_4_886 b_4 NI_4 NS_886 0 1.5204008153785182e-06
GC_4_887 b_4 NI_4 NS_887 0 3.9312423495778983e-07
GC_4_888 b_4 NI_4 NS_888 0 -1.2255152231020714e-07
GC_4_889 b_4 NI_4 NS_889 0 -2.7361002675958044e-06
GC_4_890 b_4 NI_4 NS_890 0 -1.8487251802552486e-06
GC_4_891 b_4 NI_4 NS_891 0 -4.3417375922905614e-06
GC_4_892 b_4 NI_4 NS_892 0 6.4984050247919764e-07
GC_4_893 b_4 NI_4 NS_893 0 -1.7585016188861143e-05
GC_4_894 b_4 NI_4 NS_894 0 9.5836826644337131e-06
GC_4_895 b_4 NI_4 NS_895 0 -9.3307317351278146e-06
GC_4_896 b_4 NI_4 NS_896 0 3.7420412834633494e-05
GC_4_897 b_4 NI_4 NS_897 0 -7.2143700657483774e-06
GC_4_898 b_4 NI_4 NS_898 0 3.1323471495145904e-07
GC_4_899 b_4 NI_4 NS_899 0 -1.3394815734579146e-05
GC_4_900 b_4 NI_4 NS_900 0 1.8225008014360002e-06
GC_4_901 b_4 NI_4 NS_901 0 -4.6183393508244359e-06
GC_4_902 b_4 NI_4 NS_902 0 -3.3980542949431298e-06
GC_4_903 b_4 NI_4 NS_903 0 -6.3783028251204404e-06
GC_4_904 b_4 NI_4 NS_904 0 1.0293199306953365e-06
GC_4_905 b_4 NI_4 NS_905 0 -3.0260508508823639e-06
GC_4_906 b_4 NI_4 NS_906 0 8.8999088917734460e-07
GC_4_907 b_4 NI_4 NS_907 0 -1.7736247285231777e-06
GC_4_908 b_4 NI_4 NS_908 0 -9.4941202370394659e-07
GC_4_909 b_4 NI_4 NS_909 0 -2.6169661828841579e-10
GC_4_910 b_4 NI_4 NS_910 0 4.2344984006929910e-10
GC_4_911 b_4 NI_4 NS_911 0 2.2765333610106107e-09
GC_4_912 b_4 NI_4 NS_912 0 -2.6875808605142708e-08
GC_4_913 b_4 NI_4 NS_913 0 -2.1854767172194974e-05
GC_4_914 b_4 NI_4 NS_914 0 2.4289816459749788e-07
GC_4_915 b_4 NI_4 NS_915 0 1.6216332230405142e-11
GC_4_916 b_4 NI_4 NS_916 0 -4.8482477456823267e-10
GC_4_917 b_4 NI_4 NS_917 0 3.7393775930325076e-07
GC_4_918 b_4 NI_4 NS_918 0 -1.3861912788052821e-06
GC_4_919 b_4 NI_4 NS_919 0 -1.4298846730688166e-07
GC_4_920 b_4 NI_4 NS_920 0 1.1185392352529650e-06
GC_4_921 b_4 NI_4 NS_921 0 -3.5074127154698209e-06
GC_4_922 b_4 NI_4 NS_922 0 -2.2370218340146195e-06
GC_4_923 b_4 NI_4 NS_923 0 -7.4943554678609195e-07
GC_4_924 b_4 NI_4 NS_924 0 -1.1227673776974020e-06
GC_4_925 b_4 NI_4 NS_925 0 -6.8343235483576978e-07
GC_4_926 b_4 NI_4 NS_926 0 2.6595603090851351e-06
GC_4_927 b_4 NI_4 NS_927 0 -5.0813980439902281e-06
GC_4_928 b_4 NI_4 NS_928 0 3.8742750566182634e-06
GC_4_929 b_4 NI_4 NS_929 0 9.5053017798168189e-07
GC_4_930 b_4 NI_4 NS_930 0 -1.5553106590297967e-07
GC_4_931 b_4 NI_4 NS_931 0 -2.6358677567121855e-07
GC_4_932 b_4 NI_4 NS_932 0 -5.2938841053474541e-07
GC_4_933 b_4 NI_4 NS_933 0 -1.4742657638429253e-06
GC_4_934 b_4 NI_4 NS_934 0 1.1166382189638936e-05
GC_4_935 b_4 NI_4 NS_935 0 5.7536116397122343e-06
GC_4_936 b_4 NI_4 NS_936 0 2.9700779194704775e-06
GC_4_937 b_4 NI_4 NS_937 0 7.6103126287408485e-07
GC_4_938 b_4 NI_4 NS_938 0 -4.0059626853495312e-07
GC_4_939 b_4 NI_4 NS_939 0 1.7105181073334207e-05
GC_4_940 b_4 NI_4 NS_940 0 -2.9782855486281345e-07
GC_4_941 b_4 NI_4 NS_941 0 7.0007413537231753e-07
GC_4_942 b_4 NI_4 NS_942 0 1.7703040411275750e-07
GC_4_943 b_4 NI_4 NS_943 0 6.4126716900091920e-06
GC_4_944 b_4 NI_4 NS_944 0 -4.4402806930105708e-07
GC_4_945 b_4 NI_4 NS_945 0 -8.2381908705341755e-07
GC_4_946 b_4 NI_4 NS_946 0 -1.7747643070895794e-05
GC_4_947 b_4 NI_4 NS_947 0 -2.8347586617026986e-07
GC_4_948 b_4 NI_4 NS_948 0 2.3003557029879567e-07
GC_4_949 b_4 NI_4 NS_949 0 -1.0769402728137246e-05
GC_4_950 b_4 NI_4 NS_950 0 -9.4805211249177230e-06
GC_4_951 b_4 NI_4 NS_951 0 -1.3423577506100233e-06
GC_4_952 b_4 NI_4 NS_952 0 -8.1223759872771400e-07
GC_4_953 b_4 NI_4 NS_953 0 -1.6041434634542301e-06
GC_4_954 b_4 NI_4 NS_954 0 4.5694567055229850e-07
GC_4_955 b_4 NI_4 NS_955 0 -9.3337978055074404e-06
GC_4_956 b_4 NI_4 NS_956 0 6.4384894147404959e-06
GC_4_957 b_4 NI_4 NS_957 0 6.7351370458432691e-08
GC_4_958 b_4 NI_4 NS_958 0 -3.9969578173484985e-07
GC_4_959 b_4 NI_4 NS_959 0 -7.1799745178599831e-07
GC_4_960 b_4 NI_4 NS_960 0 7.2325982005443138e-06
GC_4_961 b_4 NI_4 NS_961 0 2.0739498174393436e-06
GC_4_962 b_4 NI_4 NS_962 0 2.4611628766514453e-06
GC_4_963 b_4 NI_4 NS_963 0 6.1968367427695239e-07
GC_4_964 b_4 NI_4 NS_964 0 -2.5247692690298510e-07
GC_4_965 b_4 NI_4 NS_965 0 4.6128184160872715e-06
GC_4_966 b_4 NI_4 NS_966 0 3.3398294150878946e-07
GC_4_967 b_4 NI_4 NS_967 0 1.7628451888920533e-07
GC_4_968 b_4 NI_4 NS_968 0 5.3873509046987961e-07
GC_4_969 b_4 NI_4 NS_969 0 -7.4074208245587423e-07
GC_4_970 b_4 NI_4 NS_970 0 -4.2044547435599453e-08
GC_4_971 b_4 NI_4 NS_971 0 7.4597929506847012e-07
GC_4_972 b_4 NI_4 NS_972 0 -5.2039377330471755e-07
GC_4_973 b_4 NI_4 NS_973 0 1.8298787725929494e-06
GC_4_974 b_4 NI_4 NS_974 0 4.7566212180873274e-07
GC_4_975 b_4 NI_4 NS_975 0 1.7708201016725741e-07
GC_4_976 b_4 NI_4 NS_976 0 4.5205125323859083e-07
GC_4_977 b_4 NI_4 NS_977 0 -4.4618844941618460e-07
GC_4_978 b_4 NI_4 NS_978 0 2.3604775227973096e-07
GC_4_979 b_4 NI_4 NS_979 0 6.4977383034298413e-07
GC_4_980 b_4 NI_4 NS_980 0 -3.4554335979702546e-07
GC_4_981 b_4 NI_4 NS_981 0 1.8733452338606092e-06
GC_4_982 b_4 NI_4 NS_982 0 -2.9393847929439938e-08
GC_4_983 b_4 NI_4 NS_983 0 2.9827015766943346e-07
GC_4_984 b_4 NI_4 NS_984 0 5.0985735925117628e-07
GC_4_985 b_4 NI_4 NS_985 0 -3.1520321551798122e-07
GC_4_986 b_4 NI_4 NS_986 0 4.5596753583975247e-07
GC_4_987 b_4 NI_4 NS_987 0 5.5349955998593382e-07
GC_4_988 b_4 NI_4 NS_988 0 -4.4726733255932155e-08
GC_4_989 b_4 NI_4 NS_989 0 1.9808632497757551e-06
GC_4_990 b_4 NI_4 NS_990 0 -4.0113966041143841e-07
GC_4_991 b_4 NI_4 NS_991 0 4.1702659532878273e-07
GC_4_992 b_4 NI_4 NS_992 0 7.7175591712430932e-07
GC_4_993 b_4 NI_4 NS_993 0 5.0614553585015396e-07
GC_4_994 b_4 NI_4 NS_994 0 7.2776774131763674e-07
GC_4_995 b_4 NI_4 NS_995 0 9.0283036718147660e-07
GC_4_996 b_4 NI_4 NS_996 0 9.8988163168824922e-07
GC_4_997 b_4 NI_4 NS_997 0 1.6386468331098094e-06
GC_4_998 b_4 NI_4 NS_998 0 -9.9921089482154668e-06
GC_4_999 b_4 NI_4 NS_999 0 2.8725374011669274e-06
GC_4_1000 b_4 NI_4 NS_1000 0 -1.2252033651352955e-06
GC_4_1001 b_4 NI_4 NS_1001 0 3.1669806614815572e-08
GC_4_1002 b_4 NI_4 NS_1002 0 -4.6445308824083604e-08
GC_4_1003 b_4 NI_4 NS_1003 0 1.4054939829729767e-06
GC_4_1004 b_4 NI_4 NS_1004 0 1.6971691651276979e-07
GC_4_1005 b_4 NI_4 NS_1005 0 9.7902016590363323e-07
GC_4_1006 b_4 NI_4 NS_1006 0 -4.9521388351017388e-07
GC_4_1007 b_4 NI_4 NS_1007 0 6.9358534173974595e-07
GC_4_1008 b_4 NI_4 NS_1008 0 1.3039571994991967e-06
GC_4_1009 b_4 NI_4 NS_1009 0 1.3369614011280808e-06
GC_4_1010 b_4 NI_4 NS_1010 0 1.9875861961340982e-06
GC_4_1011 b_4 NI_4 NS_1011 0 -9.2424559965123485e-08
GC_4_1012 b_4 NI_4 NS_1012 0 -2.7737045504929095e-08
GC_4_1013 b_4 NI_4 NS_1013 0 -5.3471519390956546e-07
GC_4_1014 b_4 NI_4 NS_1014 0 1.8250407830955292e-07
GC_4_1015 b_4 NI_4 NS_1015 0 3.1922710460514613e-07
GC_4_1016 b_4 NI_4 NS_1016 0 -3.6120216504117670e-07
GC_4_1017 b_4 NI_4 NS_1017 0 1.1468241244892509e-08
GC_4_1018 b_4 NI_4 NS_1018 0 -6.0659715012515068e-07
GC_4_1019 b_4 NI_4 NS_1019 0 5.2308415641760929e-08
GC_4_1020 b_4 NI_4 NS_1020 0 1.0683060259231827e-07
GC_4_1021 b_4 NI_4 NS_1021 0 2.9594357765409567e-07
GC_4_1022 b_4 NI_4 NS_1022 0 -1.4209554253537407e-09
GC_4_1023 b_4 NI_4 NS_1023 0 -2.9859354991135366e-12
GC_4_1024 b_4 NI_4 NS_1024 0 -1.0058312362903942e-11
GC_4_1025 b_4 NI_4 NS_1025 0 9.3178043776951157e-10
GC_4_1026 b_4 NI_4 NS_1026 0 3.3553872894577571e-09
GC_4_1027 b_4 NI_4 NS_1027 0 4.4178785319363510e-05
GC_4_1028 b_4 NI_4 NS_1028 0 -2.5097414830611203e-07
GC_4_1029 b_4 NI_4 NS_1029 0 -1.3616414611152599e-11
GC_4_1030 b_4 NI_4 NS_1030 0 3.6731315089110825e-10
GC_4_1031 b_4 NI_4 NS_1031 0 9.4989296719706942e-07
GC_4_1032 b_4 NI_4 NS_1032 0 -2.0375961263284038e-07
GC_4_1033 b_4 NI_4 NS_1033 0 1.1052397143613937e-06
GC_4_1034 b_4 NI_4 NS_1034 0 -6.5609253799507365e-07
GC_4_1035 b_4 NI_4 NS_1035 0 1.6285599716196344e-06
GC_4_1036 b_4 NI_4 NS_1036 0 -3.6726495688526768e-06
GC_4_1037 b_4 NI_4 NS_1037 0 -2.3668556541845549e-06
GC_4_1038 b_4 NI_4 NS_1038 0 -1.3304942517987226e-06
GC_4_1039 b_4 NI_4 NS_1039 0 -2.0337087226444095e-07
GC_4_1040 b_4 NI_4 NS_1040 0 -2.4446335426407611e-06
GC_4_1041 b_4 NI_4 NS_1041 0 -7.1160020081714316e-06
GC_4_1042 b_4 NI_4 NS_1042 0 -2.8108035938938544e-06
GC_4_1043 b_4 NI_4 NS_1043 0 1.7245506138685559e-06
GC_4_1044 b_4 NI_4 NS_1044 0 1.3116943226209031e-06
GC_4_1045 b_4 NI_4 NS_1045 0 -1.6513642825738437e-06
GC_4_1046 b_4 NI_4 NS_1046 0 9.9670711616958754e-07
GC_4_1047 b_4 NI_4 NS_1047 0 -2.8708731157829446e-06
GC_4_1048 b_4 NI_4 NS_1048 0 -1.6219533090785700e-06
GC_4_1049 b_4 NI_4 NS_1049 0 -2.0401471303158766e-06
GC_4_1050 b_4 NI_4 NS_1050 0 2.9684645514153721e-06
GC_4_1051 b_4 NI_4 NS_1051 0 -1.1731543824776094e-06
GC_4_1052 b_4 NI_4 NS_1052 0 1.1051536084384857e-06
GC_4_1053 b_4 NI_4 NS_1053 0 -2.0979525889962789e-06
GC_4_1054 b_4 NI_4 NS_1054 0 1.5287389846010870e-06
GC_4_1055 b_4 NI_4 NS_1055 0 -9.4304098054933286e-07
GC_4_1056 b_4 NI_4 NS_1056 0 1.4308247192055752e-06
GC_4_1057 b_4 NI_4 NS_1057 0 -1.4825500403294639e-06
GC_4_1058 b_4 NI_4 NS_1058 0 1.7944073437166627e-06
GC_4_1059 b_4 NI_4 NS_1059 0 2.5486696308179273e-07
GC_4_1060 b_4 NI_4 NS_1060 0 1.3614197700271948e-06
GC_4_1061 b_4 NI_4 NS_1061 0 -8.4242882476324215e-07
GC_4_1062 b_4 NI_4 NS_1062 0 1.3601202987463379e-06
GC_4_1063 b_4 NI_4 NS_1063 0 9.0836422971755285e-07
GC_4_1064 b_4 NI_4 NS_1064 0 1.8505879666381964e-06
GC_4_1065 b_4 NI_4 NS_1065 0 -7.6710000019533483e-07
GC_4_1066 b_4 NI_4 NS_1066 0 5.7089372560201280e-07
GC_4_1067 b_4 NI_4 NS_1067 0 -8.0358978753517408e-07
GC_4_1068 b_4 NI_4 NS_1068 0 1.5919658742721013e-06
GC_4_1069 b_4 NI_4 NS_1069 0 1.2780290906950902e-06
GC_4_1070 b_4 NI_4 NS_1070 0 5.6829643318520355e-07
GC_4_1071 b_4 NI_4 NS_1071 0 -6.6681055451127382e-07
GC_4_1072 b_4 NI_4 NS_1072 0 6.5600765806854083e-07
GC_4_1073 b_4 NI_4 NS_1073 0 5.3995055796842147e-07
GC_4_1074 b_4 NI_4 NS_1074 0 1.7897672046569296e-06
GC_4_1075 b_4 NI_4 NS_1075 0 -2.5637126677758715e-07
GC_4_1076 b_4 NI_4 NS_1076 0 -3.2549822731339401e-07
GC_4_1077 b_4 NI_4 NS_1077 0 -4.7493597711810636e-07
GC_4_1078 b_4 NI_4 NS_1078 0 6.1075915571438494e-07
GC_4_1079 b_4 NI_4 NS_1079 0 1.1438101830125642e-07
GC_4_1080 b_4 NI_4 NS_1080 0 5.8917183925621722e-07
GC_4_1081 b_4 NI_4 NS_1081 0 -3.1820582687804535e-07
GC_4_1082 b_4 NI_4 NS_1082 0 4.4619737764385523e-07
GC_4_1083 b_4 NI_4 NS_1083 0 6.3948195412325663e-08
GC_4_1084 b_4 NI_4 NS_1084 0 2.2648971896906077e-07
GC_4_1085 b_4 NI_4 NS_1085 0 -6.7255786358114895e-07
GC_4_1086 b_4 NI_4 NS_1086 0 2.4745742678073282e-07
GC_4_1087 b_4 NI_4 NS_1087 0 -1.6417396177053559e-07
GC_4_1088 b_4 NI_4 NS_1088 0 5.7608783772825818e-07
GC_4_1089 b_4 NI_4 NS_1089 0 -3.0458978009299225e-07
GC_4_1090 b_4 NI_4 NS_1090 0 2.5970624013898906e-07
GC_4_1091 b_4 NI_4 NS_1091 0 -9.8777028377088580e-08
GC_4_1092 b_4 NI_4 NS_1092 0 2.0871092020471727e-07
GC_4_1093 b_4 NI_4 NS_1093 0 -7.6626077401363075e-07
GC_4_1094 b_4 NI_4 NS_1094 0 5.3649997144231695e-08
GC_4_1095 b_4 NI_4 NS_1095 0 -4.8041816276640739e-07
GC_4_1096 b_4 NI_4 NS_1096 0 4.3220651514365625e-07
GC_4_1097 b_4 NI_4 NS_1097 0 -5.3154407773876925e-07
GC_4_1098 b_4 NI_4 NS_1098 0 2.1428843814128255e-07
GC_4_1099 b_4 NI_4 NS_1099 0 -5.2281320811898626e-07
GC_4_1100 b_4 NI_4 NS_1100 0 1.4456671131073188e-07
GC_4_1101 b_4 NI_4 NS_1101 0 -1.0034207702785726e-06
GC_4_1102 b_4 NI_4 NS_1102 0 -3.4734760508778675e-07
GC_4_1103 b_4 NI_4 NS_1103 0 -1.4398171806024672e-06
GC_4_1104 b_4 NI_4 NS_1104 0 5.4841464159536037e-07
GC_4_1105 b_4 NI_4 NS_1105 0 -1.1944227485263642e-06
GC_4_1106 b_4 NI_4 NS_1106 0 1.3611361530697586e-07
GC_4_1107 b_4 NI_4 NS_1107 0 -1.4807009808724838e-06
GC_4_1108 b_4 NI_4 NS_1108 0 7.7907310722265663e-07
GC_4_1109 b_4 NI_4 NS_1109 0 -2.2610242949178185e-06
GC_4_1110 b_4 NI_4 NS_1110 0 -8.4610008406233625e-07
GC_4_1111 b_4 NI_4 NS_1111 0 5.6641170744137498e-06
GC_4_1112 b_4 NI_4 NS_1112 0 1.1197530495996505e-05
GC_4_1113 b_4 NI_4 NS_1113 0 -2.2220234365069335e-06
GC_4_1114 b_4 NI_4 NS_1114 0 3.0965161028558778e-06
GC_4_1115 b_4 NI_4 NS_1115 0 1.1650784867846797e-08
GC_4_1116 b_4 NI_4 NS_1116 0 7.3480619387371595e-08
GC_4_1117 b_4 NI_4 NS_1117 0 -1.2474042613815890e-06
GC_4_1118 b_4 NI_4 NS_1118 0 1.6458700162005787e-06
GC_4_1119 b_4 NI_4 NS_1119 0 -6.3374293559483107e-07
GC_4_1120 b_4 NI_4 NS_1120 0 1.4521163460053209e-06
GC_4_1121 b_4 NI_4 NS_1121 0 -1.6480279988565471e-06
GC_4_1122 b_4 NI_4 NS_1122 0 -1.2214488488035870e-06
GC_4_1123 b_4 NI_4 NS_1123 0 -3.3896209506688423e-06
GC_4_1124 b_4 NI_4 NS_1124 0 -1.1084108115461467e-06
GC_4_1125 b_4 NI_4 NS_1125 0 7.2036994282885228e-09
GC_4_1126 b_4 NI_4 NS_1126 0 -1.2022175787940064e-07
GC_4_1127 b_4 NI_4 NS_1127 0 6.2010494287458527e-07
GC_4_1128 b_4 NI_4 NS_1128 0 -3.6782660756879428e-07
GC_4_1129 b_4 NI_4 NS_1129 0 -4.6878158756754556e-08
GC_4_1130 b_4 NI_4 NS_1130 0 3.9701406284898583e-07
GC_4_1131 b_4 NI_4 NS_1131 0 -5.1628328869895091e-08
GC_4_1132 b_4 NI_4 NS_1132 0 2.9624337049415743e-08
GC_4_1133 b_4 NI_4 NS_1133 0 -2.7362451388276175e-07
GC_4_1134 b_4 NI_4 NS_1134 0 1.7742806421023076e-07
GC_4_1135 b_4 NI_4 NS_1135 0 -2.2776110967290941e-07
GC_4_1136 b_4 NI_4 NS_1136 0 -6.5474361094548811e-09
GC_4_1137 b_4 NI_4 NS_1137 0 -8.0171083585737576e-12
GC_4_1138 b_4 NI_4 NS_1138 0 -8.1359707567498990e-13
GC_4_1139 b_4 NI_4 NS_1139 0 -1.1403175234596856e-09
GC_4_1140 b_4 NI_4 NS_1140 0 -2.4260034849702747e-09
GC_4_1141 b_4 NI_4 NS_1141 0 -2.7457175464435992e-05
GC_4_1142 b_4 NI_4 NS_1142 0 -1.0861375771367200e-08
GC_4_1143 b_4 NI_4 NS_1143 0 1.0271926140365442e-11
GC_4_1144 b_4 NI_4 NS_1144 0 -5.9963601959515355e-11
GC_4_1145 b_4 NI_4 NS_1145 0 -6.3440476376443139e-07
GC_4_1146 b_4 NI_4 NS_1146 0 -1.0701543353309948e-06
GC_4_1147 b_4 NI_4 NS_1147 0 -1.4351549063062625e-06
GC_4_1148 b_4 NI_4 NS_1148 0 2.3181028914989654e-06
GC_4_1149 b_4 NI_4 NS_1149 0 -3.8038707942717894e-06
GC_4_1150 b_4 NI_4 NS_1150 0 2.1755687271627198e-06
GC_4_1151 b_4 NI_4 NS_1151 0 1.9264784142359761e-06
GC_4_1152 b_4 NI_4 NS_1152 0 -2.2570743537627696e-07
GC_4_1153 b_4 NI_4 NS_1153 0 1.3997880312287504e-06
GC_4_1154 b_4 NI_4 NS_1154 0 5.7146742627488937e-06
GC_4_1155 b_4 NI_4 NS_1155 0 3.7149863121614444e-06
GC_4_1156 b_4 NI_4 NS_1156 0 3.2450442881607486e-06
GC_4_1157 b_4 NI_4 NS_1157 0 -1.4756138943720208e-06
GC_4_1158 b_4 NI_4 NS_1158 0 -9.4893910359218000e-07
GC_4_1159 b_4 NI_4 NS_1159 0 9.7600713067270137e-07
GC_4_1160 b_4 NI_4 NS_1160 0 -2.1770041907657972e-06
GC_4_1161 b_4 NI_4 NS_1161 0 6.4144828046077131e-06
GC_4_1162 b_4 NI_4 NS_1162 0 8.5313663137224008e-06
GC_4_1163 b_4 NI_4 NS_1163 0 1.3417301130663200e-06
GC_4_1164 b_4 NI_4 NS_1164 0 -9.5630037099100136e-07
GC_4_1165 b_4 NI_4 NS_1165 0 1.0785532001603222e-06
GC_4_1166 b_4 NI_4 NS_1166 0 -1.8906611050305794e-06
GC_4_1167 b_4 NI_4 NS_1167 0 1.4514873974180180e-05
GC_4_1168 b_4 NI_4 NS_1168 0 -4.1895957960225396e-06
GC_4_1169 b_4 NI_4 NS_1169 0 -2.0074949579278781e-07
GC_4_1170 b_4 NI_4 NS_1170 0 6.6361973388081865e-07
GC_4_1171 b_4 NI_4 NS_1171 0 4.9434215247234649e-06
GC_4_1172 b_4 NI_4 NS_1172 0 -2.1798278523027610e-06
GC_4_1173 b_4 NI_4 NS_1173 0 -7.7225940148000669e-07
GC_4_1174 b_4 NI_4 NS_1174 0 -1.5002472206118730e-05
GC_4_1175 b_4 NI_4 NS_1175 0 -7.8154900668258182e-08
GC_4_1176 b_4 NI_4 NS_1176 0 9.5811138250109684e-07
GC_4_1177 b_4 NI_4 NS_1177 0 -7.9220417371282762e-06
GC_4_1178 b_4 NI_4 NS_1178 0 -8.5842556791360911e-06
GC_4_1179 b_4 NI_4 NS_1179 0 -6.3253181905726959e-07
GC_4_1180 b_4 NI_4 NS_1180 0 -2.1422164227371373e-06
GC_4_1181 b_4 NI_4 NS_1181 0 -1.4548574893253164e-08
GC_4_1182 b_4 NI_4 NS_1182 0 1.1898769909048904e-06
GC_4_1183 b_4 NI_4 NS_1183 0 -7.7140637643857861e-06
GC_4_1184 b_4 NI_4 NS_1184 0 1.9652432885611870e-06
GC_4_1185 b_4 NI_4 NS_1185 0 2.3903573004148092e-07
GC_4_1186 b_4 NI_4 NS_1186 0 -1.6697067604312241e-06
GC_4_1187 b_4 NI_4 NS_1187 0 1.1429563429859467e-06
GC_4_1188 b_4 NI_4 NS_1188 0 3.0633003482939170e-06
GC_4_1189 b_4 NI_4 NS_1189 0 -9.6198671061338243e-07
GC_4_1190 b_4 NI_4 NS_1190 0 2.0271686275645204e-06
GC_4_1191 b_4 NI_4 NS_1191 0 4.5490064180851997e-07
GC_4_1192 b_4 NI_4 NS_1192 0 -1.2226961084766204e-06
GC_4_1193 b_4 NI_4 NS_1193 0 3.2356356098243548e-06
GC_4_1194 b_4 NI_4 NS_1194 0 -8.8238713653327060e-07
GC_4_1195 b_4 NI_4 NS_1195 0 -1.6006250831543167e-07
GC_4_1196 b_4 NI_4 NS_1196 0 5.0797816110313857e-07
GC_4_1197 b_4 NI_4 NS_1197 0 -8.4404600459441458e-07
GC_4_1198 b_4 NI_4 NS_1198 0 -4.1916155206995494e-07
GC_4_1199 b_4 NI_4 NS_1199 0 9.8705633441011412e-07
GC_4_1200 b_4 NI_4 NS_1200 0 -1.2634882498407525e-06
GC_4_1201 b_4 NI_4 NS_1201 0 1.4385462602533911e-06
GC_4_1202 b_4 NI_4 NS_1202 0 -5.6892650051792789e-07
GC_4_1203 b_4 NI_4 NS_1203 0 -3.3376942330729331e-08
GC_4_1204 b_4 NI_4 NS_1204 0 9.4899575177168194e-08
GC_4_1205 b_4 NI_4 NS_1205 0 -5.9608936398527831e-07
GC_4_1206 b_4 NI_4 NS_1206 0 -3.3988361224577860e-07
GC_4_1207 b_4 NI_4 NS_1207 0 9.6297867942823718e-07
GC_4_1208 b_4 NI_4 NS_1208 0 -1.0755598735569859e-06
GC_4_1209 b_4 NI_4 NS_1209 0 1.3913817512972710e-06
GC_4_1210 b_4 NI_4 NS_1210 0 -1.2415260044377168e-06
GC_4_1211 b_4 NI_4 NS_1211 0 1.6086379635187078e-07
GC_4_1212 b_4 NI_4 NS_1212 0 -4.5331258641385021e-08
GC_4_1213 b_4 NI_4 NS_1213 0 -4.8805451776307642e-07
GC_4_1214 b_4 NI_4 NS_1214 0 -5.0217409879689325e-07
GC_4_1215 b_4 NI_4 NS_1215 0 1.0601472783188935e-06
GC_4_1216 b_4 NI_4 NS_1216 0 -7.9957387704323154e-07
GC_4_1217 b_4 NI_4 NS_1217 0 1.2253839711753974e-06
GC_4_1218 b_4 NI_4 NS_1218 0 -2.1157296342534620e-06
GC_4_1219 b_4 NI_4 NS_1219 0 4.9452254592013330e-07
GC_4_1220 b_4 NI_4 NS_1220 0 -2.5500871570837064e-07
GC_4_1221 b_4 NI_4 NS_1221 0 -2.4639560876884396e-07
GC_4_1222 b_4 NI_4 NS_1222 0 -9.1751326207786005e-07
GC_4_1223 b_4 NI_4 NS_1223 0 1.9158182140988802e-06
GC_4_1224 b_4 NI_4 NS_1224 0 -9.9682355436588036e-07
GC_4_1225 b_4 NI_4 NS_1225 0 -8.0875204249474102e-06
GC_4_1226 b_4 NI_4 NS_1226 0 -9.1352253382500259e-07
GC_4_1227 b_4 NI_4 NS_1227 0 -3.1590253588749079e-07
GC_4_1228 b_4 NI_4 NS_1228 0 -3.6199237965344106e-06
GC_4_1229 b_4 NI_4 NS_1229 0 -4.8932602372537297e-08
GC_4_1230 b_4 NI_4 NS_1230 0 -3.3151019374481498e-08
GC_4_1231 b_4 NI_4 NS_1231 0 -1.0395733863158447e-07
GC_4_1232 b_4 NI_4 NS_1232 0 -1.2351489720468219e-06
GC_4_1233 b_4 NI_4 NS_1233 0 -1.0202896217314086e-06
GC_4_1234 b_4 NI_4 NS_1234 0 -6.6670072313333927e-07
GC_4_1235 b_4 NI_4 NS_1235 0 1.4550422799090461e-06
GC_4_1236 b_4 NI_4 NS_1236 0 -7.5893834669965559e-07
GC_4_1237 b_4 NI_4 NS_1237 0 1.9403652199902974e-06
GC_4_1238 b_4 NI_4 NS_1238 0 -1.8687388945452176e-06
GC_4_1239 b_4 NI_4 NS_1239 0 -2.2166835352747093e-07
GC_4_1240 b_4 NI_4 NS_1240 0 3.2466687157080480e-07
GC_4_1241 b_4 NI_4 NS_1241 0 2.1427589020083006e-07
GC_4_1242 b_4 NI_4 NS_1242 0 5.2885600557671668e-07
GC_4_1243 b_4 NI_4 NS_1243 0 -1.0742530012866069e-07
GC_4_1244 b_4 NI_4 NS_1244 0 -2.8271655508753924e-07
GC_4_1245 b_4 NI_4 NS_1245 0 7.8974543148382392e-09
GC_4_1246 b_4 NI_4 NS_1246 0 -9.5823318874660567e-08
GC_4_1247 b_4 NI_4 NS_1247 0 -8.8821466961898074e-08
GC_4_1248 b_4 NI_4 NS_1248 0 4.1483568833116789e-08
GC_4_1249 b_4 NI_4 NS_1249 0 -1.2204412635757288e-07
GC_4_1250 b_4 NI_4 NS_1250 0 -5.3450897373985041e-08
GC_4_1251 b_4 NI_4 NS_1251 0 6.1486207105914618e-12
GC_4_1252 b_4 NI_4 NS_1252 0 -1.7071101681517564e-12
GC_4_1253 b_4 NI_4 NS_1253 0 3.5216396847966851e-10
GC_4_1254 b_4 NI_4 NS_1254 0 6.9300720861198271e-10
GC_4_1255 b_4 NI_4 NS_1255 0 1.3351806524440041e-05
GC_4_1256 b_4 NI_4 NS_1256 0 -5.9008757846780447e-08
GC_4_1257 b_4 NI_4 NS_1257 0 -1.4919063025654516e-11
GC_4_1258 b_4 NI_4 NS_1258 0 1.3565960991288281e-10
GC_4_1259 b_4 NI_4 NS_1259 0 3.5691506271271351e-07
GC_4_1260 b_4 NI_4 NS_1260 0 -1.8036858474540791e-07
GC_4_1261 b_4 NI_4 NS_1261 0 2.7982048521105032e-07
GC_4_1262 b_4 NI_4 NS_1262 0 -3.4839667547971915e-07
GC_4_1263 b_4 NI_4 NS_1263 0 4.9688846269635587e-07
GC_4_1264 b_4 NI_4 NS_1264 0 -1.4211337452813549e-06
GC_4_1265 b_4 NI_4 NS_1265 0 -1.1580123258173625e-06
GC_4_1266 b_4 NI_4 NS_1266 0 -4.6157856315081518e-07
GC_4_1267 b_4 NI_4 NS_1267 0 -3.3852704035540042e-07
GC_4_1268 b_4 NI_4 NS_1268 0 -6.2315320674515955e-07
GC_4_1269 b_4 NI_4 NS_1269 0 -2.5799930629420306e-06
GC_4_1270 b_4 NI_4 NS_1270 0 -6.4781485864553902e-07
GC_4_1271 b_4 NI_4 NS_1271 0 7.1553449617308034e-07
GC_4_1272 b_4 NI_4 NS_1272 0 3.5782573118853021e-07
GC_4_1273 b_4 NI_4 NS_1273 0 -7.3448887501673240e-07
GC_4_1274 b_4 NI_4 NS_1274 0 3.7214427393301138e-07
GC_4_1275 b_4 NI_4 NS_1275 0 -9.8995956692297847e-07
GC_4_1276 b_4 NI_4 NS_1276 0 5.8052943759724086e-07
GC_4_1277 b_4 NI_4 NS_1277 0 -4.3434584694885021e-07
GC_4_1278 b_4 NI_4 NS_1278 0 2.6522544642706559e-07
GC_4_1279 b_4 NI_4 NS_1279 0 -8.4585928277618491e-07
GC_4_1280 b_4 NI_4 NS_1280 0 4.5732491897679767e-07
GC_4_1281 b_4 NI_4 NS_1281 0 1.5918351607446737e-07
GC_4_1282 b_4 NI_4 NS_1282 0 1.1045476480487622e-06
GC_4_1283 b_4 NI_4 NS_1283 0 -5.9724289476574598e-07
GC_4_1284 b_4 NI_4 NS_1284 0 1.3109632785262413e-07
GC_4_1285 b_4 NI_4 NS_1285 0 -1.8767398453801223e-06
GC_4_1286 b_4 NI_4 NS_1286 0 1.2955872931369710e-06
GC_4_1287 b_4 NI_4 NS_1287 0 2.0522697849242213e-06
GC_4_1288 b_4 NI_4 NS_1288 0 2.3513000700674817e-07
GC_4_1289 b_4 NI_4 NS_1289 0 -6.8553497679832482e-07
GC_4_1290 b_4 NI_4 NS_1290 0 2.0088559092951263e-07
GC_4_1291 b_4 NI_4 NS_1291 0 9.9851537266824263e-07
GC_4_1292 b_4 NI_4 NS_1292 0 1.6701840573103374e-06
GC_4_1293 b_4 NI_4 NS_1293 0 -2.4331619858363763e-07
GC_4_1294 b_4 NI_4 NS_1294 0 -5.7760860856555964e-07
GC_4_1295 b_4 NI_4 NS_1295 0 -9.1795053977389629e-07
GC_4_1296 b_4 NI_4 NS_1296 0 4.3082205625391277e-07
GC_4_1297 b_4 NI_4 NS_1297 0 1.4279736938233729e-06
GC_4_1298 b_4 NI_4 NS_1298 0 6.8214075708794408e-07
GC_4_1299 b_4 NI_4 NS_1299 0 -3.4147117964442255e-07
GC_4_1300 b_4 NI_4 NS_1300 0 -2.1170585652679394e-07
GC_4_1301 b_4 NI_4 NS_1301 0 -2.9973029124629886e-08
GC_4_1302 b_4 NI_4 NS_1302 0 1.4218679532590951e-06
GC_4_1303 b_4 NI_4 NS_1303 0 4.6149619415076753e-07
GC_4_1304 b_4 NI_4 NS_1304 0 -7.6771759176273458e-07
GC_4_1305 b_4 NI_4 NS_1305 0 -3.5264144880214478e-07
GC_4_1306 b_4 NI_4 NS_1306 0 4.8843516868940060e-08
GC_4_1307 b_4 NI_4 NS_1307 0 3.2445627864754730e-07
GC_4_1308 b_4 NI_4 NS_1308 0 3.7912970360789417e-07
GC_4_1309 b_4 NI_4 NS_1309 0 -1.4602257803825308e-07
GC_4_1310 b_4 NI_4 NS_1310 0 -8.6161061595591514e-09
GC_4_1311 b_4 NI_4 NS_1311 0 1.4120901015838014e-07
GC_4_1312 b_4 NI_4 NS_1312 0 1.2124343992015378e-07
GC_4_1313 b_4 NI_4 NS_1313 0 -1.9293198924225985e-07
GC_4_1314 b_4 NI_4 NS_1314 0 -6.8413937050210806e-08
GC_4_1315 b_4 NI_4 NS_1315 0 4.0854706361245367e-08
GC_4_1316 b_4 NI_4 NS_1316 0 1.9500435546223626e-07
GC_4_1317 b_4 NI_4 NS_1317 0 -1.1264866092872478e-07
GC_4_1318 b_4 NI_4 NS_1318 0 1.0076529089540708e-08
GC_4_1319 b_4 NI_4 NS_1319 0 4.5458923944770705e-08
GC_4_1320 b_4 NI_4 NS_1320 0 4.5514502242422741e-09
GC_4_1321 b_4 NI_4 NS_1321 0 -2.9963274436265323e-07
GC_4_1322 b_4 NI_4 NS_1322 0 -5.1511697798452978e-08
GC_4_1323 b_4 NI_4 NS_1323 0 -9.0274597247633483e-08
GC_4_1324 b_4 NI_4 NS_1324 0 6.0417936756737288e-08
GC_4_1325 b_4 NI_4 NS_1325 0 -2.3104818327543131e-07
GC_4_1326 b_4 NI_4 NS_1326 0 8.0694595524673617e-08
GC_4_1327 b_4 NI_4 NS_1327 0 -1.3259209334879702e-07
GC_4_1328 b_4 NI_4 NS_1328 0 -7.1016518011357883e-08
GC_4_1329 b_4 NI_4 NS_1329 0 -4.3085748570716818e-07
GC_4_1330 b_4 NI_4 NS_1330 0 -5.3628430870347146e-08
GC_4_1331 b_4 NI_4 NS_1331 0 -4.1936675387714381e-07
GC_4_1332 b_4 NI_4 NS_1332 0 6.1406752469158383e-08
GC_4_1333 b_4 NI_4 NS_1333 0 -4.4043868201302893e-07
GC_4_1334 b_4 NI_4 NS_1334 0 1.4691496328729628e-07
GC_4_1335 b_4 NI_4 NS_1335 0 -5.1097823540191924e-07
GC_4_1336 b_4 NI_4 NS_1336 0 9.9964930319413576e-08
GC_4_1337 b_4 NI_4 NS_1337 0 -9.6170663476043375e-07
GC_4_1338 b_4 NI_4 NS_1338 0 -9.6201991733592270e-08
GC_4_1339 b_4 NI_4 NS_1339 0 2.6182516020345657e-06
GC_4_1340 b_4 NI_4 NS_1340 0 2.9793837837785693e-06
GC_4_1341 b_4 NI_4 NS_1341 0 -6.1475024123758474e-07
GC_4_1342 b_4 NI_4 NS_1342 0 1.0339430972069629e-06
GC_4_1343 b_4 NI_4 NS_1343 0 9.1585165321434355e-09
GC_4_1344 b_4 NI_4 NS_1344 0 2.5337436139334555e-08
GC_4_1345 b_4 NI_4 NS_1345 0 -4.6874895434752881e-07
GC_4_1346 b_4 NI_4 NS_1346 0 8.2782653536162076e-07
GC_4_1347 b_4 NI_4 NS_1347 0 8.6795545952802341e-09
GC_4_1348 b_4 NI_4 NS_1348 0 3.8300011512099672e-07
GC_4_1349 b_4 NI_4 NS_1349 0 -8.6727475750574607e-07
GC_4_1350 b_4 NI_4 NS_1350 0 -7.0681656139383884e-08
GC_4_1351 b_4 NI_4 NS_1351 0 -9.7701459086729452e-07
GC_4_1352 b_4 NI_4 NS_1352 0 -1.7981772292353577e-07
GC_4_1353 b_4 NI_4 NS_1353 0 1.0738473523203329e-07
GC_4_1354 b_4 NI_4 NS_1354 0 -1.4754532886872966e-07
GC_4_1355 b_4 NI_4 NS_1355 0 6.6801744770247203e-08
GC_4_1356 b_4 NI_4 NS_1356 0 1.4718154706392771e-08
GC_4_1357 b_4 NI_4 NS_1357 0 -6.9818551725241095e-08
GC_4_1358 b_4 NI_4 NS_1358 0 1.6103497077786523e-07
GC_4_1359 b_4 NI_4 NS_1359 0 2.7786733489996990e-08
GC_4_1360 b_4 NI_4 NS_1360 0 -4.0821854199217278e-08
GC_4_1361 b_4 NI_4 NS_1361 0 -8.1243021840519878e-08
GC_4_1362 b_4 NI_4 NS_1362 0 1.6047194731931713e-07
GC_4_1363 b_4 NI_4 NS_1363 0 5.6556664225795340e-08
GC_4_1364 b_4 NI_4 NS_1364 0 -1.6778197183112433e-08
GC_4_1365 b_4 NI_4 NS_1365 0 -1.1804175237589369e-11
GC_4_1366 b_4 NI_4 NS_1366 0 5.2790010993857104e-12
GC_4_1367 b_4 NI_4 NS_1367 0 -3.4095401817629186e-10
GC_4_1368 b_4 NI_4 NS_1368 0 -9.7317200931801163e-10
GD_4_1 b_4 NI_4 NA_1 0 5.9084076393106178e-04
GD_4_2 b_4 NI_4 NA_2 0 1.3004902192071191e-02
GD_4_3 b_4 NI_4 NA_3 0 -4.2441400590540112e-03
GD_4_4 b_4 NI_4 NA_4 0 -8.6867583427960981e-03
GD_4_5 b_4 NI_4 NA_5 0 2.6994458370821475e-05
GD_4_6 b_4 NI_4 NA_6 0 1.0031817901016784e-04
GD_4_7 b_4 NI_4 NA_7 0 1.1836190164646708e-06
GD_4_8 b_4 NI_4 NA_8 0 3.6701583821687476e-06
GD_4_9 b_4 NI_4 NA_9 0 4.7457867232243437e-07
GD_4_10 b_4 NI_4 NA_10 0 -5.5537910586247965e-06
GD_4_11 b_4 NI_4 NA_11 0 5.6258472687503064e-06
GD_4_12 b_4 NI_4 NA_12 0 -1.8573495908082893e-06
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 -1.1889664709065413e-04
GC_5_2 b_5 NI_5 NS_2 0 -2.1515751559464628e-06
GC_5_3 b_5 NI_5 NS_3 0 -2.4447829657187102e-10
GC_5_4 b_5 NI_5 NS_4 0 2.5353390384257263e-09
GC_5_5 b_5 NI_5 NS_5 0 1.5643085686690507e-06
GC_5_6 b_5 NI_5 NS_6 0 -1.5218359227371622e-06
GC_5_7 b_5 NI_5 NS_7 0 -8.9297682017459832e-09
GC_5_8 b_5 NI_5 NS_8 0 -6.1820522075631427e-06
GC_5_9 b_5 NI_5 NS_9 0 -7.6539313511896647e-06
GC_5_10 b_5 NI_5 NS_10 0 5.3261385171082713e-07
GC_5_11 b_5 NI_5 NS_11 0 -9.8452195619778207e-07
GC_5_12 b_5 NI_5 NS_12 0 -4.3923453905293837e-06
GC_5_13 b_5 NI_5 NS_13 0 -1.5585556945236749e-05
GC_5_14 b_5 NI_5 NS_14 0 -1.3013886506004499e-06
GC_5_15 b_5 NI_5 NS_15 0 -5.3235184111459471e-06
GC_5_16 b_5 NI_5 NS_16 0 1.9150004917651977e-05
GC_5_17 b_5 NI_5 NS_17 0 4.4241059733161001e-06
GC_5_18 b_5 NI_5 NS_18 0 -3.1123179387206526e-06
GC_5_19 b_5 NI_5 NS_19 0 1.2804781909340864e-07
GC_5_20 b_5 NI_5 NS_20 0 -2.5891791652787207e-06
GC_5_21 b_5 NI_5 NS_21 0 -2.4876404667236962e-05
GC_5_22 b_5 NI_5 NS_22 0 2.8210753508880433e-05
GC_5_23 b_5 NI_5 NS_23 0 2.7762971339719761e-05
GC_5_24 b_5 NI_5 NS_24 0 -8.7259228628811039e-06
GC_5_25 b_5 NI_5 NS_25 0 -7.7819274365814059e-06
GC_5_26 b_5 NI_5 NS_26 0 -4.1753177848418828e-06
GC_5_27 b_5 NI_5 NS_27 0 1.2787916911927672e-05
GC_5_28 b_5 NI_5 NS_28 0 2.6107424750830461e-05
GC_5_29 b_5 NI_5 NS_29 0 1.4270067300445181e-06
GC_5_30 b_5 NI_5 NS_30 0 -8.8305598524600137e-06
GC_5_31 b_5 NI_5 NS_31 0 -2.7324697223825537e-05
GC_5_32 b_5 NI_5 NS_32 0 5.0137306908634824e-06
GC_5_33 b_5 NI_5 NS_33 0 4.0396636342590801e-05
GC_5_34 b_5 NI_5 NS_34 0 9.6550510286998473e-06
GC_5_35 b_5 NI_5 NS_35 0 -2.8820961577319625e-06
GC_5_36 b_5 NI_5 NS_36 0 -4.3143668047876754e-06
GC_5_37 b_5 NI_5 NS_37 0 1.3053639552501346e-05
GC_5_38 b_5 NI_5 NS_38 0 1.8104097869826252e-05
GC_5_39 b_5 NI_5 NS_39 0 3.5097808609263850e-06
GC_5_40 b_5 NI_5 NS_40 0 -1.0678067996826689e-05
GC_5_41 b_5 NI_5 NS_41 0 -6.1544159323469088e-06
GC_5_42 b_5 NI_5 NS_42 0 1.0310052233501291e-06
GC_5_43 b_5 NI_5 NS_43 0 1.8592829956304333e-05
GC_5_44 b_5 NI_5 NS_44 0 4.7647989951188255e-06
GC_5_45 b_5 NI_5 NS_45 0 -1.6257210838219363e-07
GC_5_46 b_5 NI_5 NS_46 0 -4.0317313270447696e-06
GC_5_47 b_5 NI_5 NS_47 0 5.3001343913731225e-06
GC_5_48 b_5 NI_5 NS_48 0 1.3913340945965307e-05
GC_5_49 b_5 NI_5 NS_49 0 7.3647530309034177e-06
GC_5_50 b_5 NI_5 NS_50 0 -1.1146120787191955e-05
GC_5_51 b_5 NI_5 NS_51 0 -1.3430338482860120e-06
GC_5_52 b_5 NI_5 NS_52 0 1.0232543447877870e-06
GC_5_53 b_5 NI_5 NS_53 0 1.0874239404547311e-05
GC_5_54 b_5 NI_5 NS_54 0 3.8626538755829085e-06
GC_5_55 b_5 NI_5 NS_55 0 1.6867602056248018e-06
GC_5_56 b_5 NI_5 NS_56 0 -5.9600522694430144e-07
GC_5_57 b_5 NI_5 NS_57 0 5.6731243600739530e-06
GC_5_58 b_5 NI_5 NS_58 0 1.6014340974434156e-06
GC_5_59 b_5 NI_5 NS_59 0 3.3818682820134912e-06
GC_5_60 b_5 NI_5 NS_60 0 2.0535676221903238e-06
GC_5_61 b_5 NI_5 NS_61 0 1.1002372226381559e-05
GC_5_62 b_5 NI_5 NS_62 0 3.6804861048338245e-06
GC_5_63 b_5 NI_5 NS_63 0 4.8497228696269655e-06
GC_5_64 b_5 NI_5 NS_64 0 -8.6121319731254356e-08
GC_5_65 b_5 NI_5 NS_65 0 9.9794194201138728e-06
GC_5_66 b_5 NI_5 NS_66 0 -1.1587617265640389e-06
GC_5_67 b_5 NI_5 NS_67 0 8.2788149453850880e-06
GC_5_68 b_5 NI_5 NS_68 0 2.9673089861178826e-06
GC_5_69 b_5 NI_5 NS_69 0 1.9120277045620166e-05
GC_5_70 b_5 NI_5 NS_70 0 -5.6689227296960076e-06
GC_5_71 b_5 NI_5 NS_71 0 7.2485954309899656e-06
GC_5_72 b_5 NI_5 NS_72 0 -4.0295065063293499e-06
GC_5_73 b_5 NI_5 NS_73 0 1.3800813549045525e-05
GC_5_74 b_5 NI_5 NS_74 0 -1.2000538368758908e-05
GC_5_75 b_5 NI_5 NS_75 0 1.2506358383096459e-05
GC_5_76 b_5 NI_5 NS_76 0 -3.9183447949779621e-06
GC_5_77 b_5 NI_5 NS_77 0 9.3634142103169569e-06
GC_5_78 b_5 NI_5 NS_78 0 -2.6978357354144362e-05
GC_5_79 b_5 NI_5 NS_79 0 2.5168592864109854e-06
GC_5_80 b_5 NI_5 NS_80 0 -1.2425235379422644e-05
GC_5_81 b_5 NI_5 NS_81 0 -8.1224252588395234e-06
GC_5_82 b_5 NI_5 NS_82 0 -1.8906424310558306e-05
GC_5_83 b_5 NI_5 NS_83 0 -4.4970473439652277e-06
GC_5_84 b_5 NI_5 NS_84 0 -1.2065329732568956e-05
GC_5_85 b_5 NI_5 NS_85 0 5.2902140736998074e-05
GC_5_86 b_5 NI_5 NS_86 0 -8.9264414192413187e-05
GC_5_87 b_5 NI_5 NS_87 0 -9.8974233966754843e-06
GC_5_88 b_5 NI_5 NS_88 0 6.3392390148234806e-07
GC_5_89 b_5 NI_5 NS_89 0 3.8297079174503616e-07
GC_5_90 b_5 NI_5 NS_90 0 -1.3807140095383701e-07
GC_5_91 b_5 NI_5 NS_91 0 -2.6243898425164280e-06
GC_5_92 b_5 NI_5 NS_92 0 -2.3105604725278385e-06
GC_5_93 b_5 NI_5 NS_93 0 -4.4577511518001965e-06
GC_5_94 b_5 NI_5 NS_94 0 2.7145419442112930e-07
GC_5_95 b_5 NI_5 NS_95 0 -1.7068913134340521e-05
GC_5_96 b_5 NI_5 NS_96 0 9.6343678953072643e-06
GC_5_97 b_5 NI_5 NS_97 0 -8.5804545863665989e-06
GC_5_98 b_5 NI_5 NS_98 0 3.7246476925015236e-05
GC_5_99 b_5 NI_5 NS_99 0 -7.2739651809057006e-06
GC_5_100 b_5 NI_5 NS_100 0 3.7766522596988243e-07
GC_5_101 b_5 NI_5 NS_101 0 -1.3438135991974461e-05
GC_5_102 b_5 NI_5 NS_102 0 1.9879391735282895e-06
GC_5_103 b_5 NI_5 NS_103 0 -4.6768387281282922e-06
GC_5_104 b_5 NI_5 NS_104 0 -3.4323461426562934e-06
GC_5_105 b_5 NI_5 NS_105 0 -6.4511241002083884e-06
GC_5_106 b_5 NI_5 NS_106 0 1.0470458507243154e-06
GC_5_107 b_5 NI_5 NS_107 0 -3.0717704024622102e-06
GC_5_108 b_5 NI_5 NS_108 0 8.7596279999525800e-07
GC_5_109 b_5 NI_5 NS_109 0 -1.8095974786191948e-06
GC_5_110 b_5 NI_5 NS_110 0 -9.3346422712773053e-07
GC_5_111 b_5 NI_5 NS_111 0 -2.5782257563899458e-10
GC_5_112 b_5 NI_5 NS_112 0 4.1882528067564739e-10
GC_5_113 b_5 NI_5 NS_113 0 2.1382066443717849e-09
GC_5_114 b_5 NI_5 NS_114 0 -2.6515544411045013e-08
GC_5_115 b_5 NI_5 NS_115 0 -3.8127591865756122e-05
GC_5_116 b_5 NI_5 NS_116 0 2.2429767180709047e-06
GC_5_117 b_5 NI_5 NS_117 0 5.7510496873688842e-11
GC_5_118 b_5 NI_5 NS_118 0 3.0676964445858673e-09
GC_5_119 b_5 NI_5 NS_119 0 -1.9281103331311003e-06
GC_5_120 b_5 NI_5 NS_120 0 -1.7008098849606101e-06
GC_5_121 b_5 NI_5 NS_121 0 -5.6014731867516261e-06
GC_5_122 b_5 NI_5 NS_122 0 2.8809775549826579e-06
GC_5_123 b_5 NI_5 NS_123 0 -1.6609394906148689e-05
GC_5_124 b_5 NI_5 NS_124 0 1.9115780634440216e-05
GC_5_125 b_5 NI_5 NS_125 0 1.5381275932041268e-05
GC_5_126 b_5 NI_5 NS_126 0 1.0271579380547803e-05
GC_5_127 b_5 NI_5 NS_127 0 1.7283129879715551e-05
GC_5_128 b_5 NI_5 NS_128 0 2.3212258180843902e-05
GC_5_129 b_5 NI_5 NS_129 0 3.0965004130508651e-05
GC_5_130 b_5 NI_5 NS_130 0 5.3090198320120298e-06
GC_5_131 b_5 NI_5 NS_131 0 -3.3865791025794973e-06
GC_5_132 b_5 NI_5 NS_132 0 -2.1456102217143211e-06
GC_5_133 b_5 NI_5 NS_133 0 1.7199397368067215e-05
GC_5_134 b_5 NI_5 NS_134 0 -2.1238048569866466e-06
GC_5_135 b_5 NI_5 NS_135 0 1.2959164412501719e-04
GC_5_136 b_5 NI_5 NS_136 0 3.5268884941509057e-05
GC_5_137 b_5 NI_5 NS_137 0 -2.8361249489568621e-05
GC_5_138 b_5 NI_5 NS_138 0 -1.0001870664112396e-04
GC_5_139 b_5 NI_5 NS_139 0 2.5325861595112814e-05
GC_5_140 b_5 NI_5 NS_140 0 -3.1108753041936399e-05
GC_5_141 b_5 NI_5 NS_141 0 -4.1100398159582652e-05
GC_5_142 b_5 NI_5 NS_142 0 -1.6753408761562176e-04
GC_5_143 b_5 NI_5 NS_143 0 -4.1818795879431327e-05
GC_5_144 b_5 NI_5 NS_144 0 -5.5999248943759956e-06
GC_5_145 b_5 NI_5 NS_145 0 2.2902356589975465e-05
GC_5_146 b_5 NI_5 NS_146 0 -1.5132347380506316e-04
GC_5_147 b_5 NI_5 NS_147 0 -2.3194036016245897e-04
GC_5_148 b_5 NI_5 NS_148 0 1.1299732452236540e-04
GC_5_149 b_5 NI_5 NS_149 0 -3.7469245150731993e-05
GC_5_150 b_5 NI_5 NS_150 0 1.3726672460795792e-05
GC_5_151 b_5 NI_5 NS_151 0 -1.3772298123038604e-04
GC_5_152 b_5 NI_5 NS_152 0 1.2973733095056485e-04
GC_5_153 b_5 NI_5 NS_153 0 3.6014582026270066e-05
GC_5_154 b_5 NI_5 NS_154 0 4.1758562918810051e-05
GC_5_155 b_5 NI_5 NS_155 0 -3.8325642753743231e-05
GC_5_156 b_5 NI_5 NS_156 0 4.2732818851908030e-05
GC_5_157 b_5 NI_5 NS_157 0 8.7551066675110124e-05
GC_5_158 b_5 NI_5 NS_158 0 1.1830579937756195e-04
GC_5_159 b_5 NI_5 NS_159 0 2.7199706886354564e-05
GC_5_160 b_5 NI_5 NS_160 0 1.0487347192525999e-05
GC_5_161 b_5 NI_5 NS_161 0 8.6918393408963348e-05
GC_5_162 b_5 NI_5 NS_162 0 6.5387623905943581e-05
GC_5_163 b_5 NI_5 NS_163 0 2.0649678924447743e-05
GC_5_164 b_5 NI_5 NS_164 0 -5.7329131399768548e-05
GC_5_165 b_5 NI_5 NS_165 0 1.7010778322306309e-05
GC_5_166 b_5 NI_5 NS_166 0 -8.6980469626393611e-06
GC_5_167 b_5 NI_5 NS_167 0 8.3266760461515342e-06
GC_5_168 b_5 NI_5 NS_168 0 -3.3101616807591406e-05
GC_5_169 b_5 NI_5 NS_169 0 -8.8261831356155505e-06
GC_5_170 b_5 NI_5 NS_170 0 3.3237449069129020e-07
GC_5_171 b_5 NI_5 NS_171 0 -2.3513340626676673e-06
GC_5_172 b_5 NI_5 NS_172 0 8.4561586669689475e-06
GC_5_173 b_5 NI_5 NS_173 0 1.0134445593471270e-05
GC_5_174 b_5 NI_5 NS_174 0 6.1702245215249564e-06
GC_5_175 b_5 NI_5 NS_175 0 1.2106299139909123e-05
GC_5_176 b_5 NI_5 NS_176 0 -7.8948457355306812e-06
GC_5_177 b_5 NI_5 NS_177 0 -3.4457707640832506e-06
GC_5_178 b_5 NI_5 NS_178 0 -5.4105858191467699e-07
GC_5_179 b_5 NI_5 NS_179 0 2.5534799949851457e-06
GC_5_180 b_5 NI_5 NS_180 0 7.3550268394186193e-06
GC_5_181 b_5 NI_5 NS_181 0 1.3648109030606845e-05
GC_5_182 b_5 NI_5 NS_182 0 2.7056935557435033e-06
GC_5_183 b_5 NI_5 NS_183 0 4.5460336438598913e-06
GC_5_184 b_5 NI_5 NS_184 0 -1.4254847048807256e-05
GC_5_185 b_5 NI_5 NS_185 0 -5.8809752922506606e-06
GC_5_186 b_5 NI_5 NS_186 0 4.1779264621864276e-06
GC_5_187 b_5 NI_5 NS_187 0 1.0407133752414071e-05
GC_5_188 b_5 NI_5 NS_188 0 9.8673447181516309e-06
GC_5_189 b_5 NI_5 NS_189 0 1.7371589583654884e-05
GC_5_190 b_5 NI_5 NS_190 0 -4.2134201147708340e-06
GC_5_191 b_5 NI_5 NS_191 0 -9.1860417226910723e-06
GC_5_192 b_5 NI_5 NS_192 0 -1.5417465867839014e-05
GC_5_193 b_5 NI_5 NS_193 0 -3.9937499798253579e-06
GC_5_194 b_5 NI_5 NS_194 0 1.3459824227561652e-05
GC_5_195 b_5 NI_5 NS_195 0 2.1061332083120151e-05
GC_5_196 b_5 NI_5 NS_196 0 -6.9754222331097020e-07
GC_5_197 b_5 NI_5 NS_197 0 9.0885470574570329e-06
GC_5_198 b_5 NI_5 NS_198 0 -1.7352309911017163e-05
GC_5_199 b_5 NI_5 NS_199 0 1.8901206776109675e-06
GC_5_200 b_5 NI_5 NS_200 0 -1.4898986060769832e-05
GC_5_201 b_5 NI_5 NS_201 0 -1.3643861468905871e-05
GC_5_202 b_5 NI_5 NS_202 0 4.0672463723472461e-06
GC_5_203 b_5 NI_5 NS_203 0 1.3198662440719891e-08
GC_5_204 b_5 NI_5 NS_204 0 -4.9292565096098132e-08
GC_5_205 b_5 NI_5 NS_205 0 8.7094357729505977e-06
GC_5_206 b_5 NI_5 NS_206 0 1.1413293836885969e-05
GC_5_207 b_5 NI_5 NS_207 0 1.0949791557172593e-05
GC_5_208 b_5 NI_5 NS_208 0 -1.1467443916444867e-05
GC_5_209 b_5 NI_5 NS_209 0 -3.5677421690301139e-06
GC_5_210 b_5 NI_5 NS_210 0 -1.0053467973172744e-05
GC_5_211 b_5 NI_5 NS_211 0 -2.0108159777408537e-06
GC_5_212 b_5 NI_5 NS_212 0 1.3050037780383804e-05
GC_5_213 b_5 NI_5 NS_213 0 9.7275568882406164e-07
GC_5_214 b_5 NI_5 NS_214 0 -7.2791641367303127e-06
GC_5_215 b_5 NI_5 NS_215 0 7.4349155539845637e-06
GC_5_216 b_5 NI_5 NS_216 0 1.7180972443814681e-06
GC_5_217 b_5 NI_5 NS_217 0 -6.1040300134950948e-06
GC_5_218 b_5 NI_5 NS_218 0 -8.8986483549165435e-06
GC_5_219 b_5 NI_5 NS_219 0 -4.1281684490553222e-06
GC_5_220 b_5 NI_5 NS_220 0 9.6390254578565552e-06
GC_5_221 b_5 NI_5 NS_221 0 3.3246451361971314e-06
GC_5_222 b_5 NI_5 NS_222 0 6.0744664728307644e-06
GC_5_223 b_5 NI_5 NS_223 0 5.7495178745086687e-06
GC_5_224 b_5 NI_5 NS_224 0 5.2304200721594049e-07
GC_5_225 b_5 NI_5 NS_225 0 5.7042917761439440e-11
GC_5_226 b_5 NI_5 NS_226 0 1.4838831109443849e-10
GC_5_227 b_5 NI_5 NS_227 0 6.0313806619174956e-09
GC_5_228 b_5 NI_5 NS_228 0 -8.4056172822875333e-09
GC_5_229 b_5 NI_5 NS_229 0 3.0652005901740057e-04
GC_5_230 b_5 NI_5 NS_230 0 -1.4375836080391030e-05
GC_5_231 b_5 NI_5 NS_231 0 -1.2385117047136972e-09
GC_5_232 b_5 NI_5 NS_232 0 -1.9194440502993037e-08
GC_5_233 b_5 NI_5 NS_233 0 3.2004164038130290e-06
GC_5_234 b_5 NI_5 NS_234 0 -3.9681503481355950e-06
GC_5_235 b_5 NI_5 NS_235 0 -1.2573342228250492e-05
GC_5_236 b_5 NI_5 NS_236 0 -1.0250931065608287e-06
GC_5_237 b_5 NI_5 NS_237 0 3.9887653671701077e-05
GC_5_238 b_5 NI_5 NS_238 0 8.6396664766261422e-07
GC_5_239 b_5 NI_5 NS_239 0 -4.2800323533641159e-05
GC_5_240 b_5 NI_5 NS_240 0 -2.4451092254023126e-05
GC_5_241 b_5 NI_5 NS_241 0 1.1877307505924250e-06
GC_5_242 b_5 NI_5 NS_242 0 4.3284247759121258e-05
GC_5_243 b_5 NI_5 NS_243 0 1.0653262743003706e-05
GC_5_244 b_5 NI_5 NS_244 0 -4.8921231503768847e-05
GC_5_245 b_5 NI_5 NS_245 0 2.9254045420764521e-06
GC_5_246 b_5 NI_5 NS_246 0 6.2451616582240076e-06
GC_5_247 b_5 NI_5 NS_247 0 -4.5618512784543644e-05
GC_5_248 b_5 NI_5 NS_248 0 1.8884929852287794e-06
GC_5_249 b_5 NI_5 NS_249 0 1.0003123891785796e-04
GC_5_250 b_5 NI_5 NS_250 0 1.2285660411274392e-04
GC_5_251 b_5 NI_5 NS_251 0 -7.5037288390589899e-05
GC_5_252 b_5 NI_5 NS_252 0 -1.3519238234484000e-04
GC_5_253 b_5 NI_5 NS_253 0 -6.7763285286072999e-05
GC_5_254 b_5 NI_5 NS_254 0 4.9170014362576888e-05
GC_5_255 b_5 NI_5 NS_255 0 1.3378245801978103e-04
GC_5_256 b_5 NI_5 NS_256 0 -2.6374211743579703e-05
GC_5_257 b_5 NI_5 NS_257 0 -8.7278702774256256e-05
GC_5_258 b_5 NI_5 NS_258 0 -1.1628849228227016e-05
GC_5_259 b_5 NI_5 NS_259 0 -9.6762932987484436e-05
GC_5_260 b_5 NI_5 NS_260 0 2.1083572473927856e-04
GC_5_261 b_5 NI_5 NS_261 0 1.6567950605466785e-04
GC_5_262 b_5 NI_5 NS_262 0 -2.1188394429151139e-04
GC_5_263 b_5 NI_5 NS_263 0 -8.1910068389974707e-05
GC_5_264 b_5 NI_5 NS_264 0 1.9157059395536191e-05
GC_5_265 b_5 NI_5 NS_265 0 1.6054321701364379e-04
GC_5_266 b_5 NI_5 NS_266 0 4.4269398544493915e-05
GC_5_267 b_5 NI_5 NS_267 0 -8.8292491002378500e-05
GC_5_268 b_5 NI_5 NS_268 0 -7.2082536009616296e-05
GC_5_269 b_5 NI_5 NS_269 0 -8.5464952767069023e-05
GC_5_270 b_5 NI_5 NS_270 0 6.3489913137986220e-05
GC_5_271 b_5 NI_5 NS_271 0 1.4126679595945931e-04
GC_5_272 b_5 NI_5 NS_272 0 -4.6881954553281843e-05
GC_5_273 b_5 NI_5 NS_273 0 -6.6093588023825316e-05
GC_5_274 b_5 NI_5 NS_274 0 -2.4355717001953161e-05
GC_5_275 b_5 NI_5 NS_275 0 6.0401776938855225e-05
GC_5_276 b_5 NI_5 NS_276 0 1.1474581756759074e-04
GC_5_277 b_5 NI_5 NS_277 0 -2.2017764679448247e-05
GC_5_278 b_5 NI_5 NS_278 0 -1.2142962506048013e-04
GC_5_279 b_5 NI_5 NS_279 0 -4.4471483392111517e-05
GC_5_280 b_5 NI_5 NS_280 0 1.0923655437459580e-05
GC_5_281 b_5 NI_5 NS_281 0 4.7464788532059206e-05
GC_5_282 b_5 NI_5 NS_282 0 -9.9240655813282828e-06
GC_5_283 b_5 NI_5 NS_283 0 -3.2079591645760286e-05
GC_5_284 b_5 NI_5 NS_284 0 -7.5858717131385008e-06
GC_5_285 b_5 NI_5 NS_285 0 2.1298598719488319e-05
GC_5_286 b_5 NI_5 NS_286 0 -4.6121029704139652e-06
GC_5_287 b_5 NI_5 NS_287 0 -3.2316567447941033e-05
GC_5_288 b_5 NI_5 NS_288 0 -2.5188213293615734e-05
GC_5_289 b_5 NI_5 NS_289 0 1.2511323836103328e-05
GC_5_290 b_5 NI_5 NS_290 0 6.5132080002209511e-06
GC_5_291 b_5 NI_5 NS_291 0 -2.0424006351442602e-05
GC_5_292 b_5 NI_5 NS_292 0 -7.6315545719397064e-06
GC_5_293 b_5 NI_5 NS_293 0 1.3991693687049743e-05
GC_5_294 b_5 NI_5 NS_294 0 -1.2277477632724402e-05
GC_5_295 b_5 NI_5 NS_295 0 -4.1514445536045336e-05
GC_5_296 b_5 NI_5 NS_296 0 -1.6952576005547190e-05
GC_5_297 b_5 NI_5 NS_297 0 1.1564369778263144e-05
GC_5_298 b_5 NI_5 NS_298 0 -1.4313418342151018e-06
GC_5_299 b_5 NI_5 NS_299 0 -3.0401004475387423e-05
GC_5_300 b_5 NI_5 NS_300 0 5.6251336308546952e-06
GC_5_301 b_5 NI_5 NS_301 0 1.6016639662712352e-05
GC_5_302 b_5 NI_5 NS_302 0 -2.0571427143085767e-05
GC_5_303 b_5 NI_5 NS_303 0 -5.0239545299514118e-05
GC_5_304 b_5 NI_5 NS_304 0 -1.7714965386577863e-06
GC_5_305 b_5 NI_5 NS_305 0 1.1585345885533743e-05
GC_5_306 b_5 NI_5 NS_306 0 -1.1191609971557957e-05
GC_5_307 b_5 NI_5 NS_307 0 -3.2363535725972869e-05
GC_5_308 b_5 NI_5 NS_308 0 2.5180975187365517e-05
GC_5_309 b_5 NI_5 NS_309 0 1.0237907885533024e-05
GC_5_310 b_5 NI_5 NS_310 0 -3.5896465168936447e-05
GC_5_311 b_5 NI_5 NS_311 0 -3.4868718564753637e-05
GC_5_312 b_5 NI_5 NS_312 0 1.8378559938362386e-05
GC_5_313 b_5 NI_5 NS_313 0 -5.6366146617224474e-05
GC_5_314 b_5 NI_5 NS_314 0 1.3314460696518997e-04
GC_5_315 b_5 NI_5 NS_315 0 -1.5278319210330320e-05
GC_5_316 b_5 NI_5 NS_316 0 -3.1719296894040927e-05
GC_5_317 b_5 NI_5 NS_317 0 -3.7759710770529509e-07
GC_5_318 b_5 NI_5 NS_318 0 3.9613389311759361e-07
GC_5_319 b_5 NI_5 NS_319 0 -2.0157655195783879e-05
GC_5_320 b_5 NI_5 NS_320 0 3.2122140613125793e-05
GC_5_321 b_5 NI_5 NS_321 0 -1.4301666073363391e-05
GC_5_322 b_5 NI_5 NS_322 0 -3.3396349653377985e-05
GC_5_323 b_5 NI_5 NS_323 0 -6.1620332090231445e-06
GC_5_324 b_5 NI_5 NS_324 0 5.1170144430924184e-06
GC_5_325 b_5 NI_5 NS_325 0 -2.1210447911042036e-05
GC_5_326 b_5 NI_5 NS_326 0 -6.5713064447515601e-05
GC_5_327 b_5 NI_5 NS_327 0 -9.1587285794777830e-06
GC_5_328 b_5 NI_5 NS_328 0 -2.0643971600732332e-05
GC_5_329 b_5 NI_5 NS_329 0 1.5020247707457899e-05
GC_5_330 b_5 NI_5 NS_330 0 2.2754098137952523e-05
GC_5_331 b_5 NI_5 NS_331 0 -6.7861253167620815e-06
GC_5_332 b_5 NI_5 NS_332 0 2.7712147583298113e-05
GC_5_333 b_5 NI_5 NS_333 0 -1.1040554618325064e-05
GC_5_334 b_5 NI_5 NS_334 0 -2.1529685286324218e-05
GC_5_335 b_5 NI_5 NS_335 0 -1.1040049298956425e-05
GC_5_336 b_5 NI_5 NS_336 0 2.3841904655309710e-05
GC_5_337 b_5 NI_5 NS_337 0 5.1225220296293250e-06
GC_5_338 b_5 NI_5 NS_338 0 -1.5323216617572416e-05
GC_5_339 b_5 NI_5 NS_339 0 -4.7531903705875846e-10
GC_5_340 b_5 NI_5 NS_340 0 -9.1476640412662822e-10
GC_5_341 b_5 NI_5 NS_341 0 -5.5313560196141319e-08
GC_5_342 b_5 NI_5 NS_342 0 7.4254738897637690e-09
GC_5_343 b_5 NI_5 NS_343 0 -2.0465926465440562e-04
GC_5_344 b_5 NI_5 NS_344 0 -3.3255113924366404e-06
GC_5_345 b_5 NI_5 NS_345 0 1.2945496057086887e-09
GC_5_346 b_5 NI_5 NS_346 0 9.6766100896451059e-09
GC_5_347 b_5 NI_5 NS_347 0 -4.2560813252057753e-06
GC_5_348 b_5 NI_5 NS_348 0 6.2139735074423222e-06
GC_5_349 b_5 NI_5 NS_349 0 3.7169297126477360e-06
GC_5_350 b_5 NI_5 NS_350 0 -8.0226869247019894e-06
GC_5_351 b_5 NI_5 NS_351 0 2.1711134076639127e-05
GC_5_352 b_5 NI_5 NS_352 0 -8.4068450754479287e-06
GC_5_353 b_5 NI_5 NS_353 0 -2.1213740968409285e-05
GC_5_354 b_5 NI_5 NS_354 0 -1.2028648664585840e-06
GC_5_355 b_5 NI_5 NS_355 0 -2.9295847391368612e-05
GC_5_356 b_5 NI_5 NS_356 0 -2.8036650245747167e-05
GC_5_357 b_5 NI_5 NS_357 0 -4.8460987734380513e-06
GC_5_358 b_5 NI_5 NS_358 0 1.6200710300739461e-05
GC_5_359 b_5 NI_5 NS_359 0 -2.6737720054700640e-06
GC_5_360 b_5 NI_5 NS_360 0 -7.1113141233273771e-06
GC_5_361 b_5 NI_5 NS_361 0 -2.2547099050717673e-05
GC_5_362 b_5 NI_5 NS_362 0 5.7325211312431741e-06
GC_5_363 b_5 NI_5 NS_363 0 -1.8497082933064380e-04
GC_5_364 b_5 NI_5 NS_364 0 -4.4589107853631858e-05
GC_5_365 b_5 NI_5 NS_365 0 6.1993810985186491e-05
GC_5_366 b_5 NI_5 NS_366 0 1.3751678573478118e-04
GC_5_367 b_5 NI_5 NS_367 0 -3.7420883334896051e-05
GC_5_368 b_5 NI_5 NS_368 0 5.6316425798516686e-05
GC_5_369 b_5 NI_5 NS_369 0 9.5006455202844268e-05
GC_5_370 b_5 NI_5 NS_370 0 2.4592086888510807e-04
GC_5_371 b_5 NI_5 NS_371 0 7.3727691869039959e-05
GC_5_372 b_5 NI_5 NS_372 0 8.1340630329171096e-07
GC_5_373 b_5 NI_5 NS_373 0 -1.6013482313570892e-05
GC_5_374 b_5 NI_5 NS_374 0 2.6083741747888256e-04
GC_5_375 b_5 NI_5 NS_375 0 3.6487194359218118e-04
GC_5_376 b_5 NI_5 NS_376 0 -2.4275812550233797e-04
GC_5_377 b_5 NI_5 NS_377 0 6.5712946212068059e-05
GC_5_378 b_5 NI_5 NS_378 0 -2.8184590562941607e-05
GC_5_379 b_5 NI_5 NS_379 0 2.0799642420547330e-04
GC_5_380 b_5 NI_5 NS_380 0 -2.4122513466870739e-04
GC_5_381 b_5 NI_5 NS_381 0 -7.1069704680612887e-05
GC_5_382 b_5 NI_5 NS_382 0 -7.1882655589668043e-05
GC_5_383 b_5 NI_5 NS_383 0 6.4720730241308330e-05
GC_5_384 b_5 NI_5 NS_384 0 -7.5166912098191142e-05
GC_5_385 b_5 NI_5 NS_385 0 -1.7062494621390001e-04
GC_5_386 b_5 NI_5 NS_386 0 -1.8331083685746994e-04
GC_5_387 b_5 NI_5 NS_387 0 -4.8753414870632489e-05
GC_5_388 b_5 NI_5 NS_388 0 -1.9422271571646649e-05
GC_5_389 b_5 NI_5 NS_389 0 -1.4456137376859412e-04
GC_5_390 b_5 NI_5 NS_390 0 -9.5399246085555077e-05
GC_5_391 b_5 NI_5 NS_391 0 -2.7694032301989452e-05
GC_5_392 b_5 NI_5 NS_392 0 1.0380547760986706e-04
GC_5_393 b_5 NI_5 NS_393 0 -2.7258366804000391e-05
GC_5_394 b_5 NI_5 NS_394 0 1.3718071321635590e-05
GC_5_395 b_5 NI_5 NS_395 0 2.3543131378350768e-06
GC_5_396 b_5 NI_5 NS_396 0 5.0802585344004453e-05
GC_5_397 b_5 NI_5 NS_397 0 1.6821897885204081e-05
GC_5_398 b_5 NI_5 NS_398 0 -4.6940313873287393e-07
GC_5_399 b_5 NI_5 NS_399 0 1.7925272261788742e-06
GC_5_400 b_5 NI_5 NS_400 0 -1.5480347139603081e-05
GC_5_401 b_5 NI_5 NS_401 0 -1.4962445745700194e-05
GC_5_402 b_5 NI_5 NS_402 0 -1.3719794623046466e-05
GC_5_403 b_5 NI_5 NS_403 0 -1.2980299408039958e-05
GC_5_404 b_5 NI_5 NS_404 0 1.2291504479132230e-05
GC_5_405 b_5 NI_5 NS_405 0 7.7935023627879396e-06
GC_5_406 b_5 NI_5 NS_406 0 1.2794174910121825e-06
GC_5_407 b_5 NI_5 NS_407 0 -5.1334671787012359e-06
GC_5_408 b_5 NI_5 NS_408 0 -1.2739690923604260e-05
GC_5_409 b_5 NI_5 NS_409 0 -2.0684369734541903e-05
GC_5_410 b_5 NI_5 NS_410 0 -5.9679192317609380e-06
GC_5_411 b_5 NI_5 NS_411 0 1.1830376941256144e-06
GC_5_412 b_5 NI_5 NS_412 0 2.1729586492250424e-05
GC_5_413 b_5 NI_5 NS_413 0 1.2901795119742526e-05
GC_5_414 b_5 NI_5 NS_414 0 -6.8764806303115832e-06
GC_5_415 b_5 NI_5 NS_415 0 -1.7239595637413909e-05
GC_5_416 b_5 NI_5 NS_416 0 -1.6087364714276141e-05
GC_5_417 b_5 NI_5 NS_417 0 -2.7000608978044999e-05
GC_5_418 b_5 NI_5 NS_418 0 8.7818298756574216e-06
GC_5_419 b_5 NI_5 NS_419 0 2.7184780962946339e-05
GC_5_420 b_5 NI_5 NS_420 0 2.2283572700245568e-05
GC_5_421 b_5 NI_5 NS_421 0 1.1017158426387971e-05
GC_5_422 b_5 NI_5 NS_422 0 -2.1371410854884737e-05
GC_5_423 b_5 NI_5 NS_423 0 -3.0546772387422293e-05
GC_5_424 b_5 NI_5 NS_424 0 3.7146636540762667e-06
GC_5_425 b_5 NI_5 NS_425 0 -9.5336497222866023e-06
GC_5_426 b_5 NI_5 NS_426 0 3.9207841557037089e-05
GC_5_427 b_5 NI_5 NS_427 0 1.8462499023172459e-05
GC_5_428 b_5 NI_5 NS_428 0 -6.8326619094951935e-05
GC_5_429 b_5 NI_5 NS_429 0 4.3338401933859890e-05
GC_5_430 b_5 NI_5 NS_430 0 -1.7306939517286828e-05
GC_5_431 b_5 NI_5 NS_431 0 1.9831873059408375e-07
GC_5_432 b_5 NI_5 NS_432 0 -2.4930643171609978e-07
GC_5_433 b_5 NI_5 NS_433 0 -3.6889277615637413e-06
GC_5_434 b_5 NI_5 NS_434 0 -2.1088362104833448e-05
GC_5_435 b_5 NI_5 NS_435 0 -1.0619640304063651e-05
GC_5_436 b_5 NI_5 NS_436 0 1.6523074764138939e-05
GC_5_437 b_5 NI_5 NS_437 0 9.4073674995713897e-06
GC_5_438 b_5 NI_5 NS_438 0 3.1757020344530674e-05
GC_5_439 b_5 NI_5 NS_439 0 1.4489705540035967e-05
GC_5_440 b_5 NI_5 NS_440 0 -3.2770503922896179e-06
GC_5_441 b_5 NI_5 NS_441 0 -3.8741501656993795e-06
GC_5_442 b_5 NI_5 NS_442 0 1.2514849452734853e-05
GC_5_443 b_5 NI_5 NS_443 0 -1.8542557747690541e-05
GC_5_444 b_5 NI_5 NS_444 0 -3.5697562069741805e-06
GC_5_445 b_5 NI_5 NS_445 0 1.3189261521707815e-05
GC_5_446 b_5 NI_5 NS_446 0 1.3199109106000702e-05
GC_5_447 b_5 NI_5 NS_447 0 7.6293353077101078e-06
GC_5_448 b_5 NI_5 NS_448 0 -2.3004659568456430e-05
GC_5_449 b_5 NI_5 NS_449 0 -3.8543184738735028e-06
GC_5_450 b_5 NI_5 NS_450 0 -1.1714816045196064e-05
GC_5_451 b_5 NI_5 NS_451 0 -8.7383821882669537e-06
GC_5_452 b_5 NI_5 NS_452 0 -2.6220833191233551e-06
GC_5_453 b_5 NI_5 NS_453 0 5.5128509351889324e-10
GC_5_454 b_5 NI_5 NS_454 0 2.9325606221037022e-10
GC_5_455 b_5 NI_5 NS_455 0 4.2108228391939041e-08
GC_5_456 b_5 NI_5 NS_456 0 3.6979687973081052e-08
GC_5_457 b_5 NI_5 NS_457 0 -1.2879678365301597e-02
GC_5_458 b_5 NI_5 NS_458 0 1.3854981435520491e-03
GC_5_459 b_5 NI_5 NS_459 0 -2.6205840285934984e-07
GC_5_460 b_5 NI_5 NS_460 0 -3.7467072111586769e-06
GC_5_461 b_5 NI_5 NS_461 0 -2.6867049565005072e-04
GC_5_462 b_5 NI_5 NS_462 0 4.6434734670182794e-04
GC_5_463 b_5 NI_5 NS_463 0 1.3324560954779004e-03
GC_5_464 b_5 NI_5 NS_464 0 5.3750026552117352e-04
GC_5_465 b_5 NI_5 NS_465 0 -2.7601137799872538e-03
GC_5_466 b_5 NI_5 NS_466 0 -8.2597320623825881e-04
GC_5_467 b_5 NI_5 NS_467 0 3.5364628675814123e-03
GC_5_468 b_5 NI_5 NS_468 0 2.5065924206226289e-03
GC_5_469 b_5 NI_5 NS_469 0 1.1567034688187751e-03
GC_5_470 b_5 NI_5 NS_470 0 -4.2275310405896971e-03
GC_5_471 b_5 NI_5 NS_471 0 -1.7809488407363389e-03
GC_5_472 b_5 NI_5 NS_472 0 2.6938524756482214e-03
GC_5_473 b_5 NI_5 NS_473 0 -3.0415706679748621e-04
GC_5_474 b_5 NI_5 NS_474 0 -1.8023628353795466e-04
GC_5_475 b_5 NI_5 NS_475 0 3.9634827786397984e-03
GC_5_476 b_5 NI_5 NS_476 0 2.8124748378258722e-04
GC_5_477 b_5 NI_5 NS_477 0 -7.5491934513216650e-03
GC_5_478 b_5 NI_5 NS_478 0 -1.3596114662985673e-02
GC_5_479 b_5 NI_5 NS_479 0 4.4801853133997795e-03
GC_5_480 b_5 NI_5 NS_480 0 1.3516142075965857e-02
GC_5_481 b_5 NI_5 NS_481 0 6.6864812775844409e-03
GC_5_482 b_5 NI_5 NS_482 0 -4.0243778214441184e-03
GC_5_483 b_5 NI_5 NS_483 0 -1.3410293820584852e-02
GC_5_484 b_5 NI_5 NS_484 0 7.8159675612572514e-04
GC_5_485 b_5 NI_5 NS_485 0 7.8563490498532746e-03
GC_5_486 b_5 NI_5 NS_486 0 1.8570197805253192e-03
GC_5_487 b_5 NI_5 NS_487 0 1.0427284400920726e-02
GC_5_488 b_5 NI_5 NS_488 0 -1.9666894873981766e-02
GC_5_489 b_5 NI_5 NS_489 0 -1.7708792995197349e-02
GC_5_490 b_5 NI_5 NS_490 0 1.9274355532093498e-02
GC_5_491 b_5 NI_5 NS_491 0 7.6729375833858773e-03
GC_5_492 b_5 NI_5 NS_492 0 -1.4539279044187335e-03
GC_5_493 b_5 NI_5 NS_493 0 -1.5685667411793069e-02
GC_5_494 b_5 NI_5 NS_494 0 -4.6645856315018731e-03
GC_5_495 b_5 NI_5 NS_495 0 8.1074590720908602e-03
GC_5_496 b_5 NI_5 NS_496 0 7.2499065554861679e-03
GC_5_497 b_5 NI_5 NS_497 0 8.0870969212279171e-03
GC_5_498 b_5 NI_5 NS_498 0 -6.0421280239948104e-03
GC_5_499 b_5 NI_5 NS_499 0 -1.3963406797979248e-02
GC_5_500 b_5 NI_5 NS_500 0 4.6523180962944359e-03
GC_5_501 b_5 NI_5 NS_501 0 6.2461635398100186e-03
GC_5_502 b_5 NI_5 NS_502 0 2.3807834431025547e-03
GC_5_503 b_5 NI_5 NS_503 0 -6.3453822298407967e-03
GC_5_504 b_5 NI_5 NS_504 0 -1.1079792127784916e-02
GC_5_505 b_5 NI_5 NS_505 0 2.1863246186593064e-03
GC_5_506 b_5 NI_5 NS_506 0 1.1948129062760802e-02
GC_5_507 b_5 NI_5 NS_507 0 4.2064706907618977e-03
GC_5_508 b_5 NI_5 NS_508 0 -1.1782766738062396e-03
GC_5_509 b_5 NI_5 NS_509 0 -4.9335539115045891e-03
GC_5_510 b_5 NI_5 NS_510 0 1.0765974648072314e-03
GC_5_511 b_5 NI_5 NS_511 0 3.0283694698644160e-03
GC_5_512 b_5 NI_5 NS_512 0 6.9130860183737764e-04
GC_5_513 b_5 NI_5 NS_513 0 -2.2217202779697010e-03
GC_5_514 b_5 NI_5 NS_514 0 5.0249125625977391e-04
GC_5_515 b_5 NI_5 NS_515 0 3.0726777043806851e-03
GC_5_516 b_5 NI_5 NS_516 0 2.2985795667224531e-03
GC_5_517 b_5 NI_5 NS_517 0 -1.5387659365278651e-03
GC_5_518 b_5 NI_5 NS_518 0 -6.6609606018772484e-04
GC_5_519 b_5 NI_5 NS_519 0 1.8890921269302309e-03
GC_5_520 b_5 NI_5 NS_520 0 6.8214989017220163e-04
GC_5_521 b_5 NI_5 NS_521 0 -1.5634744905268954e-03
GC_5_522 b_5 NI_5 NS_522 0 1.2300996015769004e-03
GC_5_523 b_5 NI_5 NS_523 0 3.9777129314604431e-03
GC_5_524 b_5 NI_5 NS_524 0 1.4029334048311190e-03
GC_5_525 b_5 NI_5 NS_525 0 -1.5582664148642040e-03
GC_5_526 b_5 NI_5 NS_526 0 7.6117986197563422e-05
GC_5_527 b_5 NI_5 NS_527 0 2.8289093493877493e-03
GC_5_528 b_5 NI_5 NS_528 0 -6.8710722461222775e-04
GC_5_529 b_5 NI_5 NS_529 0 -1.8835386613865104e-03
GC_5_530 b_5 NI_5 NS_530 0 2.0120381834849905e-03
GC_5_531 b_5 NI_5 NS_531 0 4.9081291509083498e-03
GC_5_532 b_5 NI_5 NS_532 0 -1.8224322838858003e-04
GC_5_533 b_5 NI_5 NS_533 0 -1.6649329358349051e-03
GC_5_534 b_5 NI_5 NS_534 0 9.3127935402016456e-04
GC_5_535 b_5 NI_5 NS_535 0 3.0639848244447964e-03
GC_5_536 b_5 NI_5 NS_536 0 -2.8461931415289495e-03
GC_5_537 b_5 NI_5 NS_537 0 -1.4669285909372353e-03
GC_5_538 b_5 NI_5 NS_538 0 3.2252964315560369e-03
GC_5_539 b_5 NI_5 NS_539 0 3.7966903523395453e-03
GC_5_540 b_5 NI_5 NS_540 0 -2.9822010389922928e-03
GC_5_541 b_5 NI_5 NS_541 0 -1.8555106348092682e-03
GC_5_542 b_5 NI_5 NS_542 0 -3.8335466338367354e-03
GC_5_543 b_5 NI_5 NS_543 0 -4.1821452105082020e-04
GC_5_544 b_5 NI_5 NS_544 0 2.3792558667093044e-03
GC_5_545 b_5 NI_5 NS_545 0 -1.0537476773818887e-05
GC_5_546 b_5 NI_5 NS_546 0 -2.1101151456112947e-05
GC_5_547 b_5 NI_5 NS_547 0 8.3840691106312152e-04
GC_5_548 b_5 NI_5 NS_548 0 -3.7904942194838601e-03
GC_5_549 b_5 NI_5 NS_549 0 3.3771146867993685e-04
GC_5_550 b_5 NI_5 NS_550 0 3.3559401036911195e-03
GC_5_551 b_5 NI_5 NS_551 0 1.3516114980408969e-03
GC_5_552 b_5 NI_5 NS_552 0 -2.3818192054485521e-03
GC_5_553 b_5 NI_5 NS_553 0 2.1706665097638417e-03
GC_5_554 b_5 NI_5 NS_554 0 3.3305719674284269e-03
GC_5_555 b_5 NI_5 NS_555 0 1.1698297471202535e-03
GC_5_556 b_5 NI_5 NS_556 0 2.4039661728073787e-03
GC_5_557 b_5 NI_5 NS_557 0 -8.0769620187228397e-04
GC_5_558 b_5 NI_5 NS_558 0 -1.9803365764631633e-03
GC_5_559 b_5 NI_5 NS_559 0 3.9764634565270511e-04
GC_5_560 b_5 NI_5 NS_560 0 -2.6820418370232884e-03
GC_5_561 b_5 NI_5 NS_561 0 9.8318212604546007e-04
GC_5_562 b_5 NI_5 NS_562 0 2.7477883096377860e-03
GC_5_563 b_5 NI_5 NS_563 0 1.0389073299063309e-03
GC_5_564 b_5 NI_5 NS_564 0 -2.4201775721064485e-03
GC_5_565 b_5 NI_5 NS_565 0 -1.0840515955758212e-03
GC_5_566 b_5 NI_5 NS_566 0 1.5933774281620885e-03
GC_5_567 b_5 NI_5 NS_567 0 -1.0741032327266180e-08
GC_5_568 b_5 NI_5 NS_568 0 -2.7692023162286639e-09
GC_5_569 b_5 NI_5 NS_569 0 2.2912277515833352e-06
GC_5_570 b_5 NI_5 NS_570 0 5.4762400252556837e-07
GC_5_571 b_5 NI_5 NS_571 0 1.8114258402846400e-02
GC_5_572 b_5 NI_5 NS_572 0 6.7504951698033420e-03
GC_5_573 b_5 NI_5 NS_573 0 4.7195340056744647e-07
GC_5_574 b_5 NI_5 NS_574 0 1.4474465807824860e-06
GC_5_575 b_5 NI_5 NS_575 0 6.0855591319528462e-03
GC_5_576 b_5 NI_5 NS_576 0 1.8096362281391216e-03
GC_5_577 b_5 NI_5 NS_577 0 -6.0720623110209820e-03
GC_5_578 b_5 NI_5 NS_578 0 -6.1691308988263776e-04
GC_5_579 b_5 NI_5 NS_579 0 7.3059555360108020e-03
GC_5_580 b_5 NI_5 NS_580 0 -1.2857318021597862e-02
GC_5_581 b_5 NI_5 NS_581 0 8.4528525370748623e-03
GC_5_582 b_5 NI_5 NS_582 0 -2.4020868258508297e-04
GC_5_583 b_5 NI_5 NS_583 0 -9.6390275735754073e-03
GC_5_584 b_5 NI_5 NS_584 0 2.6170726232826115e-03
GC_5_585 b_5 NI_5 NS_585 0 -8.8462056541014373e-03
GC_5_586 b_5 NI_5 NS_586 0 -2.4392927000882001e-02
GC_5_587 b_5 NI_5 NS_587 0 -8.6515245608362996e-04
GC_5_588 b_5 NI_5 NS_588 0 4.1785645919016961e-03
GC_5_589 b_5 NI_5 NS_589 0 7.1897514053148454e-03
GC_5_590 b_5 NI_5 NS_590 0 -1.0341204426173314e-03
GC_5_591 b_5 NI_5 NS_591 0 -2.5138615464278230e-02
GC_5_592 b_5 NI_5 NS_592 0 4.8070754375990092e-03
GC_5_593 b_5 NI_5 NS_593 0 -1.9701023618046206e-02
GC_5_594 b_5 NI_5 NS_594 0 8.9743269243009718e-04
GC_5_595 b_5 NI_5 NS_595 0 1.0752501538270114e-02
GC_5_596 b_5 NI_5 NS_596 0 -2.7940137750917427e-03
GC_5_597 b_5 NI_5 NS_597 0 -4.8191051631670794e-03
GC_5_598 b_5 NI_5 NS_598 0 4.5027471493287237e-02
GC_5_599 b_5 NI_5 NS_599 0 -1.2658611388374765e-02
GC_5_600 b_5 NI_5 NS_600 0 -2.5617083899007219e-04
GC_5_601 b_5 NI_5 NS_601 0 1.5863256622517877e-02
GC_5_602 b_5 NI_5 NS_602 0 -4.0664539102301172e-03
GC_5_603 b_5 NI_5 NS_603 0 3.2252268012760092e-02
GC_5_604 b_5 NI_5 NS_604 0 1.8644568960926922e-02
GC_5_605 b_5 NI_5 NS_605 0 -1.2591689410895376e-02
GC_5_606 b_5 NI_5 NS_606 0 1.8232239084040738e-04
GC_5_607 b_5 NI_5 NS_607 0 1.7239501216885215e-02
GC_5_608 b_5 NI_5 NS_608 0 -3.5124355464666850e-02
GC_5_609 b_5 NI_5 NS_609 0 1.4036151259632836e-02
GC_5_610 b_5 NI_5 NS_610 0 4.7591218063493387e-03
GC_5_611 b_5 NI_5 NS_611 0 -1.4382232004487865e-02
GC_5_612 b_5 NI_5 NS_612 0 2.6525514398366158e-04
GC_5_613 b_5 NI_5 NS_613 0 -2.0118038005669241e-02
GC_5_614 b_5 NI_5 NS_614 0 -3.0219184026285206e-02
GC_5_615 b_5 NI_5 NS_615 0 1.0538961572883945e-02
GC_5_616 b_5 NI_5 NS_616 0 3.5722907153827124e-03
GC_5_617 b_5 NI_5 NS_617 0 -2.6760787019281366e-02
GC_5_618 b_5 NI_5 NS_618 0 1.1130945875216795e-02
GC_5_619 b_5 NI_5 NS_619 0 -1.4164601789999351e-02
GC_5_620 b_5 NI_5 NS_620 0 -2.5194349481183899e-03
GC_5_621 b_5 NI_5 NS_621 0 7.5549379428175552e-03
GC_5_622 b_5 NI_5 NS_622 0 1.5797730028683924e-03
GC_5_623 b_5 NI_5 NS_623 0 -8.4943321279293792e-04
GC_5_624 b_5 NI_5 NS_624 0 2.4400445484638173e-02
GC_5_625 b_5 NI_5 NS_625 0 -7.6205599928682510e-03
GC_5_626 b_5 NI_5 NS_626 0 2.8886133180202218e-04
GC_5_627 b_5 NI_5 NS_627 0 -5.5962845643326656e-04
GC_5_628 b_5 NI_5 NS_628 0 -5.5377893651042545e-03
GC_5_629 b_5 NI_5 NS_629 0 8.2746286078645669e-03
GC_5_630 b_5 NI_5 NS_630 0 7.0134869144217868e-03
GC_5_631 b_5 NI_5 NS_631 0 -7.1244776235215889e-04
GC_5_632 b_5 NI_5 NS_632 0 1.2089354891046790e-02
GC_5_633 b_5 NI_5 NS_633 0 -5.1470154056105690e-03
GC_5_634 b_5 NI_5 NS_634 0 -1.3515142215502854e-04
GC_5_635 b_5 NI_5 NS_635 0 -1.8292841011720048e-03
GC_5_636 b_5 NI_5 NS_636 0 -5.1716269492733313e-03
GC_5_637 b_5 NI_5 NS_637 0 9.2942858406233082e-03
GC_5_638 b_5 NI_5 NS_638 0 5.4122740160823758e-03
GC_5_639 b_5 NI_5 NS_639 0 3.5222366912643840e-03
GC_5_640 b_5 NI_5 NS_640 0 1.1687382974279023e-02
GC_5_641 b_5 NI_5 NS_641 0 -6.1347983956874259e-03
GC_5_642 b_5 NI_5 NS_642 0 1.4299471280256198e-03
GC_5_643 b_5 NI_5 NS_643 0 -2.8132859417070717e-03
GC_5_644 b_5 NI_5 NS_644 0 -7.3475993413127539e-03
GC_5_645 b_5 NI_5 NS_645 0 9.9612567433730505e-03
GC_5_646 b_5 NI_5 NS_646 0 3.3711874885421055e-03
GC_5_647 b_5 NI_5 NS_647 0 8.1789449275024868e-03
GC_5_648 b_5 NI_5 NS_648 0 1.0242403639163787e-02
GC_5_649 b_5 NI_5 NS_649 0 -6.9808965547235886e-03
GC_5_650 b_5 NI_5 NS_650 0 2.9381657992600140e-03
GC_5_651 b_5 NI_5 NS_651 0 -5.6228415414615847e-03
GC_5_652 b_5 NI_5 NS_652 0 -8.0956784923397595e-03
GC_5_653 b_5 NI_5 NS_653 0 9.8673033766100444e-03
GC_5_654 b_5 NI_5 NS_654 0 5.6094095416818512e-04
GC_5_655 b_5 NI_5 NS_655 0 -1.0918399761574738e-02
GC_5_656 b_5 NI_5 NS_656 0 1.2173665240499501e-02
GC_5_657 b_5 NI_5 NS_657 0 9.6705985847331030e-03
GC_5_658 b_5 NI_5 NS_658 0 5.0264728403737980e-03
GC_5_659 b_5 NI_5 NS_659 0 -1.9577767983728558e-05
GC_5_660 b_5 NI_5 NS_660 0 3.1186857979205405e-05
GC_5_661 b_5 NI_5 NS_661 0 -7.1178131165468414e-03
GC_5_662 b_5 NI_5 NS_662 0 4.4750771610104403e-03
GC_5_663 b_5 NI_5 NS_663 0 -7.6632721047214351e-03
GC_5_664 b_5 NI_5 NS_664 0 -5.3302256448546368e-03
GC_5_665 b_5 NI_5 NS_665 0 9.5221928859994445e-03
GC_5_666 b_5 NI_5 NS_666 0 -1.7151705510902338e-03
GC_5_667 b_5 NI_5 NS_667 0 1.2490583078224570e-02
GC_5_668 b_5 NI_5 NS_668 0 -1.3742793297989513e-03
GC_5_669 b_5 NI_5 NS_669 0 -5.0725007265825855e-03
GC_5_670 b_5 NI_5 NS_670 0 -2.7519124370864669e-03
GC_5_671 b_5 NI_5 NS_671 0 -2.2328915677616262e-03
GC_5_672 b_5 NI_5 NS_672 0 6.6013356482994088e-03
GC_5_673 b_5 NI_5 NS_673 0 8.9595363600226009e-03
GC_5_674 b_5 NI_5 NS_674 0 1.2928959390184506e-04
GC_5_675 b_5 NI_5 NS_675 0 1.2486928460366045e-02
GC_5_676 b_5 NI_5 NS_676 0 1.7755709829021036e-03
GC_5_677 b_5 NI_5 NS_677 0 -5.3764539858590461e-03
GC_5_678 b_5 NI_5 NS_678 0 4.1567506691064559e-03
GC_5_679 b_5 NI_5 NS_679 0 -1.8433718942024752e-03
GC_5_680 b_5 NI_5 NS_680 0 -5.6868607242641575e-03
GC_5_681 b_5 NI_5 NS_681 0 2.0788380545382222e-07
GC_5_682 b_5 NI_5 NS_682 0 -2.4508480559808222e-07
GC_5_683 b_5 NI_5 NS_683 0 -1.1508311415294919e-05
GC_5_684 b_5 NI_5 NS_684 0 1.8247242434575860e-05
GC_5_685 b_5 NI_5 NS_685 0 7.9886735401539961e-03
GC_5_686 b_5 NI_5 NS_686 0 -1.6009906166397658e-03
GC_5_687 b_5 NI_5 NS_687 0 -1.2329825440166125e-08
GC_5_688 b_5 NI_5 NS_688 0 -8.8365943175870924e-07
GC_5_689 b_5 NI_5 NS_689 0 1.0714030449892067e-04
GC_5_690 b_5 NI_5 NS_690 0 -5.1251764245795466e-04
GC_5_691 b_5 NI_5 NS_691 0 -1.9321159778792280e-03
GC_5_692 b_5 NI_5 NS_692 0 -5.9631983963332900e-04
GC_5_693 b_5 NI_5 NS_693 0 2.9522606672808525e-03
GC_5_694 b_5 NI_5 NS_694 0 2.2413638503497248e-03
GC_5_695 b_5 NI_5 NS_695 0 -3.5853190594994527e-03
GC_5_696 b_5 NI_5 NS_696 0 -3.0463421382723442e-03
GC_5_697 b_5 NI_5 NS_697 0 -1.6953791407142052e-03
GC_5_698 b_5 NI_5 NS_698 0 5.8334391390082027e-03
GC_5_699 b_5 NI_5 NS_699 0 4.3284002291638073e-03
GC_5_700 b_5 NI_5 NS_700 0 -2.4949667614127106e-03
GC_5_701 b_5 NI_5 NS_701 0 -1.0252446936248555e-04
GC_5_702 b_5 NI_5 NS_702 0 -9.7511075161820095e-05
GC_5_703 b_5 NI_5 NS_703 0 -4.4595020428925929e-03
GC_5_704 b_5 NI_5 NS_704 0 -9.0945608091203944e-04
GC_5_705 b_5 NI_5 NS_705 0 9.1489028587241408e-03
GC_5_706 b_5 NI_5 NS_706 0 1.7749052989247376e-02
GC_5_707 b_5 NI_5 NS_707 0 -4.0759927667455252e-03
GC_5_708 b_5 NI_5 NS_708 0 -1.7815995532837223e-02
GC_5_709 b_5 NI_5 NS_709 0 -8.2086051829402401e-03
GC_5_710 b_5 NI_5 NS_710 0 4.1974762820249393e-03
GC_5_711 b_5 NI_5 NS_711 0 1.7045924966324170e-02
GC_5_712 b_5 NI_5 NS_712 0 -4.7587338128305448e-04
GC_5_713 b_5 NI_5 NS_713 0 -9.2871624819418352e-03
GC_5_714 b_5 NI_5 NS_714 0 -3.1746354546416406e-03
GC_5_715 b_5 NI_5 NS_715 0 -1.3650848379647919e-02
GC_5_716 b_5 NI_5 NS_716 0 2.2873425818299549e-02
GC_5_717 b_5 NI_5 NS_717 0 2.2768614588535702e-02
GC_5_718 b_5 NI_5 NS_718 0 -2.2718063915562001e-02
GC_5_719 b_5 NI_5 NS_719 0 -9.2369617939143181e-03
GC_5_720 b_5 NI_5 NS_720 0 9.4042656214539378e-04
GC_5_721 b_5 NI_5 NS_721 0 1.8496822276860714e-02
GC_5_722 b_5 NI_5 NS_722 0 6.1966535518119909e-03
GC_5_723 b_5 NI_5 NS_723 0 -9.2042288301689163e-03
GC_5_724 b_5 NI_5 NS_724 0 -9.4288118152042657e-03
GC_5_725 b_5 NI_5 NS_725 0 -9.9569355470869123e-03
GC_5_726 b_5 NI_5 NS_726 0 6.4309792448890958e-03
GC_5_727 b_5 NI_5 NS_727 0 1.6827172974901664e-02
GC_5_728 b_5 NI_5 NS_728 0 -4.8950434243071172e-03
GC_5_729 b_5 NI_5 NS_729 0 -7.2263300358184823e-03
GC_5_730 b_5 NI_5 NS_730 0 -3.3851923587828758e-03
GC_5_731 b_5 NI_5 NS_731 0 6.8657296048918112e-03
GC_5_732 b_5 NI_5 NS_732 0 1.3286490716233919e-02
GC_5_733 b_5 NI_5 NS_733 0 -1.8581881524139161e-03
GC_5_734 b_5 NI_5 NS_734 0 -1.4397044103065635e-02
GC_5_735 b_5 NI_5 NS_735 0 -4.9859100078895732e-03
GC_5_736 b_5 NI_5 NS_736 0 1.0545183375540890e-03
GC_5_737 b_5 NI_5 NS_737 0 6.0007407101906390e-03
GC_5_738 b_5 NI_5 NS_738 0 -1.1126545345610764e-03
GC_5_739 b_5 NI_5 NS_739 0 -3.4683253119721469e-03
GC_5_740 b_5 NI_5 NS_740 0 -1.0780499297876050e-03
GC_5_741 b_5 NI_5 NS_741 0 2.7173467373079723e-03
GC_5_742 b_5 NI_5 NS_742 0 -5.1095685632514222e-04
GC_5_743 b_5 NI_5 NS_743 0 -3.3053412635033136e-03
GC_5_744 b_5 NI_5 NS_744 0 -2.8885150366898121e-03
GC_5_745 b_5 NI_5 NS_745 0 2.0156340107862010e-03
GC_5_746 b_5 NI_5 NS_746 0 7.7768289509255598e-04
GC_5_747 b_5 NI_5 NS_747 0 -2.0192451153385770e-03
GC_5_748 b_5 NI_5 NS_748 0 -9.6218739425117845e-04
GC_5_749 b_5 NI_5 NS_749 0 2.1198804231875317e-03
GC_5_750 b_5 NI_5 NS_750 0 -1.4705676215787074e-03
GC_5_751 b_5 NI_5 NS_751 0 -4.1910213514369625e-03
GC_5_752 b_5 NI_5 NS_752 0 -1.8092507177206196e-03
GC_5_753 b_5 NI_5 NS_753 0 2.3672939645781980e-03
GC_5_754 b_5 NI_5 NS_754 0 -3.6739647747752277e-04
GC_5_755 b_5 NI_5 NS_755 0 -3.0199644114831635e-03
GC_5_756 b_5 NI_5 NS_756 0 4.6494721848137162e-04
GC_5_757 b_5 NI_5 NS_757 0 2.7038550448384218e-03
GC_5_758 b_5 NI_5 NS_758 0 -2.7263252341181601e-03
GC_5_759 b_5 NI_5 NS_759 0 -5.0450291902992333e-03
GC_5_760 b_5 NI_5 NS_760 0 -1.2988615164204683e-04
GC_5_761 b_5 NI_5 NS_761 0 2.4275289845229501e-03
GC_5_762 b_5 NI_5 NS_762 0 -2.1667278442961120e-03
GC_5_763 b_5 NI_5 NS_763 0 -3.2524101995311627e-03
GC_5_764 b_5 NI_5 NS_764 0 2.6001223086795124e-03
GC_5_765 b_5 NI_5 NS_765 0 1.7373702900374262e-03
GC_5_766 b_5 NI_5 NS_766 0 -4.7433399597032379e-03
GC_5_767 b_5 NI_5 NS_767 0 -3.6476875627013731e-03
GC_5_768 b_5 NI_5 NS_768 0 2.5904971150401972e-03
GC_5_769 b_5 NI_5 NS_769 0 -2.8140500630920114e-03
GC_5_770 b_5 NI_5 NS_770 0 4.0553536026503049e-03
GC_5_771 b_5 NI_5 NS_771 0 -2.3077988955524218e-04
GC_5_772 b_5 NI_5 NS_772 0 -4.1951359845031145e-03
GC_5_773 b_5 NI_5 NS_773 0 -9.8757619543563190e-06
GC_5_774 b_5 NI_5 NS_774 0 7.9025157468606561e-06
GC_5_775 b_5 NI_5 NS_775 0 -1.3634151899027619e-03
GC_5_776 b_5 NI_5 NS_776 0 3.3837800922319919e-03
GC_5_777 b_5 NI_5 NS_777 0 -9.6978191554016090e-04
GC_5_778 b_5 NI_5 NS_778 0 -4.3384320358366016e-03
GC_5_779 b_5 NI_5 NS_779 0 -1.0095576378297832e-03
GC_5_780 b_5 NI_5 NS_780 0 2.2144692442646161e-03
GC_5_781 b_5 NI_5 NS_781 0 -1.6625797627074141e-03
GC_5_782 b_5 NI_5 NS_782 0 -4.4181655731749944e-03
GC_5_783 b_5 NI_5 NS_783 0 -1.4450239250894132e-03
GC_5_784 b_5 NI_5 NS_784 0 -2.4969806516489555e-03
GC_5_785 b_5 NI_5 NS_785 0 7.8582137584433766e-04
GC_5_786 b_5 NI_5 NS_786 0 2.5922239207891900e-03
GC_5_787 b_5 NI_5 NS_787 0 -6.9658839234052426e-04
GC_5_788 b_5 NI_5 NS_788 0 2.8805416794975814e-03
GC_5_789 b_5 NI_5 NS_789 0 -1.4341252988649927e-03
GC_5_790 b_5 NI_5 NS_790 0 -2.7701138494934897e-03
GC_5_791 b_5 NI_5 NS_791 0 -1.1685605982718714e-03
GC_5_792 b_5 NI_5 NS_792 0 2.6674409195710422e-03
GC_5_793 b_5 NI_5 NS_793 0 7.8095042474653166e-04
GC_5_794 b_5 NI_5 NS_794 0 -1.8732339630859263e-03
GC_5_795 b_5 NI_5 NS_795 0 2.4009828617971256e-08
GC_5_796 b_5 NI_5 NS_796 0 -6.0310105244334038e-08
GC_5_797 b_5 NI_5 NS_797 0 -9.0615469967058698e-07
GC_5_798 b_5 NI_5 NS_798 0 3.2140038270567072e-06
GC_5_799 b_5 NI_5 NS_799 0 3.0950443039044285e-03
GC_5_800 b_5 NI_5 NS_800 0 -6.1289418580224241e-04
GC_5_801 b_5 NI_5 NS_801 0 2.8121770033646162e-08
GC_5_802 b_5 NI_5 NS_802 0 -3.1528708115044329e-08
GC_5_803 b_5 NI_5 NS_803 0 2.0500773518833767e-04
GC_5_804 b_5 NI_5 NS_804 0 1.3546540150003835e-04
GC_5_805 b_5 NI_5 NS_805 0 5.6415263432640559e-04
GC_5_806 b_5 NI_5 NS_806 0 2.6382413732436175e-04
GC_5_807 b_5 NI_5 NS_807 0 3.0949151581973894e-03
GC_5_808 b_5 NI_5 NS_808 0 -2.2211775604445844e-03
GC_5_809 b_5 NI_5 NS_809 0 -1.5948050014524433e-03
GC_5_810 b_5 NI_5 NS_810 0 -2.6831568741263762e-03
GC_5_811 b_5 NI_5 NS_811 0 -2.0664405331187320e-03
GC_5_812 b_5 NI_5 NS_812 0 -3.7810168675206229e-03
GC_5_813 b_5 NI_5 NS_813 0 -4.9930248634699722e-03
GC_5_814 b_5 NI_5 NS_814 0 -1.5154929334807925e-03
GC_5_815 b_5 NI_5 NS_815 0 2.9714197086706107e-04
GC_5_816 b_5 NI_5 NS_816 0 1.9409424577538048e-04
GC_5_817 b_5 NI_5 NS_817 0 -2.8708432797730343e-03
GC_5_818 b_5 NI_5 NS_818 0 -9.4557935833778273e-04
GC_5_819 b_5 NI_5 NS_819 0 -2.2198356447053348e-02
GC_5_820 b_5 NI_5 NS_820 0 -1.0125161759749575e-02
GC_5_821 b_5 NI_5 NS_821 0 1.2231803926555148e-03
GC_5_822 b_5 NI_5 NS_822 0 2.0396448916398541e-02
GC_5_823 b_5 NI_5 NS_823 0 -5.8225964770082890e-03
GC_5_824 b_5 NI_5 NS_824 0 4.6364311842683643e-03
GC_5_825 b_5 NI_5 NS_825 0 5.8808187604699330e-03
GC_5_826 b_5 NI_5 NS_826 0 3.4493744000981631e-02
GC_5_827 b_5 NI_5 NS_827 0 8.0480772487816210e-03
GC_5_828 b_5 NI_5 NS_828 0 2.7589349738089968e-03
GC_5_829 b_5 NI_5 NS_829 0 -7.6367957292518465e-03
GC_5_830 b_5 NI_5 NS_830 0 2.9591949312289638e-02
GC_5_831 b_5 NI_5 NS_831 0 5.0679464963455052e-02
GC_5_832 b_5 NI_5 NS_832 0 -2.0315740117315708e-02
GC_5_833 b_5 NI_5 NS_833 0 7.9122592807459834e-03
GC_5_834 b_5 NI_5 NS_834 0 -1.6718962441294412e-03
GC_5_835 b_5 NI_5 NS_835 0 2.8952184632050501e-02
GC_5_836 b_5 NI_5 NS_836 0 -2.6605126129145541e-02
GC_5_837 b_5 NI_5 NS_837 0 -6.7717822711924110e-03
GC_5_838 b_5 NI_5 NS_838 0 -9.8521000534942012e-03
GC_5_839 b_5 NI_5 NS_839 0 8.4245547478698328e-03
GC_5_840 b_5 NI_5 NS_840 0 -8.0661005364070764e-03
GC_5_841 b_5 NI_5 NS_841 0 -1.9120467240054891e-02
GC_5_842 b_5 NI_5 NS_842 0 -2.5143595149441110e-02
GC_5_843 b_5 NI_5 NS_843 0 -5.4851138495895712e-03
GC_5_844 b_5 NI_5 NS_844 0 -2.8303874863051717e-03
GC_5_845 b_5 NI_5 NS_845 0 -1.7803813202940711e-02
GC_5_846 b_5 NI_5 NS_846 0 -1.3047348683002650e-02
GC_5_847 b_5 NI_5 NS_847 0 -4.7610274665251225e-03
GC_5_848 b_5 NI_5 NS_848 0 1.2568312185923518e-02
GC_5_849 b_5 NI_5 NS_849 0 -3.4539895313030031e-03
GC_5_850 b_5 NI_5 NS_850 0 1.5560260582215127e-03
GC_5_851 b_5 NI_5 NS_851 0 -6.8744300317368163e-04
GC_5_852 b_5 NI_5 NS_852 0 7.0157646284252813e-03
GC_5_853 b_5 NI_5 NS_853 0 1.8840812973413546e-03
GC_5_854 b_5 NI_5 NS_854 0 8.1060422559650478e-05
GC_5_855 b_5 NI_5 NS_855 0 3.0821856981076473e-04
GC_5_856 b_5 NI_5 NS_856 0 -1.9474452509138213e-03
GC_5_857 b_5 NI_5 NS_857 0 -1.8615158810871963e-03
GC_5_858 b_5 NI_5 NS_858 0 -1.6133456384919559e-03
GC_5_859 b_5 NI_5 NS_859 0 -2.1255689792494146e-03
GC_5_860 b_5 NI_5 NS_860 0 1.6940535978505788e-03
GC_5_861 b_5 NI_5 NS_861 0 7.6441486732342948e-04
GC_5_862 b_5 NI_5 NS_862 0 1.8569487132465409e-04
GC_5_863 b_5 NI_5 NS_863 0 -7.0068912680603475e-04
GC_5_864 b_5 NI_5 NS_864 0 -1.6760054888967197e-03
GC_5_865 b_5 NI_5 NS_865 0 -2.6855352097078546e-03
GC_5_866 b_5 NI_5 NS_866 0 -8.2394391564054239e-04
GC_5_867 b_5 NI_5 NS_867 0 -4.9849900907188009e-04
GC_5_868 b_5 NI_5 NS_868 0 2.9352188056097979e-03
GC_5_869 b_5 NI_5 NS_869 0 1.3528909986814043e-03
GC_5_870 b_5 NI_5 NS_870 0 -8.5706936164413089e-04
GC_5_871 b_5 NI_5 NS_871 0 -2.4223433396979980e-03
GC_5_872 b_5 NI_5 NS_872 0 -2.2652834660473104e-03
GC_5_873 b_5 NI_5 NS_873 0 -3.5590211421404334e-03
GC_5_874 b_5 NI_5 NS_874 0 7.4879944697761841e-04
GC_5_875 b_5 NI_5 NS_875 0 2.4605502113730074e-03
GC_5_876 b_5 NI_5 NS_876 0 3.0265645535254432e-03
GC_5_877 b_5 NI_5 NS_877 0 9.8335647735160693e-04
GC_5_878 b_5 NI_5 NS_878 0 -2.9400791209097769e-03
GC_5_879 b_5 NI_5 NS_879 0 -4.7724967855482144e-03
GC_5_880 b_5 NI_5 NS_880 0 5.7213633240375327e-05
GC_5_881 b_5 NI_5 NS_881 0 -1.7194839081914200e-03
GC_5_882 b_5 NI_5 NS_882 0 3.7113727614766913e-03
GC_5_883 b_5 NI_5 NS_883 0 -7.3866508540143636e-04
GC_5_884 b_5 NI_5 NS_884 0 1.5326963597250491e-03
GC_5_885 b_5 NI_5 NS_885 0 3.2195727075057753e-03
GC_5_886 b_5 NI_5 NS_886 0 -1.3349985164818761e-03
GC_5_887 b_5 NI_5 NS_887 0 -2.8022748169909112e-06
GC_5_888 b_5 NI_5 NS_888 0 8.9859889224592073e-06
GC_5_889 b_5 NI_5 NS_889 0 -1.8210613133963940e-03
GC_5_890 b_5 NI_5 NS_890 0 -2.5224003647436504e-03
GC_5_891 b_5 NI_5 NS_891 0 -2.4088301534687605e-03
GC_5_892 b_5 NI_5 NS_892 0 2.4933225713162236e-03
GC_5_893 b_5 NI_5 NS_893 0 1.0059037156700753e-03
GC_5_894 b_5 NI_5 NS_894 0 2.4239841643900967e-03
GC_5_895 b_5 NI_5 NS_895 0 8.4854726496080965e-04
GC_5_896 b_5 NI_5 NS_896 0 -2.6997865571465672e-03
GC_5_897 b_5 NI_5 NS_897 0 -3.0628339988005270e-04
GC_5_898 b_5 NI_5 NS_898 0 1.6736613633905092e-03
GC_5_899 b_5 NI_5 NS_899 0 -1.7824227291375022e-03
GC_5_900 b_5 NI_5 NS_900 0 -3.1430320046740709e-04
GC_5_901 b_5 NI_5 NS_901 0 1.3997488472937071e-03
GC_5_902 b_5 NI_5 NS_902 0 1.9719385380328621e-03
GC_5_903 b_5 NI_5 NS_903 0 1.0457174698470955e-03
GC_5_904 b_5 NI_5 NS_904 0 -2.2988262163664056e-03
GC_5_905 b_5 NI_5 NS_905 0 -6.9831747332173755e-04
GC_5_906 b_5 NI_5 NS_906 0 -1.4663462689947933e-03
GC_5_907 b_5 NI_5 NS_907 0 -1.3735955654334605e-03
GC_5_908 b_5 NI_5 NS_908 0 -3.1257035676522654e-04
GC_5_909 b_5 NI_5 NS_909 0 6.7938444069209254e-09
GC_5_910 b_5 NI_5 NS_910 0 -2.4700012010235619e-08
GC_5_911 b_5 NI_5 NS_911 0 -4.4377037392376030e-07
GC_5_912 b_5 NI_5 NS_912 0 1.6205767026264488e-06
GC_5_913 b_5 NI_5 NS_913 0 -1.1776549591928312e-04
GC_5_914 b_5 NI_5 NS_914 0 -2.1390371269946564e-06
GC_5_915 b_5 NI_5 NS_915 0 -2.5034434674381663e-10
GC_5_916 b_5 NI_5 NS_916 0 2.5994089614998970e-09
GC_5_917 b_5 NI_5 NS_917 0 1.6865027226507712e-06
GC_5_918 b_5 NI_5 NS_918 0 -1.5557518856712656e-06
GC_5_919 b_5 NI_5 NS_919 0 1.0498575692869478e-07
GC_5_920 b_5 NI_5 NS_920 0 -6.3346749680079760e-06
GC_5_921 b_5 NI_5 NS_921 0 -7.5924898800446669e-06
GC_5_922 b_5 NI_5 NS_922 0 2.3113153394570403e-07
GC_5_923 b_5 NI_5 NS_923 0 -1.1742330524623065e-06
GC_5_924 b_5 NI_5 NS_924 0 -4.6213210382682761e-06
GC_5_925 b_5 NI_5 NS_925 0 -1.5831640424530069e-05
GC_5_926 b_5 NI_5 NS_926 0 -1.5727952804796183e-06
GC_5_927 b_5 NI_5 NS_927 0 -6.0025257209218105e-06
GC_5_928 b_5 NI_5 NS_928 0 1.9095124188389721e-05
GC_5_929 b_5 NI_5 NS_929 0 4.6272150845831564e-06
GC_5_930 b_5 NI_5 NS_930 0 -3.0068106352501850e-06
GC_5_931 b_5 NI_5 NS_931 0 -1.4071656231230598e-08
GC_5_932 b_5 NI_5 NS_932 0 -2.6089082199603210e-06
GC_5_933 b_5 NI_5 NS_933 0 -2.5759906133282627e-05
GC_5_934 b_5 NI_5 NS_934 0 2.8490203973359023e-05
GC_5_935 b_5 NI_5 NS_935 0 2.8211387952909081e-05
GC_5_936 b_5 NI_5 NS_936 0 -8.6038967430501355e-06
GC_5_937 b_5 NI_5 NS_937 0 -8.0514516540375236e-06
GC_5_938 b_5 NI_5 NS_938 0 -4.3168391464409647e-06
GC_5_939 b_5 NI_5 NS_939 0 1.2692845785897475e-05
GC_5_940 b_5 NI_5 NS_940 0 2.6907359924712740e-05
GC_5_941 b_5 NI_5 NS_941 0 1.4541619223224465e-06
GC_5_942 b_5 NI_5 NS_942 0 -9.0171639978094192e-06
GC_5_943 b_5 NI_5 NS_943 0 -2.8297054977549664e-05
GC_5_944 b_5 NI_5 NS_944 0 4.7690830141018034e-06
GC_5_945 b_5 NI_5 NS_945 0 4.1340035815588038e-05
GC_5_946 b_5 NI_5 NS_946 0 1.0566874561950401e-05
GC_5_947 b_5 NI_5 NS_947 0 -2.9777178666927519e-06
GC_5_948 b_5 NI_5 NS_948 0 -4.5076723818426569e-06
GC_5_949 b_5 NI_5 NS_949 0 1.2968809920551739e-05
GC_5_950 b_5 NI_5 NS_950 0 1.8946404935504972e-05
GC_5_951 b_5 NI_5 NS_951 0 3.7956311228151309e-06
GC_5_952 b_5 NI_5 NS_952 0 -1.0952540284156567e-05
GC_5_953 b_5 NI_5 NS_953 0 -6.4190508555728198e-06
GC_5_954 b_5 NI_5 NS_954 0 8.3208938784613327e-07
GC_5_955 b_5 NI_5 NS_955 0 1.8890181496748065e-05
GC_5_956 b_5 NI_5 NS_956 0 5.3956719892357994e-06
GC_5_957 b_5 NI_5 NS_957 0 -7.6255255116911023e-08
GC_5_958 b_5 NI_5 NS_958 0 -4.2077103387018934e-06
GC_5_959 b_5 NI_5 NS_959 0 4.9306586447886220e-06
GC_5_960 b_5 NI_5 NS_960 0 1.4263142659157418e-05
GC_5_961 b_5 NI_5 NS_961 0 7.8225223554032850e-06
GC_5_962 b_5 NI_5 NS_962 0 -1.1202027477536485e-05
GC_5_963 b_5 NI_5 NS_963 0 -1.3847720853419338e-06
GC_5_964 b_5 NI_5 NS_964 0 9.2712256644826868e-07
GC_5_965 b_5 NI_5 NS_965 0 1.0915581787092155e-05
GC_5_966 b_5 NI_5 NS_966 0 4.0962629112943040e-06
GC_5_967 b_5 NI_5 NS_967 0 1.7204805700690176e-06
GC_5_968 b_5 NI_5 NS_968 0 -6.4492682011602175e-07
GC_5_969 b_5 NI_5 NS_969 0 5.6901265197405576e-06
GC_5_970 b_5 NI_5 NS_970 0 1.6919136190886240e-06
GC_5_971 b_5 NI_5 NS_971 0 3.4275668880499552e-06
GC_5_972 b_5 NI_5 NS_972 0 2.0300854192408932e-06
GC_5_973 b_5 NI_5 NS_973 0 1.0987680938791757e-05
GC_5_974 b_5 NI_5 NS_974 0 3.7699913596919395e-06
GC_5_975 b_5 NI_5 NS_975 0 4.8689033070844224e-06
GC_5_976 b_5 NI_5 NS_976 0 -9.2939663285077785e-08
GC_5_977 b_5 NI_5 NS_977 0 9.9989117972311659e-06
GC_5_978 b_5 NI_5 NS_978 0 -1.0950576695233314e-06
GC_5_979 b_5 NI_5 NS_979 0 8.2824376152807909e-06
GC_5_980 b_5 NI_5 NS_980 0 2.9417405406590215e-06
GC_5_981 b_5 NI_5 NS_981 0 1.9094674708988475e-05
GC_5_982 b_5 NI_5 NS_982 0 -5.5863940986972750e-06
GC_5_983 b_5 NI_5 NS_983 0 7.2293231308744144e-06
GC_5_984 b_5 NI_5 NS_984 0 -4.0341369461407490e-06
GC_5_985 b_5 NI_5 NS_985 0 1.3781905476062289e-05
GC_5_986 b_5 NI_5 NS_986 0 -1.1917593609536000e-05
GC_5_987 b_5 NI_5 NS_987 0 1.2441236848598050e-05
GC_5_988 b_5 NI_5 NS_988 0 -3.9380666699361914e-06
GC_5_989 b_5 NI_5 NS_989 0 9.3021677611912286e-06
GC_5_990 b_5 NI_5 NS_990 0 -2.6814459807702131e-05
GC_5_991 b_5 NI_5 NS_991 0 2.4411468471243563e-06
GC_5_992 b_5 NI_5 NS_992 0 -1.2372670604274647e-05
GC_5_993 b_5 NI_5 NS_993 0 -8.1267824700187677e-06
GC_5_994 b_5 NI_5 NS_994 0 -1.8722451998279471e-05
GC_5_995 b_5 NI_5 NS_995 0 -4.6961708714784151e-06
GC_5_996 b_5 NI_5 NS_996 0 -1.1981124154796818e-05
GC_5_997 b_5 NI_5 NS_997 0 5.4399747008271286e-05
GC_5_998 b_5 NI_5 NS_998 0 -8.9383189187739023e-05
GC_5_999 b_5 NI_5 NS_999 0 -9.7660143433605474e-06
GC_5_1000 b_5 NI_5 NS_1000 0 9.8738693240208092e-07
GC_5_1001 b_5 NI_5 NS_1001 0 3.8976886136704206e-07
GC_5_1002 b_5 NI_5 NS_1002 0 -1.3364777394303439e-07
GC_5_1003 b_5 NI_5 NS_1003 0 -2.5756641920700520e-06
GC_5_1004 b_5 NI_5 NS_1004 0 -2.1120215530047476e-06
GC_5_1005 b_5 NI_5 NS_1005 0 -4.3189724674128106e-06
GC_5_1006 b_5 NI_5 NS_1006 0 3.8846853618176418e-07
GC_5_1007 b_5 NI_5 NS_1007 0 -1.7308660525962059e-05
GC_5_1008 b_5 NI_5 NS_1008 0 9.7288625520407794e-06
GC_5_1009 b_5 NI_5 NS_1009 0 -8.8649401815520711e-06
GC_5_1010 b_5 NI_5 NS_1010 0 3.7519896972881330e-05
GC_5_1011 b_5 NI_5 NS_1011 0 -7.2572371004703778e-06
GC_5_1012 b_5 NI_5 NS_1012 0 3.2751357959642831e-07
GC_5_1013 b_5 NI_5 NS_1013 0 -1.3477623299685058e-05
GC_5_1014 b_5 NI_5 NS_1014 0 1.9011795167668807e-06
GC_5_1015 b_5 NI_5 NS_1015 0 -4.6310022224947511e-06
GC_5_1016 b_5 NI_5 NS_1016 0 -3.4347515913027859e-06
GC_5_1017 b_5 NI_5 NS_1017 0 -6.4037966539411824e-06
GC_5_1018 b_5 NI_5 NS_1018 0 1.0107233953113000e-06
GC_5_1019 b_5 NI_5 NS_1019 0 -3.0174082968894779e-06
GC_5_1020 b_5 NI_5 NS_1020 0 8.7541105855974870e-07
GC_5_1021 b_5 NI_5 NS_1021 0 -1.7610335328609159e-06
GC_5_1022 b_5 NI_5 NS_1022 0 -9.6128227804527740e-07
GC_5_1023 b_5 NI_5 NS_1023 0 -2.6099372611507963e-10
GC_5_1024 b_5 NI_5 NS_1024 0 4.2237635291794461e-10
GC_5_1025 b_5 NI_5 NS_1025 0 2.2554034748013341e-09
GC_5_1026 b_5 NI_5 NS_1026 0 -2.6817131746152097e-08
GC_5_1027 b_5 NI_5 NS_1027 0 -3.2388759236622915e-05
GC_5_1028 b_5 NI_5 NS_1028 0 2.2145965776025565e-06
GC_5_1029 b_5 NI_5 NS_1029 0 6.9002939971370114e-11
GC_5_1030 b_5 NI_5 NS_1030 0 3.0548434815266929e-09
GC_5_1031 b_5 NI_5 NS_1031 0 -1.7287512645275860e-06
GC_5_1032 b_5 NI_5 NS_1032 0 -1.8218260763185454e-06
GC_5_1033 b_5 NI_5 NS_1033 0 -5.3711639243487967e-06
GC_5_1034 b_5 NI_5 NS_1034 0 2.8657262423098405e-06
GC_5_1035 b_5 NI_5 NS_1035 0 -1.6530933290097456e-05
GC_5_1036 b_5 NI_5 NS_1036 0 1.8435108376158402e-05
GC_5_1037 b_5 NI_5 NS_1037 0 1.5105603169419866e-05
GC_5_1038 b_5 NI_5 NS_1038 0 9.7996894048179218e-06
GC_5_1039 b_5 NI_5 NS_1039 0 1.7319443063621244e-05
GC_5_1040 b_5 NI_5 NS_1040 0 2.2757435645912905e-05
GC_5_1041 b_5 NI_5 NS_1041 0 2.9271974718686333e-05
GC_5_1042 b_5 NI_5 NS_1042 0 4.9454578197242114e-06
GC_5_1043 b_5 NI_5 NS_1043 0 -3.0090409772668880e-06
GC_5_1044 b_5 NI_5 NS_1044 0 -1.8920180050644512e-06
GC_5_1045 b_5 NI_5 NS_1045 0 1.6961735728232527e-05
GC_5_1046 b_5 NI_5 NS_1046 0 -2.2247252949551382e-06
GC_5_1047 b_5 NI_5 NS_1047 0 1.2894021035178292e-04
GC_5_1048 b_5 NI_5 NS_1048 0 3.4692087785003753e-05
GC_5_1049 b_5 NI_5 NS_1049 0 -2.8903913355783665e-05
GC_5_1050 b_5 NI_5 NS_1050 0 -9.8807839414212338e-05
GC_5_1051 b_5 NI_5 NS_1051 0 2.4942601158106574e-05
GC_5_1052 b_5 NI_5 NS_1052 0 -3.1439987002836098e-05
GC_5_1053 b_5 NI_5 NS_1053 0 -4.1726498396969074e-05
GC_5_1054 b_5 NI_5 NS_1054 0 -1.6659245087811191e-04
GC_5_1055 b_5 NI_5 NS_1055 0 -4.1856851584360239e-05
GC_5_1056 b_5 NI_5 NS_1056 0 -4.9686691358037368e-06
GC_5_1057 b_5 NI_5 NS_1057 0 2.1526235893395072e-05
GC_5_1058 b_5 NI_5 NS_1058 0 -1.5189898289621131e-04
GC_5_1059 b_5 NI_5 NS_1059 0 -2.3067412435409638e-04
GC_5_1060 b_5 NI_5 NS_1060 0 1.1454640495307338e-04
GC_5_1061 b_5 NI_5 NS_1061 0 -3.7434567658238301e-05
GC_5_1062 b_5 NI_5 NS_1062 0 1.4285340919351651e-05
GC_5_1063 b_5 NI_5 NS_1063 0 -1.3769176255905223e-04
GC_5_1064 b_5 NI_5 NS_1064 0 1.3059703857631704e-04
GC_5_1065 b_5 NI_5 NS_1065 0 3.6482332886077584e-05
GC_5_1066 b_5 NI_5 NS_1066 0 4.1333508722116121e-05
GC_5_1067 b_5 NI_5 NS_1067 0 -3.8174269489161534e-05
GC_5_1068 b_5 NI_5 NS_1068 0 4.3297681487383522e-05
GC_5_1069 b_5 NI_5 NS_1069 0 8.7698892765724140e-05
GC_5_1070 b_5 NI_5 NS_1070 0 1.1839070577946095e-04
GC_5_1071 b_5 NI_5 NS_1071 0 2.7360737824007327e-05
GC_5_1072 b_5 NI_5 NS_1072 0 1.0188167510593487e-05
GC_5_1073 b_5 NI_5 NS_1073 0 8.7309936759315205e-05
GC_5_1074 b_5 NI_5 NS_1074 0 6.5589081583361592e-05
GC_5_1075 b_5 NI_5 NS_1075 0 2.0355450374273856e-05
GC_5_1076 b_5 NI_5 NS_1076 0 -5.7134226732691831e-05
GC_5_1077 b_5 NI_5 NS_1077 0 1.6985963752125083e-05
GC_5_1078 b_5 NI_5 NS_1078 0 -8.8834521239179430e-06
GC_5_1079 b_5 NI_5 NS_1079 0 8.5005736915284884e-06
GC_5_1080 b_5 NI_5 NS_1080 0 -3.2939544299990697e-05
GC_5_1081 b_5 NI_5 NS_1081 0 -8.8537955416307639e-06
GC_5_1082 b_5 NI_5 NS_1082 0 5.2635665046007741e-07
GC_5_1083 b_5 NI_5 NS_1083 0 -2.4130970051405349e-06
GC_5_1084 b_5 NI_5 NS_1084 0 8.5086595440983610e-06
GC_5_1085 b_5 NI_5 NS_1085 0 1.0220494071670488e-05
GC_5_1086 b_5 NI_5 NS_1086 0 6.0870241551042604e-06
GC_5_1087 b_5 NI_5 NS_1087 0 1.2161244357569573e-05
GC_5_1088 b_5 NI_5 NS_1088 0 -7.8264937820389737e-06
GC_5_1089 b_5 NI_5 NS_1089 0 -3.4879226923634435e-06
GC_5_1090 b_5 NI_5 NS_1090 0 -4.4670409547315724e-07
GC_5_1091 b_5 NI_5 NS_1091 0 2.4880910172267879e-06
GC_5_1092 b_5 NI_5 NS_1092 0 7.4079276295990581e-06
GC_5_1093 b_5 NI_5 NS_1093 0 1.3650681218737403e-05
GC_5_1094 b_5 NI_5 NS_1094 0 2.6359153981096664e-06
GC_5_1095 b_5 NI_5 NS_1095 0 4.5207268684470668e-06
GC_5_1096 b_5 NI_5 NS_1096 0 -1.4188593668369723e-05
GC_5_1097 b_5 NI_5 NS_1097 0 -5.9269932085063496e-06
GC_5_1098 b_5 NI_5 NS_1098 0 4.2582988380500010e-06
GC_5_1099 b_5 NI_5 NS_1099 0 1.0309907472409518e-05
GC_5_1100 b_5 NI_5 NS_1100 0 9.9374974623675213e-06
GC_5_1101 b_5 NI_5 NS_1101 0 1.7307650756809800e-05
GC_5_1102 b_5 NI_5 NS_1102 0 -4.2709223710566292e-06
GC_5_1103 b_5 NI_5 NS_1103 0 -9.2920994066731804e-06
GC_5_1104 b_5 NI_5 NS_1104 0 -1.5315611863387798e-05
GC_5_1105 b_5 NI_5 NS_1105 0 -4.0817827727046190e-06
GC_5_1106 b_5 NI_5 NS_1106 0 1.3516513534051377e-05
GC_5_1107 b_5 NI_5 NS_1107 0 2.0928896349612372e-05
GC_5_1108 b_5 NI_5 NS_1108 0 -5.6268434394199973e-07
GC_5_1109 b_5 NI_5 NS_1109 0 8.8751443490648215e-06
GC_5_1110 b_5 NI_5 NS_1110 0 -1.7452610544080247e-05
GC_5_1111 b_5 NI_5 NS_1111 0 2.4051623201568387e-06
GC_5_1112 b_5 NI_5 NS_1112 0 -1.3697890440136892e-05
GC_5_1113 b_5 NI_5 NS_1113 0 -1.3815629790831078e-05
GC_5_1114 b_5 NI_5 NS_1114 0 4.3768013490776305e-06
GC_5_1115 b_5 NI_5 NS_1115 0 1.5477816711465733e-08
GC_5_1116 b_5 NI_5 NS_1116 0 -4.2108817393574760e-08
GC_5_1117 b_5 NI_5 NS_1117 0 8.6211007962581327e-06
GC_5_1118 b_5 NI_5 NS_1118 0 1.1597928740736822e-05
GC_5_1119 b_5 NI_5 NS_1119 0 1.0904667048937961e-05
GC_5_1120 b_5 NI_5 NS_1120 0 -1.1278359719874704e-05
GC_5_1121 b_5 NI_5 NS_1121 0 -3.7307383214002499e-06
GC_5_1122 b_5 NI_5 NS_1122 0 -1.0216263848116271e-05
GC_5_1123 b_5 NI_5 NS_1123 0 -2.2940085956383701e-06
GC_5_1124 b_5 NI_5 NS_1124 0 1.2865967515829219e-05
GC_5_1125 b_5 NI_5 NS_1125 0 9.6691368501547296e-07
GC_5_1126 b_5 NI_5 NS_1126 0 -7.2695118225415127e-06
GC_5_1127 b_5 NI_5 NS_1127 0 7.5166615551516553e-06
GC_5_1128 b_5 NI_5 NS_1128 0 1.6931639200690833e-06
GC_5_1129 b_5 NI_5 NS_1129 0 -6.1012188469366923e-06
GC_5_1130 b_5 NI_5 NS_1130 0 -8.8953961914716168e-06
GC_5_1131 b_5 NI_5 NS_1131 0 -4.1215010615351704e-06
GC_5_1132 b_5 NI_5 NS_1132 0 9.6659601508050505e-06
GC_5_1133 b_5 NI_5 NS_1133 0 3.3268438650112730e-06
GC_5_1134 b_5 NI_5 NS_1134 0 6.0367137962417184e-06
GC_5_1135 b_5 NI_5 NS_1135 0 5.6518862078818838e-06
GC_5_1136 b_5 NI_5 NS_1136 0 5.1680465825212542e-07
GC_5_1137 b_5 NI_5 NS_1137 0 6.1804773114340677e-11
GC_5_1138 b_5 NI_5 NS_1138 0 1.4894831662766201e-10
GC_5_1139 b_5 NI_5 NS_1139 0 5.9431745329487181e-09
GC_5_1140 b_5 NI_5 NS_1140 0 -8.3385692131560821e-09
GC_5_1141 b_5 NI_5 NS_1141 0 8.4593945000548755e-05
GC_5_1142 b_5 NI_5 NS_1142 0 1.9043587625876777e-07
GC_5_1143 b_5 NI_5 NS_1143 0 2.0152904745714104e-11
GC_5_1144 b_5 NI_5 NS_1144 0 -9.4454556293862621e-10
GC_5_1145 b_5 NI_5 NS_1145 0 8.8362777003077878e-07
GC_5_1146 b_5 NI_5 NS_1146 0 5.7800682294055158e-08
GC_5_1147 b_5 NI_5 NS_1147 0 1.1605036444501343e-06
GC_5_1148 b_5 NI_5 NS_1148 0 6.9649917256652249e-08
GC_5_1149 b_5 NI_5 NS_1149 0 3.3633123224175221e-06
GC_5_1150 b_5 NI_5 NS_1150 0 -3.2270897511278628e-06
GC_5_1151 b_5 NI_5 NS_1151 0 -2.0864345922270994e-06
GC_5_1152 b_5 NI_5 NS_1152 0 -1.7323699217737436e-06
GC_5_1153 b_5 NI_5 NS_1153 0 1.9309984599618422e-06
GC_5_1154 b_5 NI_5 NS_1154 0 -2.2101001938191571e-06
GC_5_1155 b_5 NI_5 NS_1155 0 -5.8945393732665389e-06
GC_5_1156 b_5 NI_5 NS_1156 0 -7.1428808150440553e-06
GC_5_1157 b_5 NI_5 NS_1157 0 9.5034301878745669e-07
GC_5_1158 b_5 NI_5 NS_1158 0 2.2267366763210283e-06
GC_5_1159 b_5 NI_5 NS_1159 0 -2.2769834521873638e-06
GC_5_1160 b_5 NI_5 NS_1160 0 8.0128600459136622e-07
GC_5_1161 b_5 NI_5 NS_1161 0 5.8089039639728494e-07
GC_5_1162 b_5 NI_5 NS_1162 0 -4.8941802449791671e-06
GC_5_1163 b_5 NI_5 NS_1163 0 -6.4026889471751261e-06
GC_5_1164 b_5 NI_5 NS_1164 0 2.7563303125947548e-06
GC_5_1165 b_5 NI_5 NS_1165 0 -1.0161047564424483e-06
GC_5_1166 b_5 NI_5 NS_1166 0 1.6584680650572350e-06
GC_5_1167 b_5 NI_5 NS_1167 0 -3.3725642687036418e-06
GC_5_1168 b_5 NI_5 NS_1168 0 -2.5283990267920066e-06
GC_5_1169 b_5 NI_5 NS_1169 0 -2.2050141382453023e-06
GC_5_1170 b_5 NI_5 NS_1170 0 2.3624367573428191e-06
GC_5_1171 b_5 NI_5 NS_1171 0 1.5143152836767460e-06
GC_5_1172 b_5 NI_5 NS_1172 0 2.6092777460438463e-06
GC_5_1173 b_5 NI_5 NS_1173 0 -5.1177184610017399e-06
GC_5_1174 b_5 NI_5 NS_1174 0 -2.0375229565224095e-06
GC_5_1175 b_5 NI_5 NS_1175 0 -1.4942736644421925e-06
GC_5_1176 b_5 NI_5 NS_1176 0 2.2229726160365799e-06
GC_5_1177 b_5 NI_5 NS_1177 0 -4.8187213931578911e-08
GC_5_1178 b_5 NI_5 NS_1178 0 -1.0705803435921213e-06
GC_5_1179 b_5 NI_5 NS_1179 0 -2.7776412989789354e-06
GC_5_1180 b_5 NI_5 NS_1180 0 1.7676655625548331e-06
GC_5_1181 b_5 NI_5 NS_1181 0 -7.8794273890799669e-07
GC_5_1182 b_5 NI_5 NS_1182 0 2.3418921801307255e-06
GC_5_1183 b_5 NI_5 NS_1183 0 -1.0030646093228123e-06
GC_5_1184 b_5 NI_5 NS_1184 0 -1.3429446642495102e-06
GC_5_1185 b_5 NI_5 NS_1185 0 -1.8385161218631746e-06
GC_5_1186 b_5 NI_5 NS_1186 0 1.3366200313583133e-06
GC_5_1187 b_5 NI_5 NS_1187 0 5.5156955604000339e-07
GC_5_1188 b_5 NI_5 NS_1188 0 1.6537064897059237e-07
GC_5_1189 b_5 NI_5 NS_1189 0 -2.9420518113438026e-06
GC_5_1190 b_5 NI_5 NS_1190 0 3.7600509563664154e-07
GC_5_1191 b_5 NI_5 NS_1191 0 -9.6513326839409760e-07
GC_5_1192 b_5 NI_5 NS_1192 0 7.1182570839700041e-07
GC_5_1193 b_5 NI_5 NS_1193 0 -1.9725838231954989e-06
GC_5_1194 b_5 NI_5 NS_1194 0 -7.9480779743760974e-07
GC_5_1195 b_5 NI_5 NS_1195 0 -1.4687827304167386e-06
GC_5_1196 b_5 NI_5 NS_1196 0 6.2110219255598796e-07
GC_5_1197 b_5 NI_5 NS_1197 0 -1.1171949295931075e-06
GC_5_1198 b_5 NI_5 NS_1198 0 -3.9215291987900519e-07
GC_5_1199 b_5 NI_5 NS_1199 0 -2.4596159752342797e-06
GC_5_1200 b_5 NI_5 NS_1200 0 -6.3464719198008013e-07
GC_5_1201 b_5 NI_5 NS_1201 0 -3.0281906283826005e-06
GC_5_1202 b_5 NI_5 NS_1202 0 -3.1125413008622031e-07
GC_5_1203 b_5 NI_5 NS_1203 0 -2.1722949475214690e-06
GC_5_1204 b_5 NI_5 NS_1204 0 3.1827804888742888e-07
GC_5_1205 b_5 NI_5 NS_1205 0 -2.7407143734378282e-06
GC_5_1206 b_5 NI_5 NS_1206 0 3.0329373432768444e-07
GC_5_1207 b_5 NI_5 NS_1207 0 -4.2063163428023859e-06
GC_5_1208 b_5 NI_5 NS_1208 0 -7.3431075745416663e-07
GC_5_1209 b_5 NI_5 NS_1209 0 -5.6821682966511445e-06
GC_5_1210 b_5 NI_5 NS_1210 0 2.2501731868374763e-06
GC_5_1211 b_5 NI_5 NS_1211 0 -3.1748898490624498e-06
GC_5_1212 b_5 NI_5 NS_1212 0 1.8636231219688072e-06
GC_5_1213 b_5 NI_5 NS_1213 0 -4.1156147229978165e-06
GC_5_1214 b_5 NI_5 NS_1214 0 3.2996224993116206e-06
GC_5_1215 b_5 NI_5 NS_1215 0 -5.6743085523639884e-06
GC_5_1216 b_5 NI_5 NS_1216 0 1.3489552094601021e-06
GC_5_1217 b_5 NI_5 NS_1217 0 -3.5124576738228077e-06
GC_5_1218 b_5 NI_5 NS_1218 0 8.2350288171693081e-06
GC_5_1219 b_5 NI_5 NS_1219 0 -2.3080098975186840e-06
GC_5_1220 b_5 NI_5 NS_1220 0 4.5638946591091121e-06
GC_5_1221 b_5 NI_5 NS_1221 0 1.1256601544700588e-06
GC_5_1222 b_5 NI_5 NS_1222 0 5.4143284542593726e-06
GC_5_1223 b_5 NI_5 NS_1223 0 -1.8435302805147160e-06
GC_5_1224 b_5 NI_5 NS_1224 0 3.4528263916341807e-06
GC_5_1225 b_5 NI_5 NS_1225 0 -7.0146493688396952e-06
GC_5_1226 b_5 NI_5 NS_1226 0 3.7171371102132301e-05
GC_5_1227 b_5 NI_5 NS_1227 0 6.9438866436203685e-07
GC_5_1228 b_5 NI_5 NS_1228 0 2.6520874225041247e-06
GC_5_1229 b_5 NI_5 NS_1229 0 -8.4705184097565194e-08
GC_5_1230 b_5 NI_5 NS_1230 0 1.1842643871216040e-07
GC_5_1231 b_5 NI_5 NS_1231 0 -7.2474320830791814e-07
GC_5_1232 b_5 NI_5 NS_1232 0 3.4155277428189345e-06
GC_5_1233 b_5 NI_5 NS_1233 0 6.7707583142192229e-07
GC_5_1234 b_5 NI_5 NS_1234 0 8.6166755388301319e-07
GC_5_1235 b_5 NI_5 NS_1235 0 2.2818966074561194e-06
GC_5_1236 b_5 NI_5 NS_1236 0 -3.1368165094551809e-06
GC_5_1237 b_5 NI_5 NS_1237 0 -1.5493209398909649e-06
GC_5_1238 b_5 NI_5 NS_1238 0 -1.1843770573482743e-05
GC_5_1239 b_5 NI_5 NS_1239 0 2.0448389812803482e-06
GC_5_1240 b_5 NI_5 NS_1240 0 -7.3745612845071367e-07
GC_5_1241 b_5 NI_5 NS_1241 0 4.5136869169633078e-06
GC_5_1242 b_5 NI_5 NS_1242 0 -4.0126002828835334e-07
GC_5_1243 b_5 NI_5 NS_1243 0 1.2442633300173642e-06
GC_5_1244 b_5 NI_5 NS_1244 0 1.9854525450116060e-06
GC_5_1245 b_5 NI_5 NS_1245 0 1.7412906472416892e-06
GC_5_1246 b_5 NI_5 NS_1246 0 -7.6164097003040966e-07
GC_5_1247 b_5 NI_5 NS_1247 0 5.8319842415258926e-07
GC_5_1248 b_5 NI_5 NS_1248 0 5.1106052599804624e-07
GC_5_1249 b_5 NI_5 NS_1249 0 6.5667009545007142e-07
GC_5_1250 b_5 NI_5 NS_1250 0 -7.6188570425170858e-08
GC_5_1251 b_5 NI_5 NS_1251 0 2.2923100423621418e-11
GC_5_1252 b_5 NI_5 NS_1252 0 -9.3363869332698833e-11
GC_5_1253 b_5 NI_5 NS_1253 0 -1.8301880559619860e-09
GC_5_1254 b_5 NI_5 NS_1254 0 4.0621497241107225e-09
GC_5_1255 b_5 NI_5 NS_1255 0 -6.3086645279662940e-05
GC_5_1256 b_5 NI_5 NS_1256 0 3.1407867978578684e-07
GC_5_1257 b_5 NI_5 NS_1257 0 1.6213866530362793e-11
GC_5_1258 b_5 NI_5 NS_1258 0 -9.0527175141136995e-11
GC_5_1259 b_5 NI_5 NS_1259 0 -1.1178109159694303e-06
GC_5_1260 b_5 NI_5 NS_1260 0 -1.7847510948111635e-06
GC_5_1261 b_5 NI_5 NS_1261 0 -1.9986015271080415e-06
GC_5_1262 b_5 NI_5 NS_1262 0 1.9870799049704329e-06
GC_5_1263 b_5 NI_5 NS_1263 0 -9.6875187598289361e-06
GC_5_1264 b_5 NI_5 NS_1264 0 6.6933774804672807e-07
GC_5_1265 b_5 NI_5 NS_1265 0 -2.3281015655076691e-07
GC_5_1266 b_5 NI_5 NS_1266 0 3.4992261183088638e-06
GC_5_1267 b_5 NI_5 NS_1267 0 -2.1124315053196704e-06
GC_5_1268 b_5 NI_5 NS_1268 0 1.1812007203418651e-05
GC_5_1269 b_5 NI_5 NS_1269 0 6.7540161416432809e-06
GC_5_1270 b_5 NI_5 NS_1270 0 1.2474526010109672e-05
GC_5_1271 b_5 NI_5 NS_1271 0 -1.9954500394169794e-06
GC_5_1272 b_5 NI_5 NS_1272 0 -2.3039269237009676e-06
GC_5_1273 b_5 NI_5 NS_1273 0 1.6659035743044277e-06
GC_5_1274 b_5 NI_5 NS_1274 0 9.5797696227169434e-07
GC_5_1275 b_5 NI_5 NS_1275 0 7.5629424579188954e-06
GC_5_1276 b_5 NI_5 NS_1276 0 3.8828221112901028e-05
GC_5_1277 b_5 NI_5 NS_1277 0 2.3010290785898298e-05
GC_5_1278 b_5 NI_5 NS_1278 0 -1.1868416740827938e-05
GC_5_1279 b_5 NI_5 NS_1279 0 8.3672968413770518e-06
GC_5_1280 b_5 NI_5 NS_1280 0 1.6445429537527524e-06
GC_5_1281 b_5 NI_5 NS_1281 0 4.8509109833355077e-05
GC_5_1282 b_5 NI_5 NS_1282 0 -2.5181062648604696e-05
GC_5_1283 b_5 NI_5 NS_1283 0 -8.8536567940270809e-07
GC_5_1284 b_5 NI_5 NS_1284 0 -7.8651555507748873e-06
GC_5_1285 b_5 NI_5 NS_1285 0 3.4167774046203124e-05
GC_5_1286 b_5 NI_5 NS_1286 0 -7.8499469664938443e-06
GC_5_1287 b_5 NI_5 NS_1287 0 -3.8183050727541407e-05
GC_5_1288 b_5 NI_5 NS_1288 0 -5.2548380026202231e-05
GC_5_1289 b_5 NI_5 NS_1289 0 -4.5027047674618118e-06
GC_5_1290 b_5 NI_5 NS_1290 0 -4.3379498095764061e-06
GC_5_1291 b_5 NI_5 NS_1291 0 -3.9815354980797148e-05
GC_5_1292 b_5 NI_5 NS_1292 0 -2.0116802145661636e-05
GC_5_1293 b_5 NI_5 NS_1293 0 -4.8511669074329962e-06
GC_5_1294 b_5 NI_5 NS_1294 0 6.2282646849232519e-06
GC_5_1295 b_5 NI_5 NS_1295 0 -8.5210919686255102e-06
GC_5_1296 b_5 NI_5 NS_1296 0 -4.5734694863787880e-07
GC_5_1297 b_5 NI_5 NS_1297 0 -1.5552803078521248e-05
GC_5_1298 b_5 NI_5 NS_1298 0 2.4319404154174891e-05
GC_5_1299 b_5 NI_5 NS_1299 0 1.1127387886890431e-06
GC_5_1300 b_5 NI_5 NS_1300 0 2.3765188209660730e-06
GC_5_1301 b_5 NI_5 NS_1301 0 3.2444555840893669e-06
GC_5_1302 b_5 NI_5 NS_1302 0 1.8514021733069055e-05
GC_5_1303 b_5 NI_5 NS_1303 0 7.5499014163536519e-06
GC_5_1304 b_5 NI_5 NS_1304 0 -1.4049668828526414e-06
GC_5_1305 b_5 NI_5 NS_1305 0 2.9997394428970235e-06
GC_5_1306 b_5 NI_5 NS_1306 0 -5.0735584451537584e-07
GC_5_1307 b_5 NI_5 NS_1307 0 7.6482564242695034e-06
GC_5_1308 b_5 NI_5 NS_1308 0 -4.5383957103544794e-06
GC_5_1309 b_5 NI_5 NS_1309 0 -8.6323819922225607e-07
GC_5_1310 b_5 NI_5 NS_1310 0 -4.4782532919575186e-07
GC_5_1311 b_5 NI_5 NS_1311 0 -1.7220285686243629e-06
GC_5_1312 b_5 NI_5 NS_1312 0 1.8650698046659519e-07
GC_5_1313 b_5 NI_5 NS_1313 0 1.6124745586651558e-06
GC_5_1314 b_5 NI_5 NS_1314 0 -2.3833195904553990e-08
GC_5_1315 b_5 NI_5 NS_1315 0 3.7027745012660569e-06
GC_5_1316 b_5 NI_5 NS_1316 0 -9.2679739402290550e-07
GC_5_1317 b_5 NI_5 NS_1317 0 -8.7848001086322951e-08
GC_5_1318 b_5 NI_5 NS_1318 0 -3.4244846245808609e-07
GC_5_1319 b_5 NI_5 NS_1319 0 -5.7040535905980130e-07
GC_5_1320 b_5 NI_5 NS_1320 0 5.1106374703081481e-07
GC_5_1321 b_5 NI_5 NS_1321 0 2.4651881959351212e-06
GC_5_1322 b_5 NI_5 NS_1322 0 1.0968662789096046e-07
GC_5_1323 b_5 NI_5 NS_1323 0 3.4038999996556152e-06
GC_5_1324 b_5 NI_5 NS_1324 0 -2.8600674099549354e-06
GC_5_1325 b_5 NI_5 NS_1325 0 -2.6935639532301614e-07
GC_5_1326 b_5 NI_5 NS_1326 0 -4.9653644332205106e-08
GC_5_1327 b_5 NI_5 NS_1327 0 7.1909391291809887e-07
GC_5_1328 b_5 NI_5 NS_1328 0 1.0039440381761531e-06
GC_5_1329 b_5 NI_5 NS_1329 0 3.5525123624457384e-06
GC_5_1330 b_5 NI_5 NS_1330 0 3.5543547594451926e-08
GC_5_1331 b_5 NI_5 NS_1331 0 2.4198778221187198e-06
GC_5_1332 b_5 NI_5 NS_1332 0 -4.6562318473497734e-06
GC_5_1333 b_5 NI_5 NS_1333 0 4.5355979519440496e-07
GC_5_1334 b_5 NI_5 NS_1334 0 1.1318772898967800e-06
GC_5_1335 b_5 NI_5 NS_1335 0 3.6738603367761573e-06
GC_5_1336 b_5 NI_5 NS_1336 0 -6.8877976680333246e-07
GC_5_1337 b_5 NI_5 NS_1337 0 5.6188310830190173e-06
GC_5_1338 b_5 NI_5 NS_1338 0 -9.6837063983801948e-07
GC_5_1339 b_5 NI_5 NS_1339 0 -1.6176022882134558e-05
GC_5_1340 b_5 NI_5 NS_1340 0 -1.0667578796652355e-05
GC_5_1341 b_5 NI_5 NS_1341 0 9.4792211858896026e-07
GC_5_1342 b_5 NI_5 NS_1342 0 -7.4950609659774466e-06
GC_5_1343 b_5 NI_5 NS_1343 0 -6.7190881648230835e-08
GC_5_1344 b_5 NI_5 NS_1344 0 -1.4892210323190501e-07
GC_5_1345 b_5 NI_5 NS_1345 0 1.8092881233205507e-06
GC_5_1346 b_5 NI_5 NS_1346 0 -1.8934174919403702e-06
GC_5_1347 b_5 NI_5 NS_1347 0 5.4099645297281473e-07
GC_5_1348 b_5 NI_5 NS_1348 0 -3.3989041988201642e-06
GC_5_1349 b_5 NI_5 NS_1349 0 3.4155695217391424e-06
GC_5_1350 b_5 NI_5 NS_1350 0 -1.3122435379063151e-06
GC_5_1351 b_5 NI_5 NS_1351 0 4.5902932245826417e-06
GC_5_1352 b_5 NI_5 NS_1352 0 -7.9885751780107605e-07
GC_5_1353 b_5 NI_5 NS_1353 0 -1.9723755486015696e-07
GC_5_1354 b_5 NI_5 NS_1354 0 -2.0613870518459506e-07
GC_5_1355 b_5 NI_5 NS_1355 0 7.0253925868440331e-07
GC_5_1356 b_5 NI_5 NS_1356 0 1.4071776829324501e-06
GC_5_1357 b_5 NI_5 NS_1357 0 -7.0005252233569601e-07
GC_5_1358 b_5 NI_5 NS_1358 0 -1.4722237414631031e-06
GC_5_1359 b_5 NI_5 NS_1359 0 -6.2852494578832304e-07
GC_5_1360 b_5 NI_5 NS_1360 0 8.2374766447794051e-07
GC_5_1361 b_5 NI_5 NS_1361 0 2.2513794143056179e-07
GC_5_1362 b_5 NI_5 NS_1362 0 6.5418615274512713e-07
GC_5_1363 b_5 NI_5 NS_1363 0 6.0606486366309532e-07
GC_5_1364 b_5 NI_5 NS_1364 0 2.1063180908266877e-08
GC_5_1365 b_5 NI_5 NS_1365 0 1.3944022897221253e-11
GC_5_1366 b_5 NI_5 NS_1366 0 5.4831938948527919e-13
GC_5_1367 b_5 NI_5 NS_1367 0 4.3772280629553725e-10
GC_5_1368 b_5 NI_5 NS_1368 0 1.6923733613232480e-09
GD_5_1 b_5 NI_5 NA_1 0 5.3912437032568475e-06
GD_5_2 b_5 NI_5 NA_2 0 2.4210553079270388e-06
GD_5_3 b_5 NI_5 NA_3 0 1.0031817881093703e-04
GD_5_4 b_5 NI_5 NA_4 0 2.7000166674696918e-05
GD_5_5 b_5 NI_5 NA_5 0 -8.8807860850851610e-03
GD_5_6 b_5 NI_5 NA_6 0 -4.2218428274150514e-03
GD_5_7 b_5 NI_5 NA_7 0 1.2979344857305371e-02
GD_5_8 b_5 NI_5 NA_8 0 5.8608994894660622e-04
GD_5_9 b_5 NI_5 NA_9 0 4.8704189576553740e-06
GD_5_10 b_5 NI_5 NA_10 0 1.2379598094560608e-06
GD_5_11 b_5 NI_5 NA_11 0 -6.7055790994299297e-06
GD_5_12 b_5 NI_5 NA_12 0 1.0203935186402119e-05
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 -3.8126167498904904e-05
GC_6_2 b_6 NI_6 NS_2 0 2.2429781029594003e-06
GC_6_3 b_6 NI_6 NS_3 0 5.7510359651917983e-11
GC_6_4 b_6 NI_6 NS_4 0 3.0676995634755480e-09
GC_6_5 b_6 NI_6 NS_5 0 -1.9278398255944989e-06
GC_6_6 b_6 NI_6 NS_6 0 -1.7007518341002390e-06
GC_6_7 b_6 NI_6 NS_7 0 -5.6017359168061826e-06
GC_6_8 b_6 NI_6 NS_8 0 2.8809325672355818e-06
GC_6_9 b_6 NI_6 NS_9 0 -1.6609153059418861e-05
GC_6_10 b_6 NI_6 NS_10 0 1.9115492548943403e-05
GC_6_11 b_6 NI_6 NS_11 0 1.5381836614873184e-05
GC_6_12 b_6 NI_6 NS_12 0 1.0271591444337598e-05
GC_6_13 b_6 NI_6 NS_13 0 1.7283116207380704e-05
GC_6_14 b_6 NI_6 NS_14 0 2.3212335716383672e-05
GC_6_15 b_6 NI_6 NS_15 0 3.0964752020319569e-05
GC_6_16 b_6 NI_6 NS_16 0 5.3078575569417221e-06
GC_6_17 b_6 NI_6 NS_17 0 -3.3865366264644635e-06
GC_6_18 b_6 NI_6 NS_18 0 -2.1454228487573289e-06
GC_6_19 b_6 NI_6 NS_19 0 1.7199897151050782e-05
GC_6_20 b_6 NI_6 NS_20 0 -2.1239550484374399e-06
GC_6_21 b_6 NI_6 NS_21 0 1.2959269891114192e-04
GC_6_22 b_6 NI_6 NS_22 0 3.5268000057704650e-05
GC_6_23 b_6 NI_6 NS_23 0 -2.8363540471269497e-05
GC_6_24 b_6 NI_6 NS_24 0 -1.0001972403792202e-04
GC_6_25 b_6 NI_6 NS_25 0 2.5326199919349488e-05
GC_6_26 b_6 NI_6 NS_26 0 -3.1109554325742436e-05
GC_6_27 b_6 NI_6 NS_27 0 -4.1103626820163804e-05
GC_6_28 b_6 NI_6 NS_28 0 -1.6753402429527917e-04
GC_6_29 b_6 NI_6 NS_29 0 -4.1819869166084924e-05
GC_6_30 b_6 NI_6 NS_30 0 -5.5994631628349588e-06
GC_6_31 b_6 NI_6 NS_31 0 2.2900987906483162e-05
GC_6_32 b_6 NI_6 NS_32 0 -1.5132579346638524e-04
GC_6_33 b_6 NI_6 NS_33 0 -2.3194062743486644e-04
GC_6_34 b_6 NI_6 NS_34 0 1.1300294583693434e-04
GC_6_35 b_6 NI_6 NS_35 0 -3.7469906640010690e-05
GC_6_36 b_6 NI_6 NS_36 0 1.3727346542828026e-05
GC_6_37 b_6 NI_6 NS_37 0 -1.3772206217606826e-04
GC_6_38 b_6 NI_6 NS_38 0 1.2973991888027455e-04
GC_6_39 b_6 NI_6 NS_39 0 3.6015990640722157e-05
GC_6_40 b_6 NI_6 NS_40 0 4.1758736276267767e-05
GC_6_41 b_6 NI_6 NS_41 0 -3.8325873809074661e-05
GC_6_42 b_6 NI_6 NS_42 0 4.2733754272956775e-05
GC_6_43 b_6 NI_6 NS_43 0 8.7553202112611349e-05
GC_6_44 b_6 NI_6 NS_44 0 1.1830509427155053e-04
GC_6_45 b_6 NI_6 NS_45 0 2.7200342058781531e-05
GC_6_46 b_6 NI_6 NS_46 0 1.0487248295016989e-05
GC_6_47 b_6 NI_6 NS_47 0 8.6919299627232434e-05
GC_6_48 b_6 NI_6 NS_48 0 6.5387413656876116e-05
GC_6_49 b_6 NI_6 NS_49 0 2.0648990667106847e-05
GC_6_50 b_6 NI_6 NS_50 0 -5.7329957147797706e-05
GC_6_51 b_6 NI_6 NS_51 0 1.7010942654229642e-05
GC_6_52 b_6 NI_6 NS_52 0 -8.6982089229162380e-06
GC_6_53 b_6 NI_6 NS_53 0 8.3263460328043318e-06
GC_6_54 b_6 NI_6 NS_54 0 -3.3101466474613745e-05
GC_6_55 b_6 NI_6 NS_55 0 -8.8263215473903780e-06
GC_6_56 b_6 NI_6 NS_56 0 3.3245562859718456e-07
GC_6_57 b_6 NI_6 NS_57 0 -2.3512428422783518e-06
GC_6_58 b_6 NI_6 NS_58 0 8.4561786477537828e-06
GC_6_59 b_6 NI_6 NS_59 0 1.0134608961356484e-05
GC_6_60 b_6 NI_6 NS_60 0 6.1703161236356179e-06
GC_6_61 b_6 NI_6 NS_61 0 1.2106284013512765e-05
GC_6_62 b_6 NI_6 NS_62 0 -7.8947994038582263e-06
GC_6_63 b_6 NI_6 NS_63 0 -3.4458122283526067e-06
GC_6_64 b_6 NI_6 NS_64 0 -5.4102859497677728e-07
GC_6_65 b_6 NI_6 NS_65 0 2.5535456873308740e-06
GC_6_66 b_6 NI_6 NS_66 0 7.3550398515627659e-06
GC_6_67 b_6 NI_6 NS_67 0 1.3648181308741491e-05
GC_6_68 b_6 NI_6 NS_68 0 2.7057431484486200e-06
GC_6_69 b_6 NI_6 NS_69 0 4.5460300386772046e-06
GC_6_70 b_6 NI_6 NS_70 0 -1.4254775541062906e-05
GC_6_71 b_6 NI_6 NS_71 0 -5.8809803714181202e-06
GC_6_72 b_6 NI_6 NS_72 0 4.1779767899001233e-06
GC_6_73 b_6 NI_6 NS_73 0 1.0407200121259603e-05
GC_6_74 b_6 NI_6 NS_74 0 9.8673822299743229e-06
GC_6_75 b_6 NI_6 NS_75 0 1.7371591998047629e-05
GC_6_76 b_6 NI_6 NS_76 0 -4.2133716606638691e-06
GC_6_77 b_6 NI_6 NS_77 0 -9.1859937904139183e-06
GC_6_78 b_6 NI_6 NS_78 0 -1.5417368825990374e-05
GC_6_79 b_6 NI_6 NS_79 0 -3.9937397375735811e-06
GC_6_80 b_6 NI_6 NS_80 0 1.3459880288383124e-05
GC_6_81 b_6 NI_6 NS_81 0 2.1061389715988901e-05
GC_6_82 b_6 NI_6 NS_82 0 -6.9747416149329755e-07
GC_6_83 b_6 NI_6 NS_83 0 9.0884891473744352e-06
GC_6_84 b_6 NI_6 NS_84 0 -1.7352200317051005e-05
GC_6_85 b_6 NI_6 NS_85 0 1.8906782029196468e-06
GC_6_86 b_6 NI_6 NS_86 0 -1.4899320073310816e-05
GC_6_87 b_6 NI_6 NS_87 0 -1.3643677216078234e-05
GC_6_88 b_6 NI_6 NS_88 0 4.0673663154417879e-06
GC_6_89 b_6 NI_6 NS_89 0 1.3202624173125460e-08
GC_6_90 b_6 NI_6 NS_90 0 -4.9293050598111986e-08
GC_6_91 b_6 NI_6 NS_91 0 8.7095241516492612e-06
GC_6_92 b_6 NI_6 NS_92 0 1.1413353069764621e-05
GC_6_93 b_6 NI_6 NS_93 0 1.0949855281381823e-05
GC_6_94 b_6 NI_6 NS_94 0 -1.1467433621744669e-05
GC_6_95 b_6 NI_6 NS_95 0 -3.5678171995323697e-06
GC_6_96 b_6 NI_6 NS_96 0 -1.0053365775096303e-05
GC_6_97 b_6 NI_6 NS_97 0 -2.0108357603882727e-06
GC_6_98 b_6 NI_6 NS_98 0 1.3050211452451848e-05
GC_6_99 b_6 NI_6 NS_99 0 9.7274313567565796e-07
GC_6_100 b_6 NI_6 NS_100 0 -7.2791931807776694e-06
GC_6_101 b_6 NI_6 NS_101 0 7.4348969472655980e-06
GC_6_102 b_6 NI_6 NS_102 0 1.7180575561354758e-06
GC_6_103 b_6 NI_6 NS_103 0 -6.1040136152446632e-06
GC_6_104 b_6 NI_6 NS_104 0 -8.8986588350437229e-06
GC_6_105 b_6 NI_6 NS_105 0 -4.1281705029553164e-06
GC_6_106 b_6 NI_6 NS_106 0 9.6390055647591743e-06
GC_6_107 b_6 NI_6 NS_107 0 3.3246533998431558e-06
GC_6_108 b_6 NI_6 NS_108 0 6.0744635697527594e-06
GC_6_109 b_6 NI_6 NS_109 0 5.7495241645993535e-06
GC_6_110 b_6 NI_6 NS_110 0 5.2303412184843215e-07
GC_6_111 b_6 NI_6 NS_111 0 5.7042472242073175e-11
GC_6_112 b_6 NI_6 NS_112 0 1.4838931782381694e-10
GC_6_113 b_6 NI_6 NS_113 0 6.0314106867941374e-09
GC_6_114 b_6 NI_6 NS_114 0 -8.4056555786174642e-09
GC_6_115 b_6 NI_6 NS_115 0 -1.1990417440852588e-04
GC_6_116 b_6 NI_6 NS_116 0 -2.1506583358240569e-06
GC_6_117 b_6 NI_6 NS_117 0 -2.4444181352678074e-10
GC_6_118 b_6 NI_6 NS_118 0 2.5345869598460184e-09
GC_6_119 b_6 NI_6 NS_119 0 1.5459797113158055e-06
GC_6_120 b_6 NI_6 NS_120 0 -1.4954279590271684e-06
GC_6_121 b_6 NI_6 NS_121 0 -2.6328574170036756e-08
GC_6_122 b_6 NI_6 NS_122 0 -6.1347873435825482e-06
GC_6_123 b_6 NI_6 NS_123 0 -7.5890813797956327e-06
GC_6_124 b_6 NI_6 NS_124 0 6.3141463932684011e-07
GC_6_125 b_6 NI_6 NS_125 0 -9.4093704978995330e-07
GC_6_126 b_6 NI_6 NS_126 0 -4.4034014118364766e-06
GC_6_127 b_6 NI_6 NS_127 0 -1.5515996069313019e-05
GC_6_128 b_6 NI_6 NS_128 0 -1.2262225651697471e-06
GC_6_129 b_6 NI_6 NS_129 0 -5.1272327664245586e-06
GC_6_130 b_6 NI_6 NS_130 0 1.9057489030099395e-05
GC_6_131 b_6 NI_6 NS_131 0 4.3659578823061098e-06
GC_6_132 b_6 NI_6 NS_132 0 -3.1091686385509134e-06
GC_6_133 b_6 NI_6 NS_133 0 1.2739379514196837e-07
GC_6_134 b_6 NI_6 NS_134 0 -2.6189011600412056e-06
GC_6_135 b_6 NI_6 NS_135 0 -2.4695118632619753e-05
GC_6_136 b_6 NI_6 NS_136 0 2.8214913353463016e-05
GC_6_137 b_6 NI_6 NS_137 0 2.7678010805490588e-05
GC_6_138 b_6 NI_6 NS_138 0 -8.8491169767577627e-06
GC_6_139 b_6 NI_6 NS_139 0 -7.7786900857718351e-06
GC_6_140 b_6 NI_6 NS_140 0 -4.1717377847997626e-06
GC_6_141 b_6 NI_6 NS_141 0 1.2852721032089346e-05
GC_6_142 b_6 NI_6 NS_142 0 2.5989431798251348e-05
GC_6_143 b_6 NI_6 NS_143 0 1.3965872811729415e-06
GC_6_144 b_6 NI_6 NS_144 0 -8.8467713029253539e-06
GC_6_145 b_6 NI_6 NS_145 0 -2.7274070350010502e-05
GC_6_146 b_6 NI_6 NS_146 0 5.0518924522466653e-06
GC_6_147 b_6 NI_6 NS_147 0 4.0358168113828382e-05
GC_6_148 b_6 NI_6 NS_148 0 9.5136822509538962e-06
GC_6_149 b_6 NI_6 NS_149 0 -2.8939298288639839e-06
GC_6_150 b_6 NI_6 NS_150 0 -4.3230654062133983e-06
GC_6_151 b_6 NI_6 NS_151 0 1.3068135327278249e-05
GC_6_152 b_6 NI_6 NS_152 0 1.8039409574162778e-05
GC_6_153 b_6 NI_6 NS_153 0 3.4806890041344376e-06
GC_6_154 b_6 NI_6 NS_154 0 -1.0690735079403716e-05
GC_6_155 b_6 NI_6 NS_155 0 -6.1534218898160505e-06
GC_6_156 b_6 NI_6 NS_156 0 1.0246668015362979e-06
GC_6_157 b_6 NI_6 NS_157 0 1.8579425228197407e-05
GC_6_158 b_6 NI_6 NS_158 0 4.7194966317507613e-06
GC_6_159 b_6 NI_6 NS_159 0 -1.7163668492294431e-07
GC_6_160 b_6 NI_6 NS_160 0 -4.0410338058817101e-06
GC_6_161 b_6 NI_6 NS_161 0 5.3110691348675666e-06
GC_6_162 b_6 NI_6 NS_162 0 1.3887857656229515e-05
GC_6_163 b_6 NI_6 NS_163 0 7.3444730767557989e-06
GC_6_164 b_6 NI_6 NS_164 0 -1.1159205176177959e-05
GC_6_165 b_6 NI_6 NS_165 0 -1.3421714957123194e-06
GC_6_166 b_6 NI_6 NS_166 0 1.0174183700969009e-06
GC_6_167 b_6 NI_6 NS_167 0 1.0876591141454416e-05
GC_6_168 b_6 NI_6 NS_168 0 3.8402785340936240e-06
GC_6_169 b_6 NI_6 NS_169 0 1.6848232680845111e-06
GC_6_170 b_6 NI_6 NS_170 0 -6.0383776755681599e-07
GC_6_171 b_6 NI_6 NS_171 0 5.6746776763057712e-06
GC_6_172 b_6 NI_6 NS_172 0 1.5928961566815613e-06
GC_6_173 b_6 NI_6 NS_173 0 3.3876858951859986e-06
GC_6_174 b_6 NI_6 NS_174 0 2.0447825481673611e-06
GC_6_175 b_6 NI_6 NS_175 0 1.1009150710055745e-05
GC_6_176 b_6 NI_6 NS_176 0 3.6665168110645397e-06
GC_6_177 b_6 NI_6 NS_177 0 4.8524825097967841e-06
GC_6_178 b_6 NI_6 NS_178 0 -9.3154958796501975e-08
GC_6_179 b_6 NI_6 NS_179 0 9.9846404982325201e-06
GC_6_180 b_6 NI_6 NS_180 0 -1.1688009489528576e-06
GC_6_181 b_6 NI_6 NS_181 0 8.2907546430226168e-06
GC_6_182 b_6 NI_6 NS_182 0 2.9619519518434585e-06
GC_6_183 b_6 NI_6 NS_183 0 1.9135356567013588e-05
GC_6_184 b_6 NI_6 NS_184 0 -5.6872197204318334e-06
GC_6_185 b_6 NI_6 NS_185 0 7.2561490929741689e-06
GC_6_186 b_6 NI_6 NS_186 0 -4.0375692779454695e-06
GC_6_187 b_6 NI_6 NS_187 0 1.3814374772253572e-05
GC_6_188 b_6 NI_6 NS_188 0 -1.2017012419790670e-05
GC_6_189 b_6 NI_6 NS_189 0 1.2524732366842470e-05
GC_6_190 b_6 NI_6 NS_190 0 -3.9196660386618501e-06
GC_6_191 b_6 NI_6 NS_191 0 9.3874019958160737e-06
GC_6_192 b_6 NI_6 NS_192 0 -2.7008491593010351e-05
GC_6_193 b_6 NI_6 NS_193 0 2.5340509141880350e-06
GC_6_194 b_6 NI_6 NS_194 0 -1.2433576174181965e-05
GC_6_195 b_6 NI_6 NS_195 0 -8.1011422336396857e-06
GC_6_196 b_6 NI_6 NS_196 0 -1.8935729582527257e-05
GC_6_197 b_6 NI_6 NS_197 0 -4.4539207899344550e-06
GC_6_198 b_6 NI_6 NS_198 0 -1.2056802916593666e-05
GC_6_199 b_6 NI_6 NS_199 0 5.2729054732788339e-05
GC_6_200 b_6 NI_6 NS_200 0 -8.9465544404301233e-05
GC_6_201 b_6 NI_6 NS_201 0 -9.8695735230671165e-06
GC_6_202 b_6 NI_6 NS_202 0 5.5951851249645228e-07
GC_6_203 b_6 NI_6 NS_203 0 3.8236083341678917e-07
GC_6_204 b_6 NI_6 NS_204 0 -1.3957348841041311e-07
GC_6_205 b_6 NI_6 NS_205 0 -2.6066255324181425e-06
GC_6_206 b_6 NI_6 NS_206 0 -2.3472557574728509e-06
GC_6_207 b_6 NI_6 NS_207 0 -4.4561576353773485e-06
GC_6_208 b_6 NI_6 NS_208 0 2.3602466711457792e-07
GC_6_209 b_6 NI_6 NS_209 0 -1.7027355767154582e-05
GC_6_210 b_6 NI_6 NS_210 0 9.6526754645207218e-06
GC_6_211 b_6 NI_6 NS_211 0 -8.5113175886080545e-06
GC_6_212 b_6 NI_6 NS_212 0 3.7251828582572745e-05
GC_6_213 b_6 NI_6 NS_213 0 -7.2790849656625347e-06
GC_6_214 b_6 NI_6 NS_214 0 3.7957317663237260e-07
GC_6_215 b_6 NI_6 NS_215 0 -1.3447171477509145e-05
GC_6_216 b_6 NI_6 NS_216 0 1.9992894116103447e-06
GC_6_217 b_6 NI_6 NS_217 0 -4.6778654474372175e-06
GC_6_218 b_6 NI_6 NS_218 0 -3.4374763063909167e-06
GC_6_219 b_6 NI_6 NS_219 0 -6.4554994467250189e-06
GC_6_220 b_6 NI_6 NS_220 0 1.0434673451375805e-06
GC_6_221 b_6 NI_6 NS_221 0 -3.0715773509490951e-06
GC_6_222 b_6 NI_6 NS_222 0 8.7380282997168591e-07
GC_6_223 b_6 NI_6 NS_223 0 -1.8084091140574290e-06
GC_6_224 b_6 NI_6 NS_224 0 -9.3492551845693792e-07
GC_6_225 b_6 NI_6 NS_225 0 -2.5769930139644211e-10
GC_6_226 b_6 NI_6 NS_226 0 4.1862385617761563e-10
GC_6_227 b_6 NI_6 NS_227 0 2.1402111055303004e-09
GC_6_228 b_6 NI_6 NS_228 0 -2.6513263824301824e-08
GC_6_229 b_6 NI_6 NS_229 0 -2.0458585301878410e-04
GC_6_230 b_6 NI_6 NS_230 0 -3.3255724775698829e-06
GC_6_231 b_6 NI_6 NS_231 0 1.2945366104495201e-09
GC_6_232 b_6 NI_6 NS_232 0 9.6769689612394179e-09
GC_6_233 b_6 NI_6 NS_233 0 -4.2458928393087929e-06
GC_6_234 b_6 NI_6 NS_234 0 6.2176569447482565e-06
GC_6_235 b_6 NI_6 NS_235 0 3.7003799270299823e-06
GC_6_236 b_6 NI_6 NS_236 0 -8.0289276916718963e-06
GC_6_237 b_6 NI_6 NS_237 0 2.1715322490767114e-05
GC_6_238 b_6 NI_6 NS_238 0 -8.4141854411167379e-06
GC_6_239 b_6 NI_6 NS_239 0 -2.1191980736283601e-05
GC_6_240 b_6 NI_6 NS_240 0 -1.1902007288802127e-06
GC_6_241 b_6 NI_6 NS_241 0 -2.9306371123143939e-05
GC_6_242 b_6 NI_6 NS_242 0 -2.8028703547120027e-05
GC_6_243 b_6 NI_6 NS_243 0 -4.8383266125104130e-06
GC_6_244 b_6 NI_6 NS_244 0 1.6178945784831173e-05
GC_6_245 b_6 NI_6 NS_245 0 -2.6738580746843629e-06
GC_6_246 b_6 NI_6 NS_246 0 -7.1112471266582359e-06
GC_6_247 b_6 NI_6 NS_247 0 -2.2526885815362042e-05
GC_6_248 b_6 NI_6 NS_248 0 5.7341816120098449e-06
GC_6_249 b_6 NI_6 NS_249 0 -1.8493942568726518e-04
GC_6_250 b_6 NI_6 NS_250 0 -4.4593183009224079e-05
GC_6_251 b_6 NI_6 NS_251 0 6.1949165212607686e-05
GC_6_252 b_6 NI_6 NS_252 0 1.3746856757030927e-04
GC_6_253 b_6 NI_6 NS_253 0 -3.7405898064622544e-05
GC_6_254 b_6 NI_6 NS_254 0 5.6303425873817561e-05
GC_6_255 b_6 NI_6 NS_255 0 9.4942291767869671e-05
GC_6_256 b_6 NI_6 NS_256 0 2.4590670669831483e-04
GC_6_257 b_6 NI_6 NS_257 0 7.3705220794178337e-05
GC_6_258 b_6 NI_6 NS_258 0 8.1377176446628900e-07
GC_6_259 b_6 NI_6 NS_259 0 -1.6021262781592606e-05
GC_6_260 b_6 NI_6 NS_260 0 2.6079713653264403e-04
GC_6_261 b_6 NI_6 NS_261 0 3.6483923862603917e-04
GC_6_262 b_6 NI_6 NS_262 0 -2.4267030115152232e-04
GC_6_263 b_6 NI_6 NS_263 0 6.5700688792376432e-05
GC_6_264 b_6 NI_6 NS_264 0 -2.8179946309243476e-05
GC_6_265 b_6 NI_6 NS_265 0 2.0799814233101970e-04
GC_6_266 b_6 NI_6 NS_266 0 -2.4118641771770299e-04
GC_6_267 b_6 NI_6 NS_267 0 -7.1054866303209331e-05
GC_6_268 b_6 NI_6 NS_268 0 -7.1872563795687225e-05
GC_6_269 b_6 NI_6 NS_269 0 6.4713639744293268e-05
GC_6_270 b_6 NI_6 NS_270 0 -7.5159631385643411e-05
GC_6_271 b_6 NI_6 NS_271 0 -1.7059831812829158e-04
GC_6_272 b_6 NI_6 NS_272 0 -1.8330408566816754e-04
GC_6_273 b_6 NI_6 NS_273 0 -4.8748184805615901e-05
GC_6_274 b_6 NI_6 NS_274 0 -1.9418952382699223e-05
GC_6_275 b_6 NI_6 NS_275 0 -1.4455356566856845e-04
GC_6_276 b_6 NI_6 NS_276 0 -9.5394431626107823e-05
GC_6_277 b_6 NI_6 NS_277 0 -2.7691635109998453e-05
GC_6_278 b_6 NI_6 NS_278 0 1.0379604914975364e-04
GC_6_279 b_6 NI_6 NS_279 0 -2.7256719908858158e-05
GC_6_280 b_6 NI_6 NS_280 0 1.3718670016430038e-05
GC_6_281 b_6 NI_6 NS_281 0 2.3523424080992041e-06
GC_6_282 b_6 NI_6 NS_282 0 5.0801561545545480e-05
GC_6_283 b_6 NI_6 NS_283 0 1.6821087314061997e-05
GC_6_284 b_6 NI_6 NS_284 0 -4.6980927479556252e-07
GC_6_285 b_6 NI_6 NS_285 0 1.7928529627305196e-06
GC_6_286 b_6 NI_6 NS_286 0 -1.5479232675569013e-05
GC_6_287 b_6 NI_6 NS_287 0 -1.4962774714117813e-05
GC_6_288 b_6 NI_6 NS_288 0 -1.3717819235812415e-05
GC_6_289 b_6 NI_6 NS_289 0 -1.2980734800636639e-05
GC_6_290 b_6 NI_6 NS_290 0 1.2292198345894048e-05
GC_6_291 b_6 NI_6 NS_291 0 7.7931171930762812e-06
GC_6_292 b_6 NI_6 NS_292 0 1.2794676169096903e-06
GC_6_293 b_6 NI_6 NS_293 0 -5.1332453849388358e-06
GC_6_294 b_6 NI_6 NS_294 0 -1.2738560750606821e-05
GC_6_295 b_6 NI_6 NS_295 0 -2.0684795124414265e-05
GC_6_296 b_6 NI_6 NS_296 0 -5.9665468130640008e-06
GC_6_297 b_6 NI_6 NS_297 0 1.1819040472549766e-06
GC_6_298 b_6 NI_6 NS_298 0 2.1730414503038183e-05
GC_6_299 b_6 NI_6 NS_299 0 1.2900858380811721e-05
GC_6_300 b_6 NI_6 NS_300 0 -6.8760461060615192e-06
GC_6_301 b_6 NI_6 NS_301 0 -1.7239529500358760e-05
GC_6_302 b_6 NI_6 NS_302 0 -1.6085703129405644e-05
GC_6_303 b_6 NI_6 NS_303 0 -2.7001164672358822e-05
GC_6_304 b_6 NI_6 NS_304 0 8.7822995036184545e-06
GC_6_305 b_6 NI_6 NS_305 0 2.7182342780655655e-05
GC_6_306 b_6 NI_6 NS_306 0 2.2285113098474868e-05
GC_6_307 b_6 NI_6 NS_307 0 1.1015441453869381e-05
GC_6_308 b_6 NI_6 NS_308 0 -2.1370449312243821e-05
GC_6_309 b_6 NI_6 NS_309 0 -3.0546883461561383e-05
GC_6_310 b_6 NI_6 NS_310 0 3.7167535851965737e-06
GC_6_311 b_6 NI_6 NS_311 0 -9.5362996097765346e-06
GC_6_312 b_6 NI_6 NS_312 0 3.9206783737611231e-05
GC_6_313 b_6 NI_6 NS_313 0 1.8475870824928794e-05
GC_6_314 b_6 NI_6 NS_314 0 -6.8312003710643791e-05
GC_6_315 b_6 NI_6 NS_315 0 4.3335413356248404e-05
GC_6_316 b_6 NI_6 NS_316 0 -1.7301382280612726e-05
GC_6_317 b_6 NI_6 NS_317 0 1.9835697952987444e-07
GC_6_318 b_6 NI_6 NS_318 0 -2.4920152709344818e-07
GC_6_319 b_6 NI_6 NS_319 0 -3.6902306344177573e-06
GC_6_320 b_6 NI_6 NS_320 0 -2.1085259586667824e-05
GC_6_321 b_6 NI_6 NS_321 0 -1.0619037346988501e-05
GC_6_322 b_6 NI_6 NS_322 0 1.6525274164308984e-05
GC_6_323 b_6 NI_6 NS_323 0 9.4041738316938413e-06
GC_6_324 b_6 NI_6 NS_324 0 3.1755351788998414e-05
GC_6_325 b_6 NI_6 NS_325 0 1.4484099630514317e-05
GC_6_326 b_6 NI_6 NS_326 0 -3.2769465151681074e-06
GC_6_327 b_6 NI_6 NS_327 0 -3.8735042578730275e-06
GC_6_328 b_6 NI_6 NS_328 0 1.2514301901764475e-05
GC_6_329 b_6 NI_6 NS_329 0 -1.8541636231517283e-05
GC_6_330 b_6 NI_6 NS_330 0 -3.5705385275779103e-06
GC_6_331 b_6 NI_6 NS_331 0 1.3189368067071406e-05
GC_6_332 b_6 NI_6 NS_332 0 1.3199058329263715e-05
GC_6_333 b_6 NI_6 NS_333 0 7.6290957955450738e-06
GC_6_334 b_6 NI_6 NS_334 0 -2.3004370043197377e-05
GC_6_335 b_6 NI_6 NS_335 0 -3.8544197275024396e-06
GC_6_336 b_6 NI_6 NS_336 0 -1.1714514700122241e-05
GC_6_337 b_6 NI_6 NS_337 0 -8.7383925756588958e-06
GC_6_338 b_6 NI_6 NS_338 0 -2.6219006542583555e-06
GC_6_339 b_6 NI_6 NS_339 0 5.5124511635412701e-10
GC_6_340 b_6 NI_6 NS_340 0 2.9329249742701159e-10
GC_6_341 b_6 NI_6 NS_341 0 4.2110179087631447e-08
GC_6_342 b_6 NI_6 NS_342 0 3.6978461741640886e-08
GC_6_343 b_6 NI_6 NS_343 0 3.0649011568140226e-04
GC_6_344 b_6 NI_6 NS_344 0 -1.4375817923524661e-05
GC_6_345 b_6 NI_6 NS_345 0 -1.2385100341500104e-09
GC_6_346 b_6 NI_6 NS_346 0 -1.9194463860806588e-08
GC_6_347 b_6 NI_6 NS_347 0 3.1995092094640503e-06
GC_6_348 b_6 NI_6 NS_348 0 -3.9682765746908864e-06
GC_6_349 b_6 NI_6 NS_349 0 -1.2574826046013604e-05
GC_6_350 b_6 NI_6 NS_350 0 -1.0246051903399496e-06
GC_6_351 b_6 NI_6 NS_351 0 3.9886438442920930e-05
GC_6_352 b_6 NI_6 NS_352 0 8.6693123462557758e-07
GC_6_353 b_6 NI_6 NS_353 0 -4.2799425036890471e-05
GC_6_354 b_6 NI_6 NS_354 0 -2.4449725321246623e-05
GC_6_355 b_6 NI_6 NS_355 0 1.1879748166074783e-06
GC_6_356 b_6 NI_6 NS_356 0 4.3287498219921517e-05
GC_6_357 b_6 NI_6 NS_357 0 1.0659388275690759e-05
GC_6_358 b_6 NI_6 NS_358 0 -4.8918960787292568e-05
GC_6_359 b_6 NI_6 NS_359 0 2.9240468151127566e-06
GC_6_360 b_6 NI_6 NS_360 0 6.2438629693545048e-06
GC_6_361 b_6 NI_6 NS_361 0 -4.5617839235685449e-05
GC_6_362 b_6 NI_6 NS_362 0 1.8881731452199659e-06
GC_6_363 b_6 NI_6 NS_363 0 1.0003674527520744e-04
GC_6_364 b_6 NI_6 NS_364 0 1.2285988338553864e-04
GC_6_365 b_6 NI_6 NS_365 0 -7.5037904137923594e-05
GC_6_366 b_6 NI_6 NS_366 0 -1.3519685095232968e-04
GC_6_367 b_6 NI_6 NS_367 0 -6.7762987642152041e-05
GC_6_368 b_6 NI_6 NS_368 0 4.9170696746967472e-05
GC_6_369 b_6 NI_6 NS_369 0 1.3378660856916194e-04
GC_6_370 b_6 NI_6 NS_370 0 -2.6377113959114133e-05
GC_6_371 b_6 NI_6 NS_371 0 -8.7279467970655258e-05
GC_6_372 b_6 NI_6 NS_372 0 -1.1629395608239069e-05
GC_6_373 b_6 NI_6 NS_373 0 -9.6761215501000905e-05
GC_6_374 b_6 NI_6 NS_374 0 2.1083875744212584e-04
GC_6_375 b_6 NI_6 NS_375 0 1.6568017263390885e-04
GC_6_376 b_6 NI_6 NS_376 0 -2.1189014081227875e-04
GC_6_377 b_6 NI_6 NS_377 0 -8.1910387912064998e-05
GC_6_378 b_6 NI_6 NS_378 0 1.9157070531825873e-05
GC_6_379 b_6 NI_6 NS_379 0 1.6054550630096706e-04
GC_6_380 b_6 NI_6 NS_380 0 4.4267036256209022e-05
GC_6_381 b_6 NI_6 NS_381 0 -8.8293783631838947e-05
GC_6_382 b_6 NI_6 NS_382 0 -7.2083231971925536e-05
GC_6_383 b_6 NI_6 NS_383 0 -8.5464792061992634e-05
GC_6_384 b_6 NI_6 NS_384 0 6.3490320429460787e-05
GC_6_385 b_6 NI_6 NS_385 0 1.4126735068420898e-04
GC_6_386 b_6 NI_6 NS_386 0 -4.6884427786891157e-05
GC_6_387 b_6 NI_6 NS_387 0 -6.6094061620913729e-05
GC_6_388 b_6 NI_6 NS_388 0 -2.4355974498980151e-05
GC_6_389 b_6 NI_6 NS_389 0 6.0403145019141326e-05
GC_6_390 b_6 NI_6 NS_390 0 1.1474521655020386e-04
GC_6_391 b_6 NI_6 NS_391 0 -2.2018823140410008e-05
GC_6_392 b_6 NI_6 NS_392 0 -1.2143064060892460e-04
GC_6_393 b_6 NI_6 NS_393 0 -4.4471467095189203e-05
GC_6_394 b_6 NI_6 NS_394 0 1.0923645353414605e-05
GC_6_395 b_6 NI_6 NS_395 0 4.7465213375204489e-05
GC_6_396 b_6 NI_6 NS_396 0 -9.9250316061151325e-06
GC_6_397 b_6 NI_6 NS_397 0 -3.2079696418122039e-05
GC_6_398 b_6 NI_6 NS_398 0 -7.5861024012300463e-06
GC_6_399 b_6 NI_6 NS_399 0 2.1298742222753475e-05
GC_6_400 b_6 NI_6 NS_400 0 -4.6124677725614252e-06
GC_6_401 b_6 NI_6 NS_401 0 -3.2316439417008971e-05
GC_6_402 b_6 NI_6 NS_402 0 -2.5188454677234861e-05
GC_6_403 b_6 NI_6 NS_403 0 1.2511646400606411e-05
GC_6_404 b_6 NI_6 NS_404 0 6.5127529663205033e-06
GC_6_405 b_6 NI_6 NS_405 0 -2.0423934944665891e-05
GC_6_406 b_6 NI_6 NS_406 0 -7.6317417885396732e-06
GC_6_407 b_6 NI_6 NS_407 0 1.3991873400459053e-05
GC_6_408 b_6 NI_6 NS_408 0 -1.2277806987148266e-05
GC_6_409 b_6 NI_6 NS_409 0 -4.1514157232219387e-05
GC_6_410 b_6 NI_6 NS_410 0 -1.6952621529593864e-05
GC_6_411 b_6 NI_6 NS_411 0 1.1564885983757774e-05
GC_6_412 b_6 NI_6 NS_412 0 -1.4317471345907240e-06
GC_6_413 b_6 NI_6 NS_413 0 -3.0400739425575863e-05
GC_6_414 b_6 NI_6 NS_414 0 5.6250440257640977e-06
GC_6_415 b_6 NI_6 NS_415 0 1.6017175635959856e-05
GC_6_416 b_6 NI_6 NS_416 0 -2.0571747385402424e-05
GC_6_417 b_6 NI_6 NS_417 0 -5.0238950786053664e-05
GC_6_418 b_6 NI_6 NS_418 0 -1.7712107646080508e-06
GC_6_419 b_6 NI_6 NS_419 0 1.1586540402757849e-05
GC_6_420 b_6 NI_6 NS_420 0 -1.1192316510744958e-05
GC_6_421 b_6 NI_6 NS_421 0 -3.2362722016465725e-05
GC_6_422 b_6 NI_6 NS_422 0 2.5180888667828709e-05
GC_6_423 b_6 NI_6 NS_423 0 1.0238942192233166e-05
GC_6_424 b_6 NI_6 NS_424 0 -3.5897417274142958e-05
GC_6_425 b_6 NI_6 NS_425 0 -3.4867044696462863e-05
GC_6_426 b_6 NI_6 NS_426 0 1.8379101490889946e-05
GC_6_427 b_6 NI_6 NS_427 0 -5.6371127018361011e-05
GC_6_428 b_6 NI_6 NS_428 0 1.3313684165777189e-04
GC_6_429 b_6 NI_6 NS_429 0 -1.5277007312846139e-05
GC_6_430 b_6 NI_6 NS_430 0 -3.1721922232380093e-05
GC_6_431 b_6 NI_6 NS_431 0 -3.7761111382457722e-07
GC_6_432 b_6 NI_6 NS_432 0 3.9607623736698750e-07
GC_6_433 b_6 NI_6 NS_433 0 -2.0156817478431632e-05
GC_6_434 b_6 NI_6 NS_434 0 3.2120811481426594e-05
GC_6_435 b_6 NI_6 NS_435 0 -1.4301599752765425e-05
GC_6_436 b_6 NI_6 NS_436 0 -3.3397595497313907e-05
GC_6_437 b_6 NI_6 NS_437 0 -6.1607123258380034e-06
GC_6_438 b_6 NI_6 NS_438 0 5.1177451472368140e-06
GC_6_439 b_6 NI_6 NS_439 0 -2.1208239294884812e-05
GC_6_440 b_6 NI_6 NS_440 0 -6.5712465638575912e-05
GC_6_441 b_6 NI_6 NS_441 0 -9.1589658582704834e-06
GC_6_442 b_6 NI_6 NS_442 0 -2.0643900451616891e-05
GC_6_443 b_6 NI_6 NS_443 0 1.5019856418118165e-05
GC_6_444 b_6 NI_6 NS_444 0 2.2754441630860790e-05
GC_6_445 b_6 NI_6 NS_445 0 -6.7861489212176697e-06
GC_6_446 b_6 NI_6 NS_446 0 2.7711938674333513e-05
GC_6_447 b_6 NI_6 NS_447 0 -1.1040736293399200e-05
GC_6_448 b_6 NI_6 NS_448 0 -2.1529802587475341e-05
GC_6_449 b_6 NI_6 NS_449 0 -1.1040032853012634e-05
GC_6_450 b_6 NI_6 NS_450 0 2.3841805289329355e-05
GC_6_451 b_6 NI_6 NS_451 0 5.1225289505725196e-06
GC_6_452 b_6 NI_6 NS_452 0 -1.5323283156518190e-05
GC_6_453 b_6 NI_6 NS_453 0 -4.7531527344006197e-10
GC_6_454 b_6 NI_6 NS_454 0 -9.1476846523738587e-10
GC_6_455 b_6 NI_6 NS_455 0 -5.5313689758702332e-08
GC_6_456 b_6 NI_6 NS_456 0 7.4255355920546604e-09
GC_6_457 b_6 NI_6 NS_457 0 1.8114336726378237e-02
GC_6_458 b_6 NI_6 NS_458 0 6.7504950789270771e-03
GC_6_459 b_6 NI_6 NS_459 0 4.7195338559849647e-07
GC_6_460 b_6 NI_6 NS_460 0 1.4474468434174021e-06
GC_6_461 b_6 NI_6 NS_461 0 6.0855621012505454e-03
GC_6_462 b_6 NI_6 NS_462 0 1.8096380663553218e-03
GC_6_463 b_6 NI_6 NS_463 0 -6.0720566036892168e-03
GC_6_464 b_6 NI_6 NS_464 0 -6.1691169805710381e-04
GC_6_465 b_6 NI_6 NS_465 0 7.3059720479077064e-03
GC_6_466 b_6 NI_6 NS_466 0 -1.2857326416673347e-02
GC_6_467 b_6 NI_6 NS_467 0 8.4528504344314574e-03
GC_6_468 b_6 NI_6 NS_468 0 -2.4022241147047242e-04
GC_6_469 b_6 NI_6 NS_469 0 -9.6390200420795689e-03
GC_6_470 b_6 NI_6 NS_470 0 2.6170482566423084e-03
GC_6_471 b_6 NI_6 NS_471 0 -8.8462744979591855e-03
GC_6_472 b_6 NI_6 NS_472 0 -2.4392959822013820e-02
GC_6_473 b_6 NI_6 NS_473 0 -8.6513314638808137e-04
GC_6_474 b_6 NI_6 NS_474 0 4.1785829106014459e-03
GC_6_475 b_6 NI_6 NS_475 0 7.1897431411497006e-03
GC_6_476 b_6 NI_6 NS_476 0 -1.0341095893621919e-03
GC_6_477 b_6 NI_6 NS_477 0 -2.5138645072588950e-02
GC_6_478 b_6 NI_6 NS_478 0 4.8070865083379025e-03
GC_6_479 b_6 NI_6 NS_479 0 -1.9701009719807039e-02
GC_6_480 b_6 NI_6 NS_480 0 8.9744558209220253e-04
GC_6_481 b_6 NI_6 NS_481 0 1.0752500089229648e-02
GC_6_482 b_6 NI_6 NS_482 0 -2.7940120004926136e-03
GC_6_483 b_6 NI_6 NS_483 0 -4.8191103593353398e-03
GC_6_484 b_6 NI_6 NS_484 0 4.5027482262602128e-02
GC_6_485 b_6 NI_6 NS_485 0 -1.2658610976822868e-02
GC_6_486 b_6 NI_6 NS_486 0 -2.5616841623795901e-04
GC_6_487 b_6 NI_6 NS_487 0 1.5863247740453730e-02
GC_6_488 b_6 NI_6 NS_488 0 -4.0664544956435138e-03
GC_6_489 b_6 NI_6 NS_489 0 3.2252275281977195e-02
GC_6_490 b_6 NI_6 NS_490 0 1.8644583367589632e-02
GC_6_491 b_6 NI_6 NS_491 0 -1.2591689401929772e-02
GC_6_492 b_6 NI_6 NS_492 0 1.8232431906525104e-04
GC_6_493 b_6 NI_6 NS_493 0 1.7239503477483986e-02
GC_6_494 b_6 NI_6 NS_494 0 -3.5124347146081980e-02
GC_6_495 b_6 NI_6 NS_495 0 1.4036153295910738e-02
GC_6_496 b_6 NI_6 NS_496 0 4.7591216408185933e-03
GC_6_497 b_6 NI_6 NS_497 0 -1.4382232517467267e-02
GC_6_498 b_6 NI_6 NS_498 0 2.6525603918567918e-04
GC_6_499 b_6 NI_6 NS_499 0 -2.0118036411998018e-02
GC_6_500 b_6 NI_6 NS_500 0 -3.0219180480418165e-02
GC_6_501 b_6 NI_6 NS_501 0 1.0538961723180695e-02
GC_6_502 b_6 NI_6 NS_502 0 3.5722915431533422e-03
GC_6_503 b_6 NI_6 NS_503 0 -2.6760788520027837e-02
GC_6_504 b_6 NI_6 NS_504 0 1.1130949460103706e-02
GC_6_505 b_6 NI_6 NS_505 0 -1.4164599537369994e-02
GC_6_506 b_6 NI_6 NS_506 0 -2.5194340438023577e-03
GC_6_507 b_6 NI_6 NS_507 0 7.5549375462437215e-03
GC_6_508 b_6 NI_6 NS_508 0 1.5797736822532342e-03
GC_6_509 b_6 NI_6 NS_509 0 -8.4943300011940299e-04
GC_6_510 b_6 NI_6 NS_510 0 2.4400448231884354e-02
GC_6_511 b_6 NI_6 NS_511 0 -7.6205595722672066e-03
GC_6_512 b_6 NI_6 NS_512 0 2.8886210045845116e-04
GC_6_513 b_6 NI_6 NS_513 0 -5.5962819680513843e-04
GC_6_514 b_6 NI_6 NS_514 0 -5.5377887589299884e-03
GC_6_515 b_6 NI_6 NS_515 0 8.2746280902484051e-03
GC_6_516 b_6 NI_6 NS_516 0 7.0134873305525832e-03
GC_6_517 b_6 NI_6 NS_517 0 -7.1244862543303302e-04
GC_6_518 b_6 NI_6 NS_518 0 1.2089356154987857e-02
GC_6_519 b_6 NI_6 NS_519 0 -5.1470157612647106e-03
GC_6_520 b_6 NI_6 NS_520 0 -1.3515068051033914e-04
GC_6_521 b_6 NI_6 NS_521 0 -1.8292844590348980e-03
GC_6_522 b_6 NI_6 NS_522 0 -5.1716258721766781e-03
GC_6_523 b_6 NI_6 NS_523 0 9.2942847359328250e-03
GC_6_524 b_6 NI_6 NS_524 0 5.4122746528868027e-03
GC_6_525 b_6 NI_6 NS_525 0 3.5222357042379066e-03
GC_6_526 b_6 NI_6 NS_526 0 1.1687384805598805e-02
GC_6_527 b_6 NI_6 NS_527 0 -6.1347989585944819e-03
GC_6_528 b_6 NI_6 NS_528 0 1.4299478940445018e-03
GC_6_529 b_6 NI_6 NS_529 0 -2.8132867938864218e-03
GC_6_530 b_6 NI_6 NS_530 0 -7.3475979127943731e-03
GC_6_531 b_6 NI_6 NS_531 0 9.9612552254398547e-03
GC_6_532 b_6 NI_6 NS_532 0 3.3711876920198467e-03
GC_6_533 b_6 NI_6 NS_533 0 8.1789432230964746e-03
GC_6_534 b_6 NI_6 NS_534 0 1.0242406137098934e-02
GC_6_535 b_6 NI_6 NS_535 0 -6.9808979899865786e-03
GC_6_536 b_6 NI_6 NS_536 0 2.9381665597750604e-03
GC_6_537 b_6 NI_6 NS_537 0 -5.6228431035891752e-03
GC_6_538 b_6 NI_6 NS_538 0 -8.0956760510053367e-03
GC_6_539 b_6 NI_6 NS_539 0 9.8672997141965712e-03
GC_6_540 b_6 NI_6 NS_540 0 5.6094055159328809e-04
GC_6_541 b_6 NI_6 NS_541 0 -1.0918385564126758e-02
GC_6_542 b_6 NI_6 NS_542 0 1.2173680036568374e-02
GC_6_543 b_6 NI_6 NS_543 0 9.6705968610813695e-03
GC_6_544 b_6 NI_6 NS_544 0 5.0264789717576076e-03
GC_6_545 b_6 NI_6 NS_545 0 -1.9577711367124114e-05
GC_6_546 b_6 NI_6 NS_546 0 3.1186968928240080e-05
GC_6_547 b_6 NI_6 NS_547 0 -7.1178143638970419e-03
GC_6_548 b_6 NI_6 NS_548 0 4.4750802374604057e-03
GC_6_549 b_6 NI_6 NS_549 0 -7.6632719766099328e-03
GC_6_550 b_6 NI_6 NS_550 0 -5.3302228771389785e-03
GC_6_551 b_6 NI_6 NS_551 0 9.5221895684981569e-03
GC_6_552 b_6 NI_6 NS_552 0 -1.7151716787258886e-03
GC_6_553 b_6 NI_6 NS_553 0 1.2490577802569460e-02
GC_6_554 b_6 NI_6 NS_554 0 -1.3742794733717415e-03
GC_6_555 b_6 NI_6 NS_555 0 -5.0725003257807650e-03
GC_6_556 b_6 NI_6 NS_556 0 -2.7519126603801516e-03
GC_6_557 b_6 NI_6 NS_557 0 -2.2328908867392814e-03
GC_6_558 b_6 NI_6 NS_558 0 6.6013347722753595e-03
GC_6_559 b_6 NI_6 NS_559 0 8.9595364541943893e-03
GC_6_560 b_6 NI_6 NS_560 0 1.2929001117796933e-04
GC_6_561 b_6 NI_6 NS_561 0 1.2486928827837990e-02
GC_6_562 b_6 NI_6 NS_562 0 1.7755711650586708e-03
GC_6_563 b_6 NI_6 NS_563 0 -5.3764540243771194e-03
GC_6_564 b_6 NI_6 NS_564 0 4.1567508156257968e-03
GC_6_565 b_6 NI_6 NS_565 0 -1.8433719828635322e-03
GC_6_566 b_6 NI_6 NS_566 0 -5.6868606296735574e-03
GC_6_567 b_6 NI_6 NS_567 0 2.0788378680101645e-07
GC_6_568 b_6 NI_6 NS_568 0 -2.4508479457560462e-07
GC_6_569 b_6 NI_6 NS_569 0 -1.1508310640103534e-05
GC_6_570 b_6 NI_6 NS_570 0 1.8247241596861921e-05
GC_6_571 b_6 NI_6 NS_571 0 -1.2879678365302492e-02
GC_6_572 b_6 NI_6 NS_572 0 1.3854981435521057e-03
GC_6_573 b_6 NI_6 NS_573 0 -2.6205840285931289e-07
GC_6_574 b_6 NI_6 NS_574 0 -3.7467072111589030e-06
GC_6_575 b_6 NI_6 NS_575 0 -2.6867049565011604e-04
GC_6_576 b_6 NI_6 NS_576 0 4.6434734670184545e-04
GC_6_577 b_6 NI_6 NS_577 0 1.3324560954778317e-03
GC_6_578 b_6 NI_6 NS_578 0 5.3750026552126112e-04
GC_6_579 b_6 NI_6 NS_579 0 -2.7601137799872586e-03
GC_6_580 b_6 NI_6 NS_580 0 -8.2597320623793811e-04
GC_6_581 b_6 NI_6 NS_581 0 3.5364628675816283e-03
GC_6_582 b_6 NI_6 NS_582 0 2.5065924206227009e-03
GC_6_583 b_6 NI_6 NS_583 0 1.1567034688189696e-03
GC_6_584 b_6 NI_6 NS_584 0 -4.2275310405893692e-03
GC_6_585 b_6 NI_6 NS_585 0 -1.7809488407351775e-03
GC_6_586 b_6 NI_6 NS_586 0 2.6938524756479174e-03
GC_6_587 b_6 NI_6 NS_587 0 -3.0415706679788281e-04
GC_6_588 b_6 NI_6 NS_588 0 -1.8023628353797827e-04
GC_6_589 b_6 NI_6 NS_589 0 3.9634827786398704e-03
GC_6_590 b_6 NI_6 NS_590 0 2.8124748378237623e-04
GC_6_591 b_6 NI_6 NS_591 0 -7.5491934513208427e-03
GC_6_592 b_6 NI_6 NS_592 0 -1.3596114662986087e-02
GC_6_593 b_6 NI_6 NS_593 0 4.4801853133992764e-03
GC_6_594 b_6 NI_6 NS_594 0 1.3516142075965383e-02
GC_6_595 b_6 NI_6 NS_595 0 6.6864812775845666e-03
GC_6_596 b_6 NI_6 NS_596 0 -4.0243778214442945e-03
GC_6_597 b_6 NI_6 NS_597 0 -1.3410293820585199e-02
GC_6_598 b_6 NI_6 NS_598 0 7.8159675612468605e-04
GC_6_599 b_6 NI_6 NS_599 0 7.8563490498530526e-03
GC_6_600 b_6 NI_6 NS_600 0 1.8570197805252227e-03
GC_6_601 b_6 NI_6 NS_601 0 1.0427284400921158e-02
GC_6_602 b_6 NI_6 NS_602 0 -1.9666894873982640e-02
GC_6_603 b_6 NI_6 NS_603 0 -1.7708792995199098e-02
GC_6_604 b_6 NI_6 NS_604 0 1.9274355532093747e-02
GC_6_605 b_6 NI_6 NS_605 0 7.6729375833856136e-03
GC_6_606 b_6 NI_6 NS_606 0 -1.4539279044187810e-03
GC_6_607 b_6 NI_6 NS_607 0 -1.5685667411794307e-02
GC_6_608 b_6 NI_6 NS_608 0 -4.6645856315015591e-03
GC_6_609 b_6 NI_6 NS_609 0 8.1074590720908689e-03
GC_6_610 b_6 NI_6 NS_610 0 7.2499065554865556e-03
GC_6_611 b_6 NI_6 NS_611 0 8.0870969212275233e-03
GC_6_612 b_6 NI_6 NS_612 0 -6.0421280239948182e-03
GC_6_613 b_6 NI_6 NS_613 0 -1.3963406797979428e-02
GC_6_614 b_6 NI_6 NS_614 0 4.6523180962955244e-03
GC_6_615 b_6 NI_6 NS_615 0 6.2461635398100481e-03
GC_6_616 b_6 NI_6 NS_616 0 2.3807834431027711e-03
GC_6_617 b_6 NI_6 NS_617 0 -6.3453822298409727e-03
GC_6_618 b_6 NI_6 NS_618 0 -1.1079792127784103e-02
GC_6_619 b_6 NI_6 NS_619 0 2.1863246186598290e-03
GC_6_620 b_6 NI_6 NS_620 0 1.1948129062760812e-02
GC_6_621 b_6 NI_6 NS_621 0 4.2064706907619497e-03
GC_6_622 b_6 NI_6 NS_622 0 -1.1782766738060943e-03
GC_6_623 b_6 NI_6 NS_623 0 -4.9335539115042491e-03
GC_6_624 b_6 NI_6 NS_624 0 1.0765974648074038e-03
GC_6_625 b_6 NI_6 NS_625 0 3.0283694698645287e-03
GC_6_626 b_6 NI_6 NS_626 0 6.9130860183735910e-04
GC_6_627 b_6 NI_6 NS_627 0 -2.2217202779696243e-03
GC_6_628 b_6 NI_6 NS_628 0 5.0249125625974030e-04
GC_6_629 b_6 NI_6 NS_629 0 3.0726777043807167e-03
GC_6_630 b_6 NI_6 NS_630 0 2.2985795667224392e-03
GC_6_631 b_6 NI_6 NS_631 0 -1.5387659365278582e-03
GC_6_632 b_6 NI_6 NS_632 0 -6.6609606018771877e-04
GC_6_633 b_6 NI_6 NS_633 0 1.8890921269302129e-03
GC_6_634 b_6 NI_6 NS_634 0 6.8214989017222364e-04
GC_6_635 b_6 NI_6 NS_635 0 -1.5634744905268791e-03
GC_6_636 b_6 NI_6 NS_636 0 1.2300996015769425e-03
GC_6_637 b_6 NI_6 NS_637 0 3.9777129314604023e-03
GC_6_638 b_6 NI_6 NS_638 0 1.4029334048311682e-03
GC_6_639 b_6 NI_6 NS_639 0 -1.5582664148641758e-03
GC_6_640 b_6 NI_6 NS_640 0 7.6117986197686913e-05
GC_6_641 b_6 NI_6 NS_641 0 2.8289093493877714e-03
GC_6_642 b_6 NI_6 NS_642 0 -6.8710722461214296e-04
GC_6_643 b_6 NI_6 NS_643 0 -1.8835386613863484e-03
GC_6_644 b_6 NI_6 NS_644 0 2.0120381834850959e-03
GC_6_645 b_6 NI_6 NS_645 0 4.9081291509085389e-03
GC_6_646 b_6 NI_6 NS_646 0 -1.8224322838839835e-04
GC_6_647 b_6 NI_6 NS_647 0 -1.6649329358344050e-03
GC_6_648 b_6 NI_6 NS_648 0 9.3127935401977164e-04
GC_6_649 b_6 NI_6 NS_649 0 3.0639848244451745e-03
GC_6_650 b_6 NI_6 NS_650 0 -2.8461931415294174e-03
GC_6_651 b_6 NI_6 NS_651 0 -1.4669285909377561e-03
GC_6_652 b_6 NI_6 NS_652 0 3.2252964315548712e-03
GC_6_653 b_6 NI_6 NS_653 0 3.7966903523392161e-03
GC_6_654 b_6 NI_6 NS_654 0 -2.9822010389947864e-03
GC_6_655 b_6 NI_6 NS_655 0 -1.8555106347963872e-03
GC_6_656 b_6 NI_6 NS_656 0 -3.8335466338409192e-03
GC_6_657 b_6 NI_6 NS_657 0 -4.1821452105519392e-04
GC_6_658 b_6 NI_6 NS_658 0 2.3792558667108952e-03
GC_6_659 b_6 NI_6 NS_659 0 -1.0537476773856996e-05
GC_6_660 b_6 NI_6 NS_660 0 -2.1101151455955165e-05
GC_6_661 b_6 NI_6 NS_661 0 8.3840691106141748e-04
GC_6_662 b_6 NI_6 NS_662 0 -3.7904942194814180e-03
GC_6_663 b_6 NI_6 NS_663 0 3.3771146868055366e-04
GC_6_664 b_6 NI_6 NS_664 0 3.3559401036935654e-03
GC_6_665 b_6 NI_6 NS_665 0 1.3516114980381638e-03
GC_6_666 b_6 NI_6 NS_666 0 -2.3818192054469644e-03
GC_6_667 b_6 NI_6 NS_667 0 2.1706665097617436e-03
GC_6_668 b_6 NI_6 NS_668 0 3.3305719674323908e-03
GC_6_669 b_6 NI_6 NS_669 0 1.1698297471200250e-03
GC_6_670 b_6 NI_6 NS_670 0 2.4039661728071462e-03
GC_6_671 b_6 NI_6 NS_671 0 -8.0769620187296290e-04
GC_6_672 b_6 NI_6 NS_672 0 -1.9803365764637011e-03
GC_6_673 b_6 NI_6 NS_673 0 3.9764634565289062e-04
GC_6_674 b_6 NI_6 NS_674 0 -2.6820418370234818e-03
GC_6_675 b_6 NI_6 NS_675 0 9.8318212604539611e-04
GC_6_676 b_6 NI_6 NS_676 0 2.7477883096375484e-03
GC_6_677 b_6 NI_6 NS_677 0 1.0389073299063981e-03
GC_6_678 b_6 NI_6 NS_678 0 -2.4201775721065136e-03
GC_6_679 b_6 NI_6 NS_679 0 -1.0840515955757514e-03
GC_6_680 b_6 NI_6 NS_680 0 1.5933774281620492e-03
GC_6_681 b_6 NI_6 NS_681 0 -1.0741032327255962e-08
GC_6_682 b_6 NI_6 NS_682 0 -2.7692023162416547e-09
GC_6_683 b_6 NI_6 NS_683 0 2.2912277515828723e-06
GC_6_684 b_6 NI_6 NS_684 0 5.4762400252624081e-07
GC_6_685 b_6 NI_6 NS_685 0 3.0950382312358348e-03
GC_6_686 b_6 NI_6 NS_686 0 -6.1289419798521319e-04
GC_6_687 b_6 NI_6 NS_687 0 2.8121768878839131e-08
GC_6_688 b_6 NI_6 NS_688 0 -3.1528677817600243e-08
GC_6_689 b_6 NI_6 NS_689 0 2.0500748585094983e-04
GC_6_690 b_6 NI_6 NS_690 0 1.3546525477488530e-04
GC_6_691 b_6 NI_6 NS_691 0 5.6415243191910817e-04
GC_6_692 b_6 NI_6 NS_692 0 2.6382416820019744e-04
GC_6_693 b_6 NI_6 NS_693 0 3.0949145134964461e-03
GC_6_694 b_6 NI_6 NS_694 0 -2.2211768851412165e-03
GC_6_695 b_6 NI_6 NS_695 0 -1.5948048524675490e-03
GC_6_696 b_6 NI_6 NS_696 0 -2.6831565094566677e-03
GC_6_697 b_6 NI_6 NS_697 0 -2.0664402392753137e-03
GC_6_698 b_6 NI_6 NS_698 0 -3.7810164178167459e-03
GC_6_699 b_6 NI_6 NS_699 0 -4.9930244901123036e-03
GC_6_700 b_6 NI_6 NS_700 0 -1.5154927482942545e-03
GC_6_701 b_6 NI_6 NS_701 0 2.9714191439280416e-04
GC_6_702 b_6 NI_6 NS_702 0 1.9409431795050511e-04
GC_6_703 b_6 NI_6 NS_703 0 -2.8708433682436492e-03
GC_6_704 b_6 NI_6 NS_704 0 -9.4557921921435803e-04
GC_6_705 b_6 NI_6 NS_705 0 -2.2198356736887599e-02
GC_6_706 b_6 NI_6 NS_706 0 -1.0125160141378329e-02
GC_6_707 b_6 NI_6 NS_707 0 1.2231820575138205e-03
GC_6_708 b_6 NI_6 NS_708 0 2.0396448737431221e-02
GC_6_709 b_6 NI_6 NS_709 0 -5.8225961277874978e-03
GC_6_710 b_6 NI_6 NS_710 0 4.6364315826257912e-03
GC_6_711 b_6 NI_6 NS_711 0 5.8808211908528488e-03
GC_6_712 b_6 NI_6 NS_712 0 3.4493742857532289e-02
GC_6_713 b_6 NI_6 NS_713 0 8.0480773190338330e-03
GC_6_714 b_6 NI_6 NS_714 0 2.7589344816132395e-03
GC_6_715 b_6 NI_6 NS_715 0 -7.6367946407707851e-03
GC_6_716 b_6 NI_6 NS_716 0 2.9591949309510923e-02
GC_6_717 b_6 NI_6 NS_717 0 5.0679464028395106e-02
GC_6_718 b_6 NI_6 NS_718 0 -2.0315742013374386e-02
GC_6_719 b_6 NI_6 NS_719 0 7.9122593953820479e-03
GC_6_720 b_6 NI_6 NS_720 0 -1.6718964658466130e-03
GC_6_721 b_6 NI_6 NS_721 0 2.8952184056961927e-02
GC_6_722 b_6 NI_6 NS_722 0 -2.6605127391588643e-02
GC_6_723 b_6 NI_6 NS_723 0 -6.7717827268786619e-03
GC_6_724 b_6 NI_6 NS_724 0 -9.8521000025668815e-03
GC_6_725 b_6 NI_6 NS_725 0 8.4245545407999993e-03
GC_6_726 b_6 NI_6 NS_726 0 -8.0661008711107925e-03
GC_6_727 b_6 NI_6 NS_727 0 -1.9120468064156206e-02
GC_6_728 b_6 NI_6 NS_728 0 -2.5143594558669744e-02
GC_6_729 b_6 NI_6 NS_729 0 -5.4851139330865679e-03
GC_6_730 b_6 NI_6 NS_730 0 -2.8303873467052537e-03
GC_6_731 b_6 NI_6 NS_731 0 -1.7803813480559819e-02
GC_6_732 b_6 NI_6 NS_732 0 -1.3047347988247594e-02
GC_6_733 b_6 NI_6 NS_733 0 -4.7610269326944302e-03
GC_6_734 b_6 NI_6 NS_734 0 1.2568312262639526e-02
GC_6_735 b_6 NI_6 NS_735 0 -3.4539894384810407e-03
GC_6_736 b_6 NI_6 NS_736 0 1.5560262362348150e-03
GC_6_737 b_6 NI_6 NS_737 0 -6.8744234581335681e-04
GC_6_738 b_6 NI_6 NS_738 0 7.0157646921948941e-03
GC_6_739 b_6 NI_6 NS_739 0 1.8840814926340055e-03
GC_6_740 b_6 NI_6 NS_740 0 8.1060298282552100e-05
GC_6_741 b_6 NI_6 NS_741 0 3.0821871518978410e-04
GC_6_742 b_6 NI_6 NS_742 0 -1.9474453973633067e-03
GC_6_743 b_6 NI_6 NS_743 0 -1.8615157413656570e-03
GC_6_744 b_6 NI_6 NS_744 0 -1.6133457408893396e-03
GC_6_745 b_6 NI_6 NS_745 0 -2.1255689202463648e-03
GC_6_746 b_6 NI_6 NS_746 0 1.6940535316767151e-03
GC_6_747 b_6 NI_6 NS_747 0 7.6441490542901956e-04
GC_6_748 b_6 NI_6 NS_748 0 1.8569494676258749e-04
GC_6_749 b_6 NI_6 NS_749 0 -7.0068891017052899e-04
GC_6_750 b_6 NI_6 NS_750 0 -1.6760053666460058e-03
GC_6_751 b_6 NI_6 NS_751 0 -2.6855348527751056e-03
GC_6_752 b_6 NI_6 NS_752 0 -8.2394361514492246e-04
GC_6_753 b_6 NI_6 NS_753 0 -4.9849815543533745e-04
GC_6_754 b_6 NI_6 NS_754 0 2.9352185660264530e-03
GC_6_755 b_6 NI_6 NS_755 0 1.3528913556508026e-03
GC_6_756 b_6 NI_6 NS_756 0 -8.5706965935815045e-04
GC_6_757 b_6 NI_6 NS_757 0 -2.4223431242854049e-03
GC_6_758 b_6 NI_6 NS_758 0 -2.2652839991051110e-03
GC_6_759 b_6 NI_6 NS_759 0 -3.5590208528511838e-03
GC_6_760 b_6 NI_6 NS_760 0 7.4879929799389179e-04
GC_6_761 b_6 NI_6 NS_761 0 2.4605503807920157e-03
GC_6_762 b_6 NI_6 NS_762 0 3.0265640475578299e-03
GC_6_763 b_6 NI_6 NS_763 0 9.8335663828499247e-04
GC_6_764 b_6 NI_6 NS_764 0 -2.9400791630671023e-03
GC_6_765 b_6 NI_6 NS_765 0 -4.7724963150962184e-03
GC_6_766 b_6 NI_6 NS_766 0 5.7213286454470044e-05
GC_6_767 b_6 NI_6 NS_767 0 -1.7194828880382198e-03
GC_6_768 b_6 NI_6 NS_768 0 3.7113727647197681e-03
GC_6_769 b_6 NI_6 NS_769 0 -7.3866856711920408e-04
GC_6_770 b_6 NI_6 NS_770 0 1.5326975789382120e-03
GC_6_771 b_6 NI_6 NS_771 0 3.2195727687087785e-03
GC_6_772 b_6 NI_6 NS_772 0 -1.3350001774915094e-03
GC_6_773 b_6 NI_6 NS_773 0 -2.8023014575452787e-06
GC_6_774 b_6 NI_6 NS_774 0 8.9859617450905297e-06
GC_6_775 b_6 NI_6 NS_775 0 -1.8210613622819710e-03
GC_6_776 b_6 NI_6 NS_776 0 -2.5224011940836355e-03
GC_6_777 b_6 NI_6 NS_777 0 -2.4088305468615932e-03
GC_6_778 b_6 NI_6 NS_778 0 2.4933219626362391e-03
GC_6_779 b_6 NI_6 NS_779 0 1.0059044462660349e-03
GC_6_780 b_6 NI_6 NS_780 0 2.4239835194429511e-03
GC_6_781 b_6 NI_6 NS_781 0 8.4854758676541247e-04
GC_6_782 b_6 NI_6 NS_782 0 -2.6997877237450976e-03
GC_6_783 b_6 NI_6 NS_783 0 -3.0628340275732643e-04
GC_6_784 b_6 NI_6 NS_784 0 1.6736613987153562e-03
GC_6_785 b_6 NI_6 NS_785 0 -1.7824226315017089e-03
GC_6_786 b_6 NI_6 NS_786 0 -3.1430312550315115e-04
GC_6_787 b_6 NI_6 NS_787 0 1.3997487929992233e-03
GC_6_788 b_6 NI_6 NS_788 0 1.9719385103700712e-03
GC_6_789 b_6 NI_6 NS_789 0 1.0457174132094895e-03
GC_6_790 b_6 NI_6 NS_790 0 -2.2988261700395063e-03
GC_6_791 b_6 NI_6 NS_791 0 -6.9831750467137744e-04
GC_6_792 b_6 NI_6 NS_792 0 -1.4663462620118804e-03
GC_6_793 b_6 NI_6 NS_793 0 -1.3735955854149045e-03
GC_6_794 b_6 NI_6 NS_794 0 -3.1257035056182108e-04
GC_6_795 b_6 NI_6 NS_795 0 6.7938417477142257e-09
GC_6_796 b_6 NI_6 NS_796 0 -2.4700008532305917e-08
GC_6_797 b_6 NI_6 NS_797 0 -4.4377025843547366e-07
GC_6_798 b_6 NI_6 NS_798 0 1.6205765415415968e-06
GC_6_799 b_6 NI_6 NS_799 0 7.9886718564914586e-03
GC_6_800 b_6 NI_6 NS_800 0 -1.6009906145810682e-03
GC_6_801 b_6 NI_6 NS_801 0 -1.2329825278621210e-08
GC_6_802 b_6 NI_6 NS_802 0 -8.8365943549159953e-07
GC_6_803 b_6 NI_6 NS_803 0 1.0714040931158705e-04
GC_6_804 b_6 NI_6 NS_804 0 -5.1251769138420085e-04
GC_6_805 b_6 NI_6 NS_805 0 -1.9321158086619804e-03
GC_6_806 b_6 NI_6 NS_806 0 -5.9632008190260016e-04
GC_6_807 b_6 NI_6 NS_807 0 2.9522602799263277e-03
GC_6_808 b_6 NI_6 NS_808 0 2.2413628935615626e-03
GC_6_809 b_6 NI_6 NS_809 0 -3.5853198941042494e-03
GC_6_810 b_6 NI_6 NS_810 0 -3.0463419422841957e-03
GC_6_811 b_6 NI_6 NS_811 0 -1.6953804469390229e-03
GC_6_812 b_6 NI_6 NS_812 0 5.8334393047821814e-03
GC_6_813 b_6 NI_6 NS_813 0 4.3284000327929867e-03
GC_6_814 b_6 NI_6 NS_814 0 -2.4949638211468903e-03
GC_6_815 b_6 NI_6 NS_815 0 -1.0252417117198533e-04
GC_6_816 b_6 NI_6 NS_816 0 -9.7511923675885258e-05
GC_6_817 b_6 NI_6 NS_817 0 -4.4595016509466840e-03
GC_6_818 b_6 NI_6 NS_818 0 -9.0945578513100013e-04
GC_6_819 b_6 NI_6 NS_819 0 9.1489031894844020e-03
GC_6_820 b_6 NI_6 NS_820 0 1.7749054714789689e-02
GC_6_821 b_6 NI_6 NS_821 0 -4.0759917581847131e-03
GC_6_822 b_6 NI_6 NS_822 0 -1.7815996221333397e-02
GC_6_823 b_6 NI_6 NS_823 0 -8.2086049935102910e-03
GC_6_824 b_6 NI_6 NS_824 0 4.1974764955479910e-03
GC_6_825 b_6 NI_6 NS_825 0 1.7045926423172802e-02
GC_6_826 b_6 NI_6 NS_826 0 -4.7587324944727921e-04
GC_6_827 b_6 NI_6 NS_827 0 -9.2871622319565666e-03
GC_6_828 b_6 NI_6 NS_828 0 -3.1746356713083655e-03
GC_6_829 b_6 NI_6 NS_829 0 -1.3650847444386357e-02
GC_6_830 b_6 NI_6 NS_830 0 2.2873426936243200e-02
GC_6_831 b_6 NI_6 NS_831 0 2.2768615050962539e-02
GC_6_832 b_6 NI_6 NS_832 0 -2.2718066481022287e-02
GC_6_833 b_6 NI_6 NS_833 0 -9.2369617596561628e-03
GC_6_834 b_6 NI_6 NS_834 0 9.4042622161431659e-04
GC_6_835 b_6 NI_6 NS_835 0 1.8496821948025884e-02
GC_6_836 b_6 NI_6 NS_836 0 6.1966524489086711e-03
GC_6_837 b_6 NI_6 NS_837 0 -9.2042290956656121e-03
GC_6_838 b_6 NI_6 NS_838 0 -9.4288117675606926e-03
GC_6_839 b_6 NI_6 NS_839 0 -9.9569355407995441e-03
GC_6_840 b_6 NI_6 NS_840 0 6.4309790701951178e-03
GC_6_841 b_6 NI_6 NS_841 0 1.6827172549741917e-02
GC_6_842 b_6 NI_6 NS_842 0 -4.8950436122962970e-03
GC_6_843 b_6 NI_6 NS_843 0 -7.2263300997448031e-03
GC_6_844 b_6 NI_6 NS_844 0 -3.3851923813650975e-03
GC_6_845 b_6 NI_6 NS_845 0 6.8657294741519279e-03
GC_6_846 b_6 NI_6 NS_846 0 1.3286490499937905e-02
GC_6_847 b_6 NI_6 NS_847 0 -1.8581882785385891e-03
GC_6_848 b_6 NI_6 NS_848 0 -1.4397044018698350e-02
GC_6_849 b_6 NI_6 NS_849 0 -4.9859100376690429e-03
GC_6_850 b_6 NI_6 NS_850 0 1.0545183003565538e-03
GC_6_851 b_6 NI_6 NS_851 0 6.0007405862819137e-03
GC_6_852 b_6 NI_6 NS_852 0 -1.1126545524495599e-03
GC_6_853 b_6 NI_6 NS_853 0 -3.4683253358492178e-03
GC_6_854 b_6 NI_6 NS_854 0 -1.0780499139734631e-03
GC_6_855 b_6 NI_6 NS_855 0 2.7173467256017179e-03
GC_6_856 b_6 NI_6 NS_856 0 -5.1095685074015369e-04
GC_6_857 b_6 NI_6 NS_857 0 -3.3053412645821360e-03
GC_6_858 b_6 NI_6 NS_858 0 -2.8885150443896733e-03
GC_6_859 b_6 NI_6 NS_859 0 2.0156340101056048e-03
GC_6_860 b_6 NI_6 NS_860 0 7.7768287534719764e-04
GC_6_861 b_6 NI_6 NS_861 0 -2.0192451140979666e-03
GC_6_862 b_6 NI_6 NS_862 0 -9.6218740591897441e-04
GC_6_863 b_6 NI_6 NS_863 0 2.1198804241646689e-03
GC_6_864 b_6 NI_6 NS_864 0 -1.4705676416475093e-03
GC_6_865 b_6 NI_6 NS_865 0 -4.1910213329290702e-03
GC_6_866 b_6 NI_6 NS_866 0 -1.8092507381325311e-03
GC_6_867 b_6 NI_6 NS_867 0 2.3672939675763033e-03
GC_6_868 b_6 NI_6 NS_868 0 -3.6739652409029675e-04
GC_6_869 b_6 NI_6 NS_869 0 -3.0199644098802153e-03
GC_6_870 b_6 NI_6 NS_870 0 4.6494719899224359e-04
GC_6_871 b_6 NI_6 NS_871 0 2.7038550460648783e-03
GC_6_872 b_6 NI_6 NS_872 0 -2.7263252651663740e-03
GC_6_873 b_6 NI_6 NS_873 0 -5.0450291676011286e-03
GC_6_874 b_6 NI_6 NS_874 0 -1.2988616567672113e-04
GC_6_875 b_6 NI_6 NS_875 0 2.4275289959737115e-03
GC_6_876 b_6 NI_6 NS_876 0 -2.1667278959752049e-03
GC_6_877 b_6 NI_6 NS_877 0 -3.2524101807385095e-03
GC_6_878 b_6 NI_6 NS_878 0 2.6001222878699486e-03
GC_6_879 b_6 NI_6 NS_879 0 1.7373703013879420e-03
GC_6_880 b_6 NI_6 NS_880 0 -4.7433400082752316e-03
GC_6_881 b_6 NI_6 NS_881 0 -3.6476875040186317e-03
GC_6_882 b_6 NI_6 NS_882 0 2.5904971008593315e-03
GC_6_883 b_6 NI_6 NS_883 0 -2.8140501870579254e-03
GC_6_884 b_6 NI_6 NS_884 0 4.0553534120779710e-03
GC_6_885 b_6 NI_6 NS_885 0 -2.3077989557968603e-04
GC_6_886 b_6 NI_6 NS_886 0 -4.1951360849193280e-03
GC_6_887 b_6 NI_6 NS_887 0 -9.8757633350850921e-06
GC_6_888 b_6 NI_6 NS_888 0 7.9025145348525824e-06
GC_6_889 b_6 NI_6 NS_889 0 -1.3634151857812153e-03
GC_6_890 b_6 NI_6 NS_890 0 3.3837800441968188e-03
GC_6_891 b_6 NI_6 NS_891 0 -9.6978192790284936e-04
GC_6_892 b_6 NI_6 NS_892 0 -4.3384320717327141e-03
GC_6_893 b_6 NI_6 NS_893 0 -1.0095576030072948e-03
GC_6_894 b_6 NI_6 NS_894 0 2.2144692472069946e-03
GC_6_895 b_6 NI_6 NS_895 0 -1.6625797227517180e-03
GC_6_896 b_6 NI_6 NS_896 0 -4.4181655691939922e-03
GC_6_897 b_6 NI_6 NS_897 0 -1.4450239354741865e-03
GC_6_898 b_6 NI_6 NS_898 0 -2.4969806541893561e-03
GC_6_899 b_6 NI_6 NS_899 0 7.8582136017313418e-04
GC_6_900 b_6 NI_6 NS_900 0 2.5922239209250839e-03
GC_6_901 b_6 NI_6 NS_901 0 -6.9658839153502678e-04
GC_6_902 b_6 NI_6 NS_902 0 2.8805416668427936e-03
GC_6_903 b_6 NI_6 NS_903 0 -1.4341253084519639e-03
GC_6_904 b_6 NI_6 NS_904 0 -2.7701138559925145e-03
GC_6_905 b_6 NI_6 NS_905 0 -1.1685605973488871e-03
GC_6_906 b_6 NI_6 NS_906 0 2.6674409158219509e-03
GC_6_907 b_6 NI_6 NS_907 0 7.8095042677383999e-04
GC_6_908 b_6 NI_6 NS_908 0 -1.8732339653541421e-03
GC_6_909 b_6 NI_6 NS_909 0 2.4009828897753121e-08
GC_6_910 b_6 NI_6 NS_910 0 -6.0310105638829654e-08
GC_6_911 b_6 NI_6 NS_911 0 -9.0615471211111128e-07
GC_6_912 b_6 NI_6 NS_912 0 3.2140038478689535e-06
GC_6_913 b_6 NI_6 NS_913 0 -3.2390014039628252e-05
GC_6_914 b_6 NI_6 NS_914 0 2.2145968349391818e-06
GC_6_915 b_6 NI_6 NS_915 0 6.9003387352594335e-11
GC_6_916 b_6 NI_6 NS_916 0 3.0548368075514108e-09
GC_6_917 b_6 NI_6 NS_917 0 -1.7288682531183328e-06
GC_6_918 b_6 NI_6 NS_918 0 -1.8218362834602113e-06
GC_6_919 b_6 NI_6 NS_919 0 -5.3710550252048930e-06
GC_6_920 b_6 NI_6 NS_920 0 2.8657841161327751e-06
GC_6_921 b_6 NI_6 NS_921 0 -1.6530935200591124e-05
GC_6_922 b_6 NI_6 NS_922 0 1.8435252433085600e-05
GC_6_923 b_6 NI_6 NS_923 0 1.5105431235745000e-05
GC_6_924 b_6 NI_6 NS_924 0 9.7996111865068432e-06
GC_6_925 b_6 NI_6 NS_925 0 1.7319502694581448e-05
GC_6_926 b_6 NI_6 NS_926 0 2.2757394178505780e-05
GC_6_927 b_6 NI_6 NS_927 0 2.9272138518862999e-05
GC_6_928 b_6 NI_6 NS_928 0 4.9456580582277570e-06
GC_6_929 b_6 NI_6 NS_929 0 -3.0091214576145782e-06
GC_6_930 b_6 NI_6 NS_930 0 -1.8920517022208892e-06
GC_6_931 b_6 NI_6 NS_931 0 1.6961528848098054e-05
GC_6_932 b_6 NI_6 NS_932 0 -2.2247633847181243e-06
GC_6_933 b_6 NI_6 NS_933 0 1.2893963562138748e-04
GC_6_934 b_6 NI_6 NS_934 0 3.4692029990748484e-05
GC_6_935 b_6 NI_6 NS_935 0 -2.8903407554710220e-05
GC_6_936 b_6 NI_6 NS_936 0 -9.8807186007577794e-05
GC_6_937 b_6 NI_6 NS_937 0 2.4942415033236781e-05
GC_6_938 b_6 NI_6 NS_938 0 -3.1439755220338349e-05
GC_6_939 b_6 NI_6 NS_939 0 -4.1725646046785009e-05
GC_6_940 b_6 NI_6 NS_940 0 -1.6659190259712107e-04
GC_6_941 b_6 NI_6 NS_941 0 -4.1856506246658079e-05
GC_6_942 b_6 NI_6 NS_942 0 -4.9686962331088147e-06
GC_6_943 b_6 NI_6 NS_943 0 2.1526363423768432e-05
GC_6_944 b_6 NI_6 NS_944 0 -1.5189810226539369e-04
GC_6_945 b_6 NI_6 NS_945 0 -2.3067318505825529e-04
GC_6_946 b_6 NI_6 NS_946 0 1.1454500107577453e-04
GC_6_947 b_6 NI_6 NS_947 0 -3.7434333413019959e-05
GC_6_948 b_6 NI_6 NS_948 0 1.4285228464980720e-05
GC_6_949 b_6 NI_6 NS_949 0 -1.3769140869420373e-04
GC_6_950 b_6 NI_6 NS_950 0 1.3059617306283538e-04
GC_6_951 b_6 NI_6 NS_951 0 3.6482049042413936e-05
GC_6_952 b_6 NI_6 NS_952 0 4.1333283787605529e-05
GC_6_953 b_6 NI_6 NS_953 0 -3.8174085160099896e-05
GC_6_954 b_6 NI_6 NS_954 0 4.3297472102082107e-05
GC_6_955 b_6 NI_6 NS_955 0 8.7698357445220097e-05
GC_6_956 b_6 NI_6 NS_956 0 1.1839030779539430e-04
GC_6_957 b_6 NI_6 NS_957 0 2.7360612542350974e-05
GC_6_958 b_6 NI_6 NS_958 0 1.0188100382097638e-05
GC_6_959 b_6 NI_6 NS_959 0 8.7309716226071317e-05
GC_6_960 b_6 NI_6 NS_960 0 6.5588843902989925e-05
GC_6_961 b_6 NI_6 NS_961 0 2.0355359357981297e-05
GC_6_962 b_6 NI_6 NS_962 0 -5.7134032658953713e-05
GC_6_963 b_6 NI_6 NS_963 0 1.6985922200782407e-05
GC_6_964 b_6 NI_6 NS_964 0 -8.8834615292880465e-06
GC_6_965 b_6 NI_6 NS_965 0 8.5005626246362991e-06
GC_6_966 b_6 NI_6 NS_966 0 -3.2939559475869608e-05
GC_6_967 b_6 NI_6 NS_967 0 -8.8537845861441833e-06
GC_6_968 b_6 NI_6 NS_968 0 5.2634464415455461e-07
GC_6_969 b_6 NI_6 NS_969 0 -2.4131094009220924e-06
GC_6_970 b_6 NI_6 NS_970 0 8.5086288701673128e-06
GC_6_971 b_6 NI_6 NS_971 0 1.0220485698027697e-05
GC_6_972 b_6 NI_6 NS_972 0 6.0869789107552902e-06
GC_6_973 b_6 NI_6 NS_973 0 1.2161238146989670e-05
GC_6_974 b_6 NI_6 NS_974 0 -7.8265430245217932e-06
GC_6_975 b_6 NI_6 NS_975 0 -3.4879205658343131e-06
GC_6_976 b_6 NI_6 NS_976 0 -4.4672850085974351e-07
GC_6_977 b_6 NI_6 NS_977 0 2.4880740196761714e-06
GC_6_978 b_6 NI_6 NS_978 0 7.4078962050123298e-06
GC_6_979 b_6 NI_6 NS_979 0 1.3650682690915544e-05
GC_6_980 b_6 NI_6 NS_980 0 2.6358815458922924e-06
GC_6_981 b_6 NI_6 NS_981 0 4.5207259374290918e-06
GC_6_982 b_6 NI_6 NS_982 0 -1.4188658811183454e-05
GC_6_983 b_6 NI_6 NS_983 0 -5.9269896814877524e-06
GC_6_984 b_6 NI_6 NS_984 0 4.2582630527983580e-06
GC_6_985 b_6 NI_6 NS_985 0 1.0309894186695443e-05
GC_6_986 b_6 NI_6 NS_986 0 9.9374602338136075e-06
GC_6_987 b_6 NI_6 NS_987 0 1.7307677770632080e-05
GC_6_988 b_6 NI_6 NS_988 0 -4.2709456587488918e-06
GC_6_989 b_6 NI_6 NS_989 0 -9.2921107155477020e-06
GC_6_990 b_6 NI_6 NS_990 0 -1.5315722003550935e-05
GC_6_991 b_6 NI_6 NS_991 0 -4.0817827079819463e-06
GC_6_992 b_6 NI_6 NS_992 0 1.3516462742767822e-05
GC_6_993 b_6 NI_6 NS_993 0 2.0928883496707156e-05
GC_6_994 b_6 NI_6 NS_994 0 -5.6272698079524161e-07
GC_6_995 b_6 NI_6 NS_995 0 8.8752322769539971e-06
GC_6_996 b_6 NI_6 NS_996 0 -1.7452661177579576e-05
GC_6_997 b_6 NI_6 NS_997 0 2.4046519159941763e-06
GC_6_998 b_6 NI_6 NS_998 0 -1.3697816600924368e-05
GC_6_999 b_6 NI_6 NS_999 0 -1.3815730852452067e-05
GC_6_1000 b_6 NI_6 NS_1000 0 4.3766364382718171e-06
GC_6_1001 b_6 NI_6 NS_1001 0 1.5474698591371230e-08
GC_6_1002 b_6 NI_6 NS_1002 0 -4.2110169672286724e-08
GC_6_1003 b_6 NI_6 NS_1003 0 8.6210482478020084e-06
GC_6_1004 b_6 NI_6 NS_1004 0 1.1597858429387650e-05
GC_6_1005 b_6 NI_6 NS_1005 0 1.0904635273326424e-05
GC_6_1006 b_6 NI_6 NS_1006 0 -1.1278378645792159e-05
GC_6_1007 b_6 NI_6 NS_1007 0 -3.7306489925559210e-06
GC_6_1008 b_6 NI_6 NS_1008 0 -1.0216318601489494e-05
GC_6_1009 b_6 NI_6 NS_1009 0 -2.2939498007368056e-06
GC_6_1010 b_6 NI_6 NS_1010 0 1.2865849123138874e-05
GC_6_1011 b_6 NI_6 NS_1011 0 9.6692461205432523e-07
GC_6_1012 b_6 NI_6 NS_1012 0 -7.2694845896985628e-06
GC_6_1013 b_6 NI_6 NS_1013 0 7.5166670708700643e-06
GC_6_1014 b_6 NI_6 NS_1014 0 1.6932063938841812e-06
GC_6_1015 b_6 NI_6 NS_1015 0 -6.1012272786711993e-06
GC_6_1016 b_6 NI_6 NS_1016 0 -8.8953909081834784e-06
GC_6_1017 b_6 NI_6 NS_1017 0 -4.1215017348301262e-06
GC_6_1018 b_6 NI_6 NS_1018 0 9.6659695441382806e-06
GC_6_1019 b_6 NI_6 NS_1019 0 3.3268386126868005e-06
GC_6_1020 b_6 NI_6 NS_1020 0 6.0367148503069703e-06
GC_6_1021 b_6 NI_6 NS_1021 0 5.6518831888826545e-06
GC_6_1022 b_6 NI_6 NS_1022 0 5.1680977150041462e-07
GC_6_1023 b_6 NI_6 NS_1023 0 6.1805231258568372e-11
GC_6_1024 b_6 NI_6 NS_1024 0 1.4894745424933786e-10
GC_6_1025 b_6 NI_6 NS_1025 0 5.9431479387531336e-09
GC_6_1026 b_6 NI_6 NS_1026 0 -8.3385319270295699e-09
GC_6_1027 b_6 NI_6 NS_1027 0 -1.1661777288417189e-04
GC_6_1028 b_6 NI_6 NS_1028 0 -2.1401249863265484e-06
GC_6_1029 b_6 NI_6 NS_1029 0 -2.5040563395500051e-10
GC_6_1030 b_6 NI_6 NS_1030 0 2.6003943407366943e-09
GC_6_1031 b_6 NI_6 NS_1031 0 1.7091685439947068e-06
GC_6_1032 b_6 NI_6 NS_1032 0 -1.5815004738969752e-06
GC_6_1033 b_6 NI_6 NS_1033 0 1.2865051068519264e-07
GC_6_1034 b_6 NI_6 NS_1034 0 -6.3839769896420464e-06
GC_6_1035 b_6 NI_6 NS_1035 0 -7.6493576643321340e-06
GC_6_1036 b_6 NI_6 NS_1036 0 1.1913597516753361e-07
GC_6_1037 b_6 NI_6 NS_1037 0 -1.2236191159811348e-06
GC_6_1038 b_6 NI_6 NS_1038 0 -4.6177283043391817e-06
GC_6_1039 b_6 NI_6 NS_1039 0 -1.5901242919148968e-05
GC_6_1040 b_6 NI_6 NS_1040 0 -1.6609733378310446e-06
GC_6_1041 b_6 NI_6 NS_1041 0 -6.2265113072427868e-06
GC_6_1042 b_6 NI_6 NS_1042 0 1.9173247687082512e-05
GC_6_1043 b_6 NI_6 NS_1043 0 4.6915551938611535e-06
GC_6_1044 b_6 NI_6 NS_1044 0 -3.0032579975535514e-06
GC_6_1045 b_6 NI_6 NS_1045 0 -1.8663087645730341e-08
GC_6_1046 b_6 NI_6 NS_1046 0 -2.5775024901231838e-06
GC_6_1047 b_6 NI_6 NS_1047 0 -2.5961794166318029e-05
GC_6_1048 b_6 NI_6 NS_1048 0 2.8474538110682057e-05
GC_6_1049 b_6 NI_6 NS_1049 0 2.8294920597577886e-05
GC_6_1050 b_6 NI_6 NS_1050 0 -8.4647889953265115e-06
GC_6_1051 b_6 NI_6 NS_1051 0 -8.0582938112588949e-06
GC_6_1052 b_6 NI_6 NS_1052 0 -4.3213664382356313e-06
GC_6_1053 b_6 NI_6 NS_1053 0 1.2613103596079510e-05
GC_6_1054 b_6 NI_6 NS_1054 0 2.7036770171985527e-05
GC_6_1055 b_6 NI_6 NS_1055 0 1.4849126722964096e-06
GC_6_1056 b_6 NI_6 NS_1056 0 -8.9982177050187218e-06
GC_6_1057 b_6 NI_6 NS_1057 0 -2.8357601096665819e-05
GC_6_1058 b_6 NI_6 NS_1058 0 4.7238549320635328e-06
GC_6_1059 b_6 NI_6 NS_1059 0 4.1379064272345582e-05
GC_6_1060 b_6 NI_6 NS_1060 0 1.0729943250848588e-05
GC_6_1061 b_6 NI_6 NS_1061 0 -2.9667043876590270e-06
GC_6_1062 b_6 NI_6 NS_1062 0 -4.4978586788244620e-06
GC_6_1063 b_6 NI_6 NS_1063 0 1.2948378235430439e-05
GC_6_1064 b_6 NI_6 NS_1064 0 1.9022646968629201e-05
GC_6_1065 b_6 NI_6 NS_1065 0 3.8280367364778569e-06
GC_6_1066 b_6 NI_6 NS_1066 0 -1.0937998111740748e-05
GC_6_1067 b_6 NI_6 NS_1067 0 -6.4224020386920832e-06
GC_6_1068 b_6 NI_6 NS_1068 0 8.3857918304212696e-07
GC_6_1069 b_6 NI_6 NS_1069 0 1.8903998409317655e-05
GC_6_1070 b_6 NI_6 NS_1070 0 5.4505926645612402e-06
GC_6_1071 b_6 NI_6 NS_1071 0 -6.6494122269438248e-08
GC_6_1072 b_6 NI_6 NS_1072 0 -4.1973566944006327e-06
GC_6_1073 b_6 NI_6 NS_1073 0 4.9149594553846668e-06
GC_6_1074 b_6 NI_6 NS_1074 0 1.4293061413939560e-05
GC_6_1075 b_6 NI_6 NS_1075 0 7.8466195127653290e-06
GC_6_1076 b_6 NI_6 NS_1076 0 -1.1186119751575346e-05
GC_6_1077 b_6 NI_6 NS_1077 0 -1.3863433165926810e-06
GC_6_1078 b_6 NI_6 NS_1078 0 9.3337897080481712e-07
GC_6_1079 b_6 NI_6 NS_1079 0 1.0911665092781772e-05
GC_6_1080 b_6 NI_6 NS_1080 0 4.1227353916960456e-06
GC_6_1081 b_6 NI_6 NS_1081 0 1.7223613792981994e-06
GC_6_1082 b_6 NI_6 NS_1082 0 -6.3594465334000803e-07
GC_6_1083 b_6 NI_6 NS_1083 0 5.6879435933700723e-06
GC_6_1084 b_6 NI_6 NS_1084 0 1.7020791845857687e-06
GC_6_1085 b_6 NI_6 NS_1085 0 3.4205429817278347e-06
GC_6_1086 b_6 NI_6 NS_1086 0 2.0399774862907608e-06
GC_6_1087 b_6 NI_6 NS_1087 0 1.0979313633091584e-05
GC_6_1088 b_6 NI_6 NS_1088 0 3.7863783650519410e-06
GC_6_1089 b_6 NI_6 NS_1089 0 4.8656049211138141e-06
GC_6_1090 b_6 NI_6 NS_1090 0 -8.4828087272899293e-08
GC_6_1091 b_6 NI_6 NS_1091 0 9.9928712394695358e-06
GC_6_1092 b_6 NI_6 NS_1092 0 -1.0833541296705077e-06
GC_6_1093 b_6 NI_6 NS_1093 0 8.2687933830825651e-06
GC_6_1094 b_6 NI_6 NS_1094 0 2.9476690982364637e-06
GC_6_1095 b_6 NI_6 NS_1095 0 1.9077427671484480e-05
GC_6_1096 b_6 NI_6 NS_1096 0 -5.5657363812504012e-06
GC_6_1097 b_6 NI_6 NS_1097 0 7.2206796257772123e-06
GC_6_1098 b_6 NI_6 NS_1098 0 -4.0253014084250304e-06
GC_6_1099 b_6 NI_6 NS_1099 0 1.3766283004003216e-05
GC_6_1100 b_6 NI_6 NS_1100 0 -1.1899498834988411e-05
GC_6_1101 b_6 NI_6 NS_1101 0 1.2420481858672631e-05
GC_6_1102 b_6 NI_6 NS_1102 0 -3.9375949378219997e-06
GC_6_1103 b_6 NI_6 NS_1103 0 9.2733681412889165e-06
GC_6_1104 b_6 NI_6 NS_1104 0 -2.6781575840482539e-05
GC_6_1105 b_6 NI_6 NS_1105 0 2.4206615640181230e-06
GC_6_1106 b_6 NI_6 NS_1106 0 -1.2364181295033152e-05
GC_6_1107 b_6 NI_6 NS_1107 0 -8.1530766204066523e-06
GC_6_1108 b_6 NI_6 NS_1108 0 -1.8689492530204735e-05
GC_6_1109 b_6 NI_6 NS_1109 0 -4.7467508239185590e-06
GC_6_1110 b_6 NI_6 NS_1110 0 -1.1992670053146294e-05
GC_6_1111 b_6 NI_6 NS_1111 0 5.4596299462598027e-05
GC_6_1112 b_6 NI_6 NS_1112 0 -8.9145401776647150e-05
GC_6_1113 b_6 NI_6 NS_1113 0 -9.8008118809773754e-06
GC_6_1114 b_6 NI_6 NS_1114 0 1.0736441214074415e-06
GC_6_1115 b_6 NI_6 NS_1115 0 3.9043695298726725e-07
GC_6_1116 b_6 NI_6 NS_1116 0 -1.3188532085871934e-07
GC_6_1117 b_6 NI_6 NS_1117 0 -2.5976304984530379e-06
GC_6_1118 b_6 NI_6 NS_1118 0 -2.0694185365027691e-06
GC_6_1119 b_6 NI_6 NS_1119 0 -4.3215031298900231e-06
GC_6_1120 b_6 NI_6 NS_1120 0 4.2993116120447324e-07
GC_6_1121 b_6 NI_6 NS_1121 0 -1.7356641028179229e-05
GC_6_1122 b_6 NI_6 NS_1122 0 9.7071534452095301e-06
GC_6_1123 b_6 NI_6 NS_1123 0 -8.9446467764177907e-06
GC_6_1124 b_6 NI_6 NS_1124 0 3.7512034534949061e-05
GC_6_1125 b_6 NI_6 NS_1125 0 -7.2510360475887901e-06
GC_6_1126 b_6 NI_6 NS_1126 0 3.2526187699706002e-07
GC_6_1127 b_6 NI_6 NS_1127 0 -1.3466584909299749e-05
GC_6_1128 b_6 NI_6 NS_1128 0 1.8883241292653362e-06
GC_6_1129 b_6 NI_6 NS_1129 0 -4.6297892645653430e-06
GC_6_1130 b_6 NI_6 NS_1130 0 -3.4285052062641840e-06
GC_6_1131 b_6 NI_6 NS_1131 0 -6.3984881100776129e-06
GC_6_1132 b_6 NI_6 NS_1132 0 1.0147265503783984e-06
GC_6_1133 b_6 NI_6 NS_1133 0 -3.0176504634552640e-06
GC_6_1134 b_6 NI_6 NS_1134 0 8.7792927498512069e-07
GC_6_1135 b_6 NI_6 NS_1135 0 -1.7623655812769631e-06
GC_6_1136 b_6 NI_6 NS_1136 0 -9.5961619594108227e-07
GC_6_1137 b_6 NI_6 NS_1137 0 -2.6113581753263519e-10
GC_6_1138 b_6 NI_6 NS_1138 0 4.2260600042071674e-10
GC_6_1139 b_6 NI_6 NS_1139 0 2.2541531945995941e-09
GC_6_1140 b_6 NI_6 NS_1140 0 -2.6820925610107610e-08
GC_6_1141 b_6 NI_6 NS_1141 0 -6.3151412933162916e-05
GC_6_1142 b_6 NI_6 NS_1142 0 3.1403585067412944e-07
GC_6_1143 b_6 NI_6 NS_1143 0 1.6220251030239807e-11
GC_6_1144 b_6 NI_6 NS_1144 0 -9.0648929032137467e-11
GC_6_1145 b_6 NI_6 NS_1145 0 -1.1289888153428015e-06
GC_6_1146 b_6 NI_6 NS_1146 0 -1.7888653582797340e-06
GC_6_1147 b_6 NI_6 NS_1147 0 -1.9838385388868297e-06
GC_6_1148 b_6 NI_6 NS_1148 0 1.9933859812126820e-06
GC_6_1149 b_6 NI_6 NS_1149 0 -9.6952269089947112e-06
GC_6_1150 b_6 NI_6 NS_1150 0 6.8014552021125808e-07
GC_6_1151 b_6 NI_6 NS_1151 0 -2.5333326092830139e-07
GC_6_1152 b_6 NI_6 NS_1152 0 3.4894115077516193e-06
GC_6_1153 b_6 NI_6 NS_1153 0 -2.1026812363119473e-06
GC_6_1154 b_6 NI_6 NS_1154 0 1.1808591800302114e-05
GC_6_1155 b_6 NI_6 NS_1155 0 6.7560298423112776e-06
GC_6_1156 b_6 NI_6 NS_1156 0 1.2503590559757655e-05
GC_6_1157 b_6 NI_6 NS_1157 0 -1.9973642071478094e-06
GC_6_1158 b_6 NI_6 NS_1158 0 -2.3069618062119863e-06
GC_6_1159 b_6 NI_6 NS_1159 0 1.6477101230653152e-06
GC_6_1160 b_6 NI_6 NS_1160 0 9.5582671826801495e-07
GC_6_1161 b_6 NI_6 NS_1161 0 7.5392900420546464e-06
GC_6_1162 b_6 NI_6 NS_1162 0 3.8837518344663017e-05
GC_6_1163 b_6 NI_6 NS_1163 0 2.3057222990794385e-05
GC_6_1164 b_6 NI_6 NS_1164 0 -1.1826462400637680e-05
GC_6_1165 b_6 NI_6 NS_1165 0 8.3538340993670521e-06
GC_6_1166 b_6 NI_6 NS_1166 0 1.6579973739170061e-06
GC_6_1167 b_6 NI_6 NS_1167 0 4.8581027621243096e-05
GC_6_1168 b_6 NI_6 NS_1168 0 -2.5173278067035869e-05
GC_6_1169 b_6 NI_6 NS_1169 0 -8.6231395773316483e-07
GC_6_1170 b_6 NI_6 NS_1170 0 -7.8674969409597611e-06
GC_6_1171 b_6 NI_6 NS_1171 0 3.4181901326160067e-05
GC_6_1172 b_6 NI_6 NS_1172 0 -7.8071006464131126e-06
GC_6_1173 b_6 NI_6 NS_1173 0 -3.8154373975777992e-05
GC_6_1174 b_6 NI_6 NS_1174 0 -5.2649710161947765e-05
GC_6_1175 b_6 NI_6 NS_1175 0 -4.4897619856127532e-06
GC_6_1176 b_6 NI_6 NS_1176 0 -4.3444042605116283e-06
GC_6_1177 b_6 NI_6 NS_1177 0 -3.9819368876314178e-05
GC_6_1178 b_6 NI_6 NS_1178 0 -2.0163486747463217e-05
GC_6_1179 b_6 NI_6 NS_1179 0 -4.8690194217470156e-06
GC_6_1180 b_6 NI_6 NS_1180 0 6.2179226925258770e-06
GC_6_1181 b_6 NI_6 NS_1181 0 -8.5133371468909289e-06
GC_6_1182 b_6 NI_6 NS_1182 0 -4.6696384934552224e-07
GC_6_1183 b_6 NI_6 NS_1183 0 -1.5584992321711979e-05
GC_6_1184 b_6 NI_6 NS_1184 0 2.4311329281765552e-05
GC_6_1185 b_6 NI_6 NS_1185 0 1.1061832362806263e-06
GC_6_1186 b_6 NI_6 NS_1186 0 2.3729737616667780e-06
GC_6_1187 b_6 NI_6 NS_1187 0 3.2346258771617347e-06
GC_6_1188 b_6 NI_6 NS_1188 0 1.8506896686635081e-05
GC_6_1189 b_6 NI_6 NS_1189 0 7.5468318664760152e-06
GC_6_1190 b_6 NI_6 NS_1190 0 -1.3939200397056965e-06
GC_6_1191 b_6 NI_6 NS_1191 0 2.9977256910699787e-06
GC_6_1192 b_6 NI_6 NS_1192 0 -5.0827904240217004e-07
GC_6_1193 b_6 NI_6 NS_1193 0 7.6492577837805388e-06
GC_6_1194 b_6 NI_6 NS_1194 0 -4.5387660244908607e-06
GC_6_1195 b_6 NI_6 NS_1195 0 -8.6278313457471422e-07
GC_6_1196 b_6 NI_6 NS_1196 0 -4.4779093017176648e-07
GC_6_1197 b_6 NI_6 NS_1197 0 -1.7230529689529306e-06
GC_6_1198 b_6 NI_6 NS_1198 0 1.8501969406212277e-07
GC_6_1199 b_6 NI_6 NS_1199 0 1.6122466547583501e-06
GC_6_1200 b_6 NI_6 NS_1200 0 -2.6584366116477171e-08
GC_6_1201 b_6 NI_6 NS_1201 0 3.7023968946593426e-06
GC_6_1202 b_6 NI_6 NS_1202 0 -9.2832690185967241e-07
GC_6_1203 b_6 NI_6 NS_1203 0 -8.7822140152161259e-08
GC_6_1204 b_6 NI_6 NS_1204 0 -3.4286822398237045e-07
GC_6_1205 b_6 NI_6 NS_1205 0 -5.7132067385068352e-07
GC_6_1206 b_6 NI_6 NS_1206 0 5.0950831672416875e-07
GC_6_1207 b_6 NI_6 NS_1207 0 2.4653232085314253e-06
GC_6_1208 b_6 NI_6 NS_1208 0 1.0743181062394443e-07
GC_6_1209 b_6 NI_6 NS_1209 0 3.4040128523604692e-06
GC_6_1210 b_6 NI_6 NS_1210 0 -2.8619466186075492e-06
GC_6_1211 b_6 NI_6 NS_1211 0 -2.6885269055201470e-07
GC_6_1212 b_6 NI_6 NS_1212 0 -5.0646418891443384e-08
GC_6_1213 b_6 NI_6 NS_1213 0 7.1805136844512327e-07
GC_6_1214 b_6 NI_6 NS_1214 0 1.0014730984415872e-06
GC_6_1215 b_6 NI_6 NS_1215 0 3.5530355674587341e-06
GC_6_1216 b_6 NI_6 NS_1216 0 3.3901963100344677e-08
GC_6_1217 b_6 NI_6 NS_1217 0 2.4205266553042904e-06
GC_6_1218 b_6 NI_6 NS_1218 0 -4.6592145548201027e-06
GC_6_1219 b_6 NI_6 NS_1219 0 4.5470662367322989e-07
GC_6_1220 b_6 NI_6 NS_1220 0 1.1297769850676796e-06
GC_6_1221 b_6 NI_6 NS_1221 0 3.6719780320076916e-06
GC_6_1222 b_6 NI_6 NS_1222 0 -6.9208058610023915e-07
GC_6_1223 b_6 NI_6 NS_1223 0 5.6214527898206970e-06
GC_6_1224 b_6 NI_6 NS_1224 0 -9.7041518949798295e-07
GC_6_1225 b_6 NI_6 NS_1225 0 -1.6193992253940860e-05
GC_6_1226 b_6 NI_6 NS_1226 0 -1.0663704631159816e-05
GC_6_1227 b_6 NI_6 NS_1227 0 9.4554658235639142e-07
GC_6_1228 b_6 NI_6 NS_1228 0 -7.5011977205952859e-06
GC_6_1229 b_6 NI_6 NS_1229 0 -6.7320736114703037e-08
GC_6_1230 b_6 NI_6 NS_1230 0 -1.4895713747548512e-07
GC_6_1231 b_6 NI_6 NS_1231 0 1.8076654737825228e-06
GC_6_1232 b_6 NI_6 NS_1232 0 -1.8968921113492080e-06
GC_6_1233 b_6 NI_6 NS_1233 0 5.3801167530998830e-07
GC_6_1234 b_6 NI_6 NS_1234 0 -3.4001964422691600e-06
GC_6_1235 b_6 NI_6 NS_1235 0 3.4182945433875275e-06
GC_6_1236 b_6 NI_6 NS_1236 0 -1.3139500667336976e-06
GC_6_1237 b_6 NI_6 NS_1237 0 4.5934124285159817e-06
GC_6_1238 b_6 NI_6 NS_1238 0 -8.0352769388052409e-07
GC_6_1239 b_6 NI_6 NS_1239 0 -1.9741084180160554e-07
GC_6_1240 b_6 NI_6 NS_1240 0 -2.0545957757459614e-07
GC_6_1241 b_6 NI_6 NS_1241 0 7.0278600693210790e-07
GC_6_1242 b_6 NI_6 NS_1242 0 1.4079551510481559e-06
GC_6_1243 b_6 NI_6 NS_1243 0 -7.0034243446401849e-07
GC_6_1244 b_6 NI_6 NS_1244 0 -1.4717274282637138e-06
GC_6_1245 b_6 NI_6 NS_1245 0 -6.2802116210858779e-07
GC_6_1246 b_6 NI_6 NS_1246 0 8.2384067677339933e-07
GC_6_1247 b_6 NI_6 NS_1247 0 2.2514720897460290e-07
GC_6_1248 b_6 NI_6 NS_1248 0 6.5403211782103257e-07
GC_6_1249 b_6 NI_6 NS_1249 0 6.0595862787083812e-07
GC_6_1250 b_6 NI_6 NS_1250 0 2.0968784538918057e-08
GC_6_1251 b_6 NI_6 NS_1251 0 1.3952678356298665e-11
GC_6_1252 b_6 NI_6 NS_1252 0 5.3757766528821378e-13
GC_6_1253 b_6 NI_6 NS_1253 0 4.3669559151899307e-10
GC_6_1254 b_6 NI_6 NS_1254 0 1.6922264807395784e-09
GC_6_1255 b_6 NI_6 NS_1255 0 8.4580441885574267e-05
GC_6_1256 b_6 NI_6 NS_1256 0 1.9045627260079454e-07
GC_6_1257 b_6 NI_6 NS_1257 0 2.0155349797010242e-11
GC_6_1258 b_6 NI_6 NS_1258 0 -9.4458366716786394e-10
GC_6_1259 b_6 NI_6 NS_1259 0 8.8329950078659573e-07
GC_6_1260 b_6 NI_6 NS_1260 0 5.7933410032693081e-08
GC_6_1261 b_6 NI_6 NS_1261 0 1.1602010333246419e-06
GC_6_1262 b_6 NI_6 NS_1262 0 6.9968060309644224e-08
GC_6_1263 b_6 NI_6 NS_1263 0 3.3628861670148171e-06
GC_6_1264 b_6 NI_6 NS_1264 0 -3.2258609865283838e-06
GC_6_1265 b_6 NI_6 NS_1265 0 -2.0855281120377587e-06
GC_6_1266 b_6 NI_6 NS_1266 0 -1.7319080803057424e-06
GC_6_1267 b_6 NI_6 NS_1267 0 1.9313030219999392e-06
GC_6_1268 b_6 NI_6 NS_1268 0 -2.2094017217683040e-06
GC_6_1269 b_6 NI_6 NS_1269 0 -5.8922113760948743e-06
GC_6_1270 b_6 NI_6 NS_1270 0 -7.1422704868014034e-06
GC_6_1271 b_6 NI_6 NS_1271 0 9.4972546152650628e-07
GC_6_1272 b_6 NI_6 NS_1272 0 2.2263820793064395e-06
GC_6_1273 b_6 NI_6 NS_1273 0 -2.2764211064392485e-06
GC_6_1274 b_6 NI_6 NS_1274 0 8.0098709406874246e-07
GC_6_1275 b_6 NI_6 NS_1275 0 5.8207621621017356e-07
GC_6_1276 b_6 NI_6 NS_1276 0 -4.8941596542781979e-06
GC_6_1277 b_6 NI_6 NS_1277 0 -6.4023893087137282e-06
GC_6_1278 b_6 NI_6 NS_1278 0 2.7555986163904220e-06
GC_6_1279 b_6 NI_6 NS_1279 0 -1.0155998643423423e-06
GC_6_1280 b_6 NI_6 NS_1280 0 1.6581852898093884e-06
GC_6_1281 b_6 NI_6 NS_1281 0 -3.3720580419558081e-06
GC_6_1282 b_6 NI_6 NS_1282 0 -2.5292965278981153e-06
GC_6_1283 b_6 NI_6 NS_1283 0 -2.2047548846699165e-06
GC_6_1284 b_6 NI_6 NS_1284 0 2.3621389807175671e-06
GC_6_1285 b_6 NI_6 NS_1285 0 1.5152439389848234e-06
GC_6_1286 b_6 NI_6 NS_1286 0 2.6088614488997900e-06
GC_6_1287 b_6 NI_6 NS_1287 0 -5.1183458323236233e-06
GC_6_1288 b_6 NI_6 NS_1288 0 -2.0383784860213075e-06
GC_6_1289 b_6 NI_6 NS_1289 0 -1.4940205830940762e-06
GC_6_1290 b_6 NI_6 NS_1290 0 2.2226898044353675e-06
GC_6_1291 b_6 NI_6 NS_1291 0 -4.8359506912936854e-08
GC_6_1292 b_6 NI_6 NS_1292 0 -1.0715149264375543e-06
GC_6_1293 b_6 NI_6 NS_1293 0 -2.7776174406962234e-06
GC_6_1294 b_6 NI_6 NS_1294 0 1.7676086511505876e-06
GC_6_1295 b_6 NI_6 NS_1295 0 -7.8765238619305550e-07
GC_6_1296 b_6 NI_6 NS_1296 0 2.3415814563196124e-06
GC_6_1297 b_6 NI_6 NS_1297 0 -1.0034711604867534e-06
GC_6_1298 b_6 NI_6 NS_1298 0 -1.3434469428920311e-06
GC_6_1299 b_6 NI_6 NS_1299 0 -1.8384294735799558e-06
GC_6_1300 b_6 NI_6 NS_1300 0 1.3364981937370700e-06
GC_6_1301 b_6 NI_6 NS_1301 0 5.5164889569962535e-07
GC_6_1302 b_6 NI_6 NS_1302 0 1.6482326980356122e-07
GC_6_1303 b_6 NI_6 NS_1303 0 -2.9422070238049622e-06
GC_6_1304 b_6 NI_6 NS_1304 0 3.7599790525194355e-07
GC_6_1305 b_6 NI_6 NS_1305 0 -9.6502850468555684e-07
GC_6_1306 b_6 NI_6 NS_1306 0 7.1171509973821910e-07
GC_6_1307 b_6 NI_6 NS_1307 0 -1.9725521449073548e-06
GC_6_1308 b_6 NI_6 NS_1308 0 -7.9508488333266449e-07
GC_6_1309 b_6 NI_6 NS_1309 0 -1.4687383839295035e-06
GC_6_1310 b_6 NI_6 NS_1310 0 6.2098843680546771e-07
GC_6_1311 b_6 NI_6 NS_1311 0 -1.1171723959211045e-06
GC_6_1312 b_6 NI_6 NS_1312 0 -3.9225834327974472e-07
GC_6_1313 b_6 NI_6 NS_1313 0 -2.4594674717299084e-06
GC_6_1314 b_6 NI_6 NS_1314 0 -6.3473555889208913e-07
GC_6_1315 b_6 NI_6 NS_1315 0 -3.0280708493996779e-06
GC_6_1316 b_6 NI_6 NS_1316 0 -3.1143928614956113e-07
GC_6_1317 b_6 NI_6 NS_1317 0 -2.1722197722341397e-06
GC_6_1318 b_6 NI_6 NS_1318 0 3.1818642490006887e-07
GC_6_1319 b_6 NI_6 NS_1319 0 -2.7406254282083332e-06
GC_6_1320 b_6 NI_6 NS_1320 0 3.0317818988046178e-07
GC_6_1321 b_6 NI_6 NS_1321 0 -4.2061080053554374e-06
GC_6_1322 b_6 NI_6 NS_1322 0 -7.3435615652531226e-07
GC_6_1323 b_6 NI_6 NS_1323 0 -5.6819242117623174e-06
GC_6_1324 b_6 NI_6 NS_1324 0 2.2499643219191249e-06
GC_6_1325 b_6 NI_6 NS_1325 0 -3.1747527371648695e-06
GC_6_1326 b_6 NI_6 NS_1326 0 1.8635247466779249e-06
GC_6_1327 b_6 NI_6 NS_1327 0 -4.1153813581479546e-06
GC_6_1328 b_6 NI_6 NS_1328 0 3.2994553883685435e-06
GC_6_1329 b_6 NI_6 NS_1329 0 -5.6740252637713997e-06
GC_6_1330 b_6 NI_6 NS_1330 0 1.3489957159606564e-06
GC_6_1331 b_6 NI_6 NS_1331 0 -3.5119892405271267e-06
GC_6_1332 b_6 NI_6 NS_1332 0 8.2346884832062347e-06
GC_6_1333 b_6 NI_6 NS_1333 0 -2.3076937381871103e-06
GC_6_1334 b_6 NI_6 NS_1334 0 4.5638150843544540e-06
GC_6_1335 b_6 NI_6 NS_1335 0 1.1261134166295056e-06
GC_6_1336 b_6 NI_6 NS_1336 0 5.4139214768042226e-06
GC_6_1337 b_6 NI_6 NS_1337 0 -1.8428018552436910e-06
GC_6_1338 b_6 NI_6 NS_1338 0 3.4530155984992758e-06
GC_6_1339 b_6 NI_6 NS_1339 0 -7.0172872193463425e-06
GC_6_1340 b_6 NI_6 NS_1340 0 3.7168276293635202e-05
GC_6_1341 b_6 NI_6 NS_1341 0 6.9494403352830797e-07
GC_6_1342 b_6 NI_6 NS_1342 0 2.6509036898796044e-06
GC_6_1343 b_6 NI_6 NS_1343 0 -8.4712142809652004e-08
GC_6_1344 b_6 NI_6 NS_1344 0 1.1840328113808305e-07
GC_6_1345 b_6 NI_6 NS_1345 0 -7.2440145532804653e-07
GC_6_1346 b_6 NI_6 NS_1346 0 3.4149225061309473e-06
GC_6_1347 b_6 NI_6 NS_1347 0 6.7713289819938791e-07
GC_6_1348 b_6 NI_6 NS_1348 0 8.6106570699078578e-07
GC_6_1349 b_6 NI_6 NS_1349 0 2.2825499247774992e-06
GC_6_1350 b_6 NI_6 NS_1350 0 -3.1366047579595443e-06
GC_6_1351 b_6 NI_6 NS_1351 0 -1.5483035100097255e-06
GC_6_1352 b_6 NI_6 NS_1352 0 -1.1843702648401331e-05
GC_6_1353 b_6 NI_6 NS_1353 0 2.0447488873369180e-06
GC_6_1354 b_6 NI_6 NS_1354 0 -7.3740350738974669e-07
GC_6_1355 b_6 NI_6 NS_1355 0 4.5134996031002569e-06
GC_6_1356 b_6 NI_6 NS_1356 0 -4.0110313678626961e-07
GC_6_1357 b_6 NI_6 NS_1357 0 1.2442188583003029e-06
GC_6_1358 b_6 NI_6 NS_1358 0 1.9853482106865495e-06
GC_6_1359 b_6 NI_6 NS_1359 0 1.7411980788475754e-06
GC_6_1360 b_6 NI_6 NS_1360 0 -7.6164694793204105e-07
GC_6_1361 b_6 NI_6 NS_1361 0 5.8319424544753120e-07
GC_6_1362 b_6 NI_6 NS_1362 0 5.1104638665066464e-07
GC_6_1363 b_6 NI_6 NS_1363 0 6.5669154015749160e-07
GC_6_1364 b_6 NI_6 NS_1364 0 -7.6193870552889512e-08
GC_6_1365 b_6 NI_6 NS_1365 0 2.2925806713632255e-11
GC_6_1366 b_6 NI_6 NS_1366 0 -9.3367259394458185e-11
GC_6_1367 b_6 NI_6 NS_1367 0 -1.8302761542260993e-09
GC_6_1368 b_6 NI_6 NS_1368 0 4.0623342428613867e-09
GD_6_1 b_6 NI_6 NA_1 0 2.4205669908689932e-06
GD_6_2 b_6 NI_6 NA_2 0 5.6585683135627450e-06
GD_6_3 b_6 NI_6 NA_3 0 2.6994450242091276e-05
GD_6_4 b_6 NI_6 NA_4 0 1.0032020453594625e-04
GD_6_5 b_6 NI_6 NA_5 0 -4.2218527252709283e-03
GD_6_6 b_6 NI_6 NA_6 0 -8.8807860850851975e-03
GD_6_7 b_6 NI_6 NA_7 0 5.8609053537462120e-04
GD_6_8 b_6 NI_6 NA_8 0 1.2979344926715285e-02
GD_6_9 b_6 NI_6 NA_9 0 1.2382102020478832e-06
GD_6_10 b_6 NI_6 NA_10 0 4.5909852458775341e-06
GD_6_11 b_6 NI_6 NA_11 0 1.0213241742056417e-05
GD_6_12 b_6 NI_6 NA_12 0 -6.7028356753559600e-06
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 6.6651395226593446e-05
GC_7_2 b_7 NI_7 NS_2 0 2.1491723682076291e-07
GC_7_3 b_7 NI_7 NS_3 0 2.2385585951271399e-11
GC_7_4 b_7 NI_7 NS_4 0 -9.9158362627394574e-10
GC_7_5 b_7 NI_7 NS_5 0 4.2970867628739517e-07
GC_7_6 b_7 NI_7 NS_6 0 1.8577073712703544e-07
GC_7_7 b_7 NI_7 NS_7 0 6.0303233302483539e-07
GC_7_8 b_7 NI_7 NS_8 0 5.0409511194905893e-07
GC_7_9 b_7 NI_7 NS_9 0 2.9694846239807247e-06
GC_7_10 b_7 NI_7 NS_10 0 -1.5587272750997241e-06
GC_7_11 b_7 NI_7 NS_11 0 -1.1975758908224287e-06
GC_7_12 b_7 NI_7 NS_12 0 -1.1247596178524118e-06
GC_7_13 b_7 NI_7 NS_13 0 2.3738782563121335e-06
GC_7_14 b_7 NI_7 NS_14 0 -8.6541711146762024e-07
GC_7_15 b_7 NI_7 NS_15 0 -2.5702159316134982e-06
GC_7_16 b_7 NI_7 NS_16 0 -6.4135430623265797e-06
GC_7_17 b_7 NI_7 NS_17 0 1.0932674090802925e-07
GC_7_18 b_7 NI_7 NS_18 0 1.6956899406107657e-06
GC_7_19 b_7 NI_7 NS_19 0 -1.7209484488795267e-06
GC_7_20 b_7 NI_7 NS_20 0 5.0733424606346524e-07
GC_7_21 b_7 NI_7 NS_21 0 3.1297099056602458e-06
GC_7_22 b_7 NI_7 NS_22 0 -4.3417948521078290e-06
GC_7_23 b_7 NI_7 NS_23 0 -6.6647730569680949e-06
GC_7_24 b_7 NI_7 NS_24 0 1.1555774756580657e-06
GC_7_25 b_7 NI_7 NS_25 0 -4.7409987958958329e-07
GC_7_26 b_7 NI_7 NS_26 0 1.6879959829248463e-06
GC_7_27 b_7 NI_7 NS_27 0 -2.1234786770666913e-06
GC_7_28 b_7 NI_7 NS_28 0 -4.2598558761226818e-06
GC_7_29 b_7 NI_7 NS_29 0 -2.2157160029145314e-06
GC_7_30 b_7 NI_7 NS_30 0 2.1650792667727856e-06
GC_7_31 b_7 NI_7 NS_31 0 3.1625501636796751e-06
GC_7_32 b_7 NI_7 NS_32 0 3.0747064260881073e-06
GC_7_33 b_7 NI_7 NS_33 0 -6.0917990167600677e-06
GC_7_34 b_7 NI_7 NS_34 0 -4.4592809515001279e-06
GC_7_35 b_7 NI_7 NS_35 0 -1.2974854949068915e-06
GC_7_36 b_7 NI_7 NS_36 0 2.1674364872245917e-06
GC_7_37 b_7 NI_7 NS_37 0 2.8446479470887342e-07
GC_7_38 b_7 NI_7 NS_38 0 -2.8074508254494171e-06
GC_7_39 b_7 NI_7 NS_39 0 -3.1954505258888206e-06
GC_7_40 b_7 NI_7 NS_40 0 1.8332573472179427e-06
GC_7_41 b_7 NI_7 NS_41 0 -3.1171902547485514e-07
GC_7_42 b_7 NI_7 NS_42 0 2.3433549194794608e-06
GC_7_43 b_7 NI_7 NS_43 0 -1.4634075039204026e-06
GC_7_44 b_7 NI_7 NS_44 0 -2.6245710689058521e-06
GC_7_45 b_7 NI_7 NS_45 0 -1.8978822129495256e-06
GC_7_46 b_7 NI_7 NS_46 0 1.3684809820861400e-06
GC_7_47 b_7 NI_7 NS_47 0 1.1604804990486382e-06
GC_7_48 b_7 NI_7 NS_48 0 -6.4651801919968443e-07
GC_7_49 b_7 NI_7 NS_49 0 -3.5975087539003598e-06
GC_7_50 b_7 NI_7 NS_50 0 2.8531228570685067e-07
GC_7_51 b_7 NI_7 NS_51 0 -8.2535295211906401e-07
GC_7_52 b_7 NI_7 NS_52 0 7.2325695071756399e-07
GC_7_53 b_7 NI_7 NS_53 0 -1.8919627985384480e-06
GC_7_54 b_7 NI_7 NS_54 0 -1.3288986485561596e-06
GC_7_55 b_7 NI_7 NS_55 0 -1.4489681039056087e-06
GC_7_56 b_7 NI_7 NS_56 0 5.5809478590132472e-07
GC_7_57 b_7 NI_7 NS_57 0 -1.0695912189731418e-06
GC_7_58 b_7 NI_7 NS_58 0 -5.9316176529777295e-07
GC_7_59 b_7 NI_7 NS_59 0 -2.3263765873560001e-06
GC_7_60 b_7 NI_7 NS_60 0 -6.7330265383212068e-07
GC_7_61 b_7 NI_7 NS_61 0 -2.7997955960603955e-06
GC_7_62 b_7 NI_7 NS_62 0 -5.7610658089754747e-07
GC_7_63 b_7 NI_7 NS_63 0 -2.0698223915583871e-06
GC_7_64 b_7 NI_7 NS_64 0 2.3466856413826063e-07
GC_7_65 b_7 NI_7 NS_65 0 -2.5964216970808608e-06
GC_7_66 b_7 NI_7 NS_66 0 1.0337928925644831e-07
GC_7_67 b_7 NI_7 NS_67 0 -3.9140718115779829e-06
GC_7_68 b_7 NI_7 NS_68 0 -7.2803069343779683e-07
GC_7_69 b_7 NI_7 NS_69 0 -5.2745683725303073e-06
GC_7_70 b_7 NI_7 NS_70 0 1.8892502292319134e-06
GC_7_71 b_7 NI_7 NS_71 0 -2.9583282966023254e-06
GC_7_72 b_7 NI_7 NS_72 0 1.7283197517667315e-06
GC_7_73 b_7 NI_7 NS_73 0 -3.7941649358827489e-06
GC_7_74 b_7 NI_7 NS_74 0 2.9619619744595650e-06
GC_7_75 b_7 NI_7 NS_75 0 -5.2505214068579155e-06
GC_7_76 b_7 NI_7 NS_76 0 1.3684591777873211e-06
GC_7_77 b_7 NI_7 NS_77 0 -2.9715071557620697e-06
GC_7_78 b_7 NI_7 NS_78 0 7.6158271046329488e-06
GC_7_79 b_7 NI_7 NS_79 0 -1.9293754786165259e-06
GC_7_80 b_7 NI_7 NS_80 0 4.3918277104109253e-06
GC_7_81 b_7 NI_7 NS_81 0 1.5652485241654182e-06
GC_7_82 b_7 NI_7 NS_82 0 4.8415896671958495e-06
GC_7_83 b_7 NI_7 NS_83 0 -9.8516304305767552e-07
GC_7_84 b_7 NI_7 NS_84 0 3.6448228758872711e-06
GC_7_85 b_7 NI_7 NS_85 0 -1.0328830379784172e-05
GC_7_86 b_7 NI_7 NS_86 0 3.3088912137429090e-05
GC_7_87 b_7 NI_7 NS_87 0 1.3184345525628459e-06
GC_7_88 b_7 NI_7 NS_88 0 1.2141108945396767e-06
GC_7_89 b_7 NI_7 NS_89 0 -9.3725637884325672e-08
GC_7_90 b_7 NI_7 NS_90 0 8.7540936220571663e-08
GC_7_91 b_7 NI_7 NS_91 0 -3.3374053911318109e-07
GC_7_92 b_7 NI_7 NS_92 0 2.6694950287872457e-06
GC_7_93 b_7 NI_7 NS_93 0 7.2381464980109734e-07
GC_7_94 b_7 NI_7 NS_94 0 1.5751128059479532e-07
GC_7_95 b_7 NI_7 NS_95 0 3.0782521100305982e-06
GC_7_96 b_7 NI_7 NS_96 0 -2.7783598765447664e-06
GC_7_97 b_7 NI_7 NS_97 0 -1.9583289015566573e-07
GC_7_98 b_7 NI_7 NS_98 0 -1.1673005728529611e-05
GC_7_99 b_7 NI_7 NS_99 0 1.9428743350714970e-06
GC_7_100 b_7 NI_7 NS_100 0 -6.7931477102352031e-07
GC_7_101 b_7 NI_7 NS_101 0 4.3055692616212471e-06
GC_7_102 b_7 NI_7 NS_102 0 -1.7836135856419890e-07
GC_7_103 b_7 NI_7 NS_103 0 1.2120139151790877e-06
GC_7_104 b_7 NI_7 NS_104 0 1.8707239129279736e-06
GC_7_105 b_7 NI_7 NS_105 0 1.6462419048354493e-06
GC_7_106 b_7 NI_7 NS_106 0 -7.9777719050203501e-07
GC_7_107 b_7 NI_7 NS_107 0 5.9154547673270931e-07
GC_7_108 b_7 NI_7 NS_108 0 4.7809429223504250e-07
GC_7_109 b_7 NI_7 NS_109 0 6.8253522757825861e-07
GC_7_110 b_7 NI_7 NS_110 0 -9.6305426361160791e-08
GC_7_111 b_7 NI_7 NS_111 0 2.5759036258521212e-11
GC_7_112 b_7 NI_7 NS_112 0 -9.7284646978416518e-11
GC_7_113 b_7 NI_7 NS_113 0 -1.9602950447272410e-09
GC_7_114 b_7 NI_7 NS_114 0 4.2975214246468881e-09
GC_7_115 b_7 NI_7 NS_115 0 -6.1954668528806759e-05
GC_7_116 b_7 NI_7 NS_116 0 3.1010277272149012e-07
GC_7_117 b_7 NI_7 NS_117 0 1.6335111360845019e-11
GC_7_118 b_7 NI_7 NS_118 0 -8.7576778327166667e-11
GC_7_119 b_7 NI_7 NS_119 0 -1.1069939491847854e-06
GC_7_120 b_7 NI_7 NS_120 0 -1.7649929252806386e-06
GC_7_121 b_7 NI_7 NS_121 0 -1.9904427073590616e-06
GC_7_122 b_7 NI_7 NS_122 0 1.9660076452518763e-06
GC_7_123 b_7 NI_7 NS_123 0 -9.5690872219586335e-06
GC_7_124 b_7 NI_7 NS_124 0 6.6947457516555216e-07
GC_7_125 b_7 NI_7 NS_125 0 -2.0966027349281020e-07
GC_7_126 b_7 NI_7 NS_126 0 3.5162839675861130e-06
GC_7_127 b_7 NI_7 NS_127 0 -2.1093932240475288e-06
GC_7_128 b_7 NI_7 NS_128 0 1.1709180626269876e-05
GC_7_129 b_7 NI_7 NS_129 0 6.8681806977884982e-06
GC_7_130 b_7 NI_7 NS_130 0 1.2213086956571670e-05
GC_7_131 b_7 NI_7 NS_131 0 -2.0257228280576450e-06
GC_7_132 b_7 NI_7 NS_132 0 -2.2559648199057840e-06
GC_7_133 b_7 NI_7 NS_133 0 1.6633441224004873e-06
GC_7_134 b_7 NI_7 NS_134 0 1.0211503096341604e-06
GC_7_135 b_7 NI_7 NS_135 0 7.4141092589786562e-06
GC_7_136 b_7 NI_7 NS_136 0 3.8490345184527506e-05
GC_7_137 b_7 NI_7 NS_137 0 2.2911880060839566e-05
GC_7_138 b_7 NI_7 NS_138 0 -1.2059855698341216e-05
GC_7_139 b_7 NI_7 NS_139 0 8.4232931218459287e-06
GC_7_140 b_7 NI_7 NS_140 0 1.7608828801453713e-06
GC_7_141 b_7 NI_7 NS_141 0 4.7761677973413127e-05
GC_7_142 b_7 NI_7 NS_142 0 -2.5200268829866126e-05
GC_7_143 b_7 NI_7 NS_143 0 -9.4026374769014827e-07
GC_7_144 b_7 NI_7 NS_144 0 -8.0488267987794041e-06
GC_7_145 b_7 NI_7 NS_145 0 3.4272852320129750e-05
GC_7_146 b_7 NI_7 NS_146 0 -7.7701628827419183e-06
GC_7_147 b_7 NI_7 NS_147 0 -3.8695798007954010e-05
GC_7_148 b_7 NI_7 NS_148 0 -5.1800859309168322e-05
GC_7_149 b_7 NI_7 NS_149 0 -4.5827306906996563e-06
GC_7_150 b_7 NI_7 NS_150 0 -4.5466881110385093e-06
GC_7_151 b_7 NI_7 NS_151 0 -3.9429359404879865e-05
GC_7_152 b_7 NI_7 NS_152 0 -1.9669236457993503e-05
GC_7_153 b_7 NI_7 NS_153 0 -4.8828620506727606e-06
GC_7_154 b_7 NI_7 NS_154 0 6.5890061936388160e-06
GC_7_155 b_7 NI_7 NS_155 0 -8.6504788990616727e-06
GC_7_156 b_7 NI_7 NS_156 0 -6.8353874478790871e-07
GC_7_157 b_7 NI_7 NS_157 0 -1.4941086151591754e-05
GC_7_158 b_7 NI_7 NS_158 0 2.4266072002972179e-05
GC_7_159 b_7 NI_7 NS_159 0 1.0803053485065640e-06
GC_7_160 b_7 NI_7 NS_160 0 2.6351383752883833e-06
GC_7_161 b_7 NI_7 NS_161 0 3.0586501998123282e-06
GC_7_162 b_7 NI_7 NS_162 0 1.8296341364419156e-05
GC_7_163 b_7 NI_7 NS_163 0 7.7541134486955442e-06
GC_7_164 b_7 NI_7 NS_164 0 -1.6862231100172924e-06
GC_7_165 b_7 NI_7 NS_165 0 2.9848520776057727e-06
GC_7_166 b_7 NI_7 NS_166 0 -3.4525646248578768e-07
GC_7_167 b_7 NI_7 NS_167 0 7.3238406918135273e-06
GC_7_168 b_7 NI_7 NS_168 0 -4.5245365513310109e-06
GC_7_169 b_7 NI_7 NS_169 0 -8.5067708889949019e-07
GC_7_170 b_7 NI_7 NS_170 0 -5.4051518072296651e-07
GC_7_171 b_7 NI_7 NS_171 0 -1.6424475805550522e-06
GC_7_172 b_7 NI_7 NS_172 0 2.2866431246454443e-07
GC_7_173 b_7 NI_7 NS_173 0 1.5095996113746468e-06
GC_7_174 b_7 NI_7 NS_174 0 1.1390141461049452e-07
GC_7_175 b_7 NI_7 NS_175 0 3.6033404625123502e-06
GC_7_176 b_7 NI_7 NS_176 0 -8.9568462471850732e-07
GC_7_177 b_7 NI_7 NS_177 0 -7.2228808817236548e-08
GC_7_178 b_7 NI_7 NS_178 0 -3.6299637882924652e-07
GC_7_179 b_7 NI_7 NS_179 0 -5.1726466935765200e-07
GC_7_180 b_7 NI_7 NS_180 0 5.5090740117428724e-07
GC_7_181 b_7 NI_7 NS_181 0 2.4011105758347735e-06
GC_7_182 b_7 NI_7 NS_182 0 2.0003027444575224e-07
GC_7_183 b_7 NI_7 NS_183 0 3.3592392521777601e-06
GC_7_184 b_7 NI_7 NS_184 0 -2.8048521107672629e-06
GC_7_185 b_7 NI_7 NS_185 0 -2.6349845455119420e-07
GC_7_186 b_7 NI_7 NS_186 0 -4.2643787599283132e-08
GC_7_187 b_7 NI_7 NS_187 0 7.5184337178203697e-07
GC_7_188 b_7 NI_7 NS_188 0 1.0635520301885617e-06
GC_7_189 b_7 NI_7 NS_189 0 3.5136228654918580e-06
GC_7_190 b_7 NI_7 NS_190 0 7.3949176580705062e-08
GC_7_191 b_7 NI_7 NS_191 0 2.4236009488381908e-06
GC_7_192 b_7 NI_7 NS_192 0 -4.5985061226050391e-06
GC_7_193 b_7 NI_7 NS_193 0 4.5788524517994155e-07
GC_7_194 b_7 NI_7 NS_194 0 1.1656944105502196e-06
GC_7_195 b_7 NI_7 NS_195 0 3.6840047676407798e-06
GC_7_196 b_7 NI_7 NS_196 0 -6.3710032086859174e-07
GC_7_197 b_7 NI_7 NS_197 0 5.5747457580953034e-06
GC_7_198 b_7 NI_7 NS_198 0 -9.4416434491423118e-07
GC_7_199 b_7 NI_7 NS_199 0 -1.6037170782393021e-05
GC_7_200 b_7 NI_7 NS_200 0 -1.0587154011010986e-05
GC_7_201 b_7 NI_7 NS_201 0 9.9723791127887326e-07
GC_7_202 b_7 NI_7 NS_202 0 -7.4331324412775383e-06
GC_7_203 b_7 NI_7 NS_203 0 -6.5807671162971059e-08
GC_7_204 b_7 NI_7 NS_204 0 -1.4868602657859884e-07
GC_7_205 b_7 NI_7 NS_205 0 1.8273983843745492e-06
GC_7_206 b_7 NI_7 NS_206 0 -1.8611918947902145e-06
GC_7_207 b_7 NI_7 NS_207 0 5.4344727667920102e-07
GC_7_208 b_7 NI_7 NS_208 0 -3.3780247178151217e-06
GC_7_209 b_7 NI_7 NS_209 0 3.3863434938638565e-06
GC_7_210 b_7 NI_7 NS_210 0 -1.3093484481067862e-06
GC_7_211 b_7 NI_7 NS_211 0 4.5638544082905546e-06
GC_7_212 b_7 NI_7 NS_212 0 -7.9244139665554490e-07
GC_7_213 b_7 NI_7 NS_213 0 -2.0240554356759675e-07
GC_7_214 b_7 NI_7 NS_214 0 -2.0622442440132221e-07
GC_7_215 b_7 NI_7 NS_215 0 7.0565518318475020e-07
GC_7_216 b_7 NI_7 NS_216 0 1.3955197437072695e-06
GC_7_217 b_7 NI_7 NS_217 0 -7.0553670025418633e-07
GC_7_218 b_7 NI_7 NS_218 0 -1.4723664045162816e-06
GC_7_219 b_7 NI_7 NS_219 0 -6.2774322295708976e-07
GC_7_220 b_7 NI_7 NS_220 0 8.2972056091408928e-07
GC_7_221 b_7 NI_7 NS_221 0 2.2261764753178066e-07
GC_7_222 b_7 NI_7 NS_222 0 6.5380930400920033e-07
GC_7_223 b_7 NI_7 NS_223 0 5.9764910180051477e-07
GC_7_224 b_7 NI_7 NS_224 0 2.1145577749465740e-08
GC_7_225 b_7 NI_7 NS_225 0 1.4034147424980890e-11
GC_7_226 b_7 NI_7 NS_226 0 1.0178601678075054e-12
GC_7_227 b_7 NI_7 NS_227 0 4.3186556234341503e-10
GC_7_228 b_7 NI_7 NS_228 0 1.6518450780175544e-09
GC_7_229 b_7 NI_7 NS_229 0 -1.1096947632922644e-04
GC_7_230 b_7 NI_7 NS_230 0 -2.1483030788235585e-06
GC_7_231 b_7 NI_7 NS_231 0 -2.5029536456035706e-10
GC_7_232 b_7 NI_7 NS_232 0 2.6115897804582410e-09
GC_7_233 b_7 NI_7 NS_233 0 1.8723152996615109e-06
GC_7_234 b_7 NI_7 NS_234 0 -1.6074371587623970e-06
GC_7_235 b_7 NI_7 NS_235 0 3.2540198515411774e-07
GC_7_236 b_7 NI_7 NS_236 0 -6.5210480568463915e-06
GC_7_237 b_7 NI_7 NS_237 0 -7.4589938105618449e-06
GC_7_238 b_7 NI_7 NS_238 0 -4.2413629392557597e-07
GC_7_239 b_7 NI_7 NS_239 0 -1.5203206927382317e-06
GC_7_240 b_7 NI_7 NS_240 0 -4.8607526669801257e-06
GC_7_241 b_7 NI_7 NS_241 0 -1.6019418891776626e-05
GC_7_242 b_7 NI_7 NS_242 0 -2.1097785541593303e-06
GC_7_243 b_7 NI_7 NS_243 0 -7.3376609740444753e-06
GC_7_244 b_7 NI_7 NS_244 0 1.8827315790490709e-05
GC_7_245 b_7 NI_7 NS_245 0 4.9694020224546027e-06
GC_7_246 b_7 NI_7 NS_246 0 -2.7979707241907394e-06
GC_7_247 b_7 NI_7 NS_247 0 -2.3130527386348392e-07
GC_7_248 b_7 NI_7 NS_248 0 -2.4916638620577636e-06
GC_7_249 b_7 NI_7 NS_249 0 -2.6811396922216118e-05
GC_7_250 b_7 NI_7 NS_250 0 2.8304979034737248e-05
GC_7_251 b_7 NI_7 NS_251 0 2.8363182534895550e-05
GC_7_252 b_7 NI_7 NS_252 0 -7.9685184347202437e-06
GC_7_253 b_7 NI_7 NS_253 0 -8.2696309984664953e-06
GC_7_254 b_7 NI_7 NS_254 0 -4.3355266577867571e-06
GC_7_255 b_7 NI_7 NS_255 0 1.2216122407712467e-05
GC_7_256 b_7 NI_7 NS_256 0 2.7630082381633001e-05
GC_7_257 b_7 NI_7 NS_257 0 1.4665316269874782e-06
GC_7_258 b_7 NI_7 NS_258 0 -8.9517362454360325e-06
GC_7_259 b_7 NI_7 NS_259 0 -2.8979852867188356e-05
GC_7_260 b_7 NI_7 NS_260 0 4.5865772933158950e-06
GC_7_261 b_7 NI_7 NS_261 0 4.1777950415176427e-05
GC_7_262 b_7 NI_7 NS_262 0 1.1538570991021152e-05
GC_7_263 b_7 NI_7 NS_263 0 -3.0566435995561944e-06
GC_7_264 b_7 NI_7 NS_264 0 -4.4930605616670374e-06
GC_7_265 b_7 NI_7 NS_265 0 1.2853449371907263e-05
GC_7_266 b_7 NI_7 NS_266 0 1.9652908107745760e-05
GC_7_267 b_7 NI_7 NS_267 0 3.9663199709835847e-06
GC_7_268 b_7 NI_7 NS_268 0 -1.0991933395157395e-05
GC_7_269 b_7 NI_7 NS_269 0 -6.6134810366712868e-06
GC_7_270 b_7 NI_7 NS_270 0 8.3132153445807294e-07
GC_7_271 b_7 NI_7 NS_271 0 1.9091619983326353e-05
GC_7_272 b_7 NI_7 NS_272 0 5.9084922004889624e-06
GC_7_273 b_7 NI_7 NS_273 0 -5.2595700895616686e-08
GC_7_274 b_7 NI_7 NS_274 0 -4.2237277391127255e-06
GC_7_275 b_7 NI_7 NS_275 0 4.6917577039684095e-06
GC_7_276 b_7 NI_7 NS_276 0 1.4599971541569883e-05
GC_7_277 b_7 NI_7 NS_277 0 8.0921059616469052e-06
GC_7_278 b_7 NI_7 NS_278 0 -1.1172243804813273e-05
GC_7_279 b_7 NI_7 NS_279 0 -1.4419299066455765e-06
GC_7_280 b_7 NI_7 NS_280 0 9.2581086788118407e-07
GC_7_281 b_7 NI_7 NS_281 0 1.0893573744911831e-05
GC_7_282 b_7 NI_7 NS_282 0 4.3229016053897261e-06
GC_7_283 b_7 NI_7 NS_283 0 1.7169271600087595e-06
GC_7_284 b_7 NI_7 NS_284 0 -6.1401554701592235e-07
GC_7_285 b_7 NI_7 NS_285 0 5.6792606388942149e-06
GC_7_286 b_7 NI_7 NS_286 0 1.7812865326755582e-06
GC_7_287 b_7 NI_7 NS_287 0 3.3801496357575606e-06
GC_7_288 b_7 NI_7 NS_288 0 2.0631599266954777e-06
GC_7_289 b_7 NI_7 NS_289 0 1.0923423331254490e-05
GC_7_290 b_7 NI_7 NS_290 0 3.8982229304169792e-06
GC_7_291 b_7 NI_7 NS_291 0 4.8460147107683885e-06
GC_7_292 b_7 NI_7 NS_292 0 -4.9709687826177298e-08
GC_7_293 b_7 NI_7 NS_293 0 9.9733339305699591e-06
GC_7_294 b_7 NI_7 NS_294 0 -1.0087353174344295e-06
GC_7_295 b_7 NI_7 NS_295 0 8.2004983820208192e-06
GC_7_296 b_7 NI_7 NS_296 0 2.9626422923044113e-06
GC_7_297 b_7 NI_7 NS_297 0 1.9001978238327890e-05
GC_7_298 b_7 NI_7 NS_298 0 -5.4549101619188935e-06
GC_7_299 b_7 NI_7 NS_299 0 7.1770831496727890e-06
GC_7_300 b_7 NI_7 NS_300 0 -3.9934629514992428e-06
GC_7_301 b_7 NI_7 NS_301 0 1.3699651583989786e-05
GC_7_302 b_7 NI_7 NS_302 0 -1.1820624762517893e-05
GC_7_303 b_7 NI_7 NS_303 0 1.2324204653282462e-05
GC_7_304 b_7 NI_7 NS_304 0 -3.9604839339864568e-06
GC_7_305 b_7 NI_7 NS_305 0 9.1123486855265143e-06
GC_7_306 b_7 NI_7 NS_306 0 -2.6652120845181560e-05
GC_7_307 b_7 NI_7 NS_307 0 2.3022873208221930e-06
GC_7_308 b_7 NI_7 NS_308 0 -1.2345511296129843e-05
GC_7_309 b_7 NI_7 NS_309 0 -8.3181277144407404e-06
GC_7_310 b_7 NI_7 NS_310 0 -1.8540253186369953e-05
GC_7_311 b_7 NI_7 NS_311 0 -5.0234187730604801e-06
GC_7_312 b_7 NI_7 NS_312 0 -1.2083006440560419e-05
GC_7_313 b_7 NI_7 NS_313 0 5.5479944473029043e-05
GC_7_314 b_7 NI_7 NS_314 0 -8.7812850579345664e-05
GC_7_315 b_7 NI_7 NS_315 0 -1.0021971644718903e-05
GC_7_316 b_7 NI_7 NS_316 0 1.5204007518003601e-06
GC_7_317 b_7 NI_7 NS_317 0 3.9312421047716012e-07
GC_7_318 b_7 NI_7 NS_318 0 -1.2255150701407386e-07
GC_7_319 b_7 NI_7 NS_319 0 -2.7361008414823335e-06
GC_7_320 b_7 NI_7 NS_320 0 -1.8487249511656589e-06
GC_7_321 b_7 NI_7 NS_321 0 -4.3417378304751225e-06
GC_7_322 b_7 NI_7 NS_322 0 6.4984108977149633e-07
GC_7_323 b_7 NI_7 NS_323 0 -1.7585017188580527e-05
GC_7_324 b_7 NI_7 NS_324 0 9.5836826651943876e-06
GC_7_325 b_7 NI_7 NS_325 0 -9.3307328044960533e-06
GC_7_326 b_7 NI_7 NS_326 0 3.7420413713601040e-05
GC_7_327 b_7 NI_7 NS_327 0 -7.2143701029164127e-06
GC_7_328 b_7 NI_7 NS_328 0 3.1323464805898862e-07
GC_7_329 b_7 NI_7 NS_329 0 -1.3394815867343368e-05
GC_7_330 b_7 NI_7 NS_330 0 1.8225006353996621e-06
GC_7_331 b_7 NI_7 NS_331 0 -4.6183393044890613e-06
GC_7_332 b_7 NI_7 NS_332 0 -3.3980543668483128e-06
GC_7_333 b_7 NI_7 NS_333 0 -6.3783028965084890e-06
GC_7_334 b_7 NI_7 NS_334 0 1.0293198666757153e-06
GC_7_335 b_7 NI_7 NS_335 0 -3.0260508872381594e-06
GC_7_336 b_7 NI_7 NS_336 0 8.8999083430359657e-07
GC_7_337 b_7 NI_7 NS_337 0 -1.7736248050664465e-06
GC_7_338 b_7 NI_7 NS_338 0 -9.4941207327739369e-07
GC_7_339 b_7 NI_7 NS_339 0 -2.6169660456978880e-10
GC_7_340 b_7 NI_7 NS_340 0 4.2344984639673645e-10
GC_7_341 b_7 NI_7 NS_341 0 2.2765355998656356e-09
GC_7_342 b_7 NI_7 NS_342 0 -2.6875809354253909e-08
GC_7_343 b_7 NI_7 NS_343 0 -3.2372793675769435e-05
GC_7_344 b_7 NI_7 NS_344 0 2.2170624816836781e-06
GC_7_345 b_7 NI_7 NS_345 0 6.8027978620421370e-11
GC_7_346 b_7 NI_7 NS_346 0 3.0563821472967812e-09
GC_7_347 b_7 NI_7 NS_347 0 -1.7154493989158952e-06
GC_7_348 b_7 NI_7 NS_348 0 -1.8282394835220974e-06
GC_7_349 b_7 NI_7 NS_349 0 -5.3489870944485623e-06
GC_7_350 b_7 NI_7 NS_350 0 2.8545579486756558e-06
GC_7_351 b_7 NI_7 NS_351 0 -1.6536860512617667e-05
GC_7_352 b_7 NI_7 NS_352 0 1.8376536443352042e-05
GC_7_353 b_7 NI_7 NS_353 0 1.5065513794082128e-05
GC_7_354 b_7 NI_7 NS_354 0 9.7700004202360959e-06
GC_7_355 b_7 NI_7 NS_355 0 1.7310065515790403e-05
GC_7_356 b_7 NI_7 NS_356 0 2.2719511694977962e-05
GC_7_357 b_7 NI_7 NS_357 0 2.9106418238744251e-05
GC_7_358 b_7 NI_7 NS_358 0 4.9741088700431950e-06
GC_7_359 b_7 NI_7 NS_359 0 -2.9664953684222354e-06
GC_7_360 b_7 NI_7 NS_360 0 -1.8803163852775914e-06
GC_7_361 b_7 NI_7 NS_361 0 1.6935354701209207e-05
GC_7_362 b_7 NI_7 NS_362 0 -2.2272191577551574e-06
GC_7_363 b_7 NI_7 NS_363 0 1.2887339116148414e-04
GC_7_364 b_7 NI_7 NS_364 0 3.4716987891549303e-05
GC_7_365 b_7 NI_7 NS_365 0 -2.8880066770719539e-05
GC_7_366 b_7 NI_7 NS_366 0 -9.8668884724106948e-05
GC_7_367 b_7 NI_7 NS_367 0 2.4897333171307355e-05
GC_7_368 b_7 NI_7 NS_368 0 -3.1464745437285747e-05
GC_7_369 b_7 NI_7 NS_369 0 -4.1613526385584626e-05
GC_7_370 b_7 NI_7 NS_370 0 -1.6650660432456367e-04
GC_7_371 b_7 NI_7 NS_371 0 -4.1829246325416142e-05
GC_7_372 b_7 NI_7 NS_372 0 -4.8975553301523531e-06
GC_7_373 b_7 NI_7 NS_373 0 2.1413285400932403e-05
GC_7_374 b_7 NI_7 NS_374 0 -1.5190691096604676e-04
GC_7_375 b_7 NI_7 NS_375 0 -2.3047173609290730e-04
GC_7_376 b_7 NI_7 NS_376 0 1.1445427944248418e-04
GC_7_377 b_7 NI_7 NS_377 0 -3.7402325583902109e-05
GC_7_378 b_7 NI_7 NS_378 0 1.4353147909159939e-05
GC_7_379 b_7 NI_7 NS_379 0 -1.3776506643005027e-04
GC_7_380 b_7 NI_7 NS_380 0 1.3054867195267246e-04
GC_7_381 b_7 NI_7 NS_381 0 3.6495597907398555e-05
GC_7_382 b_7 NI_7 NS_382 0 4.1231367218348888e-05
GC_7_383 b_7 NI_7 NS_383 0 -3.8131821131968828e-05
GC_7_384 b_7 NI_7 NS_384 0 4.3361765599396536e-05
GC_7_385 b_7 NI_7 NS_385 0 8.7557362523959367e-05
GC_7_386 b_7 NI_7 NS_386 0 1.1842876064752804e-04
GC_7_387 b_7 NI_7 NS_387 0 2.7361988942612091e-05
GC_7_388 b_7 NI_7 NS_388 0 1.0121130071608856e-05
GC_7_389 b_7 NI_7 NS_389 0 8.7345264965090651e-05
GC_7_390 b_7 NI_7 NS_390 0 6.5655787961544002e-05
GC_7_391 b_7 NI_7 NS_391 0 2.0320869993186259e-05
GC_7_392 b_7 NI_7 NS_392 0 -5.7039458798704093e-05
GC_7_393 b_7 NI_7 NS_393 0 1.6979053458257079e-05
GC_7_394 b_7 NI_7 NS_394 0 -8.9186484557698138e-06
GC_7_395 b_7 NI_7 NS_395 0 8.5888456914327081e-06
GC_7_396 b_7 NI_7 NS_396 0 -3.2921175825737181e-05
GC_7_397 b_7 NI_7 NS_397 0 -8.8489257001714316e-06
GC_7_398 b_7 NI_7 NS_398 0 5.5973327772758237e-07
GC_7_399 b_7 NI_7 NS_399 0 -2.4313502166907265e-06
GC_7_400 b_7 NI_7 NS_400 0 8.5078727077167666e-06
GC_7_401 b_7 NI_7 NS_401 0 1.0241027934446232e-05
GC_7_402 b_7 NI_7 NS_402 0 6.0555285793864828e-06
GC_7_403 b_7 NI_7 NS_403 0 1.2188370687158073e-05
GC_7_404 b_7 NI_7 NS_404 0 -7.8214192982394923e-06
GC_7_405 b_7 NI_7 NS_405 0 -3.4896515207433228e-06
GC_7_406 b_7 NI_7 NS_406 0 -4.3242994459391390e-07
GC_7_407 b_7 NI_7 NS_407 0 2.4744439391553291e-06
GC_7_408 b_7 NI_7 NS_408 0 7.4084000170307223e-06
GC_7_409 b_7 NI_7 NS_409 0 1.3659441427521366e-05
GC_7_410 b_7 NI_7 NS_410 0 2.6169987568719063e-06
GC_7_411 b_7 NI_7 NS_411 0 4.5330381249675863e-06
GC_7_412 b_7 NI_7 NS_412 0 -1.4186449253844688e-05
GC_7_413 b_7 NI_7 NS_413 0 -5.9288383715752856e-06
GC_7_414 b_7 NI_7 NS_414 0 4.2661989006015329e-06
GC_7_415 b_7 NI_7 NS_415 0 1.0298083342534541e-05
GC_7_416 b_7 NI_7 NS_416 0 9.9363523172252303e-06
GC_7_417 b_7 NI_7 NS_417 0 1.7307571191362386e-05
GC_7_418 b_7 NI_7 NS_418 0 -4.2766747205646557e-06
GC_7_419 b_7 NI_7 NS_419 0 -9.2959986063347761e-06
GC_7_420 b_7 NI_7 NS_420 0 -1.5305295968264376e-05
GC_7_421 b_7 NI_7 NS_421 0 -4.0930024002385150e-06
GC_7_422 b_7 NI_7 NS_422 0 1.3520443357300372e-05
GC_7_423 b_7 NI_7 NS_423 0 2.0923711950966015e-05
GC_7_424 b_7 NI_7 NS_424 0 -5.4861416410453748e-07
GC_7_425 b_7 NI_7 NS_425 0 8.8628372349261842e-06
GC_7_426 b_7 NI_7 NS_426 0 -1.7438295562352121e-05
GC_7_427 b_7 NI_7 NS_427 0 2.5769557923970334e-06
GC_7_428 b_7 NI_7 NS_428 0 -1.3773219476720520e-05
GC_7_429 b_7 NI_7 NS_429 0 -1.3801271941799888e-05
GC_7_430 b_7 NI_7 NS_430 0 4.4172099355676620e-06
GC_7_431 b_7 NI_7 NS_431 0 1.6026938278347075e-08
GC_7_432 b_7 NI_7 NS_432 0 -4.1748330078890164e-08
GC_7_433 b_7 NI_7 NS_433 0 8.6200600656242058e-06
GC_7_434 b_7 NI_7 NS_434 0 1.1611776953423100e-05
GC_7_435 b_7 NI_7 NS_435 0 1.0921480498370843e-05
GC_7_436 b_7 NI_7 NS_436 0 -1.1277715889265224e-05
GC_7_437 b_7 NI_7 NS_437 0 -3.7556080862363798e-06
GC_7_438 b_7 NI_7 NS_438 0 -1.0184108583187385e-05
GC_7_439 b_7 NI_7 NS_439 0 -2.3203003839844270e-06
GC_7_440 b_7 NI_7 NS_440 0 1.2932028574310902e-05
GC_7_441 b_7 NI_7 NS_441 0 9.7592643620746211e-07
GC_7_442 b_7 NI_7 NS_442 0 -7.2834871420775187e-06
GC_7_443 b_7 NI_7 NS_443 0 7.5033886046929981e-06
GC_7_444 b_7 NI_7 NS_444 0 1.6764901263525001e-06
GC_7_445 b_7 NI_7 NS_445 0 -6.0990783078124833e-06
GC_7_446 b_7 NI_7 NS_446 0 -8.8899526074007653e-06
GC_7_447 b_7 NI_7 NS_447 0 -4.1231996937442593e-06
GC_7_448 b_7 NI_7 NS_448 0 9.6572565344449938e-06
GC_7_449 b_7 NI_7 NS_449 0 3.3299269741274347e-06
GC_7_450 b_7 NI_7 NS_450 0 6.0429561035493425e-06
GC_7_451 b_7 NI_7 NS_451 0 5.6621074359150492e-06
GC_7_452 b_7 NI_7 NS_452 0 5.1491103758648471e-07
GC_7_453 b_7 NI_7 NS_453 0 6.1217261406704931e-11
GC_7_454 b_7 NI_7 NS_454 0 1.4945694433861397e-10
GC_7_455 b_7 NI_7 NS_455 0 5.9799730470138591e-09
GC_7_456 b_7 NI_7 NS_456 0 -8.3554688903502913e-09
GC_7_457 b_7 NI_7 NS_457 0 7.9886719687266468e-03
GC_7_458 b_7 NI_7 NS_458 0 -1.6009906150823261e-03
GC_7_459 b_7 NI_7 NS_459 0 -1.2329825313203087e-08
GC_7_460 b_7 NI_7 NS_460 0 -8.8365943464764703e-07
GC_7_461 b_7 NI_7 NS_461 0 1.0714040963905273e-04
GC_7_462 b_7 NI_7 NS_462 0 -5.1251769106129259e-04
GC_7_463 b_7 NI_7 NS_463 0 -1.9321158080111735e-03
GC_7_464 b_7 NI_7 NS_464 0 -5.9632008157690084e-04
GC_7_465 b_7 NI_7 NS_465 0 2.9522602817683378e-03
GC_7_466 b_7 NI_7 NS_466 0 2.2413628932075177e-03
GC_7_467 b_7 NI_7 NS_467 0 -3.5853198938722280e-03
GC_7_468 b_7 NI_7 NS_468 0 -3.0463419434418994e-03
GC_7_469 b_7 NI_7 NS_469 0 -1.6953804455786278e-03
GC_7_470 b_7 NI_7 NS_470 0 5.8334393037870217e-03
GC_7_471 b_7 NI_7 NS_471 0 4.3284000323277711e-03
GC_7_472 b_7 NI_7 NS_472 0 -2.4949638253823044e-03
GC_7_473 b_7 NI_7 NS_473 0 -1.0252417147585616e-04
GC_7_474 b_7 NI_7 NS_474 0 -9.7511922486949928e-05
GC_7_475 b_7 NI_7 NS_475 0 -4.4595016515740311e-03
GC_7_476 b_7 NI_7 NS_476 0 -9.0945578566390946e-04
GC_7_477 b_7 NI_7 NS_477 0 9.1489031895608114e-03
GC_7_478 b_7 NI_7 NS_478 0 1.7749054711310407e-02
GC_7_479 b_7 NI_7 NS_479 0 -4.0759917605376643e-03
GC_7_480 b_7 NI_7 NS_480 0 -1.7815996220547831e-02
GC_7_481 b_7 NI_7 NS_481 0 -8.2086049937415903e-03
GC_7_482 b_7 NI_7 NS_482 0 4.1974764949610768e-03
GC_7_483 b_7 NI_7 NS_483 0 1.7045926420419414e-02
GC_7_484 b_7 NI_7 NS_484 0 -4.7587325095690757e-04
GC_7_485 b_7 NI_7 NS_485 0 -9.2871622325277261e-03
GC_7_486 b_7 NI_7 NS_486 0 -3.1746356711356018e-03
GC_7_487 b_7 NI_7 NS_487 0 -1.3650847444118451e-02
GC_7_488 b_7 NI_7 NS_488 0 2.2873426934236631e-02
GC_7_489 b_7 NI_7 NS_489 0 2.2768615047399743e-02
GC_7_490 b_7 NI_7 NS_490 0 -2.2718066479614066e-02
GC_7_491 b_7 NI_7 NS_491 0 -9.2369617601131045e-03
GC_7_492 b_7 NI_7 NS_492 0 9.4042622149346643e-04
GC_7_493 b_7 NI_7 NS_493 0 1.8496821945441961e-02
GC_7_494 b_7 NI_7 NS_494 0 6.1966524487003230e-03
GC_7_495 b_7 NI_7 NS_495 0 -9.2042290959818938e-03
GC_7_496 b_7 NI_7 NS_496 0 -9.4288117669458025e-03
GC_7_497 b_7 NI_7 NS_497 0 -9.9569355412411319e-03
GC_7_498 b_7 NI_7 NS_498 0 6.4309790696960552e-03
GC_7_499 b_7 NI_7 NS_499 0 1.6827172547774764e-02
GC_7_500 b_7 NI_7 NS_500 0 -4.8950436115088071e-03
GC_7_501 b_7 NI_7 NS_501 0 -7.2263301001000719e-03
GC_7_502 b_7 NI_7 NS_502 0 -3.3851923812586305e-03
GC_7_503 b_7 NI_7 NS_503 0 6.8657294726293385e-03
GC_7_504 b_7 NI_7 NS_504 0 1.3286490499213545e-02
GC_7_505 b_7 NI_7 NS_505 0 -1.8581882790271163e-03
GC_7_506 b_7 NI_7 NS_506 0 -1.4397044017763719e-02
GC_7_507 b_7 NI_7 NS_507 0 -4.9859100379437485e-03
GC_7_508 b_7 NI_7 NS_508 0 1.0545183001181540e-03
GC_7_509 b_7 NI_7 NS_509 0 6.0007405850145039e-03
GC_7_510 b_7 NI_7 NS_510 0 -1.1126545527218486e-03
GC_7_511 b_7 NI_7 NS_511 0 -3.4683253362858234e-03
GC_7_512 b_7 NI_7 NS_512 0 -1.0780499140241905e-03
GC_7_513 b_7 NI_7 NS_513 0 2.7173467250648019e-03
GC_7_514 b_7 NI_7 NS_514 0 -5.1095685090648527e-04
GC_7_515 b_7 NI_7 NS_515 0 -3.3053412650086182e-03
GC_7_516 b_7 NI_7 NS_516 0 -2.8885150449347230e-03
GC_7_517 b_7 NI_7 NS_517 0 2.0156340091641960e-03
GC_7_518 b_7 NI_7 NS_518 0 7.7768287470312224e-04
GC_7_519 b_7 NI_7 NS_519 0 -2.0192451145490406e-03
GC_7_520 b_7 NI_7 NS_520 0 -9.6218740624151307e-04
GC_7_521 b_7 NI_7 NS_521 0 2.1198804234619558e-03
GC_7_522 b_7 NI_7 NS_522 0 -1.4705676421229831e-03
GC_7_523 b_7 NI_7 NS_523 0 -4.1910213331247488e-03
GC_7_524 b_7 NI_7 NS_524 0 -1.8092507391981442e-03
GC_7_525 b_7 NI_7 NS_525 0 2.3672939662825270e-03
GC_7_526 b_7 NI_7 NS_526 0 -3.6739652555426171e-04
GC_7_527 b_7 NI_7 NS_527 0 -3.0199644103893878e-03
GC_7_528 b_7 NI_7 NS_528 0 4.6494719814711943e-04
GC_7_529 b_7 NI_7 NS_529 0 2.7038550449039562e-03
GC_7_530 b_7 NI_7 NS_530 0 -2.7263252666909770e-03
GC_7_531 b_7 NI_7 NS_531 0 -5.0450291670743755e-03
GC_7_532 b_7 NI_7 NS_532 0 -1.2988616762432291e-04
GC_7_533 b_7 NI_7 NS_533 0 2.4275289935295806e-03
GC_7_534 b_7 NI_7 NS_534 0 -2.1667278995723548e-03
GC_7_535 b_7 NI_7 NS_535 0 -3.2524101809915723e-03
GC_7_536 b_7 NI_7 NS_536 0 2.6001222852165681e-03
GC_7_537 b_7 NI_7 NS_537 0 1.7373702982732264e-03
GC_7_538 b_7 NI_7 NS_538 0 -4.7433400124927355e-03
GC_7_539 b_7 NI_7 NS_539 0 -3.6476875004110092e-03
GC_7_540 b_7 NI_7 NS_540 0 2.5904970938509944e-03
GC_7_541 b_7 NI_7 NS_541 0 -2.8140502655213716e-03
GC_7_542 b_7 NI_7 NS_542 0 4.0553534803892460e-03
GC_7_543 b_7 NI_7 NS_543 0 -2.3077990758292572e-04
GC_7_544 b_7 NI_7 NS_544 0 -4.1951360936145288e-03
GC_7_545 b_7 NI_7 NS_545 0 -9.8757636544501269e-06
GC_7_546 b_7 NI_7 NS_546 0 7.9025145318081258e-06
GC_7_547 b_7 NI_7 NS_547 0 -1.3634151928128525e-03
GC_7_548 b_7 NI_7 NS_548 0 3.3837800378031975e-03
GC_7_549 b_7 NI_7 NS_549 0 -9.6978193674661427e-04
GC_7_550 b_7 NI_7 NS_550 0 -4.3384320742976901e-03
GC_7_551 b_7 NI_7 NS_551 0 -1.0095575941227899e-03
GC_7_552 b_7 NI_7 NS_552 0 2.2144692343813123e-03
GC_7_553 b_7 NI_7 NS_553 0 -1.6625797156473046e-03
GC_7_554 b_7 NI_7 NS_554 0 -4.4181655959373714e-03
GC_7_555 b_7 NI_7 NS_555 0 -1.4450239319927873e-03
GC_7_556 b_7 NI_7 NS_556 0 -2.4969806502863779e-03
GC_7_557 b_7 NI_7 NS_557 0 7.8582136666740165e-04
GC_7_558 b_7 NI_7 NS_558 0 2.5922239268502865e-03
GC_7_559 b_7 NI_7 NS_559 0 -6.9658839312940007e-04
GC_7_560 b_7 NI_7 NS_560 0 2.8805416718650518e-03
GC_7_561 b_7 NI_7 NS_561 0 -1.4341253052850243e-03
GC_7_562 b_7 NI_7 NS_562 0 -2.7701138532130187e-03
GC_7_563 b_7 NI_7 NS_563 0 -1.1685605976010783e-03
GC_7_564 b_7 NI_7 NS_564 0 2.6674409169131453e-03
GC_7_565 b_7 NI_7 NS_565 0 7.8095042626851233e-04
GC_7_566 b_7 NI_7 NS_566 0 -1.8732339647521070e-03
GC_7_567 b_7 NI_7 NS_567 0 2.4009828839562907e-08
GC_7_568 b_7 NI_7 NS_568 0 -6.0310105547878327e-08
GC_7_569 b_7 NI_7 NS_569 0 -9.0615470945560529e-07
GC_7_570 b_7 NI_7 NS_570 0 3.2140038429780433e-06
GC_7_571 b_7 NI_7 NS_571 0 3.0950442684637689e-03
GC_7_572 b_7 NI_7 NS_572 0 -6.1289418565353064e-04
GC_7_573 b_7 NI_7 NS_573 0 2.8121770040342655e-08
GC_7_574 b_7 NI_7 NS_574 0 -3.1528708375438252e-08
GC_7_575 b_7 NI_7 NS_575 0 2.0500773537449369e-04
GC_7_576 b_7 NI_7 NS_576 0 1.3546540067660017e-04
GC_7_577 b_7 NI_7 NS_577 0 5.6415263403009920e-04
GC_7_578 b_7 NI_7 NS_578 0 2.6382413588216193e-04
GC_7_579 b_7 NI_7 NS_579 0 3.0949151549668013e-03
GC_7_580 b_7 NI_7 NS_580 0 -2.2211775627329808e-03
GC_7_581 b_7 NI_7 NS_581 0 -1.5948050035838408e-03
GC_7_582 b_7 NI_7 NS_582 0 -2.6831568726140829e-03
GC_7_583 b_7 NI_7 NS_583 0 -2.0664405370191857e-03
GC_7_584 b_7 NI_7 NS_584 0 -3.7810168676189805e-03
GC_7_585 b_7 NI_7 NS_585 0 -4.9930248682110937e-03
GC_7_586 b_7 NI_7 NS_586 0 -1.5154929244419533e-03
GC_7_587 b_7 NI_7 NS_587 0 2.9714197312462673e-04
GC_7_588 b_7 NI_7 NS_588 0 1.9409424377540510e-04
GC_7_589 b_7 NI_7 NS_589 0 -2.8708432790663062e-03
GC_7_590 b_7 NI_7 NS_590 0 -9.4557935639995880e-04
GC_7_591 b_7 NI_7 NS_591 0 -2.2198356450817740e-02
GC_7_592 b_7 NI_7 NS_592 0 -1.0125161751702071e-02
GC_7_593 b_7 NI_7 NS_593 0 1.2231803991193074e-03
GC_7_594 b_7 NI_7 NS_594 0 2.0396448916834346e-02
GC_7_595 b_7 NI_7 NS_595 0 -5.8225964768853526e-03
GC_7_596 b_7 NI_7 NS_596 0 4.6364311860234734e-03
GC_7_597 b_7 NI_7 NS_597 0 5.8808187670633828e-03
GC_7_598 b_7 NI_7 NS_598 0 3.4493744006799471e-02
GC_7_599 b_7 NI_7 NS_599 0 8.0480772505822865e-03
GC_7_600 b_7 NI_7 NS_600 0 2.7589349736136890e-03
GC_7_601 b_7 NI_7 NS_601 0 -7.6367957306050704e-03
GC_7_602 b_7 NI_7 NS_602 0 2.9591949318747611e-02
GC_7_603 b_7 NI_7 NS_603 0 5.0679464975272162e-02
GC_7_604 b_7 NI_7 NS_604 0 -2.0315740121607310e-02
GC_7_605 b_7 NI_7 NS_605 0 7.9122592824869085e-03
GC_7_606 b_7 NI_7 NS_606 0 -1.6718962437624119e-03
GC_7_607 b_7 NI_7 NS_607 0 2.8952184642265309e-02
GC_7_608 b_7 NI_7 NS_608 0 -2.6605126130389931e-02
GC_7_609 b_7 NI_7 NS_609 0 -6.7717822704580306e-03
GC_7_610 b_7 NI_7 NS_610 0 -9.8521000565271986e-03
GC_7_611 b_7 NI_7 NS_611 0 8.4245547512454711e-03
GC_7_612 b_7 NI_7 NS_612 0 -8.0661005349519956e-03
GC_7_613 b_7 NI_7 NS_613 0 -1.9120467233820587e-02
GC_7_614 b_7 NI_7 NS_614 0 -2.5143595159399457e-02
GC_7_615 b_7 NI_7 NS_615 0 -5.4851138485096556e-03
GC_7_616 b_7 NI_7 NS_616 0 -2.8303874885823427e-03
GC_7_617 b_7 NI_7 NS_617 0 -1.7803813193018086e-02
GC_7_618 b_7 NI_7 NS_618 0 -1.3047348691410436e-02
GC_7_619 b_7 NI_7 NS_619 0 -4.7610274735247673e-03
GC_7_620 b_7 NI_7 NS_620 0 1.2568312179295930e-02
GC_7_621 b_7 NI_7 NS_621 0 -3.4539895302149216e-03
GC_7_622 b_7 NI_7 NS_622 0 1.5560260535347045e-03
GC_7_623 b_7 NI_7 NS_623 0 -6.8744301160818852e-04
GC_7_624 b_7 NI_7 NS_624 0 7.0157646198823961e-03
GC_7_625 b_7 NI_7 NS_625 0 1.8840812938743672e-03
GC_7_626 b_7 NI_7 NS_626 0 8.1060422034459124e-05
GC_7_627 b_7 NI_7 NS_627 0 3.0821856660416725e-04
GC_7_628 b_7 NI_7 NS_628 0 -1.9474452512085389e-03
GC_7_629 b_7 NI_7 NS_629 0 -1.8615158836804292e-03
GC_7_630 b_7 NI_7 NS_630 0 -1.6133456398352728e-03
GC_7_631 b_7 NI_7 NS_631 0 -2.1255689831030998e-03
GC_7_632 b_7 NI_7 NS_632 0 1.6940535977075833e-03
GC_7_633 b_7 NI_7 NS_633 0 7.6441486570389902e-04
GC_7_634 b_7 NI_7 NS_634 0 1.8569487153379248e-04
GC_7_635 b_7 NI_7 NS_635 0 -7.0068912884497700e-04
GC_7_636 b_7 NI_7 NS_636 0 -1.6760054883672331e-03
GC_7_637 b_7 NI_7 NS_637 0 -2.6855352118105341e-03
GC_7_638 b_7 NI_7 NS_638 0 -8.2394391646450156e-04
GC_7_639 b_7 NI_7 NS_639 0 -4.9849901251835345e-04
GC_7_640 b_7 NI_7 NS_640 0 2.9352188065828711e-03
GC_7_641 b_7 NI_7 NS_641 0 1.3528909970584714e-03
GC_7_642 b_7 NI_7 NS_642 0 -8.5706936120598116e-04
GC_7_643 b_7 NI_7 NS_643 0 -2.4223433422766818e-03
GC_7_644 b_7 NI_7 NS_644 0 -2.2652834647004906e-03
GC_7_645 b_7 NI_7 NS_645 0 -3.5590211448898431e-03
GC_7_646 b_7 NI_7 NS_646 0 7.4879944628055664e-04
GC_7_647 b_7 NI_7 NS_647 0 2.4605502070294822e-03
GC_7_648 b_7 NI_7 NS_648 0 3.0265645572291468e-03
GC_7_649 b_7 NI_7 NS_649 0 9.8335647412217220e-04
GC_7_650 b_7 NI_7 NS_650 0 -2.9400791196709047e-03
GC_7_651 b_7 NI_7 NS_651 0 -4.7724967890530262e-03
GC_7_652 b_7 NI_7 NS_652 0 5.7213638812192586e-05
GC_7_653 b_7 NI_7 NS_653 0 -1.7194839186640846e-03
GC_7_654 b_7 NI_7 NS_654 0 3.7113727622575536e-03
GC_7_655 b_7 NI_7 NS_655 0 -7.3866503981761427e-04
GC_7_656 b_7 NI_7 NS_656 0 1.5326962516858823e-03
GC_7_657 b_7 NI_7 NS_657 0 3.2195727081450842e-03
GC_7_658 b_7 NI_7 NS_658 0 -1.3349984962042201e-03
GC_7_659 b_7 NI_7 NS_659 0 -2.8022744863773488e-06
GC_7_660 b_7 NI_7 NS_660 0 8.9859893355038973e-06
GC_7_661 b_7 NI_7 NS_661 0 -1.8210613106944347e-03
GC_7_662 b_7 NI_7 NS_662 0 -2.5224003501537356e-03
GC_7_663 b_7 NI_7 NS_663 0 -2.4088301415847433e-03
GC_7_664 b_7 NI_7 NS_664 0 2.4933225812579884e-03
GC_7_665 b_7 NI_7 NS_665 0 1.0059037045019317e-03
GC_7_666 b_7 NI_7 NS_666 0 2.4239841912818559e-03
GC_7_667 b_7 NI_7 NS_667 0 8.4854727983707892e-04
GC_7_668 b_7 NI_7 NS_668 0 -2.6997865154174635e-03
GC_7_669 b_7 NI_7 NS_669 0 -3.0628340201132090e-04
GC_7_670 b_7 NI_7 NS_670 0 1.6736613642944682e-03
GC_7_671 b_7 NI_7 NS_671 0 -1.7824227358932520e-03
GC_7_672 b_7 NI_7 NS_672 0 -3.1430319732621211e-04
GC_7_673 b_7 NI_7 NS_673 0 1.3997488467847605e-03
GC_7_674 b_7 NI_7 NS_674 0 1.9719385369297336e-03
GC_7_675 b_7 NI_7 NS_675 0 1.0457174689825668e-03
GC_7_676 b_7 NI_7 NS_676 0 -2.2988262166401927e-03
GC_7_677 b_7 NI_7 NS_677 0 -6.9831747326666224e-04
GC_7_678 b_7 NI_7 NS_678 0 -1.4663462692674385e-03
GC_7_679 b_7 NI_7 NS_679 0 -1.3735955652843634e-03
GC_7_680 b_7 NI_7 NS_680 0 -3.1257035693694839e-04
GC_7_681 b_7 NI_7 NS_681 0 6.7938444254092591e-09
GC_7_682 b_7 NI_7 NS_682 0 -2.4700012038159102e-08
GC_7_683 b_7 NI_7 NS_683 0 -4.4377037472335511e-07
GC_7_684 b_7 NI_7 NS_684 0 1.6205767041468295e-06
GC_7_685 b_7 NI_7 NS_685 0 -1.2879661893680934e-02
GC_7_686 b_7 NI_7 NS_686 0 1.3854988955549130e-03
GC_7_687 b_7 NI_7 NS_687 0 -2.6205633593858005e-07
GC_7_688 b_7 NI_7 NS_688 0 -3.7467198181028706e-06
GC_7_689 b_7 NI_7 NS_689 0 -2.6866989055314156e-04
GC_7_690 b_7 NI_7 NS_690 0 4.6434496467892680e-04
GC_7_691 b_7 NI_7 NS_691 0 1.3324545855155981e-03
GC_7_692 b_7 NI_7 NS_692 0 5.3749686531473473e-04
GC_7_693 b_7 NI_7 NS_693 0 -2.7601218902434522e-03
GC_7_694 b_7 NI_7 NS_694 0 -8.2597386150402288e-04
GC_7_695 b_7 NI_7 NS_695 0 3.5364630190112636e-03
GC_7_696 b_7 NI_7 NS_696 0 2.5065964003169227e-03
GC_7_697 b_7 NI_7 NS_697 0 1.1567014953989302e-03
GC_7_698 b_7 NI_7 NS_698 0 -4.2275297822350101e-03
GC_7_699 b_7 NI_7 NS_699 0 -1.7809474208909243e-03
GC_7_700 b_7 NI_7 NS_700 0 2.6938537326557425e-03
GC_7_701 b_7 NI_7 NS_701 0 -3.0415845838287475e-04
GC_7_702 b_7 NI_7 NS_702 0 -1.8023605520433862e-04
GC_7_703 b_7 NI_7 NS_703 0 3.9634813471252951e-03
GC_7_704 b_7 NI_7 NS_704 0 2.8124797281969984e-04
GC_7_705 b_7 NI_7 NS_705 0 -7.5492073290113421e-03
GC_7_706 b_7 NI_7 NS_706 0 -1.3596105032115028e-02
GC_7_707 b_7 NI_7 NS_707 0 4.4801999487899058e-03
GC_7_708 b_7 NI_7 NS_708 0 1.3516145121002989e-02
GC_7_709 b_7 NI_7 NS_709 0 6.6864828442972004e-03
GC_7_710 b_7 NI_7 NS_710 0 -4.0243772389796572e-03
GC_7_711 b_7 NI_7 NS_711 0 -1.3410282976857637e-02
GC_7_712 b_7 NI_7 NS_712 0 7.8159746019152234e-04
GC_7_713 b_7 NI_7 NS_713 0 7.8563500433258583e-03
GC_7_714 b_7 NI_7 NS_714 0 1.8570145277325496e-03
GC_7_715 b_7 NI_7 NS_715 0 1.0427285557680787e-02
GC_7_716 b_7 NI_7 NS_716 0 -1.9666904344150672e-02
GC_7_717 b_7 NI_7 NS_717 0 -1.7708800298312597e-02
GC_7_718 b_7 NI_7 NS_718 0 1.9274360121932153e-02
GC_7_719 b_7 NI_7 NS_719 0 7.6729361596684295e-03
GC_7_720 b_7 NI_7 NS_720 0 -1.4539298525646294e-03
GC_7_721 b_7 NI_7 NS_721 0 -1.5685670877969335e-02
GC_7_722 b_7 NI_7 NS_722 0 -4.6645791485753502e-03
GC_7_723 b_7 NI_7 NS_723 0 8.1074614701308161e-03
GC_7_724 b_7 NI_7 NS_724 0 7.2499038698249293e-03
GC_7_725 b_7 NI_7 NS_725 0 8.0870945772521258e-03
GC_7_726 b_7 NI_7 NS_726 0 -6.0421323777582201e-03
GC_7_727 b_7 NI_7 NS_727 0 -1.3963410688590893e-02
GC_7_728 b_7 NI_7 NS_728 0 4.6523251530976315e-03
GC_7_729 b_7 NI_7 NS_729 0 6.2461630182085509e-03
GC_7_730 b_7 NI_7 NS_730 0 2.3807828503421983e-03
GC_7_731 b_7 NI_7 NS_731 0 -6.3453899443727969e-03
GC_7_732 b_7 NI_7 NS_732 0 -1.1079783746456554e-02
GC_7_733 b_7 NI_7 NS_733 0 2.1863328123651947e-03
GC_7_734 b_7 NI_7 NS_734 0 1.1948129394737978e-02
GC_7_735 b_7 NI_7 NS_735 0 4.2064703276400483e-03
GC_7_736 b_7 NI_7 NS_736 0 -1.1782772225451279e-03
GC_7_737 b_7 NI_7 NS_737 0 -4.9335527767871562e-03
GC_7_738 b_7 NI_7 NS_738 0 1.0766011735707035e-03
GC_7_739 b_7 NI_7 NS_739 0 3.0283700722116540e-03
GC_7_740 b_7 NI_7 NS_740 0 6.9130831203059924e-04
GC_7_741 b_7 NI_7 NS_741 0 -2.2217200917590755e-03
GC_7_742 b_7 NI_7 NS_742 0 5.0249262505259811e-04
GC_7_743 b_7 NI_7 NS_743 0 3.0726777265681435e-03
GC_7_744 b_7 NI_7 NS_744 0 2.2985803293223478e-03
GC_7_745 b_7 NI_7 NS_745 0 -1.5387652809863699e-03
GC_7_746 b_7 NI_7 NS_746 0 -6.6609294789863672e-04
GC_7_747 b_7 NI_7 NS_747 0 1.8890934059918336e-03
GC_7_748 b_7 NI_7 NS_748 0 6.8215091802094937e-04
GC_7_749 b_7 NI_7 NS_749 0 -1.5634721390540408e-03
GC_7_750 b_7 NI_7 NS_750 0 1.2301006580442344e-03
GC_7_751 b_7 NI_7 NS_751 0 3.9777148057023558e-03
GC_7_752 b_7 NI_7 NS_752 0 1.4029339285898073e-03
GC_7_753 b_7 NI_7 NS_753 0 -1.5582641540631832e-03
GC_7_754 b_7 NI_7 NS_754 0 7.6118044831076411e-05
GC_7_755 b_7 NI_7 NS_755 0 2.8289105703623767e-03
GC_7_756 b_7 NI_7 NS_756 0 -6.8710742116771903e-04
GC_7_757 b_7 NI_7 NS_757 0 -1.8835368104045142e-03
GC_7_758 b_7 NI_7 NS_758 0 2.0120377226582834e-03
GC_7_759 b_7 NI_7 NS_759 0 4.9081314997195527e-03
GC_7_760 b_7 NI_7 NS_760 0 -1.8224246863975143e-04
GC_7_761 b_7 NI_7 NS_761 0 -1.6649296084399012e-03
GC_7_762 b_7 NI_7 NS_762 0 9.3127546830156763e-04
GC_7_763 b_7 NI_7 NS_763 0 3.0639871877217134e-03
GC_7_764 b_7 NI_7 NS_764 0 -2.8461960120540119e-03
GC_7_765 b_7 NI_7 NS_765 0 -1.4669304701028073e-03
GC_7_766 b_7 NI_7 NS_766 0 3.2252900410917858e-03
GC_7_767 b_7 NI_7 NS_767 0 3.7966921645121439e-03
GC_7_768 b_7 NI_7 NS_768 0 -2.9822109805926690e-03
GC_7_769 b_7 NI_7 NS_769 0 -1.8554837958068560e-03
GC_7_770 b_7 NI_7 NS_770 0 -3.8335174704752098e-03
GC_7_771 b_7 NI_7 NS_771 0 -4.1823215155716828e-04
GC_7_772 b_7 NI_7 NS_772 0 2.3792558316471351e-03
GC_7_773 b_7 NI_7 NS_773 0 -1.0537744852492320e-05
GC_7_774 b_7 NI_7 NS_774 0 -2.1100618635940101e-05
GC_7_775 b_7 NI_7 NS_775 0 8.3839973512957351e-04
GC_7_776 b_7 NI_7 NS_776 0 -3.7904895272166620e-03
GC_7_777 b_7 NI_7 NS_777 0 3.3770948816713774e-04
GC_7_778 b_7 NI_7 NS_778 0 3.3559461662644812e-03
GC_7_779 b_7 NI_7 NS_779 0 1.3516061376476706e-03
GC_7_780 b_7 NI_7 NS_780 0 -2.3818220972734333e-03
GC_7_781 b_7 NI_7 NS_781 0 2.1706557714886890e-03
GC_7_782 b_7 NI_7 NS_782 0 3.3305696475555871e-03
GC_7_783 b_7 NI_7 NS_783 0 1.1698305133410849e-03
GC_7_784 b_7 NI_7 NS_784 0 2.4039647807662296e-03
GC_7_785 b_7 NI_7 NS_785 0 -8.0769436557370062e-04
GC_7_786 b_7 NI_7 NS_786 0 -1.9803395337626233e-03
GC_7_787 b_7 NI_7 NS_787 0 3.9764806952550017e-04
GC_7_788 b_7 NI_7 NS_788 0 -2.6820412711366500e-03
GC_7_789 b_7 NI_7 NS_789 0 9.8318323283809613e-04
GC_7_790 b_7 NI_7 NS_790 0 2.7477869287563547e-03
GC_7_791 b_7 NI_7 NS_791 0 1.0389080540843193e-03
GC_7_792 b_7 NI_7 NS_792 0 -2.4201775873018898e-03
GC_7_793 b_7 NI_7 NS_793 0 -1.0840508105159909e-03
GC_7_794 b_7 NI_7 NS_794 0 1.5933775231735778e-03
GC_7_795 b_7 NI_7 NS_795 0 -1.0740497992730731e-08
GC_7_796 b_7 NI_7 NS_796 0 -2.7688799863433892e-09
GC_7_797 b_7 NI_7 NS_797 0 2.2912016356065106e-06
GC_7_798 b_7 NI_7 NS_798 0 5.4762552454809914e-07
GC_7_799 b_7 NI_7 NS_799 0 1.8114453226673231e-02
GC_7_800 b_7 NI_7 NS_800 0 6.7504807670764888e-03
GC_7_801 b_7 NI_7 NS_801 0 4.7185838901615210e-07
GC_7_802 b_7 NI_7 NS_802 0 1.4478146766472033e-06
GC_7_803 b_7 NI_7 NS_803 0 6.0855570153400792e-03
GC_7_804 b_7 NI_7 NS_804 0 1.8096281666483943e-03
GC_7_805 b_7 NI_7 NS_805 0 -6.0720763787918894e-03
GC_7_806 b_7 NI_7 NS_806 0 -6.1692308651105148e-04
GC_7_807 b_7 NI_7 NS_807 0 7.3059161917041603e-03
GC_7_808 b_7 NI_7 NS_808 0 -1.2857310792729891e-02
GC_7_809 b_7 NI_7 NS_809 0 8.4528509146803016e-03
GC_7_810 b_7 NI_7 NS_810 0 -2.4018299117496643e-04
GC_7_811 b_7 NI_7 NS_811 0 -9.6390517778220039e-03
GC_7_812 b_7 NI_7 NS_812 0 2.6170999104785943e-03
GC_7_813 b_7 NI_7 NS_813 0 -8.8461869723790026e-03
GC_7_814 b_7 NI_7 NS_814 0 -2.4392848205199959e-02
GC_7_815 b_7 NI_7 NS_815 0 -8.6514785384649647e-04
GC_7_816 b_7 NI_7 NS_816 0 4.1785438271907827e-03
GC_7_817 b_7 NI_7 NS_817 0 7.1897714477587851e-03
GC_7_818 b_7 NI_7 NS_818 0 -1.0341053058489831e-03
GC_7_819 b_7 NI_7 NS_819 0 -2.5138553899410915e-02
GC_7_820 b_7 NI_7 NS_820 0 4.8071732780239568e-03
GC_7_821 b_7 NI_7 NS_821 0 -1.9700987247524799e-02
GC_7_822 b_7 NI_7 NS_822 0 8.9735936175270507e-04
GC_7_823 b_7 NI_7 NS_823 0 1.0752518976102793e-02
GC_7_824 b_7 NI_7 NS_824 0 -2.7940112556708060e-03
GC_7_825 b_7 NI_7 NS_825 0 -4.8190401483415232e-03
GC_7_826 b_7 NI_7 NS_826 0 4.5027436449813565e-02
GC_7_827 b_7 NI_7 NS_827 0 -1.2658610064434000e-02
GC_7_828 b_7 NI_7 NS_828 0 -2.5618591238404963e-04
GC_7_829 b_7 NI_7 NS_829 0 1.5863299541746759e-02
GC_7_830 b_7 NI_7 NS_830 0 -4.0664285067586684e-03
GC_7_831 b_7 NI_7 NS_831 0 3.2252266544197356e-02
GC_7_832 b_7 NI_7 NS_832 0 1.8644473023156336e-02
GC_7_833 b_7 NI_7 NS_833 0 -1.2591686149973691e-02
GC_7_834 b_7 NI_7 NS_834 0 1.8230672190865192e-04
GC_7_835 b_7 NI_7 NS_835 0 1.7239485177595507e-02
GC_7_836 b_7 NI_7 NS_836 0 -3.5124416646108193e-02
GC_7_837 b_7 NI_7 NS_837 0 1.4036136938523633e-02
GC_7_838 b_7 NI_7 NS_838 0 4.7591239413197128e-03
GC_7_839 b_7 NI_7 NS_839 0 -1.4382230015446227e-02
GC_7_840 b_7 NI_7 NS_840 0 2.6524601856178673e-04
GC_7_841 b_7 NI_7 NS_841 0 -2.0118060730498138e-02
GC_7_842 b_7 NI_7 NS_842 0 -3.0219205214744114e-02
GC_7_843 b_7 NI_7 NS_843 0 1.0538956622975501e-02
GC_7_844 b_7 NI_7 NS_844 0 3.5722837624055735e-03
GC_7_845 b_7 NI_7 NS_845 0 -2.6760812146001480e-02
GC_7_846 b_7 NI_7 NS_846 0 1.1130911202411223e-02
GC_7_847 b_7 NI_7 NS_847 0 -1.4164619180419190e-02
GC_7_848 b_7 NI_7 NS_848 0 -2.5194117149935293e-03
GC_7_849 b_7 NI_7 NS_849 0 7.5549284906765027e-03
GC_7_850 b_7 NI_7 NS_850 0 1.5797727451596847e-03
GC_7_851 b_7 NI_7 NS_851 0 -8.4944448061915578e-04
GC_7_852 b_7 NI_7 NS_852 0 2.4400465946428952e-02
GC_7_853 b_7 NI_7 NS_853 0 -7.6205562972541715e-03
GC_7_854 b_7 NI_7 NS_854 0 2.8886852016848051e-04
GC_7_855 b_7 NI_7 NS_855 0 -5.5962406400904469e-04
GC_7_856 b_7 NI_7 NS_856 0 -5.5377854081859164e-03
GC_7_857 b_7 NI_7 NS_857 0 8.2746292920411069e-03
GC_7_858 b_7 NI_7 NS_858 0 7.0134918747095237e-03
GC_7_859 b_7 NI_7 NS_859 0 -7.1244137286421961e-04
GC_7_860 b_7 NI_7 NS_860 0 1.2089367151269084e-02
GC_7_861 b_7 NI_7 NS_861 0 -5.1470067045460768e-03
GC_7_862 b_7 NI_7 NS_862 0 -1.3514292376944683e-04
GC_7_863 b_7 NI_7 NS_863 0 -1.8292638883539870e-03
GC_7_864 b_7 NI_7 NS_864 0 -5.1716236513630713e-03
GC_7_865 b_7 NI_7 NS_865 0 9.2943102636775868e-03
GC_7_866 b_7 NI_7 NS_866 0 5.4122832503363779e-03
GC_7_867 b_7 NI_7 NS_867 0 3.5222751302210029e-03
GC_7_868 b_7 NI_7 NS_868 0 1.1687362959038510e-02
GC_7_869 b_7 NI_7 NS_869 0 -6.1347804377410295e-03
GC_7_870 b_7 NI_7 NS_870 0 1.4299338284181934e-03
GC_7_871 b_7 NI_7 NS_871 0 -2.8132644133933632e-03
GC_7_872 b_7 NI_7 NS_872 0 -7.3476306859369582e-03
GC_7_873 b_7 NI_7 NS_873 0 9.9612926012584632e-03
GC_7_874 b_7 NI_7 NS_874 0 3.3711731333915646e-03
GC_7_875 b_7 NI_7 NS_875 0 8.1789533103228066e-03
GC_7_876 b_7 NI_7 NS_876 0 1.0242331027861944e-02
GC_7_877 b_7 NI_7 NS_877 0 -6.9808873946418607e-03
GC_7_878 b_7 NI_7 NS_878 0 2.9381312540351224e-03
GC_7_879 b_7 NI_7 NS_879 0 -5.6228582438039706e-03
GC_7_880 b_7 NI_7 NS_880 0 -8.0957312219860009e-03
GC_7_881 b_7 NI_7 NS_881 0 9.8673473079405570e-03
GC_7_882 b_7 NI_7 NS_882 0 5.6089003737183705e-04
GC_7_883 b_7 NI_7 NS_883 0 -1.0918841486865930e-02
GC_7_884 b_7 NI_7 NS_884 0 1.2173852126391086e-02
GC_7_885 b_7 NI_7 NS_885 0 9.6705226780212025e-03
GC_7_886 b_7 NI_7 NS_886 0 5.0263891167489074e-03
GC_7_887 b_7 NI_7 NS_887 0 -1.9579947268598604e-05
GC_7_888 b_7 NI_7 NS_888 0 3.1186812617212807e-05
GC_7_889 b_7 NI_7 NS_889 0 -7.1178479610792961e-03
GC_7_890 b_7 NI_7 NS_890 0 4.4750313459225788e-03
GC_7_891 b_7 NI_7 NS_891 0 -7.6633160907172053e-03
GC_7_892 b_7 NI_7 NS_892 0 -5.3302499091944225e-03
GC_7_893 b_7 NI_7 NS_893 0 9.5222517408130019e-03
GC_7_894 b_7 NI_7 NS_894 0 -1.7152207801199302e-03
GC_7_895 b_7 NI_7 NS_895 0 1.2490645341647396e-02
GC_7_896 b_7 NI_7 NS_896 0 -1.3743927858503105e-03
GC_7_897 b_7 NI_7 NS_897 0 -5.0724962539625490e-03
GC_7_898 b_7 NI_7 NS_898 0 -2.7518973835840869e-03
GC_7_899 b_7 NI_7 NS_899 0 -2.2328735438328835e-03
GC_7_900 b_7 NI_7 NS_900 0 6.6013634800430208e-03
GC_7_901 b_7 NI_7 NS_901 0 8.9595183969251330e-03
GC_7_902 b_7 NI_7 NS_902 0 1.2929296960436778e-04
GC_7_903 b_7 NI_7 NS_903 0 1.2486920853853483e-02
GC_7_904 b_7 NI_7 NS_904 0 1.7755896081662643e-03
GC_7_905 b_7 NI_7 NS_905 0 -5.3764649778781162e-03
GC_7_906 b_7 NI_7 NS_906 0 4.1567513025639958e-03
GC_7_907 b_7 NI_7 NS_907 0 -1.8433858254622215e-03
GC_7_908 b_7 NI_7 NS_908 0 -5.6868622793951554e-03
GC_7_909 b_7 NI_7 NS_909 0 2.0787691739809346e-07
GC_7_910 b_7 NI_7 NS_910 0 -2.4509522319828843e-07
GC_7_911 b_7 NI_7 NS_911 0 -1.1507782431194688e-05
GC_7_912 b_7 NI_7 NS_912 0 1.8247330623001379e-05
GC_7_913 b_7 NI_7 NS_913 0 2.8651768627693445e-04
GC_7_914 b_7 NI_7 NS_914 0 -1.4350270506552367e-05
GC_7_915 b_7 NI_7 NS_915 0 -1.2376921342242152e-09
GC_7_916 b_7 NI_7 NS_916 0 -1.9231837777704744e-08
GC_7_917 b_7 NI_7 NS_917 0 2.6656320245855035e-06
GC_7_918 b_7 NI_7 NS_918 0 -3.8233433973871865e-06
GC_7_919 b_7 NI_7 NS_919 0 -1.3224305921867278e-05
GC_7_920 b_7 NI_7 NS_920 0 -5.0206337403547749e-07
GC_7_921 b_7 NI_7 NS_921 0 3.9456084961425105e-05
GC_7_922 b_7 NI_7 NS_922 0 2.7908357503413394e-06
GC_7_923 b_7 NI_7 NS_923 0 -4.1773666457286942e-05
GC_7_924 b_7 NI_7 NS_924 0 -2.3731191064838766e-05
GC_7_925 b_7 NI_7 NS_925 0 1.7633810809398323e-06
GC_7_926 b_7 NI_7 NS_926 0 4.4847668839258310e-05
GC_7_927 b_7 NI_7 NS_927 0 1.4507221166109627e-05
GC_7_928 b_7 NI_7 NS_928 0 -4.8182187556368989e-05
GC_7_929 b_7 NI_7 NS_929 0 1.9346478235648469e-06
GC_7_930 b_7 NI_7 NS_930 0 5.6524857626343941e-06
GC_7_931 b_7 NI_7 NS_931 0 -4.4992649271795452e-05
GC_7_932 b_7 NI_7 NS_932 0 1.5680700842018532e-06
GC_7_933 b_7 NI_7 NS_933 0 1.0311100325369307e-04
GC_7_934 b_7 NI_7 NS_934 0 1.2335725337815940e-04
GC_7_935 b_7 NI_7 NS_935 0 -7.5524315977935973e-05
GC_7_936 b_7 NI_7 NS_936 0 -1.3698768740620404e-04
GC_7_937 b_7 NI_7 NS_937 0 -6.7108091795825249e-05
GC_7_938 b_7 NI_7 NS_938 0 4.9269053949164518e-05
GC_7_939 b_7 NI_7 NS_939 0 1.3517316928522222e-04
GC_7_940 b_7 NI_7 NS_940 0 -2.8539512510134432e-05
GC_7_941 b_7 NI_7 NS_941 0 -8.7330355701334414e-05
GC_7_942 b_7 NI_7 NS_942 0 -1.1763765184073353e-05
GC_7_943 b_7 NI_7 NS_943 0 -9.4644587034506777e-05
GC_7_944 b_7 NI_7 NS_944 0 2.1148789540385133e-04
GC_7_945 b_7 NI_7 NS_945 0 1.6429528258992998e-04
GC_7_946 b_7 NI_7 NS_946 0 -2.1487718422095900e-04
GC_7_947 b_7 NI_7 NS_947 0 -8.1683784350939148e-05
GC_7_948 b_7 NI_7 NS_948 0 1.9188652326562081e-05
GC_7_949 b_7 NI_7 NS_949 0 1.6096945078860142e-04
GC_7_950 b_7 NI_7 NS_950 0 4.2088604141648439e-05
GC_7_951 b_7 NI_7 NS_951 0 -8.8878228100407010e-05
GC_7_952 b_7 NI_7 NS_952 0 -7.1909714164901403e-05
GC_7_953 b_7 NI_7 NS_953 0 -8.4866179909772610e-05
GC_7_954 b_7 NI_7 NS_954 0 6.3595962069746626e-05
GC_7_955 b_7 NI_7 NS_955 0 1.4068739979468782e-04
GC_7_956 b_7 NI_7 NS_956 0 -4.8520533795343081e-05
GC_7_957 b_7 NI_7 NS_957 0 -6.6207336018025197e-05
GC_7_958 b_7 NI_7 NS_958 0 -2.4251182957480047e-05
GC_7_959 b_7 NI_7 NS_959 0 6.1224274343096440e-05
GC_7_960 b_7 NI_7 NS_960 0 1.1375729329027107e-04
GC_7_961 b_7 NI_7 NS_961 0 -2.2917748245630580e-05
GC_7_962 b_7 NI_7 NS_962 0 -1.2153249742245482e-04
GC_7_963 b_7 NI_7 NS_963 0 -4.4313280200757508e-05
GC_7_964 b_7 NI_7 NS_964 0 1.0974879861682030e-05
GC_7_965 b_7 NI_7 NS_965 0 4.7535701760196880e-05
GC_7_966 b_7 NI_7 NS_966 0 -1.0608044885966874e-05
GC_7_967 b_7 NI_7 NS_967 0 -3.2085808555960550e-05
GC_7_968 b_7 NI_7 NS_968 0 -7.6434683690190206e-06
GC_7_969 b_7 NI_7 NS_969 0 2.1333627458187977e-05
GC_7_970 b_7 NI_7 NS_970 0 -4.8747025974480145e-06
GC_7_971 b_7 NI_7 NS_971 0 -3.2213267199621815e-05
GC_7_972 b_7 NI_7 NS_972 0 -2.5250971032116176e-05
GC_7_973 b_7 NI_7 NS_973 0 1.2710451725800827e-05
GC_7_974 b_7 NI_7 NS_974 0 6.1766879660438486e-06
GC_7_975 b_7 NI_7 NS_975 0 -2.0358851588991463e-05
GC_7_976 b_7 NI_7 NS_976 0 -7.7255063667743757e-06
GC_7_977 b_7 NI_7 NS_977 0 1.4086791124182231e-05
GC_7_978 b_7 NI_7 NS_978 0 -1.2504716615467309e-05
GC_7_979 b_7 NI_7 NS_979 0 -4.1281855369796972e-05
GC_7_980 b_7 NI_7 NS_980 0 -1.6953860538917358e-05
GC_7_981 b_7 NI_7 NS_981 0 1.1908060037443579e-05
GC_7_982 b_7 NI_7 NS_982 0 -1.7650834671605370e-06
GC_7_983 b_7 NI_7 NS_983 0 -3.0212165114925223e-05
GC_7_984 b_7 NI_7 NS_984 0 5.5332079997789261e-06
GC_7_985 b_7 NI_7 NS_985 0 1.6333206664474716e-05
GC_7_986 b_7 NI_7 NS_986 0 -2.0848888570423432e-05
GC_7_987 b_7 NI_7 NS_987 0 -4.9845706090843524e-05
GC_7_988 b_7 NI_7 NS_988 0 -1.6671133391349951e-06
GC_7_989 b_7 NI_7 NS_989 0 1.2248920619281750e-05
GC_7_990 b_7 NI_7 NS_990 0 -1.1718134633326208e-05
GC_7_991 b_7 NI_7 NS_991 0 -3.1907777066314714e-05
GC_7_992 b_7 NI_7 NS_992 0 2.5076448405754126e-05
GC_7_993 b_7 NI_7 NS_993 0 1.0836001333014514e-05
GC_7_994 b_7 NI_7 NS_994 0 -3.6497129460932100e-05
GC_7_995 b_7 NI_7 NS_995 0 -3.3854597455078118e-05
GC_7_996 b_7 NI_7 NS_996 0 1.8659942635077120e-05
GC_7_997 b_7 NI_7 NS_997 0 -5.9885030775016148e-05
GC_7_998 b_7 NI_7 NS_998 0 1.2846809847204567e-04
GC_7_999 b_7 NI_7 NS_999 0 -1.4510117246787896e-05
GC_7_1000 b_7 NI_7 NS_1000 0 -3.3372794892863403e-05
GC_7_1001 b_7 NI_7 NS_1001 0 -3.8792938528746117e-07
GC_7_1002 b_7 NI_7 NS_1002 0 3.6143461469026370e-07
GC_7_1003 b_7 NI_7 NS_1003 0 -1.9684608468607042e-05
GC_7_1004 b_7 NI_7 NS_1004 0 3.1288239547052376e-05
GC_7_1005 b_7 NI_7 NS_1005 0 -1.4242871887690362e-05
GC_7_1006 b_7 NI_7 NS_1006 0 -3.4197769282285746e-05
GC_7_1007 b_7 NI_7 NS_1007 0 -5.2907352216312604e-06
GC_7_1008 b_7 NI_7 NS_1008 0 5.5319735465968331e-06
GC_7_1009 b_7 NI_7 NS_1009 0 -1.9742372090908153e-05
GC_7_1010 b_7 NI_7 NS_1010 0 -6.5467166006922959e-05
GC_7_1011 b_7 NI_7 NS_1011 0 -9.2829820999748463e-06
GC_7_1012 b_7 NI_7 NS_1012 0 -2.0586456833330478e-05
GC_7_1013 b_7 NI_7 NS_1013 0 1.4777323865722815e-05
GC_7_1014 b_7 NI_7 NS_1014 0 2.2998758109211345e-05
GC_7_1015 b_7 NI_7 NS_1015 0 -6.8231215757169168e-06
GC_7_1016 b_7 NI_7 NS_1016 0 2.7592360285689858e-05
GC_7_1017 b_7 NI_7 NS_1017 0 -1.1136047147634668e-05
GC_7_1018 b_7 NI_7 NS_1018 0 -2.1577810751687306e-05
GC_7_1019 b_7 NI_7 NS_1019 0 -1.1024479616843738e-05
GC_7_1020 b_7 NI_7 NS_1020 0 2.3799265235835828e-05
GC_7_1021 b_7 NI_7 NS_1021 0 5.1499622026257970e-06
GC_7_1022 b_7 NI_7 NS_1022 0 -1.5352080954316792e-05
GC_7_1023 b_7 NI_7 NS_1023 0 -4.7263523119410147e-10
GC_7_1024 b_7 NI_7 NS_1024 0 -9.1862440894306344e-10
GC_7_1025 b_7 NI_7 NS_1025 0 -5.5412149217665357e-08
GC_7_1026 b_7 NI_7 NS_1026 0 7.6391268743933525e-09
GC_7_1027 b_7 NI_7 NS_1027 0 -2.0271400468649996e-04
GC_7_1028 b_7 NI_7 NS_1028 0 -3.3244166343622547e-06
GC_7_1029 b_7 NI_7 NS_1029 0 1.2949661017590402e-09
GC_7_1030 b_7 NI_7 NS_1030 0 9.6758912422453085e-09
GC_7_1031 b_7 NI_7 NS_1031 0 -4.1591752799954472e-06
GC_7_1032 b_7 NI_7 NS_1032 0 6.1862098487574832e-06
GC_7_1033 b_7 NI_7 NS_1033 0 3.8149385206515077e-06
GC_7_1034 b_7 NI_7 NS_1034 0 -8.1670916783080741e-06
GC_7_1035 b_7 NI_7 NS_1035 0 2.1690370378389837e-05
GC_7_1036 b_7 NI_7 NS_1036 0 -8.8399972516782730e-06
GC_7_1037 b_7 NI_7 NS_1037 0 -2.1479600659427076e-05
GC_7_1038 b_7 NI_7 NS_1038 0 -1.1874148691720609e-06
GC_7_1039 b_7 NI_7 NS_1039 0 -2.9640120231626712e-05
GC_7_1040 b_7 NI_7 NS_1040 0 -2.8295816205185402e-05
GC_7_1041 b_7 NI_7 NS_1041 0 -5.5412991136573986e-06
GC_7_1042 b_7 NI_7 NS_1042 0 1.6552014227758522e-05
GC_7_1043 b_7 NI_7 NS_1043 0 -2.4251840788861427e-06
GC_7_1044 b_7 NI_7 NS_1044 0 -7.1420356075309639e-06
GC_7_1045 b_7 NI_7 NS_1045 0 -2.2563451770829412e-05
GC_7_1046 b_7 NI_7 NS_1046 0 6.0026123011673165e-06
GC_7_1047 b_7 NI_7 NS_1047 0 -1.8565790734937138e-04
GC_7_1048 b_7 NI_7 NS_1048 0 -4.4043350375182038e-05
GC_7_1049 b_7 NI_7 NS_1049 0 6.2654400956825562e-05
GC_7_1050 b_7 NI_7 NS_1050 0 1.3744255844417037e-04
GC_7_1051 b_7 NI_7 NS_1051 0 -3.7291590688739382e-05
GC_7_1052 b_7 NI_7 NS_1052 0 5.6617736698313637e-05
GC_7_1053 b_7 NI_7 NS_1053 0 9.5234341768614714e-05
GC_7_1054 b_7 NI_7 NS_1054 0 2.4609658732078349e-04
GC_7_1055 b_7 NI_7 NS_1055 0 7.3806894495698300e-05
GC_7_1056 b_7 NI_7 NS_1056 0 4.9082517264315611e-07
GC_7_1057 b_7 NI_7 NS_1057 0 -1.5390445972806238e-05
GC_7_1058 b_7 NI_7 NS_1058 0 2.6127685585974935e-04
GC_7_1059 b_7 NI_7 NS_1059 0 3.6437419499255378e-04
GC_7_1060 b_7 NI_7 NS_1060 0 -2.4319842581219277e-04
GC_7_1061 b_7 NI_7 NS_1061 0 6.5655663044598454e-05
GC_7_1062 b_7 NI_7 NS_1062 0 -2.8529428192746581e-05
GC_7_1063 b_7 NI_7 NS_1063 0 2.0802593133119893e-04
GC_7_1064 b_7 NI_7 NS_1064 0 -2.4142800835814839e-04
GC_7_1065 b_7 NI_7 NS_1065 0 -7.1299257465787320e-05
GC_7_1066 b_7 NI_7 NS_1066 0 -7.1473438568464272e-05
GC_7_1067 b_7 NI_7 NS_1067 0 6.4494182829781936e-05
GC_7_1068 b_7 NI_7 NS_1068 0 -7.5537526523138679e-05
GC_7_1069 b_7 NI_7 NS_1069 0 -1.7050086557019500e-04
GC_7_1070 b_7 NI_7 NS_1070 0 -1.8310153492387824e-04
GC_7_1071 b_7 NI_7 NS_1071 0 -4.8839023741566287e-05
GC_7_1072 b_7 NI_7 NS_1072 0 -1.9100995783330034e-05
GC_7_1073 b_7 NI_7 NS_1073 0 -1.4492616761180904e-04
GC_7_1074 b_7 NI_7 NS_1074 0 -9.5351253982682815e-05
GC_7_1075 b_7 NI_7 NS_1075 0 -2.7319738492277388e-05
GC_7_1076 b_7 NI_7 NS_1076 0 1.0361197434905567e-04
GC_7_1077 b_7 NI_7 NS_1077 0 -2.7244445889228455e-05
GC_7_1078 b_7 NI_7 NS_1078 0 1.3907006573924486e-05
GC_7_1079 b_7 NI_7 NS_1079 0 2.1287331775480765e-06
GC_7_1080 b_7 NI_7 NS_1080 0 5.0767895602600528e-05
GC_7_1081 b_7 NI_7 NS_1081 0 1.6812848099259353e-05
GC_7_1082 b_7 NI_7 NS_1082 0 -5.9689902238830489e-07
GC_7_1083 b_7 NI_7 NS_1083 0 1.8078605032340050e-06
GC_7_1084 b_7 NI_7 NS_1084 0 -1.5453788139724473e-05
GC_7_1085 b_7 NI_7 NS_1085 0 -1.5113187630869825e-05
GC_7_1086 b_7 NI_7 NS_1086 0 -1.3588621459978819e-05
GC_7_1087 b_7 NI_7 NS_1087 0 -1.3111062826395325e-05
GC_7_1088 b_7 NI_7 NS_1088 0 1.2341203596314654e-05
GC_7_1089 b_7 NI_7 NS_1089 0 7.7832678221314426e-06
GC_7_1090 b_7 NI_7 NS_1090 0 1.2547283828992772e-06
GC_7_1091 b_7 NI_7 NS_1091 0 -5.1390800509752550e-06
GC_7_1092 b_7 NI_7 NS_1092 0 -1.2684885561812388e-05
GC_7_1093 b_7 NI_7 NS_1093 0 -2.0804835952559483e-05
GC_7_1094 b_7 NI_7 NS_1094 0 -5.8777160580149273e-06
GC_7_1095 b_7 NI_7 NS_1095 0 1.0778177822923471e-06
GC_7_1096 b_7 NI_7 NS_1096 0 2.1822125041559117e-05
GC_7_1097 b_7 NI_7 NS_1097 0 1.2864918044895715e-05
GC_7_1098 b_7 NI_7 NS_1098 0 -6.8616156202713478e-06
GC_7_1099 b_7 NI_7 NS_1099 0 -1.7284500552021679e-05
GC_7_1100 b_7 NI_7 NS_1100 0 -1.5979338378213542e-05
GC_7_1101 b_7 NI_7 NS_1101 0 -2.7118176299836404e-05
GC_7_1102 b_7 NI_7 NS_1102 0 8.8177815691255219e-06
GC_7_1103 b_7 NI_7 NS_1103 0 2.7091326238205692e-05
GC_7_1104 b_7 NI_7 NS_1104 0 2.2446901293536093e-05
GC_7_1105 b_7 NI_7 NS_1105 0 1.0942484757867851e-05
GC_7_1106 b_7 NI_7 NS_1106 0 -2.1302974384350224e-05
GC_7_1107 b_7 NI_7 NS_1107 0 -3.0617343212276214e-05
GC_7_1108 b_7 NI_7 NS_1108 0 3.9057784790851178e-06
GC_7_1109 b_7 NI_7 NS_1109 0 -9.8014536925520751e-06
GC_7_1110 b_7 NI_7 NS_1110 0 3.9251521716220126e-05
GC_7_1111 b_7 NI_7 NS_1111 0 1.9727816453762273e-05
GC_7_1112 b_7 NI_7 NS_1112 0 -6.8538574255965398e-05
GC_7_1113 b_7 NI_7 NS_1113 0 4.3399507366581652e-05
GC_7_1114 b_7 NI_7 NS_1114 0 -1.6869783563000871e-05
GC_7_1115 b_7 NI_7 NS_1115 0 2.0639886136628772e-07
GC_7_1116 b_7 NI_7 NS_1116 0 -2.4347742686430897e-07
GC_7_1117 b_7 NI_7 NS_1117 0 -3.6328458216830294e-06
GC_7_1118 b_7 NI_7 NS_1118 0 -2.0833672030216105e-05
GC_7_1119 b_7 NI_7 NS_1119 0 -1.0494375586474375e-05
GC_7_1120 b_7 NI_7 NS_1120 0 1.6698424302608068e-05
GC_7_1121 b_7 NI_7 NS_1121 0 9.1959654082619564e-06
GC_7_1122 b_7 NI_7 NS_1122 0 3.1866768303067152e-05
GC_7_1123 b_7 NI_7 NS_1123 0 1.4280791751561903e-05
GC_7_1124 b_7 NI_7 NS_1124 0 -3.0127237457371969e-06
GC_7_1125 b_7 NI_7 NS_1125 0 -3.9054310694853980e-06
GC_7_1126 b_7 NI_7 NS_1126 0 1.2499910887324246e-05
GC_7_1127 b_7 NI_7 NS_1127 0 -1.8574401774817001e-05
GC_7_1128 b_7 NI_7 NS_1128 0 -3.6262133130471213e-06
GC_7_1129 b_7 NI_7 NS_1129 0 1.3215556396738112e-05
GC_7_1130 b_7 NI_7 NS_1130 0 1.3176894838669152e-05
GC_7_1131 b_7 NI_7 NS_1131 0 7.6361533714823685e-06
GC_7_1132 b_7 NI_7 NS_1132 0 -2.3019339363699896e-05
GC_7_1133 b_7 NI_7 NS_1133 0 -3.8459159410329157e-06
GC_7_1134 b_7 NI_7 NS_1134 0 -1.1723218514196313e-05
GC_7_1135 b_7 NI_7 NS_1135 0 -8.7362090596981494e-06
GC_7_1136 b_7 NI_7 NS_1136 0 -2.6280716201934965e-06
GC_7_1137 b_7 NI_7 NS_1137 0 5.5146535151355474e-10
GC_7_1138 b_7 NI_7 NS_1138 0 2.9343934213448563e-10
GC_7_1139 b_7 NI_7 NS_1139 0 4.2107563575441155e-08
GC_7_1140 b_7 NI_7 NS_1140 0 3.6940437896542488e-08
GC_7_1141 b_7 NI_7 NS_1141 0 -1.1163639693550968e-04
GC_7_1142 b_7 NI_7 NS_1142 0 -2.1529158609325423e-06
GC_7_1143 b_7 NI_7 NS_1143 0 -2.4619850212271531e-10
GC_7_1144 b_7 NI_7 NS_1144 0 2.5690930656971654e-09
GC_7_1145 b_7 NI_7 NS_1145 0 1.8039278164080402e-06
GC_7_1146 b_7 NI_7 NS_1146 0 -1.6072975557664492e-06
GC_7_1147 b_7 NI_7 NS_1147 0 2.5854821190860310e-07
GC_7_1148 b_7 NI_7 NS_1148 0 -6.4503864097479795e-06
GC_7_1149 b_7 NI_7 NS_1149 0 -7.5446340382405190e-06
GC_7_1150 b_7 NI_7 NS_1150 0 -3.1551875981928717e-07
GC_7_1151 b_7 NI_7 NS_1151 0 -1.4480434191738478e-06
GC_7_1152 b_7 NI_7 NS_1152 0 -4.6837951379449334e-06
GC_7_1153 b_7 NI_7 NS_1153 0 -1.5899387502200874e-05
GC_7_1154 b_7 NI_7 NS_1154 0 -1.9736058720862053e-06
GC_7_1155 b_7 NI_7 NS_1155 0 -7.0460530696893739e-06
GC_7_1156 b_7 NI_7 NS_1156 0 1.8943205321235808e-05
GC_7_1157 b_7 NI_7 NS_1157 0 4.8825937107646242e-06
GC_7_1158 b_7 NI_7 NS_1158 0 -2.8766001946831069e-06
GC_7_1159 b_7 NI_7 NS_1159 0 -1.3982129493177542e-07
GC_7_1160 b_7 NI_7 NS_1160 0 -2.4404301253185935e-06
GC_7_1161 b_7 NI_7 NS_1161 0 -2.6317281638368767e-05
GC_7_1162 b_7 NI_7 NS_1162 0 2.8135823180155724e-05
GC_7_1163 b_7 NI_7 NS_1163 0 2.8104646648151496e-05
GC_7_1164 b_7 NI_7 NS_1164 0 -7.9688315628009592e-06
GC_7_1165 b_7 NI_7 NS_1165 0 -8.0936115926343451e-06
GC_7_1166 b_7 NI_7 NS_1166 0 -4.2239601673955717e-06
GC_7_1167 b_7 NI_7 NS_1167 0 1.2266612638138046e-05
GC_7_1168 b_7 NI_7 NS_1168 0 2.7177892606694895e-05
GC_7_1169 b_7 NI_7 NS_1169 0 1.4632391604845172e-06
GC_7_1170 b_7 NI_7 NS_1170 0 -8.8115826059505750e-06
GC_7_1171 b_7 NI_7 NS_1171 0 -2.8379259351131009e-05
GC_7_1172 b_7 NI_7 NS_1172 0 4.7636960372265209e-06
GC_7_1173 b_7 NI_7 NS_1173 0 4.1223375313077263e-05
GC_7_1174 b_7 NI_7 NS_1174 0 1.0997306867440748e-05
GC_7_1175 b_7 NI_7 NS_1175 0 -2.9904643389602631e-06
GC_7_1176 b_7 NI_7 NS_1176 0 -4.3573148071414628e-06
GC_7_1177 b_7 NI_7 NS_1177 0 1.2935785684589371e-05
GC_7_1178 b_7 NI_7 NS_1178 0 1.9156001207509449e-05
GC_7_1179 b_7 NI_7 NS_1179 0 3.7957745673785355e-06
GC_7_1180 b_7 NI_7 NS_1180 0 -1.0819255556157442e-05
GC_7_1181 b_7 NI_7 NS_1181 0 -6.4497759543350755e-06
GC_7_1182 b_7 NI_7 NS_1182 0 9.6990788131141518e-07
GC_7_1183 b_7 NI_7 NS_1183 0 1.8939860646024079e-05
GC_7_1184 b_7 NI_7 NS_1184 0 5.5256304868785442e-06
GC_7_1185 b_7 NI_7 NS_1185 0 -1.0369489323891904e-07
GC_7_1186 b_7 NI_7 NS_1186 0 -4.1120694707765907e-06
GC_7_1187 b_7 NI_7 NS_1187 0 4.9329507778730780e-06
GC_7_1188 b_7 NI_7 NS_1188 0 1.4409307396633269e-05
GC_7_1189 b_7 NI_7 NS_1189 0 7.8206607248193119e-06
GC_7_1190 b_7 NI_7 NS_1190 0 -1.1148679788740902e-05
GC_7_1191 b_7 NI_7 NS_1191 0 -1.4169787281153302e-06
GC_7_1192 b_7 NI_7 NS_1192 0 9.8983545243840466e-07
GC_7_1193 b_7 NI_7 NS_1193 0 1.0881123907507149e-05
GC_7_1194 b_7 NI_7 NS_1194 0 4.1883216325746677e-06
GC_7_1195 b_7 NI_7 NS_1195 0 1.6989713673346718e-06
GC_7_1196 b_7 NI_7 NS_1196 0 -5.8201958867956544e-07
GC_7_1197 b_7 NI_7 NS_1197 0 5.6739379829910310e-06
GC_7_1198 b_7 NI_7 NS_1198 0 1.7280443514878534e-06
GC_7_1199 b_7 NI_7 NS_1199 0 3.3535644690499060e-06
GC_7_1200 b_7 NI_7 NS_1200 0 2.0815595639321636e-06
GC_7_1201 b_7 NI_7 NS_1201 0 1.0938037475103444e-05
GC_7_1202 b_7 NI_7 NS_1202 0 3.8462781645269213e-06
GC_7_1203 b_7 NI_7 NS_1203 0 4.8353425294567808e-06
GC_7_1204 b_7 NI_7 NS_1204 0 -4.4521362005255232e-08
GC_7_1205 b_7 NI_7 NS_1205 0 9.9616049377974596e-06
GC_7_1206 b_7 NI_7 NS_1206 0 -1.0482433375817011e-06
GC_7_1207 b_7 NI_7 NS_1207 0 8.1946746009049546e-06
GC_7_1208 b_7 NI_7 NS_1208 0 2.9799204274174188e-06
GC_7_1209 b_7 NI_7 NS_1209 0 1.9009426411275722e-05
GC_7_1210 b_7 NI_7 NS_1210 0 -5.5028971455175079e-06
GC_7_1211 b_7 NI_7 NS_1211 0 7.1831605069952093e-06
GC_7_1212 b_7 NI_7 NS_1212 0 -3.9855819824283925e-06
GC_7_1213 b_7 NI_7 NS_1213 0 1.3697382057704088e-05
GC_7_1214 b_7 NI_7 NS_1214 0 -1.1862009083210408e-05
GC_7_1215 b_7 NI_7 NS_1215 0 1.2345387697564614e-05
GC_7_1216 b_7 NI_7 NS_1216 0 -3.9388171235161860e-06
GC_7_1217 b_7 NI_7 NS_1217 0 9.1353069521369579e-06
GC_7_1218 b_7 NI_7 NS_1218 0 -2.6714433579846839e-05
GC_7_1219 b_7 NI_7 NS_1219 0 2.3416330847424886e-06
GC_7_1220 b_7 NI_7 NS_1220 0 -1.2350035947062383e-05
GC_7_1221 b_7 NI_7 NS_1221 0 -8.3090397673216526e-06
GC_7_1222 b_7 NI_7 NS_1222 0 -1.8612842055953615e-05
GC_7_1223 b_7 NI_7 NS_1223 0 -4.9202386355055419e-06
GC_7_1224 b_7 NI_7 NS_1224 0 -1.2088815843512124e-05
GC_7_1225 b_7 NI_7 NS_1225 0 5.4869187739346475e-05
GC_7_1226 b_7 NI_7 NS_1226 0 -8.7931493178793033e-05
GC_7_1227 b_7 NI_7 NS_1227 0 -1.0053081732229120e-05
GC_7_1228 b_7 NI_7 NS_1228 0 1.3554292903216014e-06
GC_7_1229 b_7 NI_7 NS_1229 0 3.9049610945211509e-07
GC_7_1230 b_7 NI_7 NS_1230 0 -1.2503196806407838e-07
GC_7_1231 b_7 NI_7 NS_1231 0 -2.7269127430624630e-06
GC_7_1232 b_7 NI_7 NS_1232 0 -1.9374888782496428e-06
GC_7_1233 b_7 NI_7 NS_1233 0 -4.4052555975202703e-06
GC_7_1234 b_7 NI_7 NS_1234 0 5.8881531256116932e-07
GC_7_1235 b_7 NI_7 NS_1235 0 -1.7470998453955830e-05
GC_7_1236 b_7 NI_7 NS_1236 0 9.5706307876778435e-06
GC_7_1237 b_7 NI_7 NS_1237 0 -9.2073300580411771e-06
GC_7_1238 b_7 NI_7 NS_1238 0 3.7347453100437351e-05
GC_7_1239 b_7 NI_7 NS_1239 0 -7.2389889907515128e-06
GC_7_1240 b_7 NI_7 NS_1240 0 3.3305386412017822e-07
GC_7_1241 b_7 NI_7 NS_1241 0 -1.3385051466923471e-05
GC_7_1242 b_7 NI_7 NS_1242 0 1.8624029378737059e-06
GC_7_1243 b_7 NI_7 NS_1243 0 -4.6430382324341595e-06
GC_7_1244 b_7 NI_7 NS_1244 0 -3.3916905392890218e-06
GC_7_1245 b_7 NI_7 NS_1245 0 -6.3994044318039111e-06
GC_7_1246 b_7 NI_7 NS_1246 0 1.0401449190034506e-06
GC_7_1247 b_7 NI_7 NS_1247 0 -3.0542884809419204e-06
GC_7_1248 b_7 NI_7 NS_1248 0 8.8891070214620291e-07
GC_7_1249 b_7 NI_7 NS_1249 0 -1.7965416932669041e-06
GC_7_1250 b_7 NI_7 NS_1250 0 -9.3478377772190305e-07
GC_7_1251 b_7 NI_7 NS_1251 0 -2.6064286911257407e-10
GC_7_1252 b_7 NI_7 NS_1252 0 4.2284174144260723e-10
GC_7_1253 b_7 NI_7 NS_1253 0 2.3336442188220084e-09
GC_7_1254 b_7 NI_7 NS_1254 0 -2.6682895717797015e-08
GC_7_1255 b_7 NI_7 NS_1255 0 -3.7757921460742810e-05
GC_7_1256 b_7 NI_7 NS_1256 0 2.2260818083806183e-06
GC_7_1257 b_7 NI_7 NS_1257 0 6.0497545363514610e-11
GC_7_1258 b_7 NI_7 NS_1258 0 3.0748155239702773e-09
GC_7_1259 b_7 NI_7 NS_1259 0 -1.9314697076780545e-06
GC_7_1260 b_7 NI_7 NS_1260 0 -1.7211198478621709e-06
GC_7_1261 b_7 NI_7 NS_1261 0 -5.6037063437306761e-06
GC_7_1262 b_7 NI_7 NS_1262 0 2.9249833771394349e-06
GC_7_1263 b_7 NI_7 NS_1263 0 -1.6662618290814859e-05
GC_7_1264 b_7 NI_7 NS_1264 0 1.9136410413034691e-05
GC_7_1265 b_7 NI_7 NS_1265 0 1.5401447135650260e-05
GC_7_1266 b_7 NI_7 NS_1266 0 1.0211362674985730e-05
GC_7_1267 b_7 NI_7 NS_1267 0 1.7356967279616526e-05
GC_7_1268 b_7 NI_7 NS_1268 0 2.3278421578562231e-05
GC_7_1269 b_7 NI_7 NS_1269 0 3.0898154232792304e-05
GC_7_1270 b_7 NI_7 NS_1270 0 5.3461790024660126e-06
GC_7_1271 b_7 NI_7 NS_1271 0 -3.3856270489429286e-06
GC_7_1272 b_7 NI_7 NS_1272 0 -2.1458326046312767e-06
GC_7_1273 b_7 NI_7 NS_1273 0 1.7190876278937259e-05
GC_7_1274 b_7 NI_7 NS_1274 0 -2.2223174124944080e-06
GC_7_1275 b_7 NI_7 NS_1275 0 1.2979334008016638e-04
GC_7_1276 b_7 NI_7 NS_1276 0 3.5245891749625550e-05
GC_7_1277 b_7 NI_7 NS_1277 0 -2.8532252445843134e-05
GC_7_1278 b_7 NI_7 NS_1278 0 -9.9831816067458658e-05
GC_7_1279 b_7 NI_7 NS_1279 0 2.5236659748344874e-05
GC_7_1280 b_7 NI_7 NS_1280 0 -3.1266673944117678e-05
GC_7_1281 b_7 NI_7 NS_1281 0 -4.0929319729151487e-05
GC_7_1282 b_7 NI_7 NS_1282 0 -1.6750257995001988e-04
GC_7_1283 b_7 NI_7 NS_1283 0 -4.1821228562941846e-05
GC_7_1284 b_7 NI_7 NS_1284 0 -5.3848006591397321e-06
GC_7_1285 b_7 NI_7 NS_1285 0 2.2549793276932343e-05
GC_7_1286 b_7 NI_7 NS_1286 0 -1.5151993535901580e-04
GC_7_1287 b_7 NI_7 NS_1287 0 -2.3148577820084846e-04
GC_7_1288 b_7 NI_7 NS_1288 0 1.1299683140589735e-04
GC_7_1289 b_7 NI_7 NS_1289 0 -3.7411182816105100e-05
GC_7_1290 b_7 NI_7 NS_1290 0 1.3952070823890971e-05
GC_7_1291 b_7 NI_7 NS_1291 0 -1.3781868033183495e-04
GC_7_1292 b_7 NI_7 NS_1292 0 1.2973370306020021e-04
GC_7_1293 b_7 NI_7 NS_1293 0 3.6131599498458664e-05
GC_7_1294 b_7 NI_7 NS_1294 0 4.1461236747296763e-05
GC_7_1295 b_7 NI_7 NS_1295 0 -3.8173652273211418e-05
GC_7_1296 b_7 NI_7 NS_1296 0 4.2970717763319250e-05
GC_7_1297 b_7 NI_7 NS_1297 0 8.7353505230339500e-05
GC_7_1298 b_7 NI_7 NS_1298 0 1.1821521585201738e-04
GC_7_1299 b_7 NI_7 NS_1299 0 2.7244713867421040e-05
GC_7_1300 b_7 NI_7 NS_1300 0 1.0262297459645668e-05
GC_7_1301 b_7 NI_7 NS_1301 0 8.7157827232716469e-05
GC_7_1302 b_7 NI_7 NS_1302 0 6.5380834701498107e-05
GC_7_1303 b_7 NI_7 NS_1303 0 2.0401052229024294e-05
GC_7_1304 b_7 NI_7 NS_1304 0 -5.7168348439270240e-05
GC_7_1305 b_7 NI_7 NS_1305 0 1.7001785073818202e-05
GC_7_1306 b_7 NI_7 NS_1306 0 -8.8439364054528390e-06
GC_7_1307 b_7 NI_7 NS_1307 0 8.4707962066571547e-06
GC_7_1308 b_7 NI_7 NS_1308 0 -3.3126354410214759e-05
GC_7_1309 b_7 NI_7 NS_1309 0 -8.8428232886016357e-06
GC_7_1310 b_7 NI_7 NS_1310 0 4.1504040673076701e-07
GC_7_1311 b_7 NI_7 NS_1311 0 -2.4023068832751112e-06
GC_7_1312 b_7 NI_7 NS_1312 0 8.4362071701720902e-06
GC_7_1313 b_7 NI_7 NS_1313 0 1.0207724208982013e-05
GC_7_1314 b_7 NI_7 NS_1314 0 6.0581943458280696e-06
GC_7_1315 b_7 NI_7 NS_1315 0 1.2154855319677452e-05
GC_7_1316 b_7 NI_7 NS_1316 0 -7.9359486673449747e-06
GC_7_1317 b_7 NI_7 NS_1317 0 -3.4649639534594267e-06
GC_7_1318 b_7 NI_7 NS_1318 0 -5.2259517237718180e-07
GC_7_1319 b_7 NI_7 NS_1319 0 2.5131877691080356e-06
GC_7_1320 b_7 NI_7 NS_1320 0 7.3270592462035804e-06
GC_7_1321 b_7 NI_7 NS_1321 0 1.3691620767097522e-05
GC_7_1322 b_7 NI_7 NS_1322 0 2.6181488638458732e-06
GC_7_1323 b_7 NI_7 NS_1323 0 4.5508817033720822e-06
GC_7_1324 b_7 NI_7 NS_1324 0 -1.4312593646279994e-05
GC_7_1325 b_7 NI_7 NS_1325 0 -5.8920273870422509e-06
GC_7_1326 b_7 NI_7 NS_1326 0 4.1741015812914718e-06
GC_7_1327 b_7 NI_7 NS_1327 0 1.0370342285339246e-05
GC_7_1328 b_7 NI_7 NS_1328 0 9.8155148068158105e-06
GC_7_1329 b_7 NI_7 NS_1329 0 1.7399290098632861e-05
GC_7_1330 b_7 NI_7 NS_1330 0 -4.2746509593381250e-06
GC_7_1331 b_7 NI_7 NS_1331 0 -9.2261092185140607e-06
GC_7_1332 b_7 NI_7 NS_1332 0 -1.5489846052182506e-05
GC_7_1333 b_7 NI_7 NS_1333 0 -4.0027577145914625e-06
GC_7_1334 b_7 NI_7 NS_1334 0 1.3420113206249407e-05
GC_7_1335 b_7 NI_7 NS_1335 0 2.1008720405523626e-05
GC_7_1336 b_7 NI_7 NS_1336 0 -7.6338685055023717e-07
GC_7_1337 b_7 NI_7 NS_1337 0 9.1217831177996009e-06
GC_7_1338 b_7 NI_7 NS_1338 0 -1.7455390506289775e-05
GC_7_1339 b_7 NI_7 NS_1339 0 1.4586364471653288e-06
GC_7_1340 b_7 NI_7 NS_1340 0 -1.4427293917210993e-05
GC_7_1341 b_7 NI_7 NS_1341 0 -1.3809195165323541e-05
GC_7_1342 b_7 NI_7 NS_1342 0 3.9887245742760243e-06
GC_7_1343 b_7 NI_7 NS_1343 0 9.7963032623357995e-09
GC_7_1344 b_7 NI_7 NS_1344 0 -4.8131391559212176e-08
GC_7_1345 b_7 NI_7 NS_1345 0 8.6298054466204885e-06
GC_7_1346 b_7 NI_7 NS_1346 0 1.1373549836496001e-05
GC_7_1347 b_7 NI_7 NS_1347 0 1.0873482556395874e-05
GC_7_1348 b_7 NI_7 NS_1348 0 -1.1464245838685777e-05
GC_7_1349 b_7 NI_7 NS_1349 0 -3.5306899584765455e-06
GC_7_1350 b_7 NI_7 NS_1350 0 -1.0164960324094669e-05
GC_7_1351 b_7 NI_7 NS_1351 0 -2.0124957282058730e-06
GC_7_1352 b_7 NI_7 NS_1352 0 1.2870399101246870e-05
GC_7_1353 b_7 NI_7 NS_1353 0 9.7605855869441400e-07
GC_7_1354 b_7 NI_7 NS_1354 0 -7.2620161752454795e-06
GC_7_1355 b_7 NI_7 NS_1355 0 7.4715758891157469e-06
GC_7_1356 b_7 NI_7 NS_1356 0 1.7440661053029410e-06
GC_7_1357 b_7 NI_7 NS_1357 0 -6.1165749899623893e-06
GC_7_1358 b_7 NI_7 NS_1358 0 -8.8986352361987920e-06
GC_7_1359 b_7 NI_7 NS_1359 0 -4.1366734644223145e-06
GC_7_1360 b_7 NI_7 NS_1360 0 9.6569030664131112e-06
GC_7_1361 b_7 NI_7 NS_1361 0 3.3152442455471658e-06
GC_7_1362 b_7 NI_7 NS_1362 0 6.0578135977629411e-06
GC_7_1363 b_7 NI_7 NS_1363 0 5.7049729867959353e-06
GC_7_1364 b_7 NI_7 NS_1364 0 5.2025366586525471e-07
GC_7_1365 b_7 NI_7 NS_1365 0 5.9120086526750252e-11
GC_7_1366 b_7 NI_7 NS_1366 0 1.4784861258780921e-10
GC_7_1367 b_7 NI_7 NS_1367 0 5.9030635419650698e-09
GC_7_1368 b_7 NI_7 NS_1368 0 -8.4601890096564254e-09
GD_7_1 b_7 NI_7 NA_1 0 -3.6529881690054974e-06
GD_7_2 b_7 NI_7 NA_2 0 1.0039623194473853e-05
GD_7_3 b_7 NI_7 NA_3 0 3.6701583809694909e-06
GD_7_4 b_7 NI_7 NA_4 0 1.1832478313857063e-06
GD_7_5 b_7 NI_7 NA_5 0 1.2979344923422039e-02
GD_7_6 b_7 NI_7 NA_6 0 5.8608994903672012e-04
GD_7_7 b_7 NI_7 NA_7 0 -8.8807956671789218e-03
GD_7_8 b_7 NI_7 NA_8 0 -4.2218338451908890e-03
GD_7_9 b_7 NI_7 NA_9 0 1.0377477818751231e-04
GD_7_10 b_7 NI_7 NA_10 0 2.6586126149279830e-05
GD_7_11 b_7 NI_7 NA_11 0 3.8645531634321120e-06
GD_7_12 b_7 NI_7 NA_12 0 2.4546229136042892e-06
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 -6.2021606735053564e-05
GC_8_2 b_8 NI_8 NS_2 0 3.1006125883025785e-07
GC_8_3 b_8 NI_8 NS_3 0 1.6341724892600710e-11
GC_8_4 b_8 NI_8 NS_4 0 -8.7701452471505683e-11
GC_8_5 b_8 NI_8 NS_5 0 -1.1181523833905403e-06
GC_8_6 b_8 NI_8 NS_6 0 -1.7690613015523843e-06
GC_8_7 b_8 NI_8 NS_7 0 -1.9757191082043876e-06
GC_8_8 b_8 NI_8 NS_8 0 1.9724312632021317e-06
GC_8_9 b_8 NI_8 NS_9 0 -9.5765574579279052e-06
GC_8_10 b_8 NI_8 NS_10 0 6.8033994375168141e-07
GC_8_11 b_8 NI_8 NS_11 0 -2.2987516139215162e-07
GC_8_12 b_8 NI_8 NS_12 0 3.5063276175490505e-06
GC_8_13 b_8 NI_8 NS_13 0 -2.0994403960259778e-06
GC_8_14 b_8 NI_8 NS_14 0 1.1705850578815898e-05
GC_8_15 b_8 NI_8 NS_15 0 6.8703437366734034e-06
GC_8_16 b_8 NI_8 NS_16 0 1.2241237468902691e-05
GC_8_17 b_8 NI_8 NS_17 0 -2.0277601719459714e-06
GC_8_18 b_8 NI_8 NS_18 0 -2.2588466572051667e-06
GC_8_19 b_8 NI_8 NS_19 0 1.6453766908037431e-06
GC_8_20 b_8 NI_8 NS_20 0 1.0187558204593194e-06
GC_8_21 b_8 NI_8 NS_21 0 7.3910964400549810e-06
GC_8_22 b_8 NI_8 NS_22 0 3.8498697766008035e-05
GC_8_23 b_8 NI_8 NS_23 0 2.2957030175483857e-05
GC_8_24 b_8 NI_8 NS_24 0 -1.2018259277374009e-05
GC_8_25 b_8 NI_8 NS_25 0 8.4099922233912676e-06
GC_8_26 b_8 NI_8 NS_26 0 1.7737163421784163e-06
GC_8_27 b_8 NI_8 NS_27 0 4.7831229696265145e-05
GC_8_28 b_8 NI_8 NS_28 0 -2.5191938241218791e-05
GC_8_29 b_8 NI_8 NS_29 0 -9.1802548293805272e-07
GC_8_30 b_8 NI_8 NS_30 0 -8.0507006407735592e-06
GC_8_31 b_8 NI_8 NS_31 0 3.4285625162713150e-05
GC_8_32 b_8 NI_8 NS_32 0 -7.7290006507951425e-06
GC_8_33 b_8 NI_8 NS_33 0 -3.8666315683691805e-05
GC_8_34 b_8 NI_8 NS_34 0 -5.1897453529178027e-05
GC_8_35 b_8 NI_8 NS_35 0 -4.5703061466470291e-06
GC_8_36 b_8 NI_8 NS_36 0 -4.5524709166990571e-06
GC_8_37 b_8 NI_8 NS_37 0 -3.9431758241153251e-05
GC_8_38 b_8 NI_8 NS_38 0 -1.9713943832070499e-05
GC_8_39 b_8 NI_8 NS_39 0 -4.8992939421782573e-06
GC_8_40 b_8 NI_8 NS_40 0 6.5785874555566327e-06
GC_8_41 b_8 NI_8 NS_41 0 -8.6427713688287946e-06
GC_8_42 b_8 NI_8 NS_42 0 -6.9219423033174982e-07
GC_8_43 b_8 NI_8 NS_43 0 -1.4971140805398893e-05
GC_8_44 b_8 NI_8 NS_44 0 2.4256379860371842e-05
GC_8_45 b_8 NI_8 NS_45 0 1.0744569679965700e-06
GC_8_46 b_8 NI_8 NS_46 0 2.6313437291496218e-06
GC_8_47 b_8 NI_8 NS_47 0 3.0498344198908487e-06
GC_8_48 b_8 NI_8 NS_48 0 1.8288496687766076e-05
GC_8_49 b_8 NI_8 NS_49 0 7.7498847463466521e-06
GC_8_50 b_8 NI_8 NS_50 0 -1.6761118287953399e-06
GC_8_51 b_8 NI_8 NS_51 0 2.9830305144710833e-06
GC_8_52 b_8 NI_8 NS_52 0 -3.4643478506601707e-07
GC_8_53 b_8 NI_8 NS_53 0 7.3243714717085940e-06
GC_8_54 b_8 NI_8 NS_54 0 -4.5247775712160395e-06
GC_8_55 b_8 NI_8 NS_55 0 -8.5040185247327499e-07
GC_8_56 b_8 NI_8 NS_56 0 -5.4040926398284354e-07
GC_8_57 b_8 NI_8 NS_57 0 -1.6433415732347617e-06
GC_8_58 b_8 NI_8 NS_58 0 2.2712849584384373e-07
GC_8_59 b_8 NI_8 NS_59 0 1.5096346114262030e-06
GC_8_60 b_8 NI_8 NS_60 0 1.1119782353376017e-07
GC_8_61 b_8 NI_8 NS_61 0 3.6029693279540004e-06
GC_8_62 b_8 NI_8 NS_62 0 -8.9726919190041775e-07
GC_8_63 b_8 NI_8 NS_63 0 -7.2239894776202718e-08
GC_8_64 b_8 NI_8 NS_64 0 -3.6343529785073757e-07
GC_8_65 b_8 NI_8 NS_65 0 -5.1807647677127100e-07
GC_8_66 b_8 NI_8 NS_66 0 5.4927162261811462e-07
GC_8_67 b_8 NI_8 NS_67 0 2.4014189943212754e-06
GC_8_68 b_8 NI_8 NS_68 0 1.9776742954056247e-07
GC_8_69 b_8 NI_8 NS_69 0 3.3593890252048213e-06
GC_8_70 b_8 NI_8 NS_70 0 -2.8068096152642622e-06
GC_8_71 b_8 NI_8 NS_71 0 -2.6297108066394321e-07
GC_8_72 b_8 NI_8 NS_72 0 -4.3648211821428127e-08
GC_8_73 b_8 NI_8 NS_73 0 7.5092993295866917e-07
GC_8_74 b_8 NI_8 NS_74 0 1.0610002796827943e-06
GC_8_75 b_8 NI_8 NS_75 0 3.5142730470775680e-06
GC_8_76 b_8 NI_8 NS_76 0 7.2317612413715887e-08
GC_8_77 b_8 NI_8 NS_77 0 2.4243650827701264e-06
GC_8_78 b_8 NI_8 NS_78 0 -4.6016400843597716e-06
GC_8_79 b_8 NI_8 NS_79 0 4.5912071532479023e-07
GC_8_80 b_8 NI_8 NS_80 0 1.1635563823075015e-06
GC_8_81 b_8 NI_8 NS_81 0 3.6822512841017166e-06
GC_8_82 b_8 NI_8 NS_82 0 -6.4052576650703278e-07
GC_8_83 b_8 NI_8 NS_83 0 5.5776194162597510e-06
GC_8_84 b_8 NI_8 NS_84 0 -9.4618052309093366e-07
GC_8_85 b_8 NI_8 NS_85 0 -1.6056023736853449e-05
GC_8_86 b_8 NI_8 NS_86 0 -1.0583746476577342e-05
GC_8_87 b_8 NI_8 NS_87 0 9.9492189482262888e-07
GC_8_88 b_8 NI_8 NS_88 0 -7.4396810500744624e-06
GC_8_89 b_8 NI_8 NS_89 0 -6.5942239962936902e-08
GC_8_90 b_8 NI_8 NS_90 0 -1.4872747453038400e-07
GC_8_91 b_8 NI_8 NS_91 0 1.8258064703679051e-06
GC_8_92 b_8 NI_8 NS_92 0 -1.8648483167661215e-06
GC_8_93 b_8 NI_8 NS_93 0 5.4044585703445990e-07
GC_8_94 b_8 NI_8 NS_94 0 -3.3794469469994227e-06
GC_8_95 b_8 NI_8 NS_95 0 3.3892711249337286e-06
GC_8_96 b_8 NI_8 NS_96 0 -1.3110545856615481e-06
GC_8_97 b_8 NI_8 NS_97 0 4.5672114750636040e-06
GC_8_98 b_8 NI_8 NS_98 0 -7.9721144051775361e-07
GC_8_99 b_8 NI_8 NS_99 0 -2.0258029898138505e-07
GC_8_100 b_8 NI_8 NS_100 0 -2.0551905961445139e-07
GC_8_101 b_8 NI_8 NS_101 0 7.0588785971767428e-07
GC_8_102 b_8 NI_8 NS_102 0 1.3963578036073434e-06
GC_8_103 b_8 NI_8 NS_103 0 -7.0583214309674747e-07
GC_8_104 b_8 NI_8 NS_104 0 -1.4718781177947233e-06
GC_8_105 b_8 NI_8 NS_105 0 -6.2724991724620084e-07
GC_8_106 b_8 NI_8 NS_106 0 8.2981064818168461e-07
GC_8_107 b_8 NI_8 NS_107 0 2.2262539144369858e-07
GC_8_108 b_8 NI_8 NS_108 0 6.5365102637855797e-07
GC_8_109 b_8 NI_8 NS_109 0 5.9754309503493592e-07
GC_8_110 b_8 NI_8 NS_110 0 2.1049186414085253e-08
GC_8_111 b_8 NI_8 NS_111 0 1.4042915235816373e-11
GC_8_112 b_8 NI_8 NS_112 0 1.0067978772828576e-12
GC_8_113 b_8 NI_8 NS_113 0 4.3083056118656987e-10
GC_8_114 b_8 NI_8 NS_114 0 1.6517097585592210e-09
GC_8_115 b_8 NI_8 NS_115 0 6.6701478702326392e-05
GC_8_116 b_8 NI_8 NS_116 0 2.1487602561808342e-07
GC_8_117 b_8 NI_8 NS_117 0 2.2380666884705768e-11
GC_8_118 b_8 NI_8 NS_118 0 -9.9152097981121332e-10
GC_8_119 b_8 NI_8 NS_119 0 4.3114285984214290e-07
GC_8_120 b_8 NI_8 NS_120 0 1.8615280312004883e-07
GC_8_121 b_8 NI_8 NS_121 0 6.0533479245496665e-07
GC_8_122 b_8 NI_8 NS_122 0 5.0362649972884689e-07
GC_8_123 b_8 NI_8 NS_123 0 2.9724322721516425e-06
GC_8_124 b_8 NI_8 NS_124 0 -1.5630093061709232e-06
GC_8_125 b_8 NI_8 NS_125 0 -1.1990741804850255e-06
GC_8_126 b_8 NI_8 NS_126 0 -1.1274223693487281e-06
GC_8_127 b_8 NI_8 NS_127 0 2.3740969869189682e-06
GC_8_128 b_8 NI_8 NS_128 0 -8.7014418839566818e-07
GC_8_129 b_8 NI_8 NS_129 0 -2.5791878926801263e-06
GC_8_130 b_8 NI_8 NS_130 0 -6.4188238359351265e-06
GC_8_131 b_8 NI_8 NS_131 0 1.1120470018854172e-07
GC_8_132 b_8 NI_8 NS_132 0 1.6980774846763208e-06
GC_8_133 b_8 NI_8 NS_133 0 -1.7225279931433457e-06
GC_8_134 b_8 NI_8 NS_134 0 5.0765358392714987e-07
GC_8_135 b_8 NI_8 NS_135 0 3.1223259564598447e-06
GC_8_136 b_8 NI_8 NS_136 0 -4.3467314955875459e-06
GC_8_137 b_8 NI_8 NS_137 0 -6.6651214357343690e-06
GC_8_138 b_8 NI_8 NS_138 0 1.1614615577668215e-06
GC_8_139 b_8 NI_8 NS_139 0 -4.7510519303260580e-07
GC_8_140 b_8 NI_8 NS_140 0 1.6872444372266646e-06
GC_8_141 b_8 NI_8 NS_141 0 -2.1293703716488189e-06
GC_8_142 b_8 NI_8 NS_142 0 -4.2560135982618052e-06
GC_8_143 b_8 NI_8 NS_143 0 -2.2153025138672841e-06
GC_8_144 b_8 NI_8 NS_144 0 2.1659200774326960e-06
GC_8_145 b_8 NI_8 NS_145 0 3.1593365913160003e-06
GC_8_146 b_8 NI_8 NS_146 0 3.0711649292284910e-06
GC_8_147 b_8 NI_8 NS_147 0 -6.0923058511645008e-06
GC_8_148 b_8 NI_8 NS_148 0 -4.4508806379831469e-06
GC_8_149 b_8 NI_8 NS_149 0 -1.2975247120999128e-06
GC_8_150 b_8 NI_8 NS_150 0 2.1675953995370491e-06
GC_8_151 b_8 NI_8 NS_151 0 2.8169733745596119e-07
GC_8_152 b_8 NI_8 NS_152 0 -2.8035792199559832e-06
GC_8_153 b_8 NI_8 NS_153 0 -3.1939608038239276e-06
GC_8_154 b_8 NI_8 NS_154 0 1.8340038055049179e-06
GC_8_155 b_8 NI_8 NS_155 0 -3.1234084960689102e-07
GC_8_156 b_8 NI_8 NS_156 0 2.3430257675488221e-06
GC_8_157 b_8 NI_8 NS_157 0 -1.4637158301739735e-06
GC_8_158 b_8 NI_8 NS_158 0 -2.6210655510492688e-06
GC_8_159 b_8 NI_8 NS_159 0 -1.8974250033340522e-06
GC_8_160 b_8 NI_8 NS_160 0 1.3687528370010508e-06
GC_8_161 b_8 NI_8 NS_161 0 1.1585941289080486e-06
GC_8_162 b_8 NI_8 NS_162 0 -6.4540638095425139e-07
GC_8_163 b_8 NI_8 NS_163 0 -3.5960771508100279e-06
GC_8_164 b_8 NI_8 NS_164 0 2.8645283265555657e-07
GC_8_165 b_8 NI_8 NS_165 0 -8.2546485919302936e-07
GC_8_166 b_8 NI_8 NS_166 0 7.2322598123757943e-07
GC_8_167 b_8 NI_8 NS_167 0 -1.8925801891011071e-06
GC_8_168 b_8 NI_8 NS_168 0 -1.3277337261992181e-06
GC_8_169 b_8 NI_8 NS_169 0 -1.4489411158612972e-06
GC_8_170 b_8 NI_8 NS_170 0 5.5829929489541187e-07
GC_8_171 b_8 NI_8 NS_171 0 -1.0698697945744048e-06
GC_8_172 b_8 NI_8 NS_172 0 -5.9277169872623101e-07
GC_8_173 b_8 NI_8 NS_173 0 -2.3266421240768062e-06
GC_8_174 b_8 NI_8 NS_174 0 -6.7325062334453606e-07
GC_8_175 b_8 NI_8 NS_175 0 -2.8005573602142289e-06
GC_8_176 b_8 NI_8 NS_176 0 -5.7579635065162049e-07
GC_8_177 b_8 NI_8 NS_177 0 -2.0701484255780899e-06
GC_8_178 b_8 NI_8 NS_178 0 2.3474578307455500e-07
GC_8_179 b_8 NI_8 NS_179 0 -2.5970652556167733e-06
GC_8_180 b_8 NI_8 NS_180 0 1.0366537599693077e-07
GC_8_181 b_8 NI_8 NS_181 0 -3.9148789821076441e-06
GC_8_182 b_8 NI_8 NS_182 0 -7.2842870175883121e-07
GC_8_183 b_8 NI_8 NS_183 0 -5.2762866338299168e-06
GC_8_184 b_8 NI_8 NS_184 0 1.8897598182887802e-06
GC_8_185 b_8 NI_8 NS_185 0 -2.9592147848470277e-06
GC_8_186 b_8 NI_8 NS_186 0 1.7284775866503526e-06
GC_8_187 b_8 NI_8 NS_187 0 -3.7956745639874173e-06
GC_8_188 b_8 NI_8 NS_188 0 2.9627449302113527e-06
GC_8_189 b_8 NI_8 NS_189 0 -5.2520804080494296e-06
GC_8_190 b_8 NI_8 NS_190 0 1.3679659336618500e-06
GC_8_191 b_8 NI_8 NS_191 0 -2.9739725693452381e-06
GC_8_192 b_8 NI_8 NS_192 0 7.6177906178030104e-06
GC_8_193 b_8 NI_8 NS_193 0 -1.9309245794914865e-06
GC_8_194 b_8 NI_8 NS_194 0 4.3923521415424183e-06
GC_8_195 b_8 NI_8 NS_195 0 1.5636686497098740e-06
GC_8_196 b_8 NI_8 NS_196 0 4.8436713794079585e-06
GC_8_197 b_8 NI_8 NS_197 0 -9.8795386638447127e-07
GC_8_198 b_8 NI_8 NS_198 0 3.6442595552559610e-06
GC_8_199 b_8 NI_8 NS_199 0 -1.0320720630421068e-05
GC_8_200 b_8 NI_8 NS_200 0 3.3102409889430702e-05
GC_8_201 b_8 NI_8 NS_201 0 1.3164927833764437e-06
GC_8_202 b_8 NI_8 NS_202 0 1.2184840768364405e-06
GC_8_203 b_8 NI_8 NS_203 0 -9.3710834065955694e-08
GC_8_204 b_8 NI_8 NS_204 0 8.7633969048653555e-08
GC_8_205 b_8 NI_8 NS_205 0 -3.3515210262058317e-07
GC_8_206 b_8 NI_8 NS_206 0 2.6717604987726500e-06
GC_8_207 b_8 NI_8 NS_207 0 7.2368361113139429e-07
GC_8_208 b_8 NI_8 NS_208 0 1.5966468684301533e-07
GC_8_209 b_8 NI_8 NS_209 0 3.0760810477641118e-06
GC_8_210 b_8 NI_8 NS_210 0 -2.7795578509055835e-06
GC_8_211 b_8 NI_8 NS_211 0 -1.9947428618217774e-07
GC_8_212 b_8 NI_8 NS_212 0 -1.1674120017937913e-05
GC_8_213 b_8 NI_8 NS_213 0 1.9433166998062350e-06
GC_8_214 b_8 NI_8 NS_214 0 -6.7943785955979901e-07
GC_8_215 b_8 NI_8 NS_215 0 4.3063509523488301e-06
GC_8_216 b_8 NI_8 NS_216 0 -1.7890106489573844e-07
GC_8_217 b_8 NI_8 NS_217 0 1.2121027942105582e-06
GC_8_218 b_8 NI_8 NS_218 0 1.8711460144681166e-06
GC_8_219 b_8 NI_8 NS_219 0 1.6466082897143810e-06
GC_8_220 b_8 NI_8 NS_220 0 -7.9762654538069011e-07
GC_8_221 b_8 NI_8 NS_221 0 5.9154025877315865e-07
GC_8_222 b_8 NI_8 NS_222 0 4.7824092161486622e-07
GC_8_223 b_8 NI_8 NS_223 0 6.8251383705154019e-07
GC_8_224 b_8 NI_8 NS_224 0 -9.6216812545433910e-08
GC_8_225 b_8 NI_8 NS_225 0 2.5753545760960377e-11
GC_8_226 b_8 NI_8 NS_226 0 -9.7279592873187154e-11
GC_8_227 b_8 NI_8 NS_227 0 -1.9600542294593044e-09
GC_8_228 b_8 NI_8 NS_228 0 4.2972487710579606e-09
GC_8_229 b_8 NI_8 NS_229 0 -3.2373977337425789e-05
GC_8_230 b_8 NI_8 NS_230 0 2.2170617398789061e-06
GC_8_231 b_8 NI_8 NS_231 0 6.8028427126293341e-11
GC_8_232 b_8 NI_8 NS_232 0 3.0563739672171638e-09
GC_8_233 b_8 NI_8 NS_233 0 -1.7156139982086798e-06
GC_8_234 b_8 NI_8 NS_234 0 -1.8282680237076224e-06
GC_8_235 b_8 NI_8 NS_235 0 -5.3488497316932639e-06
GC_8_236 b_8 NI_8 NS_236 0 2.8545827564616671e-06
GC_8_237 b_8 NI_8 NS_237 0 -1.6536988260264160e-05
GC_8_238 b_8 NI_8 NS_238 0 1.8376723758867093e-05
GC_8_239 b_8 NI_8 NS_239 0 1.5065179779432959e-05
GC_8_240 b_8 NI_8 NS_240 0 9.7699986544503514e-06
GC_8_241 b_8 NI_8 NS_241 0 1.7310031908075085e-05
GC_8_242 b_8 NI_8 NS_242 0 2.2719453567803186e-05
GC_8_243 b_8 NI_8 NS_243 0 2.9106631708776806e-05
GC_8_244 b_8 NI_8 NS_244 0 4.9748903172865757e-06
GC_8_245 b_8 NI_8 NS_245 0 -2.9665367336013985e-06
GC_8_246 b_8 NI_8 NS_246 0 -1.8804713539111336e-06
GC_8_247 b_8 NI_8 NS_247 0 1.6935044223643993e-05
GC_8_248 b_8 NI_8 NS_248 0 -2.2271406612322304e-06
GC_8_249 b_8 NI_8 NS_249 0 1.2887258600352908e-04
GC_8_250 b_8 NI_8 NS_250 0 3.4717434655312075e-05
GC_8_251 b_8 NI_8 NS_251 0 -2.8878620456250753e-05
GC_8_252 b_8 NI_8 NS_252 0 -9.8668107722263575e-05
GC_8_253 b_8 NI_8 NS_253 0 2.4897077674231659e-05
GC_8_254 b_8 NI_8 NS_254 0 -3.1464183790394452e-05
GC_8_255 b_8 NI_8 NS_255 0 -4.1611411743458107e-05
GC_8_256 b_8 NI_8 NS_256 0 -1.6650642318829462e-04
GC_8_257 b_8 NI_8 NS_257 0 -4.1828489446790585e-05
GC_8_258 b_8 NI_8 NS_258 0 -4.8978468111330464e-06
GC_8_259 b_8 NI_8 NS_259 0 2.1414128756167459e-05
GC_8_260 b_8 NI_8 NS_260 0 -1.5190517227923084e-04
GC_8_261 b_8 NI_8 NS_261 0 -2.3047124271565446e-04
GC_8_262 b_8 NI_8 NS_262 0 1.1445044845436983e-04
GC_8_263 b_8 NI_8 NS_263 0 -3.7401825748035043e-05
GC_8_264 b_8 NI_8 NS_264 0 1.4352682093440199e-05
GC_8_265 b_8 NI_8 NS_265 0 -1.3776551196360831e-04
GC_8_266 b_8 NI_8 NS_266 0 1.3054679569781544e-04
GC_8_267 b_8 NI_8 NS_267 0 3.6494591253322858e-05
GC_8_268 b_8 NI_8 NS_268 0 4.1231203437896011e-05
GC_8_269 b_8 NI_8 NS_269 0 -3.8131630707688927e-05
GC_8_270 b_8 NI_8 NS_270 0 4.3361081045850004e-05
GC_8_271 b_8 NI_8 NS_271 0 8.7555844314140302e-05
GC_8_272 b_8 NI_8 NS_272 0 1.1842919293832428e-04
GC_8_273 b_8 NI_8 NS_273 0 2.7361530685580764e-05
GC_8_274 b_8 NI_8 NS_274 0 1.0121201737672454e-05
GC_8_275 b_8 NI_8 NS_275 0 8.7344637251898869e-05
GC_8_276 b_8 NI_8 NS_276 0 6.5655939896238903e-05
GC_8_277 b_8 NI_8 NS_277 0 2.0321378146137156e-05
GC_8_278 b_8 NI_8 NS_278 0 -5.7038888509518223e-05
GC_8_279 b_8 NI_8 NS_279 0 1.6978946298417043e-05
GC_8_280 b_8 NI_8 NS_280 0 -8.9185276916070482e-06
GC_8_281 b_8 NI_8 NS_281 0 8.5891152829056381e-06
GC_8_282 b_8 NI_8 NS_282 0 -3.2921322821813578e-05
GC_8_283 b_8 NI_8 NS_283 0 -8.8488157050203741e-06
GC_8_284 b_8 NI_8 NS_284 0 5.5965388694198801e-07
GC_8_285 b_8 NI_8 NS_285 0 -2.4314155309708924e-06
GC_8_286 b_8 NI_8 NS_286 0 8.5078379753188616e-06
GC_8_287 b_8 NI_8 NS_287 0 1.0240904457618469e-05
GC_8_288 b_8 NI_8 NS_288 0 6.0554414451221057e-06
GC_8_289 b_8 NI_8 NS_289 0 1.2188371322591714e-05
GC_8_290 b_8 NI_8 NS_290 0 -7.8214804293912399e-06
GC_8_291 b_8 NI_8 NS_291 0 -3.4896271688717365e-06
GC_8_292 b_8 NI_8 NS_292 0 -4.3246146588597668e-07
GC_8_293 b_8 NI_8 NS_293 0 2.4743816315827772e-06
GC_8_294 b_8 NI_8 NS_294 0 7.4083949194489401e-06
GC_8_295 b_8 NI_8 NS_295 0 1.3659374209138464e-05
GC_8_296 b_8 NI_8 NS_296 0 2.6169682058911768e-06
GC_8_297 b_8 NI_8 NS_297 0 4.5330463493605632e-06
GC_8_298 b_8 NI_8 NS_298 0 -1.4186507098728478e-05
GC_8_299 b_8 NI_8 NS_299 0 -5.9288335650460138e-06
GC_8_300 b_8 NI_8 NS_300 0 4.2661558160660471e-06
GC_8_301 b_8 NI_8 NS_301 0 1.0298030473444926e-05
GC_8_302 b_8 NI_8 NS_302 0 9.9363433278093851e-06
GC_8_303 b_8 NI_8 NS_303 0 1.7307569962841289e-05
GC_8_304 b_8 NI_8 NS_304 0 -4.2766878177167002e-06
GC_8_305 b_8 NI_8 NS_305 0 -9.2960035563669747e-06
GC_8_306 b_8 NI_8 NS_306 0 -1.5305389764069588e-05
GC_8_307 b_8 NI_8 NS_307 0 -4.0930062175161154e-06
GC_8_308 b_8 NI_8 NS_308 0 1.3520391623851333e-05
GC_8_309 b_8 NI_8 NS_309 0 2.0923680867374372e-05
GC_8_310 b_8 NI_8 NS_310 0 -5.4865029872128641e-07
GC_8_311 b_8 NI_8 NS_311 0 8.8629081181941437e-06
GC_8_312 b_8 NI_8 NS_312 0 -1.7438354234438960e-05
GC_8_313 b_8 NI_8 NS_313 0 2.5763866611130719e-06
GC_8_314 b_8 NI_8 NS_314 0 -1.3772995331204317e-05
GC_8_315 b_8 NI_8 NS_315 0 -1.3801385147929991e-05
GC_8_316 b_8 NI_8 NS_316 0 4.4170656762483018e-06
GC_8_317 b_8 NI_8 NS_317 0 1.6023760120314050e-08
GC_8_318 b_8 NI_8 NS_318 0 -4.1749247038077964e-08
GC_8_319 b_8 NI_8 NS_319 0 8.6200011835323138e-06
GC_8_320 b_8 NI_8 NS_320 0 1.1611709540868862e-05
GC_8_321 b_8 NI_8 NS_321 0 1.0921436716279523e-05
GC_8_322 b_8 NI_8 NS_322 0 -1.1277737524549733e-05
GC_8_323 b_8 NI_8 NS_323 0 -3.7555133256338342e-06
GC_8_324 b_8 NI_8 NS_324 0 -1.0184188809217565e-05
GC_8_325 b_8 NI_8 NS_325 0 -2.3202504973889939e-06
GC_8_326 b_8 NI_8 NS_326 0 1.2931865048131915e-05
GC_8_327 b_8 NI_8 NS_327 0 9.7593852904956323e-07
GC_8_328 b_8 NI_8 NS_328 0 -7.2834606985686015e-06
GC_8_329 b_8 NI_8 NS_329 0 7.5034051036803983e-06
GC_8_330 b_8 NI_8 NS_330 0 1.6765299762800522e-06
GC_8_331 b_8 NI_8 NS_331 0 -6.0990911004070706e-06
GC_8_332 b_8 NI_8 NS_332 0 -8.8899452328550399e-06
GC_8_333 b_8 NI_8 NS_333 0 -4.1232006303653826e-06
GC_8_334 b_8 NI_8 NS_334 0 9.6572720631975889e-06
GC_8_335 b_8 NI_8 NS_335 0 3.3299191854629409e-06
GC_8_336 b_8 NI_8 NS_336 0 6.0429585603993354e-06
GC_8_337 b_8 NI_8 NS_337 0 5.6621019731116777e-06
GC_8_338 b_8 NI_8 NS_338 0 5.1491841621574102e-07
GC_8_339 b_8 NI_8 NS_339 0 6.1218441300162927e-11
GC_8_340 b_8 NI_8 NS_340 0 1.4945626116593220e-10
GC_8_341 b_8 NI_8 NS_341 0 5.9799306355330419e-09
GC_8_342 b_8 NI_8 NS_342 0 -8.3554324562227200e-09
GC_8_343 b_8 NI_8 NS_343 0 -1.0995071593363421e-04
GC_8_344 b_8 NI_8 NS_344 0 -2.1492391062527274e-06
GC_8_345 b_8 NI_8 NS_345 0 -2.5033374423560352e-10
GC_8_346 b_8 NI_8 NS_346 0 2.6123671577754751e-09
GC_8_347 b_8 NI_8 NS_347 0 1.8909814804427741e-06
GC_8_348 b_8 NI_8 NS_348 0 -1.6338261323707834e-06
GC_8_349 b_8 NI_8 NS_349 0 3.4328427680563642e-07
GC_8_350 b_8 NI_8 NS_350 0 -6.5685023373413638e-06
GC_8_351 b_8 NI_8 NS_351 0 -7.5232096050962672e-06
GC_8_352 b_8 NI_8 NS_352 0 -5.2405397712347920e-07
GC_8_353 b_8 NI_8 NS_353 0 -1.5644385723909789e-06
GC_8_354 b_8 NI_8 NS_354 0 -4.8503530140566803e-06
GC_8_355 b_8 NI_8 NS_355 0 -1.6089131236244526e-05
GC_8_356 b_8 NI_8 NS_356 0 -2.1861621814160747e-06
GC_8_357 b_8 NI_8 NS_357 0 -7.5367525524654000e-06
GC_8_358 b_8 NI_8 NS_358 0 1.8919009563555713e-05
GC_8_359 b_8 NI_8 NS_359 0 5.0282697868662988e-06
GC_8_360 b_8 NI_8 NS_360 0 -2.8006236751205509e-06
GC_8_361 b_8 NI_8 NS_361 0 -2.3106458747657329e-07
GC_8_362 b_8 NI_8 NS_362 0 -2.4616852107808365e-06
GC_8_363 b_8 NI_8 NS_363 0 -2.6994514413638635e-05
GC_8_364 b_8 NI_8 NS_364 0 2.8300303688318277e-05
GC_8_365 b_8 NI_8 NS_365 0 2.8448289021857441e-05
GC_8_366 b_8 NI_8 NS_366 0 -7.8440798653694632e-06
GC_8_367 b_8 NI_8 NS_367 0 -8.2731828788077668e-06
GC_8_368 b_8 NI_8 NS_368 0 -4.3391055889547900e-06
GC_8_369 b_8 NI_8 NS_369 0 1.2150359881480514e-05
GC_8_370 b_8 NI_8 NS_370 0 2.7749141253524124e-05
GC_8_371 b_8 NI_8 NS_371 0 1.4969706146806489e-06
GC_8_372 b_8 NI_8 NS_372 0 -8.9353113195543254e-06
GC_8_373 b_8 NI_8 NS_373 0 -2.9031331281288270e-05
GC_8_374 b_8 NI_8 NS_374 0 4.5480857394694135e-06
GC_8_375 b_8 NI_8 NS_375 0 4.1816723861543067e-05
GC_8_376 b_8 NI_8 NS_376 0 1.1681510531873194e-05
GC_8_377 b_8 NI_8 NS_377 0 -3.0448948219637981e-06
GC_8_378 b_8 NI_8 NS_378 0 -4.4842327319119856e-06
GC_8_379 b_8 NI_8 NS_379 0 1.2838681870413446e-05
GC_8_380 b_8 NI_8 NS_380 0 1.9718562859981764e-05
GC_8_381 b_8 NI_8 NS_381 0 3.9956457988626063e-06
GC_8_382 b_8 NI_8 NS_382 0 -1.0979149477818060e-05
GC_8_383 b_8 NI_8 NS_383 0 -6.6146714666948186e-06
GC_8_384 b_8 NI_8 NS_384 0 8.3775244381893879e-07
GC_8_385 b_8 NI_8 NS_385 0 1.9105218500751744e-05
GC_8_386 b_8 NI_8 NS_386 0 5.9545118531729413e-06
GC_8_387 b_8 NI_8 NS_387 0 -4.3481236042559753e-08
GC_8_388 b_8 NI_8 NS_388 0 -4.2143336088428541e-06
GC_8_389 b_8 NI_8 NS_389 0 4.6805663505283409e-06
GC_8_390 b_8 NI_8 NS_390 0 1.4625900374383416e-05
GC_8_391 b_8 NI_8 NS_391 0 8.1127083732355065e-06
GC_8_392 b_8 NI_8 NS_392 0 -1.1159021566279000e-05
GC_8_393 b_8 NI_8 NS_393 0 -1.4428375570273185e-06
GC_8_394 b_8 NI_8 NS_394 0 9.3170779297651210e-07
GC_8_395 b_8 NI_8 NS_395 0 1.0891210589817904e-05
GC_8_396 b_8 NI_8 NS_396 0 4.3456004040947175e-06
GC_8_397 b_8 NI_8 NS_397 0 1.7188897594320207e-06
GC_8_398 b_8 NI_8 NS_398 0 -6.0609920065333681e-07
GC_8_399 b_8 NI_8 NS_399 0 5.6777116727859837e-06
GC_8_400 b_8 NI_8 NS_400 0 1.7899370616409791e-06
GC_8_401 b_8 NI_8 NS_401 0 3.3742922933278677e-06
GC_8_402 b_8 NI_8 NS_402 0 2.0720323011922782e-06
GC_8_403 b_8 NI_8 NS_403 0 1.0916608312203075e-05
GC_8_404 b_8 NI_8 NS_404 0 3.9123303383116289e-06
GC_8_405 b_8 NI_8 NS_405 0 4.8432409649530370e-06
GC_8_406 b_8 NI_8 NS_406 0 -4.2628886166095313e-08
GC_8_407 b_8 NI_8 NS_407 0 9.9680750076085025e-06
GC_8_408 b_8 NI_8 NS_408 0 -9.9862876900387255e-07
GC_8_409 b_8 NI_8 NS_409 0 8.1884656224278131e-06
GC_8_410 b_8 NI_8 NS_410 0 2.9679944269843811e-06
GC_8_411 b_8 NI_8 NS_411 0 1.8986720032126656e-05
GC_8_412 b_8 NI_8 NS_412 0 -5.4365284664606446e-06
GC_8_413 b_8 NI_8 NS_413 0 7.1694241678354561e-06
GC_8_414 b_8 NI_8 NS_414 0 -3.9853757715760395e-06
GC_8_415 b_8 NI_8 NS_415 0 1.3685887058883454e-05
GC_8_416 b_8 NI_8 NS_416 0 -1.1804061819722942e-05
GC_8_417 b_8 NI_8 NS_417 0 1.2305622481603828e-05
GC_8_418 b_8 NI_8 NS_418 0 -3.9592531329760032e-06
GC_8_419 b_8 NI_8 NS_419 0 9.0879427380302472e-06
GC_8_420 b_8 NI_8 NS_420 0 -2.6621762682054804e-05
GC_8_421 b_8 NI_8 NS_421 0 2.2848314801757932e-06
GC_8_422 b_8 NI_8 NS_422 0 -1.2337140601772232e-05
GC_8_423 b_8 NI_8 NS_423 0 -8.3397818234636159e-06
GC_8_424 b_8 NI_8 NS_424 0 -1.8510652810791159e-05
GC_8_425 b_8 NI_8 NS_425 0 -5.0670738844842952e-06
GC_8_426 b_8 NI_8 NS_426 0 -1.2091739298219231e-05
GC_8_427 b_8 NI_8 NS_427 0 5.5654557816156790e-05
GC_8_428 b_8 NI_8 NS_428 0 -8.7608658594514623e-05
GC_8_429 b_8 NI_8 NS_429 0 -1.0050338716018578e-05
GC_8_430 b_8 NI_8 NS_430 0 1.5956330416666998e-06
GC_8_431 b_8 NI_8 NS_431 0 3.9373700602922472e-07
GC_8_432 b_8 NI_8 NS_432 0 -1.2103089213046396e-07
GC_8_433 b_8 NI_8 NS_433 0 -2.7541899515870780e-06
GC_8_434 b_8 NI_8 NS_434 0 -1.8116239241423931e-06
GC_8_435 b_8 NI_8 NS_435 0 -4.3434373575026019e-06
GC_8_436 b_8 NI_8 NS_436 0 6.8569502514683423e-07
GC_8_437 b_8 NI_8 NS_437 0 -1.7627012006832803e-05
GC_8_438 b_8 NI_8 NS_438 0 9.5650461593923458e-06
GC_8_439 b_8 NI_8 NS_439 0 -9.4006803689285239e-06
GC_8_440 b_8 NI_8 NS_440 0 3.7414742800988149e-05
GC_8_441 b_8 NI_8 NS_441 0 -7.2091675842040575e-06
GC_8_442 b_8 NI_8 NS_442 0 3.1130495402704615e-07
GC_8_443 b_8 NI_8 NS_443 0 -1.3385611199619336e-05
GC_8_444 b_8 NI_8 NS_444 0 1.8110375252004105e-06
GC_8_445 b_8 NI_8 NS_445 0 -4.6173103193827154e-06
GC_8_446 b_8 NI_8 NS_446 0 -3.3928410486765216e-06
GC_8_447 b_8 NI_8 NS_447 0 -6.3738660673577197e-06
GC_8_448 b_8 NI_8 NS_448 0 1.0329454905662900e-06
GC_8_449 b_8 NI_8 NS_449 0 -3.0262565554308511e-06
GC_8_450 b_8 NI_8 NS_450 0 8.9218043005674206e-07
GC_8_451 b_8 NI_8 NS_451 0 -1.7748342711559983e-06
GC_8_452 b_8 NI_8 NS_452 0 -9.4793262689217010e-07
GC_8_453 b_8 NI_8 NS_453 0 -2.6182135252001881e-10
GC_8_454 b_8 NI_8 NS_454 0 4.2365472539275098e-10
GC_8_455 b_8 NI_8 NS_455 0 2.2745886103270986e-09
GC_8_456 b_8 NI_8 NS_456 0 -2.6878267994866984e-08
GC_8_457 b_8 NI_8 NS_457 0 3.0950393739609121e-03
GC_8_458 b_8 NI_8 NS_458 0 -6.1289419952542960e-04
GC_8_459 b_8 NI_8 NS_459 0 2.8121768806274474e-08
GC_8_460 b_8 NI_8 NS_460 0 -3.1528675830433718e-08
GC_8_461 b_8 NI_8 NS_461 0 2.0500749013526636e-04
GC_8_462 b_8 NI_8 NS_462 0 1.3546525854947404e-04
GC_8_463 b_8 NI_8 NS_463 0 5.6415244013022291e-04
GC_8_464 b_8 NI_8 NS_464 0 2.6382417189227647e-04
GC_8_465 b_8 NI_8 NS_465 0 3.0949145364878527e-03
GC_8_466 b_8 NI_8 NS_466 0 -2.2211768907149276e-03
GC_8_467 b_8 NI_8 NS_467 0 -1.5948048505893503e-03
GC_8_468 b_8 NI_8 NS_468 0 -2.6831565243659963e-03
GC_8_469 b_8 NI_8 NS_469 0 -2.0664402239951906e-03
GC_8_470 b_8 NI_8 NS_470 0 -3.7810164315909009e-03
GC_8_471 b_8 NI_8 NS_471 0 -4.9930245005376638e-03
GC_8_472 b_8 NI_8 NS_472 0 -1.5154927975483919e-03
GC_8_473 b_8 NI_8 NS_473 0 2.9714191235064865e-04
GC_8_474 b_8 NI_8 NS_474 0 1.9409433219026896e-04
GC_8_475 b_8 NI_8 NS_475 0 -2.8708433759163355e-03
GC_8_476 b_8 NI_8 NS_476 0 -9.4557922468997484e-04
GC_8_477 b_8 NI_8 NS_477 0 -2.2198356738005930e-02
GC_8_478 b_8 NI_8 NS_478 0 -1.0125160180584833e-02
GC_8_479 b_8 NI_8 NS_479 0 1.2231820315885117e-03
GC_8_480 b_8 NI_8 NS_480 0 2.0396448747319079e-02
GC_8_481 b_8 NI_8 NS_481 0 -5.8225961304134892e-03
GC_8_482 b_8 NI_8 NS_482 0 4.6364315762052284e-03
GC_8_483 b_8 NI_8 NS_483 0 5.8808211604887356e-03
GC_8_484 b_8 NI_8 NS_484 0 3.4493742840412150e-02
GC_8_485 b_8 NI_8 NS_485 0 8.0480773127163206e-03
GC_8_486 b_8 NI_8 NS_486 0 2.7589344833169756e-03
GC_8_487 b_8 NI_8 NS_487 0 -7.6367946363373913e-03
GC_8_488 b_8 NI_8 NS_488 0 2.9591949287605196e-02
GC_8_489 b_8 NI_8 NS_489 0 5.0679463987695517e-02
GC_8_490 b_8 NI_8 NS_490 0 -2.0315742000687084e-02
GC_8_491 b_8 NI_8 NS_491 0 7.9122593904820022e-03
GC_8_492 b_8 NI_8 NS_492 0 -1.6718964677352804e-03
GC_8_493 b_8 NI_8 NS_493 0 2.8952184028047650e-02
GC_8_494 b_8 NI_8 NS_494 0 -2.6605127397770930e-02
GC_8_495 b_8 NI_8 NS_495 0 -6.7717827315056977e-03
GC_8_496 b_8 NI_8 NS_496 0 -9.8520999961726977e-03
GC_8_497 b_8 NI_8 NS_497 0 8.4245545368217545e-03
GC_8_498 b_8 NI_8 NS_498 0 -8.0661008778074826e-03
GC_8_499 b_8 NI_8 NS_499 0 -1.9120468089075335e-02
GC_8_500 b_8 NI_8 NS_500 0 -2.5143594553950769e-02
GC_8_501 b_8 NI_8 NS_501 0 -5.4851139375878344e-03
GC_8_502 b_8 NI_8 NS_502 0 -2.8303873464306118e-03
GC_8_503 b_8 NI_8 NS_503 0 -1.7803813497061571e-02
GC_8_504 b_8 NI_8 NS_504 0 -1.3047348001991631e-02
GC_8_505 b_8 NI_8 NS_505 0 -4.7610269419565525e-03
GC_8_506 b_8 NI_8 NS_506 0 1.2568312272645444e-02
GC_8_507 b_8 NI_8 NS_507 0 -3.4539894410605594e-03
GC_8_508 b_8 NI_8 NS_508 0 1.5560262320147864e-03
GC_8_509 b_8 NI_8 NS_509 0 -6.8744236182587105e-04
GC_8_510 b_8 NI_8 NS_510 0 7.0157646830849435e-03
GC_8_511 b_8 NI_8 NS_511 0 1.8840814867831794e-03
GC_8_512 b_8 NI_8 NS_512 0 8.1060295412666483e-05
GC_8_513 b_8 NI_8 NS_513 0 3.0821870820571073e-04
GC_8_514 b_8 NI_8 NS_514 0 -1.9474454026678183e-03
GC_8_515 b_8 NI_8 NS_515 0 -1.8615157448309979e-03
GC_8_516 b_8 NI_8 NS_516 0 -1.6133457519509977e-03
GC_8_517 b_8 NI_8 NS_517 0 -2.1255689319405195e-03
GC_8_518 b_8 NI_8 NS_518 0 1.6940535150088063e-03
GC_8_519 b_8 NI_8 NS_519 0 7.6441489964923851e-04
GC_8_520 b_8 NI_8 NS_520 0 1.8569493778374007e-04
GC_8_521 b_8 NI_8 NS_521 0 -7.0068892034165736e-04
GC_8_522 b_8 NI_8 NS_522 0 -1.6760053809953097e-03
GC_8_523 b_8 NI_8 NS_523 0 -2.6855348489639910e-03
GC_8_524 b_8 NI_8 NS_524 0 -8.2394364030572331e-04
GC_8_525 b_8 NI_8 NS_525 0 -4.9849817671180935e-04
GC_8_526 b_8 NI_8 NS_526 0 2.9352185203747475e-03
GC_8_527 b_8 NI_8 NS_527 0 1.3528913475371119e-03
GC_8_528 b_8 NI_8 NS_528 0 -8.5706968791956096e-04
GC_8_529 b_8 NI_8 NS_529 0 -2.4223431553966794e-03
GC_8_530 b_8 NI_8 NS_530 0 -2.2652840568361432e-03
GC_8_531 b_8 NI_8 NS_531 0 -3.5590208310841056e-03
GC_8_532 b_8 NI_8 NS_532 0 7.4879921067956545e-04
GC_8_533 b_8 NI_8 NS_533 0 2.4605502179886464e-03
GC_8_534 b_8 NI_8 NS_534 0 3.0265639065871308e-03
GC_8_535 b_8 NI_8 NS_535 0 9.8335651397548165e-04
GC_8_536 b_8 NI_8 NS_536 0 -2.9400792738963023e-03
GC_8_537 b_8 NI_8 NS_537 0 -4.7724965772711417e-03
GC_8_538 b_8 NI_8 NS_538 0 5.7213344778377536e-05
GC_8_539 b_8 NI_8 NS_539 0 -1.7194831375916303e-03
GC_8_540 b_8 NI_8 NS_540 0 3.7113726641357613e-03
GC_8_541 b_8 NI_8 NS_541 0 -7.3866808123181310e-04
GC_8_542 b_8 NI_8 NS_542 0 1.5326979983791332e-03
GC_8_543 b_8 NI_8 NS_543 0 3.2195725990708450e-03
GC_8_544 b_8 NI_8 NS_544 0 -1.3349998191154707e-03
GC_8_545 b_8 NI_8 NS_545 0 -2.8022973719014715e-06
GC_8_546 b_8 NI_8 NS_546 0 8.9859681681350464e-06
GC_8_547 b_8 NI_8 NS_547 0 -1.8210614205990429e-03
GC_8_548 b_8 NI_8 NS_548 0 -2.5224010433460703e-03
GC_8_549 b_8 NI_8 NS_549 0 -2.4088305332291343e-03
GC_8_550 b_8 NI_8 NS_550 0 2.4933220795179773e-03
GC_8_551 b_8 NI_8 NS_551 0 1.0059043253014639e-03
GC_8_552 b_8 NI_8 NS_552 0 2.4239834981763667e-03
GC_8_553 b_8 NI_8 NS_553 0 8.4854741839266010e-04
GC_8_554 b_8 NI_8 NS_554 0 -2.6997877006754720e-03
GC_8_555 b_8 NI_8 NS_555 0 -3.0628339353289791e-04
GC_8_556 b_8 NI_8 NS_556 0 1.6736613910303226e-03
GC_8_557 b_8 NI_8 NS_557 0 -1.7824226170147987e-03
GC_8_558 b_8 NI_8 NS_558 0 -3.1430315347359054e-04
GC_8_559 b_8 NI_8 NS_559 0 1.3997487969889296e-03
GC_8_560 b_8 NI_8 NS_560 0 1.9719385196850510e-03
GC_8_561 b_8 NI_8 NS_561 0 1.0457174220960381e-03
GC_8_562 b_8 NI_8 NS_562 0 -2.2988261674234353e-03
GC_8_563 b_8 NI_8 NS_563 0 -6.9831750493555068e-04
GC_8_564 b_8 NI_8 NS_564 0 -1.4663462588842982e-03
GC_8_565 b_8 NI_8 NS_565 0 -1.3735955868205236e-03
GC_8_566 b_8 NI_8 NS_566 0 -3.1257034853934335e-04
GC_8_567 b_8 NI_8 NS_567 0 6.7938416485404856e-09
GC_8_568 b_8 NI_8 NS_568 0 -2.4700008421933044e-08
GC_8_569 b_8 NI_8 NS_569 0 -4.4377025486000772e-07
GC_8_570 b_8 NI_8 NS_570 0 1.6205765284906624e-06
GC_8_571 b_8 NI_8 NS_571 0 7.9886735402679415e-03
GC_8_572 b_8 NI_8 NS_572 0 -1.6009906166401828e-03
GC_8_573 b_8 NI_8 NS_573 0 -1.2329825440157035e-08
GC_8_574 b_8 NI_8 NS_574 0 -8.8365943175808645e-07
GC_8_575 b_8 NI_8 NS_575 0 1.0714030449848763e-04
GC_8_576 b_8 NI_8 NS_576 0 -5.1251764245770735e-04
GC_8_577 b_8 NI_8 NS_577 0 -1.9321159778798245e-03
GC_8_578 b_8 NI_8 NS_578 0 -5.9631983963260346e-04
GC_8_579 b_8 NI_8 NS_579 0 2.9522606672810988e-03
GC_8_580 b_8 NI_8 NS_580 0 2.2413638503522757e-03
GC_8_581 b_8 NI_8 NS_581 0 -3.5853190594977813e-03
GC_8_582 b_8 NI_8 NS_582 0 -3.0463421382719083e-03
GC_8_583 b_8 NI_8 NS_583 0 -1.6953791407125316e-03
GC_8_584 b_8 NI_8 NS_584 0 5.8334391390102132e-03
GC_8_585 b_8 NI_8 NS_585 0 4.3284002291705736e-03
GC_8_586 b_8 NI_8 NS_586 0 -2.4949667614146062e-03
GC_8_587 b_8 NI_8 NS_587 0 -1.0252446936462651e-04
GC_8_588 b_8 NI_8 NS_588 0 -9.7511075161960906e-05
GC_8_589 b_8 NI_8 NS_589 0 -4.4595020428920577e-03
GC_8_590 b_8 NI_8 NS_590 0 -9.0945608091324605e-04
GC_8_591 b_8 NI_8 NS_591 0 9.1489028587293311e-03
GC_8_592 b_8 NI_8 NS_592 0 1.7749052989245624e-02
GC_8_593 b_8 NI_8 NS_593 0 -4.0759927667480536e-03
GC_8_594 b_8 NI_8 NS_594 0 -1.7815995532840231e-02
GC_8_595 b_8 NI_8 NS_595 0 -8.2086051829395861e-03
GC_8_596 b_8 NI_8 NS_596 0 4.1974762820242125e-03
GC_8_597 b_8 NI_8 NS_597 0 1.7045924966324344e-02
GC_8_598 b_8 NI_8 NS_598 0 -4.7587338128790482e-04
GC_8_599 b_8 NI_8 NS_599 0 -9.2871624819425552e-03
GC_8_600 b_8 NI_8 NS_600 0 -3.1746354546422903e-03
GC_8_601 b_8 NI_8 NS_601 0 -1.3650848379645064e-02
GC_8_602 b_8 NI_8 NS_602 0 2.2873425818298224e-02
GC_8_603 b_8 NI_8 NS_603 0 2.2768614588530869e-02
GC_8_604 b_8 NI_8 NS_604 0 -2.2718063915565488e-02
GC_8_605 b_8 NI_8 NS_605 0 -9.2369617939145974e-03
GC_8_606 b_8 NI_8 NS_606 0 9.4042656214467137e-04
GC_8_607 b_8 NI_8 NS_607 0 1.8496822276858445e-02
GC_8_608 b_8 NI_8 NS_608 0 6.1966535518084634e-03
GC_8_609 b_8 NI_8 NS_609 0 -9.2042288301700612e-03
GC_8_610 b_8 NI_8 NS_610 0 -9.4288118152040246e-03
GC_8_611 b_8 NI_8 NS_611 0 -9.9569355470867805e-03
GC_8_612 b_8 NI_8 NS_612 0 6.4309792448879804e-03
GC_8_613 b_8 NI_8 NS_613 0 1.6827172974898424e-02
GC_8_614 b_8 NI_8 NS_614 0 -4.8950434243086169e-03
GC_8_615 b_8 NI_8 NS_615 0 -7.2263300358190747e-03
GC_8_616 b_8 NI_8 NS_616 0 -3.3851923587831872e-03
GC_8_617 b_8 NI_8 NS_617 0 6.8657296048905189e-03
GC_8_618 b_8 NI_8 NS_618 0 1.3286490716231204e-02
GC_8_619 b_8 NI_8 NS_619 0 -1.8581881524156229e-03
GC_8_620 b_8 NI_8 NS_620 0 -1.4397044103064804e-02
GC_8_621 b_8 NI_8 NS_621 0 -4.9859100078897467e-03
GC_8_622 b_8 NI_8 NS_622 0 1.0545183375534992e-03
GC_8_623 b_8 NI_8 NS_623 0 6.0007407101891471e-03
GC_8_624 b_8 NI_8 NS_624 0 -1.1126545345625960e-03
GC_8_625 b_8 NI_8 NS_625 0 -3.4683253119726933e-03
GC_8_626 b_8 NI_8 NS_626 0 -1.0780499297880798e-03
GC_8_627 b_8 NI_8 NS_627 0 2.7173467373073912e-03
GC_8_628 b_8 NI_8 NS_628 0 -5.1095685632588728e-04
GC_8_629 b_8 NI_8 NS_629 0 -3.3053412635033852e-03
GC_8_630 b_8 NI_8 NS_630 0 -2.8885150366910208e-03
GC_8_631 b_8 NI_8 NS_631 0 2.0156340107854321e-03
GC_8_632 b_8 NI_8 NS_632 0 7.7768289509063261e-04
GC_8_633 b_8 NI_8 NS_633 0 -2.0192451153389552e-03
GC_8_634 b_8 NI_8 NS_634 0 -9.6218739425217288e-04
GC_8_635 b_8 NI_8 NS_635 0 2.1198804231868235e-03
GC_8_636 b_8 NI_8 NS_636 0 -1.4705676215802503e-03
GC_8_637 b_8 NI_8 NS_637 0 -4.1910213514362686e-03
GC_8_638 b_8 NI_8 NS_638 0 -1.8092507177228112e-03
GC_8_639 b_8 NI_8 NS_639 0 2.3672939645769807e-03
GC_8_640 b_8 NI_8 NS_640 0 -3.6739647748164003e-04
GC_8_641 b_8 NI_8 NS_641 0 -3.0199644114835412e-03
GC_8_642 b_8 NI_8 NS_642 0 4.6494721847906780e-04
GC_8_643 b_8 NI_8 NS_643 0 2.7038550448367804e-03
GC_8_644 b_8 NI_8 NS_644 0 -2.7263252341225177e-03
GC_8_645 b_8 NI_8 NS_645 0 -5.0450291902971534e-03
GC_8_646 b_8 NI_8 NS_646 0 -1.2988615164676403e-04
GC_8_647 b_8 NI_8 NS_647 0 2.4275289845173973e-03
GC_8_648 b_8 NI_8 NS_648 0 -2.1667278443055775e-03
GC_8_649 b_8 NI_8 NS_649 0 -3.2524101995323198e-03
GC_8_650 b_8 NI_8 NS_650 0 2.6001223086727374e-03
GC_8_651 b_8 NI_8 NS_651 0 1.7373702900279843e-03
GC_8_652 b_8 NI_8 NS_652 0 -4.7433399597123001e-03
GC_8_653 b_8 NI_8 NS_653 0 -3.6476875626992597e-03
GC_8_654 b_8 NI_8 NS_654 0 2.5904971150212189e-03
GC_8_655 b_8 NI_8 NS_655 0 -2.8140500630967550e-03
GC_8_656 b_8 NI_8 NS_656 0 4.0553536027748572e-03
GC_8_657 b_8 NI_8 NS_657 0 -2.3077988958867244e-04
GC_8_658 b_8 NI_8 NS_658 0 -4.1951359845090680e-03
GC_8_659 b_8 NI_8 NS_659 0 -9.8757619549949480e-06
GC_8_660 b_8 NI_8 NS_660 0 7.9025157473182216e-06
GC_8_661 b_8 NI_8 NS_661 0 -1.3634151899217524e-03
GC_8_662 b_8 NI_8 NS_662 0 3.3837800922299796e-03
GC_8_663 b_8 NI_8 NS_663 0 -9.6978191555531826e-04
GC_8_664 b_8 NI_8 NS_664 0 -4.3384320358296844e-03
GC_8_665 b_8 NI_8 NS_665 0 -1.0095576378361584e-03
GC_8_666 b_8 NI_8 NS_666 0 2.2144692442420465e-03
GC_8_667 b_8 NI_8 NS_667 0 -1.6625797627306824e-03
GC_8_668 b_8 NI_8 NS_668 0 -4.4181655732026355e-03
GC_8_669 b_8 NI_8 NS_669 0 -1.4450239250864095e-03
GC_8_670 b_8 NI_8 NS_670 0 -2.4969806516492487e-03
GC_8_671 b_8 NI_8 NS_671 0 7.8582137585162264e-04
GC_8_672 b_8 NI_8 NS_672 0 2.5922239207866972e-03
GC_8_673 b_8 NI_8 NS_673 0 -6.9658839234052242e-04
GC_8_674 b_8 NI_8 NS_674 0 2.8805416795000495e-03
GC_8_675 b_8 NI_8 NS_675 0 -1.4341252988631936e-03
GC_8_676 b_8 NI_8 NS_676 0 -2.7701138494921739e-03
GC_8_677 b_8 NI_8 NS_677 0 -1.1685605982721130e-03
GC_8_678 b_8 NI_8 NS_678 0 2.6674409195717578e-03
GC_8_679 b_8 NI_8 NS_679 0 7.8095042474608843e-04
GC_8_680 b_8 NI_8 NS_680 0 -1.8732339630854883e-03
GC_8_681 b_8 NI_8 NS_681 0 2.4009828617911146e-08
GC_8_682 b_8 NI_8 NS_682 0 -6.0310105244241711e-08
GC_8_683 b_8 NI_8 NS_683 0 -9.0615469966806918e-07
GC_8_684 b_8 NI_8 NS_684 0 3.2140038270521549e-06
GC_8_685 b_8 NI_8 NS_685 0 1.8114567005801815e-02
GC_8_686 b_8 NI_8 NS_686 0 6.7504806025154964e-03
GC_8_687 b_8 NI_8 NS_687 0 4.7185836069516976e-07
GC_8_688 b_8 NI_8 NS_688 0 1.4478151636763948e-06
GC_8_689 b_8 NI_8 NS_689 0 6.0855591005714244e-03
GC_8_690 b_8 NI_8 NS_690 0 1.8096298210349112e-03
GC_8_691 b_8 NI_8 NS_691 0 -6.0720721250795738e-03
GC_8_692 b_8 NI_8 NS_692 0 -6.1692266232205788e-04
GC_8_693 b_8 NI_8 NS_693 0 7.3059225391114381e-03
GC_8_694 b_8 NI_8 NS_694 0 -1.2857317154663782e-02
GC_8_695 b_8 NI_8 NS_695 0 8.4528484243338968e-03
GC_8_696 b_8 NI_8 NS_696 0 -2.4018652754418288e-04
GC_8_697 b_8 NI_8 NS_697 0 -9.6390501120530801e-03
GC_8_698 b_8 NI_8 NS_698 0 2.6170982247285422e-03
GC_8_699 b_8 NI_8 NS_699 0 -8.8461812087119469e-03
GC_8_700 b_8 NI_8 NS_700 0 -2.4392856975309209e-02
GC_8_701 b_8 NI_8 NS_701 0 -8.6515044653776105e-04
GC_8_702 b_8 NI_8 NS_702 0 4.1785449310926493e-03
GC_8_703 b_8 NI_8 NS_703 0 7.1897718051335798e-03
GC_8_704 b_8 NI_8 NS_704 0 -1.0341103952601766e-03
GC_8_705 b_8 NI_8 NS_705 0 -2.5138546567629309e-02
GC_8_706 b_8 NI_8 NS_706 0 4.8071402859125962e-03
GC_8_707 b_8 NI_8 NS_707 0 -1.9701012755014635e-02
GC_8_708 b_8 NI_8 NS_708 0 8.9736691668779438e-04
GC_8_709 b_8 NI_8 NS_709 0 1.0752513754578766e-02
GC_8_710 b_8 NI_8 NS_710 0 -2.7940165215852145e-03
GC_8_711 b_8 NI_8 NS_711 0 -4.8190716048252596e-03
GC_8_712 b_8 NI_8 NS_712 0 4.5027441171719258e-02
GC_8_713 b_8 NI_8 NS_713 0 -1.2658612248359759e-02
GC_8_714 b_8 NI_8 NS_714 0 -2.5617947332229969e-04
GC_8_715 b_8 NI_8 NS_715 0 1.5863284155668685e-02
GC_8_716 b_8 NI_8 NS_716 0 -4.0664340075453132e-03
GC_8_717 b_8 NI_8 NS_717 0 3.2252270959104011e-02
GC_8_718 b_8 NI_8 NS_718 0 1.8644499190453443e-02
GC_8_719 b_8 NI_8 NS_719 0 -1.2591686761975701e-02
GC_8_720 b_8 NI_8 NS_720 0 1.8230894509173965e-04
GC_8_721 b_8 NI_8 NS_721 0 1.7239482835202321e-02
GC_8_722 b_8 NI_8 NS_722 0 -3.5124406903729213e-02
GC_8_723 b_8 NI_8 NS_723 0 1.4036138781539512e-02
GC_8_724 b_8 NI_8 NS_724 0 4.7591252687124511e-03
GC_8_725 b_8 NI_8 NS_725 0 -1.4382231800877056e-02
GC_8_726 b_8 NI_8 NS_726 0 2.6524685794230554e-04
GC_8_727 b_8 NI_8 NS_727 0 -2.0118060379307190e-02
GC_8_728 b_8 NI_8 NS_728 0 -3.0219199028764330e-02
GC_8_729 b_8 NI_8 NS_729 0 1.0538956644360272e-02
GC_8_730 b_8 NI_8 NS_730 0 3.5722847305821514e-03
GC_8_731 b_8 NI_8 NS_731 0 -2.6760815132980294e-02
GC_8_732 b_8 NI_8 NS_732 0 1.1130913452571545e-02
GC_8_733 b_8 NI_8 NS_733 0 -1.4164618207772449e-02
GC_8_734 b_8 NI_8 NS_734 0 -2.5194096411398220e-03
GC_8_735 b_8 NI_8 NS_735 0 7.5549272706518667e-03
GC_8_736 b_8 NI_8 NS_736 0 1.5797729130261440e-03
GC_8_737 b_8 NI_8 NS_737 0 -8.4944731518353121e-04
GC_8_738 b_8 NI_8 NS_738 0 2.4400469191153695e-02
GC_8_739 b_8 NI_8 NS_739 0 -7.6205569716152506e-03
GC_8_740 b_8 NI_8 NS_740 0 2.8886983252414682e-04
GC_8_741 b_8 NI_8 NS_741 0 -5.5962504512421525e-04
GC_8_742 b_8 NI_8 NS_742 0 -5.5377839281866093e-03
GC_8_743 b_8 NI_8 NS_743 0 8.2746273789274325e-03
GC_8_744 b_8 NI_8 NS_744 0 7.0134928176374834e-03
GC_8_745 b_8 NI_8 NS_745 0 -7.1244355817878639e-04
GC_8_746 b_8 NI_8 NS_746 0 1.2089369788618886e-02
GC_8_747 b_8 NI_8 NS_747 0 -5.1470074791830295e-03
GC_8_748 b_8 NI_8 NS_748 0 -1.3514154647299473e-04
GC_8_749 b_8 NI_8 NS_749 0 -1.8292647115747520e-03
GC_8_750 b_8 NI_8 NS_750 0 -5.1716218544947384e-03
GC_8_751 b_8 NI_8 NS_751 0 9.2943083015114766e-03
GC_8_752 b_8 NI_8 NS_752 0 5.4122839655795073e-03
GC_8_753 b_8 NI_8 NS_753 0 3.5222729478646118e-03
GC_8_754 b_8 NI_8 NS_754 0 1.1687365551177276e-02
GC_8_755 b_8 NI_8 NS_755 0 -6.1347816103370844e-03
GC_8_756 b_8 NI_8 NS_756 0 1.4299348373071877e-03
GC_8_757 b_8 NI_8 NS_757 0 -2.8132663170310017e-03
GC_8_758 b_8 NI_8 NS_758 0 -7.3476287237787393e-03
GC_8_759 b_8 NI_8 NS_759 0 9.9612900654835329e-03
GC_8_760 b_8 NI_8 NS_760 0 3.3711728791321113e-03
GC_8_761 b_8 NI_8 NS_761 0 8.1789495854196169e-03
GC_8_762 b_8 NI_8 NS_762 0 1.0242334458720135e-02
GC_8_763 b_8 NI_8 NS_763 0 -6.9808900504393879e-03
GC_8_764 b_8 NI_8 NS_764 0 2.9381319797196896e-03
GC_8_765 b_8 NI_8 NS_765 0 -5.6228617171210716e-03
GC_8_766 b_8 NI_8 NS_766 0 -8.0957277121284713e-03
GC_8_767 b_8 NI_8 NS_767 0 9.8673412515032314e-03
GC_8_768 b_8 NI_8 NS_768 0 5.6088812580202749e-04
GC_8_769 b_8 NI_8 NS_769 0 -1.0918819997454685e-02
GC_8_770 b_8 NI_8 NS_770 0 1.2173881006687115e-02
GC_8_771 b_8 NI_8 NS_771 0 9.6705177685815370e-03
GC_8_772 b_8 NI_8 NS_772 0 5.0263989767186310e-03
GC_8_773 b_8 NI_8 NS_773 0 -1.9579885699650408e-05
GC_8_774 b_8 NI_8 NS_774 0 3.1187022397705047e-05
GC_8_775 b_8 NI_8 NS_775 0 -7.1178510223327525e-03
GC_8_776 b_8 NI_8 NS_776 0 4.4750362695304587e-03
GC_8_777 b_8 NI_8 NS_777 0 -7.6633166386158311e-03
GC_8_778 b_8 NI_8 NS_778 0 -5.3302450813859171e-03
GC_8_779 b_8 NI_8 NS_779 0 9.5222462116369335e-03
GC_8_780 b_8 NI_8 NS_780 0 -1.7152235683940242e-03
GC_8_781 b_8 NI_8 NS_781 0 1.2490636106863164e-02
GC_8_782 b_8 NI_8 NS_782 0 -1.3743942467495569e-03
GC_8_783 b_8 NI_8 NS_783 0 -5.0724955014212238e-03
GC_8_784 b_8 NI_8 NS_784 0 -2.7518977121305322e-03
GC_8_785 b_8 NI_8 NS_785 0 -2.2328721640273914e-03
GC_8_786 b_8 NI_8 NS_786 0 6.6013620628640564e-03
GC_8_787 b_8 NI_8 NS_787 0 8.9595185100321550e-03
GC_8_788 b_8 NI_8 NS_788 0 1.2929372909398451e-04
GC_8_789 b_8 NI_8 NS_789 0 1.2486921492142457e-02
GC_8_790 b_8 NI_8 NS_790 0 1.7755899763808724e-03
GC_8_791 b_8 NI_8 NS_791 0 -5.3764650581168702e-03
GC_8_792 b_8 NI_8 NS_792 0 4.1567515639541492e-03
GC_8_793 b_8 NI_8 NS_793 0 -1.8433859898151835e-03
GC_8_794 b_8 NI_8 NS_794 0 -5.6868621120399528e-03
GC_8_795 b_8 NI_8 NS_795 0 2.0787688272159232e-07
GC_8_796 b_8 NI_8 NS_796 0 -2.4509520313848799e-07
GC_8_797 b_8 NI_8 NS_797 0 -1.1507780990062321e-05
GC_8_798 b_8 NI_8 NS_798 0 1.8247329090741684e-05
GC_8_799 b_8 NI_8 NS_799 0 -1.2879661893672375e-02
GC_8_800 b_8 NI_8 NS_800 0 1.3854988955547467e-03
GC_8_801 b_8 NI_8 NS_801 0 -2.6205633593861669e-07
GC_8_802 b_8 NI_8 NS_802 0 -3.7467198181023349e-06
GC_8_803 b_8 NI_8 NS_803 0 -2.6866989055310844e-04
GC_8_804 b_8 NI_8 NS_804 0 4.6434496467886164e-04
GC_8_805 b_8 NI_8 NS_805 0 1.3324545855156662e-03
GC_8_806 b_8 NI_8 NS_806 0 5.3749686531459812e-04
GC_8_807 b_8 NI_8 NS_807 0 -2.7601218902436569e-03
GC_8_808 b_8 NI_8 NS_808 0 -8.2597386150437980e-04
GC_8_809 b_8 NI_8 NS_809 0 3.5364630190110316e-03
GC_8_810 b_8 NI_8 NS_810 0 2.5065964003169335e-03
GC_8_811 b_8 NI_8 NS_811 0 1.1567014953984948e-03
GC_8_812 b_8 NI_8 NS_812 0 -4.2275297822352590e-03
GC_8_813 b_8 NI_8 NS_813 0 -1.7809474208916719e-03
GC_8_814 b_8 NI_8 NS_814 0 2.6938537326562715e-03
GC_8_815 b_8 NI_8 NS_815 0 -3.0415845838269634e-04
GC_8_816 b_8 NI_8 NS_816 0 -1.8023605520436339e-04
GC_8_817 b_8 NI_8 NS_817 0 3.9634813471252136e-03
GC_8_818 b_8 NI_8 NS_818 0 2.8124797281994248e-04
GC_8_819 b_8 NI_8 NS_819 0 -7.5492073290123101e-03
GC_8_820 b_8 NI_8 NS_820 0 -1.3596105032114487e-02
GC_8_821 b_8 NI_8 NS_821 0 4.4801999487905477e-03
GC_8_822 b_8 NI_8 NS_822 0 1.3516145121003542e-02
GC_8_823 b_8 NI_8 NS_823 0 6.6864828442970833e-03
GC_8_824 b_8 NI_8 NS_824 0 -4.0243772389794187e-03
GC_8_825 b_8 NI_8 NS_825 0 -1.3410282976857067e-02
GC_8_826 b_8 NI_8 NS_826 0 7.8159746019269057e-04
GC_8_827 b_8 NI_8 NS_827 0 7.8563500433261272e-03
GC_8_828 b_8 NI_8 NS_828 0 1.8570145277325880e-03
GC_8_829 b_8 NI_8 NS_829 0 1.0427285557680681e-02
GC_8_830 b_8 NI_8 NS_830 0 -1.9666904344149860e-02
GC_8_831 b_8 NI_8 NS_831 0 -1.7708800298311352e-02
GC_8_832 b_8 NI_8 NS_832 0 1.9274360121931688e-02
GC_8_833 b_8 NI_8 NS_833 0 7.6729361596686351e-03
GC_8_834 b_8 NI_8 NS_834 0 -1.4539298525646338e-03
GC_8_835 b_8 NI_8 NS_835 0 -1.5685670877968981e-02
GC_8_836 b_8 NI_8 NS_836 0 -4.6645791485753684e-03
GC_8_837 b_8 NI_8 NS_837 0 8.1074614701309253e-03
GC_8_838 b_8 NI_8 NS_838 0 7.2499038698248643e-03
GC_8_839 b_8 NI_8 NS_839 0 8.0870945772520565e-03
GC_8_840 b_8 NI_8 NS_840 0 -6.0421323777580995e-03
GC_8_841 b_8 NI_8 NS_841 0 -1.3963410688590370e-02
GC_8_842 b_8 NI_8 NS_842 0 4.6523251530979472e-03
GC_8_843 b_8 NI_8 NS_843 0 6.2461630182086992e-03
GC_8_844 b_8 NI_8 NS_844 0 2.3807828503422963e-03
GC_8_845 b_8 NI_8 NS_845 0 -6.3453899443722947e-03
GC_8_846 b_8 NI_8 NS_846 0 -1.1079783746455747e-02
GC_8_847 b_8 NI_8 NS_847 0 2.1863328123657472e-03
GC_8_848 b_8 NI_8 NS_848 0 1.1948129394737579e-02
GC_8_849 b_8 NI_8 NS_849 0 4.2064703276402200e-03
GC_8_850 b_8 NI_8 NS_850 0 -1.1782772225449151e-03
GC_8_851 b_8 NI_8 NS_851 0 -4.9335527767862099e-03
GC_8_852 b_8 NI_8 NS_852 0 1.0766011735708762e-03
GC_8_853 b_8 NI_8 NS_853 0 3.0283700722119979e-03
GC_8_854 b_8 NI_8 NS_854 0 6.9130831203057322e-04
GC_8_855 b_8 NI_8 NS_855 0 -2.2217200917586262e-03
GC_8_856 b_8 NI_8 NS_856 0 5.0249262505258445e-04
GC_8_857 b_8 NI_8 NS_857 0 3.0726777265686436e-03
GC_8_858 b_8 NI_8 NS_858 0 2.2985803293225746e-03
GC_8_859 b_8 NI_8 NS_859 0 -1.5387652809854622e-03
GC_8_860 b_8 NI_8 NS_860 0 -6.6609294789864528e-04
GC_8_861 b_8 NI_8 NS_861 0 1.8890934059922553e-03
GC_8_862 b_8 NI_8 NS_862 0 6.8215091802090579e-04
GC_8_863 b_8 NI_8 NS_863 0 -1.5634721390533862e-03
GC_8_864 b_8 NI_8 NS_864 0 1.2301006580441097e-03
GC_8_865 b_8 NI_8 NS_865 0 3.9777148057030592e-03
GC_8_866 b_8 NI_8 NS_866 0 1.4029339285902298e-03
GC_8_867 b_8 NI_8 NS_867 0 -1.5582641540616048e-03
GC_8_868 b_8 NI_8 NS_868 0 7.6118044830969183e-05
GC_8_869 b_8 NI_8 NS_869 0 2.8289105703632410e-03
GC_8_870 b_8 NI_8 NS_870 0 -6.8710742116767393e-04
GC_8_871 b_8 NI_8 NS_871 0 -1.8835368104026945e-03
GC_8_872 b_8 NI_8 NS_872 0 2.0120377226579239e-03
GC_8_873 b_8 NI_8 NS_873 0 4.9081314997214973e-03
GC_8_874 b_8 NI_8 NS_874 0 -1.8224246863871897e-04
GC_8_875 b_8 NI_8 NS_875 0 -1.6649296084358578e-03
GC_8_876 b_8 NI_8 NS_876 0 9.3127546829911614e-04
GC_8_877 b_8 NI_8 NS_877 0 3.0639871877246399e-03
GC_8_878 b_8 NI_8 NS_878 0 -2.8461960120548780e-03
GC_8_879 b_8 NI_8 NS_879 0 -1.4669304700996267e-03
GC_8_880 b_8 NI_8 NS_880 0 3.2252900410869494e-03
GC_8_881 b_8 NI_8 NS_881 0 3.7966921645209827e-03
GC_8_882 b_8 NI_8 NS_882 0 -2.9822109805940984e-03
GC_8_883 b_8 NI_8 NS_883 0 -1.8554837958402789e-03
GC_8_884 b_8 NI_8 NS_884 0 -3.8335174704312676e-03
GC_8_885 b_8 NI_8 NS_885 0 -4.1823215155975898e-04
GC_8_886 b_8 NI_8 NS_886 0 2.3792558316308799e-03
GC_8_887 b_8 NI_8 NS_887 0 -1.0537744852849971e-05
GC_8_888 b_8 NI_8 NS_888 0 -2.1100618636202589e-05
GC_8_889 b_8 NI_8 NS_889 0 8.3839973512547989e-04
GC_8_890 b_8 NI_8 NS_890 0 -3.7904895272260247e-03
GC_8_891 b_8 NI_8 NS_891 0 3.3770948815916901e-04
GC_8_892 b_8 NI_8 NS_892 0 3.3559461662604284e-03
GC_8_893 b_8 NI_8 NS_893 0 1.3516061376521488e-03
GC_8_894 b_8 NI_8 NS_894 0 -2.3818220972844045e-03
GC_8_895 b_8 NI_8 NS_895 0 2.1706557714867118e-03
GC_8_896 b_8 NI_8 NS_896 0 3.3305696475383643e-03
GC_8_897 b_8 NI_8 NS_897 0 1.1698305133423109e-03
GC_8_898 b_8 NI_8 NS_898 0 2.4039647807666126e-03
GC_8_899 b_8 NI_8 NS_899 0 -8.0769436557031878e-04
GC_8_900 b_8 NI_8 NS_900 0 -1.9803395337621558e-03
GC_8_901 b_8 NI_8 NS_901 0 3.9764806952519545e-04
GC_8_902 b_8 NI_8 NS_902 0 -2.6820412711356942e-03
GC_8_903 b_8 NI_8 NS_903 0 9.8318323283865558e-04
GC_8_904 b_8 NI_8 NS_904 0 2.7477869287570482e-03
GC_8_905 b_8 NI_8 NS_905 0 1.0389080540841799e-03
GC_8_906 b_8 NI_8 NS_906 0 -2.4201775873016278e-03
GC_8_907 b_8 NI_8 NS_907 0 -1.0840508105161789e-03
GC_8_908 b_8 NI_8 NS_908 0 1.5933775231737305e-03
GC_8_909 b_8 NI_8 NS_909 0 -1.0740497992758794e-08
GC_8_910 b_8 NI_8 NS_910 0 -2.7688799863077662e-09
GC_8_911 b_8 NI_8 NS_911 0 2.2912016356077380e-06
GC_8_912 b_8 NI_8 NS_912 0 5.4762552454626479e-07
GC_8_913 b_8 NI_8 NS_913 0 -2.0263978959497164e-04
GC_8_914 b_8 NI_8 NS_914 0 -3.3244770580887213e-06
GC_8_915 b_8 NI_8 NS_915 0 1.2949514347684918e-09
GC_8_916 b_8 NI_8 NS_916 0 9.6762516394614759e-09
GC_8_917 b_8 NI_8 NS_917 0 -4.1489186934185022e-06
GC_8_918 b_8 NI_8 NS_918 0 6.1899606364191407e-06
GC_8_919 b_8 NI_8 NS_919 0 3.7984389964344715e-06
GC_8_920 b_8 NI_8 NS_920 0 -8.1732080675593972e-06
GC_8_921 b_8 NI_8 NS_921 0 2.1694994526689994e-05
GC_8_922 b_8 NI_8 NS_922 0 -8.8474234081945088e-06
GC_8_923 b_8 NI_8 NS_923 0 -2.1457575816303565e-05
GC_8_924 b_8 NI_8 NS_924 0 -1.1750497251475479e-06
GC_8_925 b_8 NI_8 NS_925 0 -2.9650349565696568e-05
GC_8_926 b_8 NI_8 NS_926 0 -2.8288020150552899e-05
GC_8_927 b_8 NI_8 NS_927 0 -5.5338663623915590e-06
GC_8_928 b_8 NI_8 NS_928 0 1.6528857182116637e-05
GC_8_929 b_8 NI_8 NS_929 0 -2.4253069455863856e-06
GC_8_930 b_8 NI_8 NS_930 0 -7.1416266789651466e-06
GC_8_931 b_8 NI_8 NS_931 0 -2.2543152931313911e-05
GC_8_932 b_8 NI_8 NS_932 0 6.0040565127403742e-06
GC_8_933 b_8 NI_8 NS_933 0 -1.8562630889099288e-04
GC_8_934 b_8 NI_8 NS_934 0 -4.4048562243151554e-05
GC_8_935 b_8 NI_8 NS_935 0 6.2607981732097084e-05
GC_8_936 b_8 NI_8 NS_936 0 1.3739430783483750e-04
GC_8_937 b_8 NI_8 NS_937 0 -3.7276502025937504e-05
GC_8_938 b_8 NI_8 NS_938 0 5.6604129431917104e-05
GC_8_939 b_8 NI_8 NS_939 0 9.5167641815725680e-05
GC_8_940 b_8 NI_8 NS_940 0 2.4608315006538429e-04
GC_8_941 b_8 NI_8 NS_941 0 7.3783611508786840e-05
GC_8_942 b_8 NI_8 NS_942 0 4.9169710703277518e-07
GC_8_943 b_8 NI_8 NS_943 0 -1.5399677886208805e-05
GC_8_944 b_8 NI_8 NS_944 0 2.6123482057269633e-04
GC_8_945 b_8 NI_8 NS_945 0 3.6434226013785947e-04
GC_8_946 b_8 NI_8 NS_946 0 -2.4310564074796038e-04
GC_8_947 b_8 NI_8 NS_947 0 6.5642862591407122e-05
GC_8_948 b_8 NI_8 NS_948 0 -2.8524093067524448e-05
GC_8_949 b_8 NI_8 NS_949 0 2.0802916538170590e-04
GC_8_950 b_8 NI_8 NS_950 0 -2.4138717484776921e-04
GC_8_951 b_8 NI_8 NS_951 0 -7.1282968464158613e-05
GC_8_952 b_8 NI_8 NS_952 0 -7.1463391602007755e-05
GC_8_953 b_8 NI_8 NS_953 0 6.4487018005666708e-05
GC_8_954 b_8 NI_8 NS_954 0 -7.5529272524564006e-05
GC_8_955 b_8 NI_8 NS_955 0 -1.7047211860671968e-04
GC_8_956 b_8 NI_8 NS_956 0 -1.8309631756382227e-04
GC_8_957 b_8 NI_8 NS_957 0 -4.8833092916089128e-05
GC_8_958 b_8 NI_8 NS_958 0 -1.9097917633156334e-05
GC_8_959 b_8 NI_8 NS_959 0 -1.4491742005655648e-04
GC_8_960 b_8 NI_8 NS_960 0 -9.5347160781365198e-05
GC_8_961 b_8 NI_8 NS_961 0 -2.7318507039288470e-05
GC_8_962 b_8 NI_8 NS_962 0 1.0360166169695989e-04
GC_8_963 b_8 NI_8 NS_963 0 -2.7242627853902513e-05
GC_8_964 b_8 NI_8 NS_964 0 1.3907339616565447e-05
GC_8_965 b_8 NI_8 NS_965 0 2.1261998392705783e-06
GC_8_966 b_8 NI_8 NS_966 0 5.0767019159586139e-05
GC_8_967 b_8 NI_8 NS_967 0 1.6811820751146959e-05
GC_8_968 b_8 NI_8 NS_968 0 -5.9722058568306759e-07
GC_8_969 b_8 NI_8 NS_969 0 1.8082668265285781e-06
GC_8_970 b_8 NI_8 NS_970 0 -1.5452703181528105e-05
GC_8_971 b_8 NI_8 NS_971 0 -1.5113316323330106e-05
GC_8_972 b_8 NI_8 NS_972 0 -1.3586603058080352e-05
GC_8_973 b_8 NI_8 NS_973 0 -1.3111587980283550e-05
GC_8_974 b_8 NI_8 NS_974 0 1.2341874062829316e-05
GC_8_975 b_8 NI_8 NS_975 0 7.7827988741129232e-06
GC_8_976 b_8 NI_8 NS_976 0 1.2547798721960272e-06
GC_8_977 b_8 NI_8 NS_977 0 -5.1388161435772339e-06
GC_8_978 b_8 NI_8 NS_978 0 -1.2683796997653751e-05
GC_8_979 b_8 NI_8 NS_979 0 -2.0805170007314526e-05
GC_8_980 b_8 NI_8 NS_980 0 -5.8763634648152639e-06
GC_8_981 b_8 NI_8 NS_981 0 1.0765921816599176e-06
GC_8_982 b_8 NI_8 NS_982 0 2.1822935208224944e-05
GC_8_983 b_8 NI_8 NS_983 0 1.2863938194178024e-05
GC_8_984 b_8 NI_8 NS_984 0 -6.8611685094012434e-06
GC_8_985 b_8 NI_8 NS_985 0 -1.7284415364374476e-05
GC_8_986 b_8 NI_8 NS_986 0 -1.5977691551219602e-05
GC_8_987 b_8 NI_8 NS_987 0 -2.7118723729779611e-05
GC_8_988 b_8 NI_8 NS_988 0 8.8182333474247121e-06
GC_8_989 b_8 NI_8 NS_989 0 2.7088817181866661e-05
GC_8_990 b_8 NI_8 NS_990 0 2.2448437556517351e-05
GC_8_991 b_8 NI_8 NS_991 0 1.0940730049857574e-05
GC_8_992 b_8 NI_8 NS_992 0 -2.1302015660056294e-05
GC_8_993 b_8 NI_8 NS_993 0 -3.0617479261810375e-05
GC_8_994 b_8 NI_8 NS_994 0 3.9079185133662579e-06
GC_8_995 b_8 NI_8 NS_995 0 -9.8041550045064697e-06
GC_8_996 b_8 NI_8 NS_996 0 3.9250454701359517e-05
GC_8_997 b_8 NI_8 NS_997 0 1.9741558437129688e-05
GC_8_998 b_8 NI_8 NS_998 0 -6.8523955460159160e-05
GC_8_999 b_8 NI_8 NS_999 0 4.3396467817959388e-05
GC_8_1000 b_8 NI_8 NS_1000 0 -1.6864135444615440e-05
GC_8_1001 b_8 NI_8 NS_1001 0 2.0643862856190492e-07
GC_8_1002 b_8 NI_8 NS_1002 0 -2.4337060907185706e-07
GC_8_1003 b_8 NI_8 NS_1003 0 -3.6341732550855647e-06
GC_8_1004 b_8 NI_8 NS_1004 0 -2.0830499348737116e-05
GC_8_1005 b_8 NI_8 NS_1005 0 -1.0493728467903484e-05
GC_8_1006 b_8 NI_8 NS_1006 0 1.6700697593232182e-05
GC_8_1007 b_8 NI_8 NS_1007 0 9.1927184657161584e-06
GC_8_1008 b_8 NI_8 NS_1008 0 3.1865117875289405e-05
GC_8_1009 b_8 NI_8 NS_1009 0 1.4275084753521822e-05
GC_8_1010 b_8 NI_8 NS_1010 0 -3.0125596276665742e-06
GC_8_1011 b_8 NI_8 NS_1011 0 -3.9047791468473868e-06
GC_8_1012 b_8 NI_8 NS_1012 0 1.2499363418251357e-05
GC_8_1013 b_8 NI_8 NS_1013 0 -1.8573493390745919e-05
GC_8_1014 b_8 NI_8 NS_1014 0 -3.6270077995313427e-06
GC_8_1015 b_8 NI_8 NS_1015 0 1.3215675947501705e-05
GC_8_1016 b_8 NI_8 NS_1016 0 1.3176842436105989e-05
GC_8_1017 b_8 NI_8 NS_1017 0 7.6359154068555492e-06
GC_8_1018 b_8 NI_8 NS_1018 0 -2.3019061748253623e-05
GC_8_1019 b_8 NI_8 NS_1019 0 -3.8460161729591072e-06
GC_8_1020 b_8 NI_8 NS_1020 0 -1.1722919458781826e-05
GC_8_1021 b_8 NI_8 NS_1021 0 -8.7362188733566225e-06
GC_8_1022 b_8 NI_8 NS_1022 0 -2.6278895744239882e-06
GC_8_1023 b_8 NI_8 NS_1023 0 5.5142537620782349e-10
GC_8_1024 b_8 NI_8 NS_1024 0 2.9347519149004545e-10
GC_8_1025 b_8 NI_8 NS_1025 0 4.2109510425955247e-08
GC_8_1026 b_8 NI_8 NS_1026 0 3.6939225733299100e-08
GC_8_1027 b_8 NI_8 NS_1027 0 2.8654995698615496e-04
GC_8_1028 b_8 NI_8 NS_1028 0 -1.4350321387929055e-05
GC_8_1029 b_8 NI_8 NS_1029 0 -1.2377044728537847e-09
GC_8_1030 b_8 NI_8 NS_1030 0 -1.9231747111375378e-08
GC_8_1031 b_8 NI_8 NS_1031 0 2.6665543881225675e-06
GC_8_1032 b_8 NI_8 NS_1032 0 -3.8232153812273274e-06
GC_8_1033 b_8 NI_8 NS_1033 0 -1.3223098695309602e-05
GC_8_1034 b_8 NI_8 NS_1034 0 -5.0242656034074541e-07
GC_8_1035 b_8 NI_8 NS_1035 0 3.9458280946503665e-05
GC_8_1036 b_8 NI_8 NS_1036 0 2.7880676543603577e-06
GC_8_1037 b_8 NI_8 NS_1037 0 -4.1775291701129227e-05
GC_8_1038 b_8 NI_8 NS_1038 0 -2.3733018972232800e-05
GC_8_1039 b_8 NI_8 NS_1039 0 1.7634788560392442e-06
GC_8_1040 b_8 NI_8 NS_1040 0 4.4845308389430388e-05
GC_8_1041 b_8 NI_8 NS_1041 0 1.4501520867389134e-05
GC_8_1042 b_8 NI_8 NS_1042 0 -4.8185833736733671e-05
GC_8_1043 b_8 NI_8 NS_1043 0 1.9359368719542762e-06
GC_8_1044 b_8 NI_8 NS_1044 0 5.6539835963371172e-06
GC_8_1045 b_8 NI_8 NS_1045 0 -4.4994174966999991e-05
GC_8_1046 b_8 NI_8 NS_1046 0 1.5684404230233881e-06
GC_8_1047 b_8 NI_8 NS_1047 0 1.0310756940268780e-04
GC_8_1048 b_8 NI_8 NS_1048 0 1.2335556499039102e-04
GC_8_1049 b_8 NI_8 NS_1049 0 -7.5525462111720085e-05
GC_8_1050 b_8 NI_8 NS_1050 0 -1.3698528309213142e-04
GC_8_1051 b_8 NI_8 NS_1051 0 -6.7109340518288558e-05
GC_8_1052 b_8 NI_8 NS_1052 0 4.9269291354921667e-05
GC_8_1053 b_8 NI_8 NS_1053 0 1.3517087394796109e-04
GC_8_1054 b_8 NI_8 NS_1054 0 -2.8537419852872702e-05
GC_8_1055 b_8 NI_8 NS_1055 0 -8.7330926140934348e-05
GC_8_1056 b_8 NI_8 NS_1056 0 -1.1763161500026704e-05
GC_8_1057 b_8 NI_8 NS_1057 0 -9.4647115795001087e-05
GC_8_1058 b_8 NI_8 NS_1058 0 2.1148781098384706e-04
GC_8_1059 b_8 NI_8 NS_1059 0 1.6429617485191900e-04
GC_8_1060 b_8 NI_8 NS_1060 0 -2.1487400993235053e-04
GC_8_1061 b_8 NI_8 NS_1061 0 -8.1684433961676421e-05
GC_8_1062 b_8 NI_8 NS_1062 0 1.9189092970388975e-05
GC_8_1063 b_8 NI_8 NS_1063 0 1.6096905530590838e-04
GC_8_1064 b_8 NI_8 NS_1064 0 4.2091213339643925e-05
GC_8_1065 b_8 NI_8 NS_1065 0 -8.8878044917091814e-05
GC_8_1066 b_8 NI_8 NS_1066 0 -7.1909596345738475e-05
GC_8_1067 b_8 NI_8 NS_1067 0 -8.4867036666413123e-05
GC_8_1068 b_8 NI_8 NS_1068 0 6.3596360809027260e-05
GC_8_1069 b_8 NI_8 NS_1069 0 1.4068805365759842e-04
GC_8_1070 b_8 NI_8 NS_1070 0 -4.8518768468088255e-05
GC_8_1071 b_8 NI_8 NS_1071 0 -6.6207483136975493e-05
GC_8_1072 b_8 NI_8 NS_1072 0 -2.4250999834822550e-05
GC_8_1073 b_8 NI_8 NS_1073 0 6.1223508913151292e-05
GC_8_1074 b_8 NI_8 NS_1074 0 1.1375862030114167e-04
GC_8_1075 b_8 NI_8 NS_1075 0 -2.2917088757141184e-05
GC_8_1076 b_8 NI_8 NS_1076 0 -1.2153227375113717e-04
GC_8_1077 b_8 NI_8 NS_1077 0 -4.4313564863393921e-05
GC_8_1078 b_8 NI_8 NS_1078 0 1.0975035201206493e-05
GC_8_1079 b_8 NI_8 NS_1079 0 4.7535486310875600e-05
GC_8_1080 b_8 NI_8 NS_1080 0 -1.0607214547266121e-05
GC_8_1081 b_8 NI_8 NS_1081 0 -3.2085902565533673e-05
GC_8_1082 b_8 NI_8 NS_1082 0 -7.6432278987721291e-06
GC_8_1083 b_8 NI_8 NS_1083 0 2.1333531471393259e-05
GC_8_1084 b_8 NI_8 NS_1084 0 -4.8743867331635505e-06
GC_8_1085 b_8 NI_8 NS_1085 0 -3.2213590322390706e-05
GC_8_1086 b_8 NI_8 NS_1086 0 -2.5250789823510624e-05
GC_8_1087 b_8 NI_8 NS_1087 0 1.2710109989460640e-05
GC_8_1088 b_8 NI_8 NS_1088 0 6.1771582786577833e-06
GC_8_1089 b_8 NI_8 NS_1089 0 -2.0359017708097009e-05
GC_8_1090 b_8 NI_8 NS_1090 0 -7.7253059720013616e-06
GC_8_1091 b_8 NI_8 NS_1091 0 1.4086578557226464e-05
GC_8_1092 b_8 NI_8 NS_1092 0 -1.2504410484793152e-05
GC_8_1093 b_8 NI_8 NS_1093 0 -4.1282285724556979e-05
GC_8_1094 b_8 NI_8 NS_1094 0 -1.6953796465321113e-05
GC_8_1095 b_8 NI_8 NS_1095 0 1.1907503991685504e-05
GC_8_1096 b_8 NI_8 NS_1096 0 -1.7646397811920671e-06
GC_8_1097 b_8 NI_8 NS_1097 0 -3.0212458392454516e-05
GC_8_1098 b_8 NI_8 NS_1098 0 5.5333503025385340e-06
GC_8_1099 b_8 NI_8 NS_1099 0 1.6332647742549352e-05
GC_8_1100 b_8 NI_8 NS_1100 0 -2.0848592978186665e-05
GC_8_1101 b_8 NI_8 NS_1101 0 -4.9846288356704498e-05
GC_8_1102 b_8 NI_8 NS_1102 0 -1.6673747788869696e-06
GC_8_1103 b_8 NI_8 NS_1103 0 1.2247659390690761e-05
GC_8_1104 b_8 NI_8 NS_1104 0 -1.1717555102861194e-05
GC_8_1105 b_8 NI_8 NS_1105 0 -3.1908583761631001e-05
GC_8_1106 b_8 NI_8 NS_1106 0 2.5076450436115475e-05
GC_8_1107 b_8 NI_8 NS_1107 0 1.0834703177704058e-05
GC_8_1108 b_8 NI_8 NS_1108 0 -3.6496291435002898e-05
GC_8_1109 b_8 NI_8 NS_1109 0 -3.3856382108538925e-05
GC_8_1110 b_8 NI_8 NS_1110 0 1.8659163397347846e-05
GC_8_1111 b_8 NI_8 NS_1111 0 -5.9880020774058210e-05
GC_8_1112 b_8 NI_8 NS_1112 0 1.2847674757906813e-04
GC_8_1113 b_8 NI_8 NS_1113 0 -1.4511897522659640e-05
GC_8_1114 b_8 NI_8 NS_1114 0 -3.3369944397924357e-05
GC_8_1115 b_8 NI_8 NS_1115 0 -3.8791639206730819e-07
GC_8_1116 b_8 NI_8 NS_1116 0 3.6149793850014854e-07
GC_8_1117 b_8 NI_8 NS_1117 0 -1.9685611879734677e-05
GC_8_1118 b_8 NI_8 NS_1118 0 3.1289659838221054e-05
GC_8_1119 b_8 NI_8 NS_1119 0 -1.4243119455904397e-05
GC_8_1120 b_8 NI_8 NS_1120 0 -3.4196322991136830e-05
GC_8_1121 b_8 NI_8 NS_1121 0 -5.2921625695160794e-06
GC_8_1122 b_8 NI_8 NS_1122 0 5.5312271491263271e-06
GC_8_1123 b_8 NI_8 NS_1123 0 -1.9744697329038625e-05
GC_8_1124 b_8 NI_8 NS_1124 0 -6.5467807952850540e-05
GC_8_1125 b_8 NI_8 NS_1125 0 -9.2827090506347975e-06
GC_8_1126 b_8 NI_8 NS_1126 0 -2.0586529693136940e-05
GC_8_1127 b_8 NI_8 NS_1127 0 1.4777871120015963e-05
GC_8_1128 b_8 NI_8 NS_1128 0 2.2998461966872429e-05
GC_8_1129 b_8 NI_8 NS_1129 0 -6.8230585923624628e-06
GC_8_1130 b_8 NI_8 NS_1130 0 2.7592666584731985e-05
GC_8_1131 b_8 NI_8 NS_1131 0 -1.1135794100712403e-05
GC_8_1132 b_8 NI_8 NS_1132 0 -2.1577734007364729e-05
GC_8_1133 b_8 NI_8 NS_1133 0 -1.1024480342705268e-05
GC_8_1134 b_8 NI_8 NS_1134 0 2.3799332207989203e-05
GC_8_1135 b_8 NI_8 NS_1135 0 5.1499148640833058e-06
GC_8_1136 b_8 NI_8 NS_1136 0 -1.5352049697044919e-05
GC_8_1137 b_8 NI_8 NS_1137 0 -4.7264158081685744e-10
GC_8_1138 b_8 NI_8 NS_1138 0 -9.1861920799933504e-10
GC_8_1139 b_8 NI_8 NS_1139 0 -5.5411894674668220e-08
GC_8_1140 b_8 NI_8 NS_1140 0 7.6386876647011339e-09
GC_8_1141 b_8 NI_8 NS_1141 0 -3.7756391871103982e-05
GC_8_1142 b_8 NI_8 NS_1142 0 2.2260817075739207e-06
GC_8_1143 b_8 NI_8 NS_1143 0 6.0497149223470972e-11
GC_8_1144 b_8 NI_8 NS_1144 0 3.0748226804822342e-09
GC_8_1145 b_8 NI_8 NS_1145 0 -1.9312553788781967e-06
GC_8_1146 b_8 NI_8 NS_1146 0 -1.7210839038780306e-06
GC_8_1147 b_8 NI_8 NS_1147 0 -5.6039610010442510e-06
GC_8_1148 b_8 NI_8 NS_1148 0 2.9249093454314825e-06
GC_8_1149 b_8 NI_8 NS_1149 0 -1.6662516292489261e-05
GC_8_1150 b_8 NI_8 NS_1150 0 1.9136220370374334e-05
GC_8_1151 b_8 NI_8 NS_1151 0 1.5401881014966517e-05
GC_8_1152 b_8 NI_8 NS_1152 0 1.0211461398455346e-05
GC_8_1153 b_8 NI_8 NS_1153 0 1.7356900880623746e-05
GC_8_1154 b_8 NI_8 NS_1154 0 2.3278497621310958e-05
GC_8_1155 b_8 NI_8 NS_1155 0 3.0897957746955270e-05
GC_8_1156 b_8 NI_8 NS_1156 0 5.3455189796430821e-06
GC_8_1157 b_8 NI_8 NS_1157 0 -3.3855510187371696e-06
GC_8_1158 b_8 NI_8 NS_1158 0 -2.1457354663976872e-06
GC_8_1159 b_8 NI_8 NS_1159 0 1.7191263830246175e-05
GC_8_1160 b_8 NI_8 NS_1160 0 -2.2223426361086429e-06
GC_8_1161 b_8 NI_8 NS_1161 0 1.2979417142367240e-04
GC_8_1162 b_8 NI_8 NS_1162 0 3.5245573480030410e-05
GC_8_1163 b_8 NI_8 NS_1163 0 -2.8533563717444207e-05
GC_8_1164 b_8 NI_8 NS_1164 0 -9.9832745627814417e-05
GC_8_1165 b_8 NI_8 NS_1165 0 2.5236941474946682e-05
GC_8_1166 b_8 NI_8 NS_1166 0 -3.1267144760796609e-05
GC_8_1167 b_8 NI_8 NS_1167 0 -4.0931240468894415e-05
GC_8_1168 b_8 NI_8 NS_1168 0 -1.6750291936513058e-04
GC_8_1169 b_8 NI_8 NS_1169 0 -4.1821888622372055e-05
GC_8_1170 b_8 NI_8 NS_1170 0 -5.3846160829576467e-06
GC_8_1171 b_8 NI_8 NS_1171 0 2.2549193408801328e-05
GC_8_1172 b_8 NI_8 NS_1172 0 -1.5152140035318152e-04
GC_8_1173 b_8 NI_8 NS_1173 0 -2.3148655017453344e-04
GC_8_1174 b_8 NI_8 NS_1174 0 1.1299995515101988e-04
GC_8_1175 b_8 NI_8 NS_1175 0 -3.7411587434928932e-05
GC_8_1176 b_8 NI_8 NS_1176 0 1.3952381998874301e-05
GC_8_1177 b_8 NI_8 NS_1177 0 -1.3781859765216794e-04
GC_8_1178 b_8 NI_8 NS_1178 0 1.2973527900085770e-04
GC_8_1179 b_8 NI_8 NS_1179 0 3.6132290534197814e-05
GC_8_1180 b_8 NI_8 NS_1180 0 4.1461477430130405e-05
GC_8_1181 b_8 NI_8 NS_1181 0 -3.8173872362586758e-05
GC_8_1182 b_8 NI_8 NS_1182 0 4.2971182494963476e-05
GC_8_1183 b_8 NI_8 NS_1183 0 8.7354662017498076e-05
GC_8_1184 b_8 NI_8 NS_1184 0 1.1821532104391714e-04
GC_8_1185 b_8 NI_8 NS_1185 0 2.7245014195505222e-05
GC_8_1186 b_8 NI_8 NS_1186 0 1.0262329164276097e-05
GC_8_1187 b_8 NI_8 NS_1187 0 8.7158310875612275e-05
GC_8_1188 b_8 NI_8 NS_1188 0 6.5380985997332623e-05
GC_8_1189 b_8 NI_8 NS_1189 0 2.0400950361572127e-05
GC_8_1190 b_8 NI_8 NS_1190 0 -5.7168781413733753e-05
GC_8_1191 b_8 NI_8 NS_1191 0 1.7001878493688136e-05
GC_8_1192 b_8 NI_8 NS_1192 0 -8.8439669638912617e-06
GC_8_1193 b_8 NI_8 NS_1193 0 8.4707453697210840e-06
GC_8_1194 b_8 NI_8 NS_1194 0 -3.3126325394680921e-05
GC_8_1195 b_8 NI_8 NS_1195 0 -8.8428601452833150e-06
GC_8_1196 b_8 NI_8 NS_1196 0 4.1505779436667061e-07
GC_8_1197 b_8 NI_8 NS_1197 0 -2.4022625298636524e-06
GC_8_1198 b_8 NI_8 NS_1198 0 8.4362264964340588e-06
GC_8_1199 b_8 NI_8 NS_1199 0 1.0207782696765641e-05
GC_8_1200 b_8 NI_8 NS_1200 0 6.0582490740494106e-06
GC_8_1201 b_8 NI_8 NS_1201 0 1.2154867902044382e-05
GC_8_1202 b_8 NI_8 NS_1202 0 -7.9359206600484449e-06
GC_8_1203 b_8 NI_8 NS_1203 0 -3.4649718930736680e-06
GC_8_1204 b_8 NI_8 NS_1204 0 -5.2258141259734934e-07
GC_8_1205 b_8 NI_8 NS_1205 0 2.5132155698399814e-06
GC_8_1206 b_8 NI_8 NS_1206 0 7.3270775928101046e-06
GC_8_1207 b_8 NI_8 NS_1207 0 1.3691636060807475e-05
GC_8_1208 b_8 NI_8 NS_1208 0 2.6181825641814769e-06
GC_8_1209 b_8 NI_8 NS_1209 0 4.5508831592651572e-06
GC_8_1210 b_8 NI_8 NS_1210 0 -1.4312547741740658e-05
GC_8_1211 b_8 NI_8 NS_1211 0 -5.8920327246913536e-06
GC_8_1212 b_8 NI_8 NS_1212 0 4.1741261851831963e-06
GC_8_1213 b_8 NI_8 NS_1213 0 1.0370350850772177e-05
GC_8_1214 b_8 NI_8 NS_1214 0 9.8155496072678491e-06
GC_8_1215 b_8 NI_8 NS_1215 0 1.7399257289212665e-05
GC_8_1216 b_8 NI_8 NS_1216 0 -4.2746276365949648e-06
GC_8_1217 b_8 NI_8 NS_1217 0 -9.2261139275781287e-06
GC_8_1218 b_8 NI_8 NS_1218 0 -1.5489745384488846e-05
GC_8_1219 b_8 NI_8 NS_1219 0 -4.0027773149285502e-06
GC_8_1220 b_8 NI_8 NS_1220 0 1.3420164125150623e-05
GC_8_1221 b_8 NI_8 NS_1221 0 2.1008731990474588e-05
GC_8_1222 b_8 NI_8 NS_1222 0 -7.6329687167041995e-07
GC_8_1223 b_8 NI_8 NS_1223 0 9.1216893504250140e-06
GC_8_1224 b_8 NI_8 NS_1224 0 -1.7455303668587114e-05
GC_8_1225 b_8 NI_8 NS_1225 0 1.4592429711582379e-06
GC_8_1226 b_8 NI_8 NS_1226 0 -1.4427431703523901e-05
GC_8_1227 b_8 NI_8 NS_1227 0 -1.3809057314624412e-05
GC_8_1228 b_8 NI_8 NS_1228 0 3.9888871008426278e-06
GC_8_1229 b_8 NI_8 NS_1229 0 9.7996655669670197e-09
GC_8_1230 b_8 NI_8 NS_1230 0 -4.8130847716981762e-08
GC_8_1231 b_8 NI_8 NS_1231 0 8.6298604282273227e-06
GC_8_1232 b_8 NI_8 NS_1232 0 1.1373623758222542e-05
GC_8_1233 b_8 NI_8 NS_1233 0 1.0873521995687701e-05
GC_8_1234 b_8 NI_8 NS_1234 0 -1.1464211290275302e-05
GC_8_1235 b_8 NI_8 NS_1235 0 -3.5307947619133511e-06
GC_8_1236 b_8 NI_8 NS_1236 0 -1.0164884438304782e-05
GC_8_1237 b_8 NI_8 NS_1237 0 -2.0125585453491757e-06
GC_8_1238 b_8 NI_8 NS_1238 0 1.2870550434852327e-05
GC_8_1239 b_8 NI_8 NS_1239 0 9.7604671977918774e-07
GC_8_1240 b_8 NI_8 NS_1240 0 -7.2620465123909737e-06
GC_8_1241 b_8 NI_8 NS_1241 0 7.4715658936411900e-06
GC_8_1242 b_8 NI_8 NS_1242 0 1.7440199310608921e-06
GC_8_1243 b_8 NI_8 NS_1243 0 -6.1165637470310682e-06
GC_8_1244 b_8 NI_8 NS_1244 0 -8.8986432282096503e-06
GC_8_1245 b_8 NI_8 NS_1245 0 -4.1366754343019081e-06
GC_8_1246 b_8 NI_8 NS_1246 0 9.6568905634304888e-06
GC_8_1247 b_8 NI_8 NS_1247 0 3.3152497347851341e-06
GC_8_1248 b_8 NI_8 NS_1248 0 6.0578125844080528e-06
GC_8_1249 b_8 NI_8 NS_1249 0 5.7049765271323486e-06
GC_8_1250 b_8 NI_8 NS_1250 0 5.2024817074559932e-07
GC_8_1251 b_8 NI_8 NS_1251 0 5.9119923053433540e-11
GC_8_1252 b_8 NI_8 NS_1252 0 1.4784982398809792e-10
GC_8_1253 b_8 NI_8 NS_1253 0 5.9030987044447657e-09
GC_8_1254 b_8 NI_8 NS_1254 0 -8.4602316835034514e-09
GC_8_1255 b_8 NI_8 NS_1255 0 -1.1277210571164117e-04
GC_8_1256 b_8 NI_8 NS_1256 0 -2.1518465391430158e-06
GC_8_1257 b_8 NI_8 NS_1257 0 -2.4613967138594873e-10
GC_8_1258 b_8 NI_8 NS_1258 0 2.5681352464362858e-09
GC_8_1259 b_8 NI_8 NS_1259 0 1.7816033195415925e-06
GC_8_1260 b_8 NI_8 NS_1260 0 -1.5815620934369930e-06
GC_8_1261 b_8 NI_8 NS_1261 0 2.3533685098906571e-07
GC_8_1262 b_8 NI_8 NS_1262 0 -6.4013236614646681e-06
GC_8_1263 b_8 NI_8 NS_1263 0 -7.4872987811586628e-06
GC_8_1264 b_8 NI_8 NS_1264 0 -2.0463961889487827e-07
GC_8_1265 b_8 NI_8 NS_1265 0 -1.3991987584388467e-06
GC_8_1266 b_8 NI_8 NS_1266 0 -4.6879150878122451e-06
GC_8_1267 b_8 NI_8 NS_1267 0 -1.5829941643410426e-05
GC_8_1268 b_8 NI_8 NS_1268 0 -1.8864567049861178e-06
GC_8_1269 b_8 NI_8 NS_1269 0 -6.8244337422190106e-06
GC_8_1270 b_8 NI_8 NS_1270 0 1.8864266590807079e-05
GC_8_1271 b_8 NI_8 NS_1271 0 4.8188264980690278e-06
GC_8_1272 b_8 NI_8 NS_1272 0 -2.8796975156571342e-06
GC_8_1273 b_8 NI_8 NS_1273 0 -1.3563216791106904e-07
GC_8_1274 b_8 NI_8 NS_1274 0 -2.4716414690498366e-06
GC_8_1275 b_8 NI_8 NS_1275 0 -2.6117097750493078e-05
GC_8_1276 b_8 NI_8 NS_1276 0 2.8150832255690094e-05
GC_8_1277 b_8 NI_8 NS_1277 0 2.8021136231863245e-05
GC_8_1278 b_8 NI_8 NS_1278 0 -8.1067139245559339e-06
GC_8_1279 b_8 NI_8 NS_1279 0 -8.0870808053768235e-06
GC_8_1280 b_8 NI_8 NS_1280 0 -4.2194541638630087e-06
GC_8_1281 b_8 NI_8 NS_1281 0 1.2345315656051745e-05
GC_8_1282 b_8 NI_8 NS_1282 0 2.7049491894651860e-05
GC_8_1283 b_8 NI_8 NS_1283 0 1.4325014300217808e-06
GC_8_1284 b_8 NI_8 NS_1284 0 -8.8303089192727698e-06
GC_8_1285 b_8 NI_8 NS_1285 0 -2.8319562928779509e-05
GC_8_1286 b_8 NI_8 NS_1286 0 4.8085423178444807e-06
GC_8_1287 b_8 NI_8 NS_1287 0 4.1184590059823326e-05
GC_8_1288 b_8 NI_8 NS_1288 0 1.0835845381587623e-05
GC_8_1289 b_8 NI_8 NS_1289 0 -3.0015681861006591e-06
GC_8_1290 b_8 NI_8 NS_1290 0 -4.3670101579512199e-06
GC_8_1291 b_8 NI_8 NS_1291 0 1.2955898723477088e-05
GC_8_1292 b_8 NI_8 NS_1292 0 1.9080714701910552e-05
GC_8_1293 b_8 NI_8 NS_1293 0 3.7635943990905342e-06
GC_8_1294 b_8 NI_8 NS_1294 0 -1.0833681912729364e-05
GC_8_1295 b_8 NI_8 NS_1295 0 -6.4466352983320422e-06
GC_8_1296 b_8 NI_8 NS_1296 0 9.6349171493023189e-07
GC_8_1297 b_8 NI_8 NS_1297 0 1.8926188289802662e-05
GC_8_1298 b_8 NI_8 NS_1298 0 5.4714303584915011e-06
GC_8_1299 b_8 NI_8 NS_1299 0 -1.1342488410580564e-07
GC_8_1300 b_8 NI_8 NS_1300 0 -4.1223382492154442e-06
GC_8_1301 b_8 NI_8 NS_1301 0 4.9483402453835254e-06
GC_8_1302 b_8 NI_8 NS_1302 0 1.4379801008978800e-05
GC_8_1303 b_8 NI_8 NS_1303 0 7.7968519737610811e-06
GC_8_1304 b_8 NI_8 NS_1304 0 -1.1164421203486066e-05
GC_8_1305 b_8 NI_8 NS_1305 0 -1.4154739430628652e-06
GC_8_1306 b_8 NI_8 NS_1306 0 9.8362926384220544e-07
GC_8_1307 b_8 NI_8 NS_1307 0 1.0884949636821620e-05
GC_8_1308 b_8 NI_8 NS_1308 0 4.1621731883249348e-06
GC_8_1309 b_8 NI_8 NS_1309 0 1.6970822711982690e-06
GC_8_1310 b_8 NI_8 NS_1310 0 -5.9090571147146150e-07
GC_8_1311 b_8 NI_8 NS_1311 0 5.6760840621048531e-06
GC_8_1312 b_8 NI_8 NS_1312 0 1.7180060549263473e-06
GC_8_1313 b_8 NI_8 NS_1313 0 3.3604894116279094e-06
GC_8_1314 b_8 NI_8 NS_1314 0 2.0717604943095358e-06
GC_8_1315 b_8 NI_8 NS_1315 0 1.0946296522207245e-05
GC_8_1316 b_8 NI_8 NS_1316 0 3.8300822011537315e-06
GC_8_1317 b_8 NI_8 NS_1317 0 4.8385991636535200e-06
GC_8_1318 b_8 NI_8 NS_1318 0 -5.2549255875003505e-08
GC_8_1319 b_8 NI_8 NS_1319 0 9.9675844057918320e-06
GC_8_1320 b_8 NI_8 NS_1320 0 -1.0598260901373119e-06
GC_8_1321 b_8 NI_8 NS_1321 0 8.2081792726570390e-06
GC_8_1322 b_8 NI_8 NS_1322 0 2.9740305938449879e-06
GC_8_1323 b_8 NI_8 NS_1323 0 1.9026488801342413e-05
GC_8_1324 b_8 NI_8 NS_1324 0 -5.5233826700775598e-06
GC_8_1325 b_8 NI_8 NS_1325 0 7.1917045387677425e-06
GC_8_1326 b_8 NI_8 NS_1326 0 -3.9943585183203122e-06
GC_8_1327 b_8 NI_8 NS_1327 0 1.3712813829442569e-05
GC_8_1328 b_8 NI_8 NS_1328 0 -1.1879978991914875e-05
GC_8_1329 b_8 NI_8 NS_1329 0 1.2365923659688710e-05
GC_8_1330 b_8 NI_8 NS_1330 0 -3.9393634434835419e-06
GC_8_1331 b_8 NI_8 NS_1331 0 9.1636805235329453e-06
GC_8_1332 b_8 NI_8 NS_1332 0 -2.6747063145897131e-05
GC_8_1333 b_8 NI_8 NS_1333 0 2.3618350267170941e-06
GC_8_1334 b_8 NI_8 NS_1334 0 -1.2358489071141205e-05
GC_8_1335 b_8 NI_8 NS_1335 0 -8.2831501532549523e-06
GC_8_1336 b_8 NI_8 NS_1336 0 -1.8645470554644219e-05
GC_8_1337 b_8 NI_8 NS_1337 0 -4.8702697771926353e-06
GC_8_1338 b_8 NI_8 NS_1338 0 -1.2077489762471531e-05
GC_8_1339 b_8 NI_8 NS_1339 0 5.4674641234461239e-05
GC_8_1340 b_8 NI_8 NS_1340 0 -8.8166250192615536e-05
GC_8_1341 b_8 NI_8 NS_1341 0 -1.0018834925856701e-05
GC_8_1342 b_8 NI_8 NS_1342 0 1.2701493750540271e-06
GC_8_1343 b_8 NI_8 NS_1343 0 3.8983285761869105e-07
GC_8_1344 b_8 NI_8 NS_1344 0 -1.2677289880177168e-07
GC_8_1345 b_8 NI_8 NS_1345 0 -2.7052832013480451e-06
GC_8_1346 b_8 NI_8 NS_1346 0 -1.9795986780020301e-06
GC_8_1347 b_8 NI_8 NS_1347 0 -4.4027981764321661e-06
GC_8_1348 b_8 NI_8 NS_1348 0 5.4784792973552464e-07
GC_8_1349 b_8 NI_8 NS_1349 0 -1.7423549724911309e-05
GC_8_1350 b_8 NI_8 NS_1350 0 9.5920509430284303e-06
GC_8_1351 b_8 NI_8 NS_1351 0 -9.1285279011593974e-06
GC_8_1352 b_8 NI_8 NS_1352 0 3.7355109248173222e-05
GC_8_1353 b_8 NI_8 NS_1353 0 -7.2451099212066974e-06
GC_8_1354 b_8 NI_8 NS_1354 0 3.3527615753167200e-07
GC_8_1355 b_8 NI_8 NS_1355 0 -1.3395935016514739e-05
GC_8_1356 b_8 NI_8 NS_1356 0 1.8751237910408046e-06
GC_8_1357 b_8 NI_8 NS_1357 0 -4.6442423183911403e-06
GC_8_1358 b_8 NI_8 NS_1358 0 -3.3978549498137963e-06
GC_8_1359 b_8 NI_8 NS_1359 0 -6.4046490468495180e-06
GC_8_1360 b_8 NI_8 NS_1360 0 1.0361836058757347e-06
GC_8_1361 b_8 NI_8 NS_1361 0 -3.0540566734107449e-06
GC_8_1362 b_8 NI_8 NS_1362 0 8.8642146114897057e-07
GC_8_1363 b_8 NI_8 NS_1363 0 -1.7952292829302740e-06
GC_8_1364 b_8 NI_8 NS_1364 0 -9.3643236874938301e-07
GC_8_1365 b_8 NI_8 NS_1365 0 -2.6050215081606893e-10
GC_8_1366 b_8 NI_8 NS_1366 0 4.2261538496435519e-10
GC_8_1367 b_8 NI_8 NS_1367 0 2.3349527041952712e-09
GC_8_1368 b_8 NI_8 NS_1368 0 -2.6679273514400198e-08
GD_8_1 b_8 NI_8 NA_1 0 1.0048973518774349e-05
GD_8_2 b_8 NI_8 NA_2 0 -3.6554694745798796e-06
GD_8_3 b_8 NI_8 NA_3 0 1.1836175979128544e-06
GD_8_4 b_8 NI_8 NA_4 0 3.4014534725073670e-06
GD_8_5 b_8 NI_8 NA_5 0 5.8609049333635207e-04
GD_8_6 b_8 NI_8 NA_6 0 1.2979344857305277e-02
GD_8_7 b_8 NI_8 NA_7 0 -4.2218420257787055e-03
GD_8_8 b_8 NI_8 NA_8 0 -8.8807956671788472e-03
GD_8_9 b_8 NI_8 NA_9 0 2.6580147436795455e-05
GD_8_10 b_8 NI_8 NA_10 0 1.0377146040001880e-04
GD_8_11 b_8 NI_8 NA_11 0 2.4542719891741668e-06
GD_8_12 b_8 NI_8 NA_12 0 4.1424656148419589e-06
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 1.3443288105640183e-05
GC_9_2 b_9 NI_9 NS_2 0 -5.8799870897186008e-08
GC_9_3 b_9 NI_9 NS_3 0 -1.4953997577932542e-11
GC_9_4 b_9 NI_9 NS_4 0 1.3605229700660727e-10
GC_9_5 b_9 NI_9 NS_5 0 3.6053355832456307e-07
GC_9_6 b_9 NI_9 NS_6 0 -1.8115037978823280e-07
GC_9_7 b_9 NI_9 NS_7 0 2.8267807135251116e-07
GC_9_8 b_9 NI_9 NS_8 0 -3.5350016201938407e-07
GC_9_9 b_9 NI_9 NS_9 0 4.9947343648778873e-07
GC_9_10 b_9 NI_9 NS_10 0 -1.4260700516352356e-06
GC_9_11 b_9 NI_9 NS_11 0 -1.1620830464528767e-06
GC_9_12 b_9 NI_9 NS_12 0 -4.7166457270345969e-07
GC_9_13 b_9 NI_9 NS_13 0 -3.4835190386945136e-07
GC_9_14 b_9 NI_9 NS_14 0 -6.2923198620062392e-07
GC_9_15 b_9 NI_9 NS_15 0 -2.5926061590113599e-06
GC_9_16 b_9 NI_9 NS_16 0 -6.4982327807015144e-07
GC_9_17 b_9 NI_9 NS_17 0 7.1999379628723664e-07
GC_9_18 b_9 NI_9 NS_18 0 3.6092310204909843e-07
GC_9_19 b_9 NI_9 NS_19 0 -7.3896660251085077e-07
GC_9_20 b_9 NI_9 NS_20 0 3.6755298553610357e-07
GC_9_21 b_9 NI_9 NS_21 0 -1.0208056174360422e-06
GC_9_22 b_9 NI_9 NS_22 0 5.9502482497461916e-07
GC_9_23 b_9 NI_9 NS_23 0 -4.1423525915172778e-07
GC_9_24 b_9 NI_9 NS_24 0 2.6100158427881656e-07
GC_9_25 b_9 NI_9 NS_25 0 -8.5708678366132292e-07
GC_9_26 b_9 NI_9 NS_26 0 4.4785382869254763e-07
GC_9_27 b_9 NI_9 NS_27 0 1.5654084253933593e-07
GC_9_28 b_9 NI_9 NS_28 0 1.1343653630107352e-06
GC_9_29 b_9 NI_9 NS_29 0 -5.9604689793783865e-07
GC_9_30 b_9 NI_9 NS_30 0 1.1950662215163326e-07
GC_9_31 b_9 NI_9 NS_31 0 -1.9175645799222253e-06
GC_9_32 b_9 NI_9 NS_32 0 1.2778549763932725e-06
GC_9_33 b_9 NI_9 NS_33 0 2.0881310633907457e-06
GC_9_34 b_9 NI_9 NS_34 0 2.7546863674275794e-07
GC_9_35 b_9 NI_9 NS_35 0 -6.8903145771085362e-07
GC_9_36 b_9 NI_9 NS_36 0 1.8923877332695052e-07
GC_9_37 b_9 NI_9 NS_37 0 9.8702541651856936e-07
GC_9_38 b_9 NI_9 NS_38 0 1.7040542666912704e-06
GC_9_39 b_9 NI_9 NS_39 0 -2.2913288399007661e-07
GC_9_40 b_9 NI_9 NS_40 0 -5.8920985370547803e-07
GC_9_41 b_9 NI_9 NS_41 0 -9.2846687238369818e-07
GC_9_42 b_9 NI_9 NS_42 0 4.1750095216738921e-07
GC_9_43 b_9 NI_9 NS_43 0 1.4336542094725202e-06
GC_9_44 b_9 NI_9 NS_44 0 7.1202838526139603e-07
GC_9_45 b_9 NI_9 NS_45 0 -3.3623676587888357e-07
GC_9_46 b_9 NI_9 NS_46 0 -2.1999177429467350e-07
GC_9_47 b_9 NI_9 NS_47 0 -5.1611154446394795e-08
GC_9_48 b_9 NI_9 NS_48 0 1.4321515496982831e-06
GC_9_49 b_9 NI_9 NS_49 0 4.8239746296067749e-07
GC_9_50 b_9 NI_9 NS_50 0 -7.6567487829049584e-07
GC_9_51 b_9 NI_9 NS_51 0 -3.5368855309321490e-07
GC_9_52 b_9 NI_9 NS_52 0 4.3186416799472187e-08
GC_9_53 b_9 NI_9 NS_53 0 3.2325024081410439e-07
GC_9_54 b_9 NI_9 NS_54 0 3.8951590294835251e-07
GC_9_55 b_9 NI_9 NS_55 0 -1.4421295037810203e-07
GC_9_56 b_9 NI_9 NS_56 0 -1.1106861819191322e-08
GC_9_57 b_9 NI_9 NS_57 0 1.4081967171401353e-07
GC_9_58 b_9 NI_9 NS_58 0 1.2556217329354836e-07
GC_9_59 b_9 NI_9 NS_59 0 -1.9026591599783155e-07
GC_9_60 b_9 NI_9 NS_60 0 -6.9780405291561863e-08
GC_9_61 b_9 NI_9 NS_61 0 3.9138880911898756e-08
GC_9_62 b_9 NI_9 NS_62 0 1.9887754419401708e-07
GC_9_63 b_9 NI_9 NS_63 0 -1.1141302976486070e-07
GC_9_64 b_9 NI_9 NS_64 0 9.4556837721573476e-09
GC_9_65 b_9 NI_9 NS_65 0 4.6234685749202573e-08
GC_9_66 b_9 NI_9 NS_66 0 7.7272943687127683e-09
GC_9_67 b_9 NI_9 NS_67 0 -2.9801153955216022e-07
GC_9_68 b_9 NI_9 NS_68 0 -5.3663285406499936e-08
GC_9_69 b_9 NI_9 NS_69 0 -9.1173201304983047e-08
GC_9_70 b_9 NI_9 NS_70 0 6.3261696460813621e-08
GC_9_71 b_9 NI_9 NS_71 0 -2.3127801741821089e-07
GC_9_72 b_9 NI_9 NS_72 0 7.8911521342620918e-08
GC_9_73 b_9 NI_9 NS_73 0 -1.3267285859459863e-07
GC_9_74 b_9 NI_9 NS_74 0 -6.8277936408681370e-08
GC_9_75 b_9 NI_9 NS_75 0 -4.3132369328655996e-07
GC_9_76 b_9 NI_9 NS_76 0 -5.7064505942510917e-08
GC_9_77 b_9 NI_9 NS_77 0 -4.2194781187280593e-07
GC_9_78 b_9 NI_9 NS_78 0 6.4454330674229473e-08
GC_9_79 b_9 NI_9 NS_79 0 -4.4334313557731583e-07
GC_9_80 b_9 NI_9 NS_80 0 1.4505056046240379e-07
GC_9_81 b_9 NI_9 NS_81 0 -5.1253938629023087e-07
GC_9_82 b_9 NI_9 NS_82 0 1.0381961058999553e-07
GC_9_83 b_9 NI_9 NS_83 0 -9.6705488514418127e-07
GC_9_84 b_9 NI_9 NS_84 0 -9.9959444515414835e-08
GC_9_85 b_9 NI_9 NS_85 0 2.6356991364168811e-06
GC_9_86 b_9 NI_9 NS_86 0 3.0027987809367931e-06
GC_9_87 b_9 NI_9 NS_87 0 -6.1775287196411023e-07
GC_9_88 b_9 NI_9 NS_88 0 1.0421155073609758e-06
GC_9_89 b_9 NI_9 NS_89 0 9.1780819392393332e-09
GC_9_90 b_9 NI_9 NS_90 0 2.5495436908622825e-08
GC_9_91 b_9 NI_9 NS_91 0 -4.7283713333114220e-07
GC_9_92 b_9 NI_9 NS_92 0 8.3077593631522014e-07
GC_9_93 b_9 NI_9 NS_93 0 9.5158816962991784e-09
GC_9_94 b_9 NI_9 NS_94 0 3.8773704411418864e-07
GC_9_95 b_9 NI_9 NS_95 0 -8.7248194685360789e-07
GC_9_96 b_9 NI_9 NS_96 0 -7.3606251122581511e-08
GC_9_97 b_9 NI_9 NS_97 0 -9.8320782969149662e-07
GC_9_98 b_9 NI_9 NS_98 0 -1.8084375269293860e-07
GC_9_99 b_9 NI_9 NS_99 0 1.0885131908241360e-07
GC_9_100 b_9 NI_9 NS_100 0 -1.4767351158519386e-07
GC_9_101 b_9 NI_9 NS_101 0 6.7365811192392759e-08
GC_9_102 b_9 NI_9 NS_102 0 1.3222898135337727e-08
GC_9_103 b_9 NI_9 NS_103 0 -6.9919566890869133e-08
GC_9_104 b_9 NI_9 NS_104 0 1.6104206303808446e-07
GC_9_105 b_9 NI_9 NS_105 0 2.8981720799672074e-08
GC_9_106 b_9 NI_9 NS_106 0 -4.0222870968357580e-08
GC_9_107 b_9 NI_9 NS_107 0 -8.1261282781496373e-08
GC_9_108 b_9 NI_9 NS_108 0 1.6009598723984954e-07
GC_9_109 b_9 NI_9 NS_109 0 5.6392814277291463e-08
GC_9_110 b_9 NI_9 NS_110 0 -1.6240567997002957e-08
GC_9_111 b_9 NI_9 NS_111 0 -1.1754944103217100e-11
GC_9_112 b_9 NI_9 NS_112 0 5.1377514848256476e-12
GC_9_113 b_9 NI_9 NS_113 0 -3.4035806327184368e-10
GC_9_114 b_9 NI_9 NS_114 0 -9.7344865412090831e-10
GC_9_115 b_9 NI_9 NS_115 0 -2.7509041501259305e-05
GC_9_116 b_9 NI_9 NS_116 0 -1.0597401274346783e-08
GC_9_117 b_9 NI_9 NS_117 0 1.0238697292720393e-11
GC_9_118 b_9 NI_9 NS_118 0 -5.9557113996745083e-11
GC_9_119 b_9 NI_9 NS_119 0 -6.3653752079486505e-07
GC_9_120 b_9 NI_9 NS_120 0 -1.0748116880182433e-06
GC_9_121 b_9 NI_9 NS_121 0 -1.4323577862559950e-06
GC_9_122 b_9 NI_9 NS_122 0 2.3248331677632947e-06
GC_9_123 b_9 NI_9 NS_123 0 -3.8131170164671199e-06
GC_9_124 b_9 NI_9 NS_124 0 2.1795976655387724e-06
GC_9_125 b_9 NI_9 NS_125 0 1.9255578571279110e-06
GC_9_126 b_9 NI_9 NS_126 0 -2.3465996891319070e-07
GC_9_127 b_9 NI_9 NS_127 0 1.4104640050251622e-06
GC_9_128 b_9 NI_9 NS_128 0 5.7203967553550945e-06
GC_9_129 b_9 NI_9 NS_129 0 3.7052085437973222e-06
GC_9_130 b_9 NI_9 NS_130 0 3.2538153353741458e-06
GC_9_131 b_9 NI_9 NS_131 0 -1.4742178717705602e-06
GC_9_132 b_9 NI_9 NS_132 0 -9.4918361300826419e-07
GC_9_133 b_9 NI_9 NS_133 0 9.7320412656241526e-07
GC_9_134 b_9 NI_9 NS_134 0 -2.1860351980158695e-06
GC_9_135 b_9 NI_9 NS_135 0 6.4354354597529846e-06
GC_9_136 b_9 NI_9 NS_136 0 8.5306894820026987e-06
GC_9_137 b_9 NI_9 NS_137 0 1.3303275548184223e-06
GC_9_138 b_9 NI_9 NS_138 0 -9.3980216222904945e-07
GC_9_139 b_9 NI_9 NS_139 0 1.0706359832758976e-06
GC_9_140 b_9 NI_9 NS_140 0 -1.9034741543419507e-06
GC_9_141 b_9 NI_9 NS_141 0 1.4528577445566961e-05
GC_9_142 b_9 NI_9 NS_142 0 -4.1922166893907221e-06
GC_9_143 b_9 NI_9 NS_143 0 -2.0125785544217147e-07
GC_9_144 b_9 NI_9 NS_144 0 6.7953589914870321e-07
GC_9_145 b_9 NI_9 NS_145 0 4.9185661972159806e-06
GC_9_146 b_9 NI_9 NS_146 0 -2.1983603756059665e-06
GC_9_147 b_9 NI_9 NS_147 0 -7.4680005137058598e-07
GC_9_148 b_9 NI_9 NS_148 0 -1.4996597882376163e-05
GC_9_149 b_9 NI_9 NS_149 0 -7.6214280688737954e-08
GC_9_150 b_9 NI_9 NS_150 0 9.7377499067124864e-07
GC_9_151 b_9 NI_9 NS_151 0 -7.9309419669178937e-06
GC_9_152 b_9 NI_9 NS_152 0 -8.5785576627352393e-06
GC_9_153 b_9 NI_9 NS_153 0 -6.2159029843692804e-07
GC_9_154 b_9 NI_9 NS_154 0 -2.1586658901070517e-06
GC_9_155 b_9 NI_9 NS_155 0 -8.3445024485419509e-09
GC_9_156 b_9 NI_9 NS_156 0 1.2073979760631016e-06
GC_9_157 b_9 NI_9 NS_157 0 -7.7192702802343068e-06
GC_9_158 b_9 NI_9 NS_158 0 1.9618087267764367e-06
GC_9_159 b_9 NI_9 NS_159 0 2.4500579579279699e-07
GC_9_160 b_9 NI_9 NS_160 0 -1.6819728413700786e-06
GC_9_161 b_9 NI_9 NS_161 0 1.1609021714110457e-06
GC_9_162 b_9 NI_9 NS_162 0 3.0678712733372934e-06
GC_9_163 b_9 NI_9 NS_163 0 -9.7673159367573392e-07
GC_9_164 b_9 NI_9 NS_164 0 2.0311448235076107e-06
GC_9_165 b_9 NI_9 NS_165 0 4.5640961975192305e-07
GC_9_166 b_9 NI_9 NS_166 0 -1.2309820271306373e-06
GC_9_167 b_9 NI_9 NS_167 0 3.2453607655045493e-06
GC_9_168 b_9 NI_9 NS_168 0 -8.8264228614508933e-07
GC_9_169 b_9 NI_9 NS_169 0 -1.6148353808492859e-07
GC_9_170 b_9 NI_9 NS_170 0 5.1316774169435726e-07
GC_9_171 b_9 NI_9 NS_171 0 -8.4629489634126805e-07
GC_9_172 b_9 NI_9 NS_172 0 -4.1984251888026910e-07
GC_9_173 b_9 NI_9 NS_173 0 9.9342089208378645e-07
GC_9_174 b_9 NI_9 NS_174 0 -1.2690023742496305e-06
GC_9_175 b_9 NI_9 NS_175 0 1.4441165221188879e-06
GC_9_176 b_9 NI_9 NS_176 0 -5.7046178189623110e-07
GC_9_177 b_9 NI_9 NS_177 0 -3.4130250200412914e-08
GC_9_178 b_9 NI_9 NS_178 0 9.6986922138785384e-08
GC_9_179 b_9 NI_9 NS_179 0 -5.9769283658525600e-07
GC_9_180 b_9 NI_9 NS_180 0 -3.4061504945716134e-07
GC_9_181 b_9 NI_9 NS_181 0 9.6765048353396503e-07
GC_9_182 b_9 NI_9 NS_182 0 -1.0810577660503904e-06
GC_9_183 b_9 NI_9 NS_183 0 1.3955346878365327e-06
GC_9_184 b_9 NI_9 NS_184 0 -1.2449194612721241e-06
GC_9_185 b_9 NI_9 NS_185 0 1.6144601941838522e-07
GC_9_186 b_9 NI_9 NS_186 0 -4.3249508155555168e-08
GC_9_187 b_9 NI_9 NS_187 0 -4.8924574449405043e-07
GC_9_188 b_9 NI_9 NS_188 0 -5.0362527561337153e-07
GC_9_189 b_9 NI_9 NS_189 0 1.0632979176975084e-06
GC_9_190 b_9 NI_9 NS_190 0 -8.0455049044801761e-07
GC_9_191 b_9 NI_9 NS_191 0 1.2280666749253875e-06
GC_9_192 b_9 NI_9 NS_192 0 -2.1206296040261025e-06
GC_9_193 b_9 NI_9 NS_193 0 4.9662065287750082e-07
GC_9_194 b_9 NI_9 NS_194 0 -2.5357201552570170e-07
GC_9_195 b_9 NI_9 NS_195 0 -2.4768517647682729e-07
GC_9_196 b_9 NI_9 NS_196 0 -9.1985226106190023e-07
GC_9_197 b_9 NI_9 NS_197 0 1.9186422021518583e-06
GC_9_198 b_9 NI_9 NS_198 0 -1.0012952206130707e-06
GC_9_199 b_9 NI_9 NS_199 0 -8.0998522776597096e-06
GC_9_200 b_9 NI_9 NS_200 0 -9.1472711760878546e-07
GC_9_201 b_9 NI_9 NS_201 0 -3.1607454298192634e-07
GC_9_202 b_9 NI_9 NS_202 0 -3.6265016944833296e-06
GC_9_203 b_9 NI_9 NS_203 0 -4.9018367158752116e-08
GC_9_204 b_9 NI_9 NS_204 0 -3.3203233017048538e-08
GC_9_205 b_9 NI_9 NS_205 0 -1.0293853396408418e-07
GC_9_206 b_9 NI_9 NS_206 0 -1.2361537897729638e-06
GC_9_207 b_9 NI_9 NS_207 0 -1.0227385934227153e-06
GC_9_208 b_9 NI_9 NS_208 0 -6.6783781207249377e-07
GC_9_209 b_9 NI_9 NS_209 0 1.4569278564815715e-06
GC_9_210 b_9 NI_9 NS_210 0 -7.6152617148752209e-07
GC_9_211 b_9 NI_9 NS_211 0 1.9436982745095111e-06
GC_9_212 b_9 NI_9 NS_212 0 -1.8722493517157300e-06
GC_9_213 b_9 NI_9 NS_213 0 -2.2230882704067001e-07
GC_9_214 b_9 NI_9 NS_214 0 3.2515851532252425e-07
GC_9_215 b_9 NI_9 NS_215 0 2.1538427757620612e-07
GC_9_216 b_9 NI_9 NS_216 0 5.2991347841554957e-07
GC_9_217 b_9 NI_9 NS_217 0 -1.0774247839097116e-07
GC_9_218 b_9 NI_9 NS_218 0 -2.8383124767849572e-07
GC_9_219 b_9 NI_9 NS_219 0 8.1696263497221109e-09
GC_9_220 b_9 NI_9 NS_220 0 -9.6164285617463144e-08
GC_9_221 b_9 NI_9 NS_221 0 -8.8650152560124967e-08
GC_9_222 b_9 NI_9 NS_222 0 4.2005177065652079e-08
GC_9_223 b_9 NI_9 NS_223 0 -1.2200379165747208e-07
GC_9_224 b_9 NI_9 NS_224 0 -5.3538923601376014e-08
GC_9_225 b_9 NI_9 NS_225 0 6.1367862149726440e-12
GC_9_226 b_9 NI_9 NS_226 0 -1.6271098060728268e-12
GC_9_227 b_9 NI_9 NS_227 0 3.5453273490338349e-10
GC_9_228 b_9 NI_9 NS_228 0 6.9229772964763057e-10
GC_9_229 b_9 NI_9 NS_229 0 4.4178795684001749e-05
GC_9_230 b_9 NI_9 NS_230 0 -2.5097412377992475e-07
GC_9_231 b_9 NI_9 NS_231 0 -1.3616422025879731e-11
GC_9_232 b_9 NI_9 NS_232 0 3.6731332412081374e-10
GC_9_233 b_9 NI_9 NS_233 0 9.4989300685535022e-07
GC_9_234 b_9 NI_9 NS_234 0 -2.0375955111976366e-07
GC_9_235 b_9 NI_9 NS_235 0 1.1052398088627723e-06
GC_9_236 b_9 NI_9 NS_236 0 -6.5609246529680960e-07
GC_9_237 b_9 NI_9 NS_237 0 1.6285602842958124e-06
GC_9_238 b_9 NI_9 NS_238 0 -3.6726495806254725e-06
GC_9_239 b_9 NI_9 NS_239 0 -2.3668555925980252e-06
GC_9_240 b_9 NI_9 NS_240 0 -1.3304944402519044e-06
GC_9_241 b_9 NI_9 NS_241 0 -2.0337063718207329e-07
GC_9_242 b_9 NI_9 NS_242 0 -2.4446336769977197e-06
GC_9_243 b_9 NI_9 NS_243 0 -7.1160019719866585e-06
GC_9_244 b_9 NI_9 NS_244 0 -2.8108042995810801e-06
GC_9_245 b_9 NI_9 NS_245 0 1.7245505252153352e-06
GC_9_246 b_9 NI_9 NS_246 0 1.3116945066209572e-06
GC_9_247 b_9 NI_9 NS_247 0 -1.6513643830306775e-06
GC_9_248 b_9 NI_9 NS_248 0 9.9670700378047566e-07
GC_9_249 b_9 NI_9 NS_249 0 -2.8708730768596750e-06
GC_9_250 b_9 NI_9 NS_250 0 -1.6219539826659549e-06
GC_9_251 b_9 NI_9 NS_251 0 -2.0401476060170159e-06
GC_9_252 b_9 NI_9 NS_252 0 2.9684647092301637e-06
GC_9_253 b_9 NI_9 NS_253 0 -1.1731544647535430e-06
GC_9_254 b_9 NI_9 NS_254 0 1.1051534896602003e-06
GC_9_255 b_9 NI_9 NS_255 0 -2.0979531877650831e-06
GC_9_256 b_9 NI_9 NS_256 0 1.5287389605739853e-06
GC_9_257 b_9 NI_9 NS_257 0 -9.4304101600369787e-07
GC_9_258 b_9 NI_9 NS_258 0 1.4308248299770105e-06
GC_9_259 b_9 NI_9 NS_259 0 -1.4825500990005666e-06
GC_9_260 b_9 NI_9 NS_260 0 1.7944073236540046e-06
GC_9_261 b_9 NI_9 NS_261 0 2.5486686778649822e-07
GC_9_262 b_9 NI_9 NS_262 0 1.3614198122281310e-06
GC_9_263 b_9 NI_9 NS_263 0 -8.4242883864902722e-07
GC_9_264 b_9 NI_9 NS_264 0 1.3601202593294448e-06
GC_9_265 b_9 NI_9 NS_265 0 9.0836400857927974e-07
GC_9_266 b_9 NI_9 NS_266 0 1.8505877418538279e-06
GC_9_267 b_9 NI_9 NS_267 0 -7.6710009486430729e-07
GC_9_268 b_9 NI_9 NS_268 0 5.7089375890636244e-07
GC_9_269 b_9 NI_9 NS_269 0 -8.0358978940475844e-07
GC_9_270 b_9 NI_9 NS_270 0 1.5919657524836671e-06
GC_9_271 b_9 NI_9 NS_271 0 1.2780286724795963e-06
GC_9_272 b_9 NI_9 NS_272 0 5.6829633813621685e-07
GC_9_273 b_9 NI_9 NS_273 0 -6.6681064550050625e-07
GC_9_274 b_9 NI_9 NS_274 0 6.5600762888398781e-07
GC_9_275 b_9 NI_9 NS_275 0 5.3995016983139459e-07
GC_9_276 b_9 NI_9 NS_276 0 1.7897668104848913e-06
GC_9_277 b_9 NI_9 NS_277 0 -2.5637152330405241e-07
GC_9_278 b_9 NI_9 NS_278 0 -3.2549791864812406e-07
GC_9_279 b_9 NI_9 NS_279 0 -4.7493611474476153e-07
GC_9_280 b_9 NI_9 NS_280 0 6.1075910422362933e-07
GC_9_281 b_9 NI_9 NS_281 0 1.1438063911167653e-07
GC_9_282 b_9 NI_9 NS_282 0 5.8917196424294711e-07
GC_9_283 b_9 NI_9 NS_283 0 -3.1820591341298959e-07
GC_9_284 b_9 NI_9 NS_284 0 4.4619744445507084e-07
GC_9_285 b_9 NI_9 NS_285 0 6.3948100415971505e-08
GC_9_286 b_9 NI_9 NS_286 0 2.2648976554529192e-07
GC_9_287 b_9 NI_9 NS_287 0 -6.7255796203573621e-07
GC_9_288 b_9 NI_9 NS_288 0 2.4745739739571638e-07
GC_9_289 b_9 NI_9 NS_289 0 -1.6417411176369926e-07
GC_9_290 b_9 NI_9 NS_290 0 5.7608780980563412e-07
GC_9_291 b_9 NI_9 NS_291 0 -3.0458984364724658e-07
GC_9_292 b_9 NI_9 NS_292 0 2.5970620496187350e-07
GC_9_293 b_9 NI_9 NS_293 0 -9.8777150532304568e-08
GC_9_294 b_9 NI_9 NS_294 0 2.0871083552509503e-07
GC_9_295 b_9 NI_9 NS_295 0 -7.6626087129431231e-07
GC_9_296 b_9 NI_9 NS_296 0 5.3649739826905492e-08
GC_9_297 b_9 NI_9 NS_297 0 -4.8041861954514509e-07
GC_9_298 b_9 NI_9 NS_298 0 4.3220631802454338e-07
GC_9_299 b_9 NI_9 NS_299 0 -5.3154429467134208e-07
GC_9_300 b_9 NI_9 NS_300 0 2.1428835224888006e-07
GC_9_301 b_9 NI_9 NS_301 0 -5.2281359921034082e-07
GC_9_302 b_9 NI_9 NS_302 0 1.4456661915265831e-07
GC_9_303 b_9 NI_9 NS_303 0 -1.0034209549637761e-06
GC_9_304 b_9 NI_9 NS_304 0 -3.4734795182094431e-07
GC_9_305 b_9 NI_9 NS_305 0 -1.4398179657191318e-06
GC_9_306 b_9 NI_9 NS_306 0 5.4841448493411644e-07
GC_9_307 b_9 NI_9 NS_307 0 -1.1944231084813713e-06
GC_9_308 b_9 NI_9 NS_308 0 1.3611333129640828e-07
GC_9_309 b_9 NI_9 NS_309 0 -1.4807018692410524e-06
GC_9_310 b_9 NI_9 NS_310 0 7.7907298742270473e-07
GC_9_311 b_9 NI_9 NS_311 0 -2.2610248475722297e-06
GC_9_312 b_9 NI_9 NS_312 0 -8.4610142913005654e-07
GC_9_313 b_9 NI_9 NS_313 0 5.6641223691681325e-06
GC_9_314 b_9 NI_9 NS_314 0 1.1197537795626094e-05
GC_9_315 b_9 NI_9 NS_315 0 -2.2220260962417380e-06
GC_9_316 b_9 NI_9 NS_316 0 3.0965170372212685e-06
GC_9_317 b_9 NI_9 NS_317 0 1.1650741949773095e-08
GC_9_318 b_9 NI_9 NS_318 0 7.3480689517925553e-08
GC_9_319 b_9 NI_9 NS_319 0 -1.2474057164821637e-06
GC_9_320 b_9 NI_9 NS_320 0 1.6458709990692271e-06
GC_9_321 b_9 NI_9 NS_321 0 -6.3374339417576425e-07
GC_9_322 b_9 NI_9 NS_322 0 1.4521176135929733e-06
GC_9_323 b_9 NI_9 NS_323 0 -1.6480293500927779e-06
GC_9_324 b_9 NI_9 NS_324 0 -1.2214497713782069e-06
GC_9_325 b_9 NI_9 NS_325 0 -3.3896234629898350e-06
GC_9_326 b_9 NI_9 NS_326 0 -1.1084113492027153e-06
GC_9_327 b_9 NI_9 NS_327 0 7.2039000991249942e-09
GC_9_328 b_9 NI_9 NS_328 0 -1.2022193290901058e-07
GC_9_329 b_9 NI_9 NS_329 0 6.2010527540438070e-07
GC_9_330 b_9 NI_9 NS_330 0 -3.6782706016118710e-07
GC_9_331 b_9 NI_9 NS_331 0 -4.6877957500379864e-08
GC_9_332 b_9 NI_9 NS_332 0 3.9701416846657599e-07
GC_9_333 b_9 NI_9 NS_333 0 -5.1628189339466620e-08
GC_9_334 b_9 NI_9 NS_334 0 2.9624232625932148e-08
GC_9_335 b_9 NI_9 NS_335 0 -2.7362447046820943e-07
GC_9_336 b_9 NI_9 NS_336 0 1.7742808204169281e-07
GC_9_337 b_9 NI_9 NS_337 0 -2.2776107167544963e-07
GC_9_338 b_9 NI_9 NS_338 0 -6.5474208636738993e-09
GC_9_339 b_9 NI_9 NS_339 0 -8.0170684652538464e-12
GC_9_340 b_9 NI_9 NS_340 0 -8.1359251355369492e-13
GC_9_341 b_9 NI_9 NS_341 0 -1.1403179256331059e-09
GC_9_342 b_9 NI_9 NS_342 0 -2.4260026294868639e-09
GC_9_343 b_9 NI_9 NS_343 0 -2.1854898732474392e-05
GC_9_344 b_9 NI_9 NS_344 0 2.4289032973213134e-07
GC_9_345 b_9 NI_9 NS_345 0 1.6216453969519895e-11
GC_9_346 b_9 NI_9 NS_346 0 -4.8482518114008598e-10
GC_9_347 b_9 NI_9 NS_347 0 3.7396392858632240e-07
GC_9_348 b_9 NI_9 NS_348 0 -1.3861162159127028e-06
GC_9_349 b_9 NI_9 NS_349 0 -1.4309825013009588e-07
GC_9_350 b_9 NI_9 NS_350 0 1.1186852052612925e-06
GC_9_351 b_9 NI_9 NS_351 0 -3.5071057701088160e-06
GC_9_352 b_9 NI_9 NS_352 0 -2.2368600656703287e-06
GC_9_353 b_9 NI_9 NS_353 0 -7.4899833313653614e-07
GC_9_354 b_9 NI_9 NS_354 0 -1.1228906775896887e-06
GC_9_355 b_9 NI_9 NS_355 0 -6.8318292371929336e-07
GC_9_356 b_9 NI_9 NS_356 0 2.6597428435692792e-06
GC_9_357 b_9 NI_9 NS_357 0 -5.0808555857082102e-06
GC_9_358 b_9 NI_9 NS_358 0 3.8731932358232743e-06
GC_9_359 b_9 NI_9 NS_359 0 9.5027397168952903e-07
GC_9_360 b_9 NI_9 NS_360 0 -1.5539847574673620e-07
GC_9_361 b_9 NI_9 NS_361 0 -2.6330610442856616e-07
GC_9_362 b_9 NI_9 NS_362 0 -5.2973856950195683e-07
GC_9_363 b_9 NI_9 NS_363 0 -1.4734358493286304e-06
GC_9_364 b_9 NI_9 NS_364 0 1.1165100596554298e-05
GC_9_365 b_9 NI_9 NS_365 0 5.7514567106243325e-06
GC_9_366 b_9 NI_9 NS_366 0 2.9696708376758333e-06
GC_9_367 b_9 NI_9 NS_367 0 7.6119639712926821e-07
GC_9_368 b_9 NI_9 NS_368 0 -4.0129844906631020e-07
GC_9_369 b_9 NI_9 NS_369 0 1.7102520244720120e-05
GC_9_370 b_9 NI_9 NS_370 0 -2.9720721131103616e-07
GC_9_371 b_9 NI_9 NS_371 0 6.9918255923296377e-07
GC_9_372 b_9 NI_9 NS_372 0 1.7754998557778110e-07
GC_9_373 b_9 NI_9 NS_373 0 6.4112249157174576e-06
GC_9_374 b_9 NI_9 NS_374 0 -4.4582134042783782e-07
GC_9_375 b_9 NI_9 NS_375 0 -8.2285114090937986e-07
GC_9_376 b_9 NI_9 NS_376 0 -1.7742557716688296e-05
GC_9_377 b_9 NI_9 NS_377 0 -2.8404103725428003e-07
GC_9_378 b_9 NI_9 NS_378 0 2.3076338376262813e-07
GC_9_379 b_9 NI_9 NS_379 0 -1.0767534489955630e-05
GC_9_380 b_9 NI_9 NS_380 0 -9.4785272528542896e-06
GC_9_381 b_9 NI_9 NS_381 0 -1.3407981958788556e-06
GC_9_382 b_9 NI_9 NS_382 0 -8.1236646810183990e-07
GC_9_383 b_9 NI_9 NS_383 0 -1.6041529792509986e-06
GC_9_384 b_9 NI_9 NS_384 0 4.5798622339895924e-07
GC_9_385 b_9 NI_9 NS_385 0 -9.3315599801851511e-06
GC_9_386 b_9 NI_9 NS_386 0 6.4364183886657689e-06
GC_9_387 b_9 NI_9 NS_387 0 6.8137731897704617e-08
GC_9_388 b_9 NI_9 NS_388 0 -4.0002747660681432e-07
GC_9_389 b_9 NI_9 NS_389 0 -7.1694151964072380e-07
GC_9_390 b_9 NI_9 NS_390 0 7.2315348962583244e-06
GC_9_391 b_9 NI_9 NS_391 0 2.0724142548992154e-06
GC_9_392 b_9 NI_9 NS_392 0 2.4601628466824145e-06
GC_9_393 b_9 NI_9 NS_393 0 6.1987265103713370e-07
GC_9_394 b_9 NI_9 NS_394 0 -2.5283369524835602e-07
GC_9_395 b_9 NI_9 NS_395 0 4.6121022659590204e-06
GC_9_396 b_9 NI_9 NS_396 0 3.3416392066753116e-07
GC_9_397 b_9 NI_9 NS_397 0 1.7600765258883748e-07
GC_9_398 b_9 NI_9 NS_398 0 5.3884837203498792e-07
GC_9_399 b_9 NI_9 NS_399 0 -7.4062783721250376e-07
GC_9_400 b_9 NI_9 NS_400 0 -4.2130513619078304e-08
GC_9_401 b_9 NI_9 NS_401 0 7.4630740639294666e-07
GC_9_402 b_9 NI_9 NS_402 0 -5.2040151645226151e-07
GC_9_403 b_9 NI_9 NS_403 0 1.8297456256238587e-06
GC_9_404 b_9 NI_9 NS_404 0 4.7558623902812081e-07
GC_9_405 b_9 NI_9 NS_405 0 1.7694711048210702e-07
GC_9_406 b_9 NI_9 NS_406 0 4.5204846932911299e-07
GC_9_407 b_9 NI_9 NS_407 0 -4.4611008130127161e-07
GC_9_408 b_9 NI_9 NS_408 0 2.3590853143460953e-07
GC_9_409 b_9 NI_9 NS_409 0 6.5001245338525778e-07
GC_9_410 b_9 NI_9 NS_410 0 -3.4566542368453864e-07
GC_9_411 b_9 NI_9 NS_411 0 1.8731754233544094e-06
GC_9_412 b_9 NI_9 NS_412 0 -2.9453286952382257e-08
GC_9_413 b_9 NI_9 NS_413 0 2.9821068831595968e-07
GC_9_414 b_9 NI_9 NS_414 0 5.0989368271927119e-07
GC_9_415 b_9 NI_9 NS_415 0 -3.1510375946607055e-07
GC_9_416 b_9 NI_9 NS_416 0 4.5573825887026289e-07
GC_9_417 b_9 NI_9 NS_417 0 5.5362650114166634e-07
GC_9_418 b_9 NI_9 NS_418 0 -4.4921605099371550e-08
GC_9_419 b_9 NI_9 NS_419 0 1.9806826658144210e-06
GC_9_420 b_9 NI_9 NS_420 0 -4.0116437661049557e-07
GC_9_421 b_9 NI_9 NS_421 0 4.1707470766635933e-07
GC_9_422 b_9 NI_9 NS_422 0 7.7173705481067036e-07
GC_9_423 b_9 NI_9 NS_423 0 5.0608697489766856e-07
GC_9_424 b_9 NI_9 NS_424 0 7.2744455312879661e-07
GC_9_425 b_9 NI_9 NS_425 0 9.0286786407057327e-07
GC_9_426 b_9 NI_9 NS_426 0 9.8962637239520543e-07
GC_9_427 b_9 NI_9 NS_427 0 1.6379038704215743e-06
GC_9_428 b_9 NI_9 NS_428 0 -9.9914033300695327e-06
GC_9_429 b_9 NI_9 NS_429 0 2.8722353464853756e-06
GC_9_430 b_9 NI_9 NS_430 0 -1.2252754867813451e-06
GC_9_431 b_9 NI_9 NS_431 0 3.1662832373194620e-08
GC_9_432 b_9 NI_9 NS_432 0 -4.6443104871015184e-08
GC_9_433 b_9 NI_9 NS_433 0 1.4053604831410736e-06
GC_9_434 b_9 NI_9 NS_434 0 1.6962628084612953e-07
GC_9_435 b_9 NI_9 NS_435 0 9.7886695774623555e-07
GC_9_436 b_9 NI_9 NS_436 0 -4.9524041064724348e-07
GC_9_437 b_9 NI_9 NS_437 0 6.9365257574961086e-07
GC_9_438 b_9 NI_9 NS_438 0 1.3037929226879007e-06
GC_9_439 b_9 NI_9 NS_439 0 1.3369678947941026e-06
GC_9_440 b_9 NI_9 NS_440 0 1.9872992037663219e-06
GC_9_441 b_9 NI_9 NS_441 0 -9.2422196943509684e-08
GC_9_442 b_9 NI_9 NS_442 0 -2.7687535711030998e-08
GC_9_443 b_9 NI_9 NS_443 0 -5.3468576582525898e-07
GC_9_444 b_9 NI_9 NS_444 0 1.8254488528542636e-07
GC_9_445 b_9 NI_9 NS_445 0 3.1918830969756021e-07
GC_9_446 b_9 NI_9 NS_446 0 -3.6116517032264078e-07
GC_9_447 b_9 NI_9 NS_447 0 1.1497614511805630e-08
GC_9_448 b_9 NI_9 NS_448 0 -6.0654804995361749e-07
GC_9_449 b_9 NI_9 NS_449 0 5.2303457259013476e-08
GC_9_450 b_9 NI_9 NS_450 0 1.0683489480045981e-07
GC_9_451 b_9 NI_9 NS_451 0 2.9593182741829641e-07
GC_9_452 b_9 NI_9 NS_452 0 -1.4168002860403877e-09
GC_9_453 b_9 NI_9 NS_453 0 -2.9849938308970166e-12
GC_9_454 b_9 NI_9 NS_454 0 -1.0058647753224846e-11
GC_9_455 b_9 NI_9 NS_455 0 9.3171479535378291e-10
GC_9_456 b_9 NI_9 NS_456 0 3.3553250630638974e-09
GC_9_457 b_9 NI_9 NS_457 0 -1.1661778302065817e-04
GC_9_458 b_9 NI_9 NS_458 0 -2.1401248505867823e-06
GC_9_459 b_9 NI_9 NS_459 0 -2.5040564412715954e-10
GC_9_460 b_9 NI_9 NS_460 0 2.6003939918206516e-09
GC_9_461 b_9 NI_9 NS_461 0 1.7091685665453935e-06
GC_9_462 b_9 NI_9 NS_462 0 -1.5815005182495531e-06
GC_9_463 b_9 NI_9 NS_463 0 1.2865051683781640e-07
GC_9_464 b_9 NI_9 NS_464 0 -6.3839770610676897e-06
GC_9_465 b_9 NI_9 NS_465 0 -7.6493577515423871e-06
GC_9_466 b_9 NI_9 NS_466 0 1.1913581114464483e-07
GC_9_467 b_9 NI_9 NS_467 0 -1.2236192411484646e-06
GC_9_468 b_9 NI_9 NS_468 0 -4.6177282954810212e-06
GC_9_469 b_9 NI_9 NS_469 0 -1.5901243080749650e-05
GC_9_470 b_9 NI_9 NS_470 0 -1.6609734490879161e-06
GC_9_471 b_9 NI_9 NS_471 0 -6.2265117659788633e-06
GC_9_472 b_9 NI_9 NS_472 0 1.9173247926651815e-05
GC_9_473 b_9 NI_9 NS_473 0 4.6915553437265260e-06
GC_9_474 b_9 NI_9 NS_474 0 -3.0032580134002338e-06
GC_9_475 b_9 NI_9 NS_475 0 -1.8663119248296669e-08
GC_9_476 b_9 NI_9 NS_476 0 -2.5775023834896314e-06
GC_9_477 b_9 NI_9 NS_477 0 -2.5961794562826505e-05
GC_9_478 b_9 NI_9 NS_478 0 2.8474538387377566e-05
GC_9_479 b_9 NI_9 NS_479 0 2.8294920892963469e-05
GC_9_480 b_9 NI_9 NS_480 0 -8.4647888184151018e-06
GC_9_481 b_9 NI_9 NS_481 0 -8.0582938353138106e-06
GC_9_482 b_9 NI_9 NS_482 0 -4.3213663683899916e-06
GC_9_483 b_9 NI_9 NS_483 0 1.2613103686100237e-05
GC_9_484 b_9 NI_9 NS_484 0 2.7036770502370558e-05
GC_9_485 b_9 NI_9 NS_485 0 1.4849127229805651e-06
GC_9_486 b_9 NI_9 NS_486 0 -8.9982176694789761e-06
GC_9_487 b_9 NI_9 NS_487 0 -2.8357601326713517e-05
GC_9_488 b_9 NI_9 NS_488 0 4.7238550692924535e-06
GC_9_489 b_9 NI_9 NS_489 0 4.1379064735050014e-05
GC_9_490 b_9 NI_9 NS_490 0 1.0729943473584398e-05
GC_9_491 b_9 NI_9 NS_491 0 -2.9667043454258169e-06
GC_9_492 b_9 NI_9 NS_492 0 -4.4978586251299466e-06
GC_9_493 b_9 NI_9 NS_493 0 1.2948378520570635e-05
GC_9_494 b_9 NI_9 NS_494 0 1.9022647176987082e-05
GC_9_495 b_9 NI_9 NS_495 0 3.8280368170438073e-06
GC_9_496 b_9 NI_9 NS_496 0 -1.0937998168637503e-05
GC_9_497 b_9 NI_9 NS_497 0 -6.4224019961541911e-06
GC_9_498 b_9 NI_9 NS_498 0 8.3857926901689193e-07
GC_9_499 b_9 NI_9 NS_499 0 1.8903998674643618e-05
GC_9_500 b_9 NI_9 NS_500 0 5.4505926039620434e-06
GC_9_501 b_9 NI_9 NS_501 0 -6.6494082866221717e-08
GC_9_502 b_9 NI_9 NS_502 0 -4.1973567158909876e-06
GC_9_503 b_9 NI_9 NS_503 0 4.9149595692373307e-06
GC_9_504 b_9 NI_9 NS_504 0 1.4293061416919800e-05
GC_9_505 b_9 NI_9 NS_505 0 7.8466195086564772e-06
GC_9_506 b_9 NI_9 NS_506 0 -1.1186119796747859e-05
GC_9_507 b_9 NI_9 NS_507 0 -1.3863433137528415e-06
GC_9_508 b_9 NI_9 NS_508 0 9.3337898051206076e-07
GC_9_509 b_9 NI_9 NS_509 0 1.0911665112220343e-05
GC_9_510 b_9 NI_9 NS_510 0 4.1227354150807296e-06
GC_9_511 b_9 NI_9 NS_511 0 1.7223613756476202e-06
GC_9_512 b_9 NI_9 NS_512 0 -6.3594465397310470e-07
GC_9_513 b_9 NI_9 NS_513 0 5.6879435487659679e-06
GC_9_514 b_9 NI_9 NS_514 0 1.7020791844560968e-06
GC_9_515 b_9 NI_9 NS_515 0 3.4205428388003651e-06
GC_9_516 b_9 NI_9 NS_516 0 2.0399774964475659e-06
GC_9_517 b_9 NI_9 NS_517 0 1.0979313467998457e-05
GC_9_518 b_9 NI_9 NS_518 0 3.7863786081901621e-06
GC_9_519 b_9 NI_9 NS_519 0 4.8656048834225336e-06
GC_9_520 b_9 NI_9 NS_520 0 -8.4827933837615759e-08
GC_9_521 b_9 NI_9 NS_521 0 9.9928712433075556e-06
GC_9_522 b_9 NI_9 NS_522 0 -1.0833538917868623e-06
GC_9_523 b_9 NI_9 NS_523 0 8.2687932540773924e-06
GC_9_524 b_9 NI_9 NS_524 0 2.9476693696081700e-06
GC_9_525 b_9 NI_9 NS_525 0 1.9077427817696007e-05
GC_9_526 b_9 NI_9 NS_526 0 -5.5657359092692164e-06
GC_9_527 b_9 NI_9 NS_527 0 7.2206796978539004e-06
GC_9_528 b_9 NI_9 NS_528 0 -4.0253011929362216e-06
GC_9_529 b_9 NI_9 NS_529 0 1.3766283198274183e-05
GC_9_530 b_9 NI_9 NS_530 0 -1.1899498487496275e-05
GC_9_531 b_9 NI_9 NS_531 0 1.2420481781473196e-05
GC_9_532 b_9 NI_9 NS_532 0 -3.9375945850844199e-06
GC_9_533 b_9 NI_9 NS_533 0 9.2733685431114432e-06
GC_9_534 b_9 NI_9 NS_534 0 -2.6781575306624002e-05
GC_9_535 b_9 NI_9 NS_535 0 2.4206615914407541e-06
GC_9_536 b_9 NI_9 NS_536 0 -1.2364180937979078e-05
GC_9_537 b_9 NI_9 NS_537 0 -8.1530762071980207e-06
GC_9_538 b_9 NI_9 NS_538 0 -1.8689491930181899e-05
GC_9_539 b_9 NI_9 NS_539 0 -4.7467512267207724e-06
GC_9_540 b_9 NI_9 NS_540 0 -1.1992669038126259e-05
GC_9_541 b_9 NI_9 NS_541 0 5.4596306723404281e-05
GC_9_542 b_9 NI_9 NS_542 0 -8.9145409232708458e-05
GC_9_543 b_9 NI_9 NS_543 0 -9.8008101984038443e-06
GC_9_544 b_9 NI_9 NS_544 0 1.0736449619741642e-06
GC_9_545 b_9 NI_9 NS_545 0 3.9043698492123622e-07
GC_9_546 b_9 NI_9 NS_546 0 -1.3188534147017998e-07
GC_9_547 b_9 NI_9 NS_547 0 -2.5976297935706871e-06
GC_9_548 b_9 NI_9 NS_548 0 -2.0694179712826741e-06
GC_9_549 b_9 NI_9 NS_549 0 -4.3215022066526412e-06
GC_9_550 b_9 NI_9 NS_550 0 4.2993150424804491e-07
GC_9_551 b_9 NI_9 NS_551 0 -1.7356641889474463e-05
GC_9_552 b_9 NI_9 NS_552 0 9.7071549881443079e-06
GC_9_553 b_9 NI_9 NS_553 0 -8.9446470999051620e-06
GC_9_554 b_9 NI_9 NS_554 0 3.7512037428891810e-05
GC_9_555 b_9 NI_9 NS_555 0 -7.2510362631633152e-06
GC_9_556 b_9 NI_9 NS_556 0 3.2526170065847205e-07
GC_9_557 b_9 NI_9 NS_557 0 -1.3466585570689415e-05
GC_9_558 b_9 NI_9 NS_558 0 1.8883237991796121e-06
GC_9_559 b_9 NI_9 NS_559 0 -4.6297889952712540e-06
GC_9_560 b_9 NI_9 NS_560 0 -3.4285053279269003e-06
GC_9_561 b_9 NI_9 NS_561 0 -6.3984880348800768e-06
GC_9_562 b_9 NI_9 NS_562 0 1.0147261805602514e-06
GC_9_563 b_9 NI_9 NS_563 0 -3.0176502765898911e-06
GC_9_564 b_9 NI_9 NS_564 0 8.7792916866856218e-07
GC_9_565 b_9 NI_9 NS_565 0 -1.7623654016110022e-06
GC_9_566 b_9 NI_9 NS_566 0 -9.5961627021492046e-07
GC_9_567 b_9 NI_9 NS_567 0 -2.6113573579157479e-10
GC_9_568 b_9 NI_9 NS_568 0 4.2260594913912326e-10
GC_9_569 b_9 NI_9 NS_569 0 2.2541520937246249e-09
GC_9_570 b_9 NI_9 NS_570 0 -2.6820923586890135e-08
GC_9_571 b_9 NI_9 NS_571 0 -3.2388760432905883e-05
GC_9_572 b_9 NI_9 NS_572 0 2.2145965300072115e-06
GC_9_573 b_9 NI_9 NS_573 0 6.9002925163924588e-11
GC_9_574 b_9 NI_9 NS_574 0 3.0548437001222061e-09
GC_9_575 b_9 NI_9 NS_575 0 -1.7287506039242528e-06
GC_9_576 b_9 NI_9 NS_576 0 -1.8218257444491899e-06
GC_9_577 b_9 NI_9 NS_577 0 -5.3711626207452347e-06
GC_9_578 b_9 NI_9 NS_578 0 2.8657252689747377e-06
GC_9_579 b_9 NI_9 NS_579 0 -1.6530934996843210e-05
GC_9_580 b_9 NI_9 NS_580 0 1.8435105761179463e-05
GC_9_581 b_9 NI_9 NS_581 0 1.5105602032401550e-05
GC_9_582 b_9 NI_9 NS_582 0 9.7996907872192122e-06
GC_9_583 b_9 NI_9 NS_583 0 1.7319442701253400e-05
GC_9_584 b_9 NI_9 NS_584 0 2.2757437399213378e-05
GC_9_585 b_9 NI_9 NS_585 0 2.9271979069670892e-05
GC_9_586 b_9 NI_9 NS_586 0 4.9454582772709867e-06
GC_9_587 b_9 NI_9 NS_587 0 -3.0090421016496078e-06
GC_9_588 b_9 NI_9 NS_588 0 -1.8920185912856242e-06
GC_9_589 b_9 NI_9 NS_589 0 1.6961736740189606e-05
GC_9_590 b_9 NI_9 NS_590 0 -2.2247267278919457e-06
GC_9_591 b_9 NI_9 NS_591 0 1.2894021431622874e-04
GC_9_592 b_9 NI_9 NS_592 0 3.4692077894225310e-05
GC_9_593 b_9 NI_9 NS_593 0 -2.8903922018055944e-05
GC_9_594 b_9 NI_9 NS_594 0 -9.8807837123790837e-05
GC_9_595 b_9 NI_9 NS_595 0 2.4942598695925002e-05
GC_9_596 b_9 NI_9 NS_596 0 -3.1439987842384161e-05
GC_9_597 b_9 NI_9 NS_597 0 -4.1726504239161669e-05
GC_9_598 b_9 NI_9 NS_598 0 -1.6659244514828447e-04
GC_9_599 b_9 NI_9 NS_599 0 -4.1856850868705463e-05
GC_9_600 b_9 NI_9 NS_600 0 -4.9686677977864620e-06
GC_9_601 b_9 NI_9 NS_601 0 2.1526232502915683e-05
GC_9_602 b_9 NI_9 NS_602 0 -1.5189898123168553e-04
GC_9_603 b_9 NI_9 NS_603 0 -2.3067411876468731e-04
GC_9_604 b_9 NI_9 NS_604 0 1.1454640770787045e-04
GC_9_605 b_9 NI_9 NS_605 0 -3.7434566688128722e-05
GC_9_606 b_9 NI_9 NS_606 0 1.4285340975099009e-05
GC_9_607 b_9 NI_9 NS_607 0 -1.3769176199644482e-04
GC_9_608 b_9 NI_9 NS_608 0 1.3059703587333312e-04
GC_9_609 b_9 NI_9 NS_609 0 3.6482331662122002e-05
GC_9_610 b_9 NI_9 NS_610 0 4.1333509032768396e-05
GC_9_611 b_9 NI_9 NS_611 0 -3.8174270410810061e-05
GC_9_612 b_9 NI_9 NS_612 0 4.3297680902104925e-05
GC_9_613 b_9 NI_9 NS_613 0 8.7698891157245531e-05
GC_9_614 b_9 NI_9 NS_614 0 1.1839070798980718e-04
GC_9_615 b_9 NI_9 NS_615 0 2.7360737653951375e-05
GC_9_616 b_9 NI_9 NS_616 0 1.0188167964850283e-05
GC_9_617 b_9 NI_9 NS_617 0 8.7309935113577867e-05
GC_9_618 b_9 NI_9 NS_618 0 6.5589082832175646e-05
GC_9_619 b_9 NI_9 NS_619 0 2.0355451241530548e-05
GC_9_620 b_9 NI_9 NS_620 0 -5.7134225715262953e-05
GC_9_621 b_9 NI_9 NS_621 0 1.6985963393561223e-05
GC_9_622 b_9 NI_9 NS_622 0 -8.8834518135941345e-06
GC_9_623 b_9 NI_9 NS_623 0 8.5005733406582173e-06
GC_9_624 b_9 NI_9 NS_624 0 -3.2939542780647770e-05
GC_9_625 b_9 NI_9 NS_625 0 -8.8537955425135874e-06
GC_9_626 b_9 NI_9 NS_626 0 5.2635716465858812e-07
GC_9_627 b_9 NI_9 NS_627 0 -2.4130971291846179e-06
GC_9_628 b_9 NI_9 NS_628 0 8.5086601830865723e-06
GC_9_629 b_9 NI_9 NS_629 0 1.0220493472574464e-05
GC_9_630 b_9 NI_9 NS_630 0 6.0870248624688566e-06
GC_9_631 b_9 NI_9 NS_631 0 1.2161244014823160e-05
GC_9_632 b_9 NI_9 NS_632 0 -7.8264921759856182e-06
GC_9_633 b_9 NI_9 NS_633 0 -3.4879227353677047e-06
GC_9_634 b_9 NI_9 NS_634 0 -4.4670318540650901e-07
GC_9_635 b_9 NI_9 NS_635 0 2.4880913836327634e-06
GC_9_636 b_9 NI_9 NS_636 0 7.4079290134155306e-06
GC_9_637 b_9 NI_9 NS_637 0 1.3650681219149200e-05
GC_9_638 b_9 NI_9 NS_638 0 2.6359170589941569e-06
GC_9_639 b_9 NI_9 NS_639 0 4.5207284179634278e-06
GC_9_640 b_9 NI_9 NS_640 0 -1.4188592293305564e-05
GC_9_641 b_9 NI_9 NS_641 0 -5.9269927649049638e-06
GC_9_642 b_9 NI_9 NS_642 0 4.2582991545093231e-06
GC_9_643 b_9 NI_9 NS_643 0 1.0309907770102586e-05
GC_9_644 b_9 NI_9 NS_644 0 9.9374981340138197e-06
GC_9_645 b_9 NI_9 NS_645 0 1.7307649562928716e-05
GC_9_646 b_9 NI_9 NS_646 0 -4.2709215632801583e-06
GC_9_647 b_9 NI_9 NS_647 0 -9.2920986707348909e-06
GC_9_648 b_9 NI_9 NS_648 0 -1.5315608286741339e-05
GC_9_649 b_9 NI_9 NS_649 0 -4.0817829305535955e-06
GC_9_650 b_9 NI_9 NS_650 0 1.3516515957847885e-05
GC_9_651 b_9 NI_9 NS_651 0 2.0928899522477301e-05
GC_9_652 b_9 NI_9 NS_652 0 -5.6268005154632278e-07
GC_9_653 b_9 NI_9 NS_653 0 8.8751455370818254e-06
GC_9_654 b_9 NI_9 NS_654 0 -1.7452600515066196e-05
GC_9_655 b_9 NI_9 NS_655 0 2.4051299250993507e-06
GC_9_656 b_9 NI_9 NS_656 0 -1.3697913930405423e-05
GC_9_657 b_9 NI_9 NS_657 0 -1.3815613859654376e-05
GC_9_658 b_9 NI_9 NS_658 0 4.3767964278833732e-06
GC_9_659 b_9 NI_9 NS_659 0 1.5477831196422835e-08
GC_9_660 b_9 NI_9 NS_660 0 -4.2109256663345421e-08
GC_9_661 b_9 NI_9 NS_661 0 8.6211060295431295e-06
GC_9_662 b_9 NI_9 NS_662 0 1.1597923913333124e-05
GC_9_663 b_9 NI_9 NS_663 0 1.0904668398954424e-05
GC_9_664 b_9 NI_9 NS_664 0 -1.1278364353956019e-05
GC_9_665 b_9 NI_9 NS_665 0 -3.7307316839072155e-06
GC_9_666 b_9 NI_9 NS_666 0 -1.0216259524811392e-05
GC_9_667 b_9 NI_9 NS_667 0 -2.2939949886592665e-06
GC_9_668 b_9 NI_9 NS_668 0 1.2865967174373309e-05
GC_9_669 b_9 NI_9 NS_669 0 9.6691381603179502e-07
GC_9_670 b_9 NI_9 NS_670 0 -7.2695105745486640e-06
GC_9_671 b_9 NI_9 NS_671 0 7.5166616339804521e-06
GC_9_672 b_9 NI_9 NS_672 0 1.6931670838971702e-06
GC_9_673 b_9 NI_9 NS_673 0 -6.1012196703864415e-06
GC_9_674 b_9 NI_9 NS_674 0 -8.8953956299886921e-06
GC_9_675 b_9 NI_9 NS_675 0 -4.1215008365320700e-06
GC_9_676 b_9 NI_9 NS_676 0 9.6659608582363802e-06
GC_9_677 b_9 NI_9 NS_677 0 3.3268437505141390e-06
GC_9_678 b_9 NI_9 NS_678 0 6.0367139269211145e-06
GC_9_679 b_9 NI_9 NS_679 0 5.6518861150013398e-06
GC_9_680 b_9 NI_9 NS_680 0 5.1680476187365464e-07
GC_9_681 b_9 NI_9 NS_681 0 6.1804623632451914e-11
GC_9_682 b_9 NI_9 NS_682 0 1.4894796998841887e-10
GC_9_683 b_9 NI_9 NS_683 0 5.9431741637554039e-09
GC_9_684 b_9 NI_9 NS_684 0 -8.3385682064926886e-09
GC_9_685 b_9 NI_9 NS_685 0 2.8654994119341019e-04
GC_9_686 b_9 NI_9 NS_686 0 -1.4350321247396221e-05
GC_9_687 b_9 NI_9 NS_687 0 -1.2377044373114563e-09
GC_9_688 b_9 NI_9 NS_688 0 -1.9231747128620347e-08
GC_9_689 b_9 NI_9 NS_689 0 2.6665546215097546e-06
GC_9_690 b_9 NI_9 NS_690 0 -3.8232154413187678e-06
GC_9_691 b_9 NI_9 NS_691 0 -1.3223098338896242e-05
GC_9_692 b_9 NI_9 NS_692 0 -5.0242681726712457e-07
GC_9_693 b_9 NI_9 NS_693 0 3.9458281226396019e-05
GC_9_694 b_9 NI_9 NS_694 0 2.7880663837424910e-06
GC_9_695 b_9 NI_9 NS_695 0 -4.1775292498016617e-05
GC_9_696 b_9 NI_9 NS_696 0 -2.3733019495907081e-05
GC_9_697 b_9 NI_9 NS_697 0 1.7634779645238484e-06
GC_9_698 b_9 NI_9 NS_698 0 4.4845306801638146e-05
GC_9_699 b_9 NI_9 NS_699 0 1.4501516010159368e-05
GC_9_700 b_9 NI_9 NS_700 0 -4.8185831961484243e-05
GC_9_701 b_9 NI_9 NS_701 0 1.9359386009817131e-06
GC_9_702 b_9 NI_9 NS_702 0 5.6539834944217649e-06
GC_9_703 b_9 NI_9 NS_703 0 -4.4994174996811817e-05
GC_9_704 b_9 NI_9 NS_704 0 1.5684412844049175e-06
GC_9_705 b_9 NI_9 NS_705 0 1.0310756751002312e-04
GC_9_706 b_9 NI_9 NS_706 0 1.2335556679895349e-04
GC_9_707 b_9 NI_9 NS_707 0 -7.5525460511100667e-05
GC_9_708 b_9 NI_9 NS_708 0 -1.3698528238335791e-04
GC_9_709 b_9 NI_9 NS_709 0 -6.7109340630338522e-05
GC_9_710 b_9 NI_9 NS_710 0 4.9269291713957249e-05
GC_9_711 b_9 NI_9 NS_711 0 1.3517087455393762e-04
GC_9_712 b_9 NI_9 NS_712 0 -2.8537418236659638e-05
GC_9_713 b_9 NI_9 NS_713 0 -8.7330925850784825e-05
GC_9_714 b_9 NI_9 NS_714 0 -1.1763161385983049e-05
GC_9_715 b_9 NI_9 NS_715 0 -9.4647116517989136e-05
GC_9_716 b_9 NI_9 NS_716 0 2.1148781166705378e-04
GC_9_717 b_9 NI_9 NS_717 0 1.6429617662777781e-04
GC_9_718 b_9 NI_9 NS_718 0 -2.1487400936091161e-04
GC_9_719 b_9 NI_9 NS_719 0 -8.1684433830341862e-05
GC_9_720 b_9 NI_9 NS_720 0 1.9189093155368882e-05
GC_9_721 b_9 NI_9 NS_721 0 1.6096905621929843e-04
GC_9_722 b_9 NI_9 NS_722 0 4.2091214227818306e-05
GC_9_723 b_9 NI_9 NS_723 0 -8.8878044591827137e-05
GC_9_724 b_9 NI_9 NS_724 0 -7.1909596477119791e-05
GC_9_725 b_9 NI_9 NS_725 0 -8.4867036650296648e-05
GC_9_726 b_9 NI_9 NS_726 0 6.3596361194763232e-05
GC_9_727 b_9 NI_9 NS_727 0 1.4068805490001222e-04
GC_9_728 b_9 NI_9 NS_728 0 -4.8518768208045298e-05
GC_9_729 b_9 NI_9 NS_729 0 -6.6207482886684264e-05
GC_9_730 b_9 NI_9 NS_730 0 -2.4250999784955779e-05
GC_9_731 b_9 NI_9 NS_731 0 6.1223509819438707e-05
GC_9_732 b_9 NI_9 NS_732 0 1.1375862113409609e-04
GC_9_733 b_9 NI_9 NS_733 0 -2.2917088222844084e-05
GC_9_734 b_9 NI_9 NS_734 0 -1.2153227439627769e-04
GC_9_735 b_9 NI_9 NS_735 0 -4.4313564574161660e-05
GC_9_736 b_9 NI_9 NS_736 0 1.0975035360452003e-05
GC_9_737 b_9 NI_9 NS_737 0 4.7535487241914023e-05
GC_9_738 b_9 NI_9 NS_738 0 -1.0607214805147562e-05
GC_9_739 b_9 NI_9 NS_739 0 -3.2085902361709370e-05
GC_9_740 b_9 NI_9 NS_740 0 -7.6432280925047340e-06
GC_9_741 b_9 NI_9 NS_741 0 2.1333531667399173e-05
GC_9_742 b_9 NI_9 NS_742 0 -4.8743868926557540e-06
GC_9_743 b_9 NI_9 NS_743 0 -3.2213590106332131e-05
GC_9_744 b_9 NI_9 NS_744 0 -2.5250789836834344e-05
GC_9_745 b_9 NI_9 NS_745 0 1.2710110264235127e-05
GC_9_746 b_9 NI_9 NS_746 0 6.1771582056737315e-06
GC_9_747 b_9 NI_9 NS_747 0 -2.0359017600187088e-05
GC_9_748 b_9 NI_9 NS_748 0 -7.7253059824133583e-06
GC_9_749 b_9 NI_9 NS_749 0 1.4086578732068812e-05
GC_9_750 b_9 NI_9 NS_750 0 -1.2504410464230536e-05
GC_9_751 b_9 NI_9 NS_751 0 -4.1282285568715805e-05
GC_9_752 b_9 NI_9 NS_752 0 -1.6953796259810693e-05
GC_9_753 b_9 NI_9 NS_753 0 1.1907504429253589e-05
GC_9_754 b_9 NI_9 NS_754 0 -1.7646396340481041e-06
GC_9_755 b_9 NI_9 NS_755 0 -3.0212458185786954e-05
GC_9_756 b_9 NI_9 NS_756 0 5.5333503981953081e-06
GC_9_757 b_9 NI_9 NS_757 0 1.6332648134970693e-05
GC_9_758 b_9 NI_9 NS_758 0 -2.0848592863771101e-05
GC_9_759 b_9 NI_9 NS_759 0 -4.9846288199787694e-05
GC_9_760 b_9 NI_9 NS_760 0 -1.6673744434439334e-06
GC_9_761 b_9 NI_9 NS_761 0 1.2247660070390668e-05
GC_9_762 b_9 NI_9 NS_762 0 -1.1717554861033940e-05
GC_9_763 b_9 NI_9 NS_763 0 -3.1908583509642189e-05
GC_9_764 b_9 NI_9 NS_764 0 2.5076450782497340e-05
GC_9_765 b_9 NI_9 NS_765 0 1.0834703979254268e-05
GC_9_766 b_9 NI_9 NS_766 0 -3.6496291107583871e-05
GC_9_767 b_9 NI_9 NS_767 0 -3.3856381860245982e-05
GC_9_768 b_9 NI_9 NS_768 0 1.8659164687801176e-05
GC_9_769 b_9 NI_9 NS_769 0 -5.9880013340861418e-05
GC_9_770 b_9 NI_9 NS_770 0 1.2847674079849642e-04
GC_9_771 b_9 NI_9 NS_771 0 -1.4511895179767261e-05
GC_9_772 b_9 NI_9 NS_772 0 -3.3369944737033570e-05
GC_9_773 b_9 NI_9 NS_773 0 -3.8791635358639323e-07
GC_9_774 b_9 NI_9 NS_774 0 3.6149788086291819e-07
GC_9_775 b_9 NI_9 NS_775 0 -1.9685610970556193e-05
GC_9_776 b_9 NI_9 NS_776 0 3.1289659338478825e-05
GC_9_777 b_9 NI_9 NS_777 0 -1.4243119222898966e-05
GC_9_778 b_9 NI_9 NS_778 0 -3.4196323239830453e-05
GC_9_779 b_9 NI_9 NS_779 0 -5.2921636740680719e-06
GC_9_780 b_9 NI_9 NS_780 0 5.5312280427685286e-06
GC_9_781 b_9 NI_9 NS_781 0 -1.9744698216205799e-05
GC_9_782 b_9 NI_9 NS_782 0 -6.5467805116979557e-05
GC_9_783 b_9 NI_9 NS_783 0 -9.2827092835254154e-06
GC_9_784 b_9 NI_9 NS_784 0 -2.0586529974831130e-05
GC_9_785 b_9 NI_9 NS_785 0 1.4777870461459807e-05
GC_9_786 b_9 NI_9 NS_786 0 2.2998461536047660e-05
GC_9_787 b_9 NI_9 NS_787 0 -6.8230582173235474e-06
GC_9_788 b_9 NI_9 NS_788 0 2.7592666302804021e-05
GC_9_789 b_9 NI_9 NS_789 0 -1.1135794198431711e-05
GC_9_790 b_9 NI_9 NS_790 0 -2.1577734503456304e-05
GC_9_791 b_9 NI_9 NS_791 0 -1.1024480213497236e-05
GC_9_792 b_9 NI_9 NS_792 0 2.3799332084794695e-05
GC_9_793 b_9 NI_9 NS_793 0 5.1499150393213775e-06
GC_9_794 b_9 NI_9 NS_794 0 -1.5352049763299690e-05
GC_9_795 b_9 NI_9 NS_795 0 -4.7264134361070035e-10
GC_9_796 b_9 NI_9 NS_796 0 -9.1861893162232335e-10
GC_9_797 b_9 NI_9 NS_797 0 -5.5411895922706338e-08
GC_9_798 b_9 NI_9 NS_798 0 7.6386903231283359e-09
GC_9_799 b_9 NI_9 NS_799 0 -2.0271395629829937e-04
GC_9_800 b_9 NI_9 NS_800 0 -3.3244175924956220e-06
GC_9_801 b_9 NI_9 NS_801 0 1.2949636216449736e-09
GC_9_802 b_9 NI_9 NS_802 0 9.6759077370154610e-09
GC_9_803 b_9 NI_9 NS_803 0 -4.1591754547047806e-06
GC_9_804 b_9 NI_9 NS_804 0 6.1862101862746297e-06
GC_9_805 b_9 NI_9 NS_805 0 3.8149382468788006e-06
GC_9_806 b_9 NI_9 NS_806 0 -8.1670905625712377e-06
GC_9_807 b_9 NI_9 NS_807 0 2.1690372977876439e-05
GC_9_808 b_9 NI_9 NS_808 0 -8.8399936853455309e-06
GC_9_809 b_9 NI_9 NS_809 0 -2.1479597125376220e-05
GC_9_810 b_9 NI_9 NS_810 0 -1.1874160555393425e-06
GC_9_811 b_9 NI_9 NS_811 0 -2.9640112064710980e-05
GC_9_812 b_9 NI_9 NS_812 0 -2.8295816058086235e-05
GC_9_813 b_9 NI_9 NS_813 0 -5.5412967258959538e-06
GC_9_814 b_9 NI_9 NS_814 0 1.6551987631820488e-05
GC_9_815 b_9 NI_9 NS_815 0 -2.4251880926817803e-06
GC_9_816 b_9 NI_9 NS_816 0 -7.1420268227042728e-06
GC_9_817 b_9 NI_9 NS_817 0 -2.2563456823229988e-05
GC_9_818 b_9 NI_9 NS_818 0 6.0026112560841037e-06
GC_9_819 b_9 NI_9 NS_819 0 -1.8565791723484809e-04
GC_9_820 b_9 NI_9 NS_820 0 -4.4043359180835937e-05
GC_9_821 b_9 NI_9 NS_821 0 6.2654398652927293e-05
GC_9_822 b_9 NI_9 NS_822 0 1.3744256670250067e-04
GC_9_823 b_9 NI_9 NS_823 0 -3.7291592346985894e-05
GC_9_824 b_9 NI_9 NS_824 0 5.6617736579859759e-05
GC_9_825 b_9 NI_9 NS_825 0 9.5234335804650312e-05
GC_9_826 b_9 NI_9 NS_826 0 2.4609659172899323e-04
GC_9_827 b_9 NI_9 NS_827 0 7.3806894491534246e-05
GC_9_828 b_9 NI_9 NS_828 0 4.9082670123317865e-07
GC_9_829 b_9 NI_9 NS_829 0 -1.5390450466594070e-05
GC_9_830 b_9 NI_9 NS_830 0 2.6127685596432742e-04
GC_9_831 b_9 NI_9 NS_831 0 3.6437419922651391e-04
GC_9_832 b_9 NI_9 NS_832 0 -2.4319841990975348e-04
GC_9_833 b_9 NI_9 NS_833 0 6.5655663518363850e-05
GC_9_834 b_9 NI_9 NS_834 0 -2.8529427648368521e-05
GC_9_835 b_9 NI_9 NS_835 0 2.0802593282129869e-04
GC_9_836 b_9 NI_9 NS_836 0 -2.4142800817523056e-04
GC_9_837 b_9 NI_9 NS_837 0 -7.1299257933555383e-05
GC_9_838 b_9 NI_9 NS_838 0 -7.1473439059096370e-05
GC_9_839 b_9 NI_9 NS_839 0 6.4494182101323667e-05
GC_9_840 b_9 NI_9 NS_840 0 -7.5537527403650909e-05
GC_9_841 b_9 NI_9 NS_841 0 -1.7050086732385352e-04
GC_9_842 b_9 NI_9 NS_842 0 -1.8310153275563076e-04
GC_9_843 b_9 NI_9 NS_843 0 -4.8839023883619615e-05
GC_9_844 b_9 NI_9 NS_844 0 -1.9100995302381975e-05
GC_9_845 b_9 NI_9 NS_845 0 -1.4492616903145106e-04
GC_9_846 b_9 NI_9 NS_846 0 -9.5351252515488732e-05
GC_9_847 b_9 NI_9 NS_847 0 -2.7319737386285937e-05
GC_9_848 b_9 NI_9 NS_848 0 1.0361197516217643e-04
GC_9_849 b_9 NI_9 NS_849 0 -2.7244445933269340e-05
GC_9_850 b_9 NI_9 NS_850 0 1.3907007011413342e-05
GC_9_851 b_9 NI_9 NS_851 0 2.1287337531585146e-06
GC_9_852 b_9 NI_9 NS_852 0 5.0767896369590149e-05
GC_9_853 b_9 NI_9 NS_853 0 1.6812848385784751e-05
GC_9_854 b_9 NI_9 NS_854 0 -5.9689891335742856e-07
GC_9_855 b_9 NI_9 NS_855 0 1.8078608279852651e-06
GC_9_856 b_9 NI_9 NS_856 0 -1.5453788161766764e-05
GC_9_857 b_9 NI_9 NS_857 0 -1.5113187240414338e-05
GC_9_858 b_9 NI_9 NS_858 0 -1.3588621551507399e-05
GC_9_859 b_9 NI_9 NS_859 0 -1.3111062599273459e-05
GC_9_860 b_9 NI_9 NS_860 0 1.2341202908884042e-05
GC_9_861 b_9 NI_9 NS_861 0 7.7832677419489880e-06
GC_9_862 b_9 NI_9 NS_862 0 1.2547280385262837e-06
GC_9_863 b_9 NI_9 NS_863 0 -5.1390801744667134e-06
GC_9_864 b_9 NI_9 NS_864 0 -1.2684886035808820e-05
GC_9_865 b_9 NI_9 NS_865 0 -2.0804835573902417e-05
GC_9_866 b_9 NI_9 NS_866 0 -5.8777168802151124e-06
GC_9_867 b_9 NI_9 NS_867 0 1.0778170013178657e-06
GC_9_868 b_9 NI_9 NS_868 0 2.1822123226377052e-05
GC_9_869 b_9 NI_9 NS_869 0 1.2864917405110838e-05
GC_9_870 b_9 NI_9 NS_870 0 -6.8616166917291685e-06
GC_9_871 b_9 NI_9 NS_871 0 -1.7284502591349766e-05
GC_9_872 b_9 NI_9 NS_872 0 -1.5979339663017199e-05
GC_9_873 b_9 NI_9 NS_873 0 -2.7118177652407545e-05
GC_9_874 b_9 NI_9 NS_874 0 8.8177797173729246e-06
GC_9_875 b_9 NI_9 NS_875 0 2.7091322514565258e-05
GC_9_876 b_9 NI_9 NS_876 0 2.2446901713034642e-05
GC_9_877 b_9 NI_9 NS_877 0 1.0942483284829456e-05
GC_9_878 b_9 NI_9 NS_878 0 -2.1302974664990888e-05
GC_9_879 b_9 NI_9 NS_879 0 -3.0617345600692943e-05
GC_9_880 b_9 NI_9 NS_880 0 3.9057790333557822e-06
GC_9_881 b_9 NI_9 NS_881 0 -9.8014557642786325e-06
GC_9_882 b_9 NI_9 NS_882 0 3.9251519218311006e-05
GC_9_883 b_9 NI_9 NS_883 0 1.9727815383755191e-05
GC_9_884 b_9 NI_9 NS_884 0 -6.8538563139313921e-05
GC_9_885 b_9 NI_9 NS_885 0 4.3399502764889287e-05
GC_9_886 b_9 NI_9 NS_886 0 -1.6869780486635635e-05
GC_9_887 b_9 NI_9 NS_887 0 2.0639883388727416e-07
GC_9_888 b_9 NI_9 NS_888 0 -2.4347731128300852e-07
GC_9_889 b_9 NI_9 NS_889 0 -3.6328478973457061e-06
GC_9_890 b_9 NI_9 NS_890 0 -2.0833670420738715e-05
GC_9_891 b_9 NI_9 NS_891 0 -1.0494376367860393e-05
GC_9_892 b_9 NI_9 NS_892 0 1.6698425758771590e-05
GC_9_893 b_9 NI_9 NS_893 0 9.1959643311532291e-06
GC_9_894 b_9 NI_9 NS_894 0 3.1866766130015869e-05
GC_9_895 b_9 NI_9 NS_895 0 1.4280789164291849e-05
GC_9_896 b_9 NI_9 NS_896 0 -3.0127252865069539e-06
GC_9_897 b_9 NI_9 NS_897 0 -3.9054310069770812e-06
GC_9_898 b_9 NI_9 NS_898 0 1.2499911281703533e-05
GC_9_899 b_9 NI_9 NS_899 0 -1.8574401620682487e-05
GC_9_900 b_9 NI_9 NS_900 0 -3.6262128898118571e-06
GC_9_901 b_9 NI_9 NS_901 0 1.3215555748716720e-05
GC_9_902 b_9 NI_9 NS_902 0 1.3176894543390360e-05
GC_9_903 b_9 NI_9 NS_903 0 7.6361524721940174e-06
GC_9_904 b_9 NI_9 NS_904 0 -2.3019338603021633e-05
GC_9_905 b_9 NI_9 NS_905 0 -3.8459167588114109e-06
GC_9_906 b_9 NI_9 NS_906 0 -1.1723218562468101e-05
GC_9_907 b_9 NI_9 NS_907 0 -8.7362100402485138e-06
GC_9_908 b_9 NI_9 NS_908 0 -2.6280717205871715e-06
GC_9_909 b_9 NI_9 NS_909 0 5.5146430931088508e-10
GC_9_910 b_9 NI_9 NS_910 0 2.9343860916888240e-10
GC_9_911 b_9 NI_9 NS_911 0 4.2107599594299634e-08
GC_9_912 b_9 NI_9 NS_912 0 3.6940438347326653e-08
GC_9_913 b_9 NI_9 NS_913 0 -1.4190176474161331e-02
GC_9_914 b_9 NI_9 NS_914 0 1.3879312341883402e-03
GC_9_915 b_9 NI_9 NS_915 0 -2.6214184849954014e-07
GC_9_916 b_9 NI_9 NS_916 0 -3.7469278865740603e-06
GC_9_917 b_9 NI_9 NS_917 0 -2.9950674534552830e-04
GC_9_918 b_9 NI_9 NS_918 0 4.7112893106086818e-04
GC_9_919 b_9 NI_9 NS_919 0 1.2936046057261958e-03
GC_9_920 b_9 NI_9 NS_920 0 5.6342157087523937e-04
GC_9_921 b_9 NI_9 NS_921 0 -2.7928160469021918e-03
GC_9_922 b_9 NI_9 NS_922 0 -7.1086069176877465e-04
GC_9_923 b_9 NI_9 NS_923 0 3.5977253048659328e-03
GC_9_924 b_9 NI_9 NS_924 0 2.5454524034539084e-03
GC_9_925 b_9 NI_9 NS_925 0 1.1770634223605939e-03
GC_9_926 b_9 NI_9 NS_926 0 -4.1367913016178504e-03
GC_9_927 b_9 NI_9 NS_927 0 -1.5549027037856109e-03
GC_9_928 b_9 NI_9 NS_928 0 2.7530000456521962e-03
GC_9_929 b_9 NI_9 NS_929 0 -3.5992331282820242e-04
GC_9_930 b_9 NI_9 NS_930 0 -2.1737589242779612e-04
GC_9_931 b_9 NI_9 NS_931 0 4.0014065019016026e-03
GC_9_932 b_9 NI_9 NS_932 0 2.5737097308870980e-04
GC_9_933 b_9 NI_9 NS_933 0 -7.3983847206872087e-03
GC_9_934 b_9 NI_9 NS_934 0 -1.3542082509394066e-02
GC_9_935 b_9 NI_9 NS_935 0 4.4843114449703864e-03
GC_9_936 b_9 NI_9 NS_936 0 1.3402112655174981e-02
GC_9_937 b_9 NI_9 NS_937 0 6.7170369768760506e-03
GC_9_938 b_9 NI_9 NS_938 0 -4.0292270424362592e-03
GC_9_939 b_9 NI_9 NS_939 0 -1.3321389325133588e-02
GC_9_940 b_9 NI_9 NS_940 0 6.8614134659124987e-04
GC_9_941 b_9 NI_9 NS_941 0 7.8581326391371671e-03
GC_9_942 b_9 NI_9 NS_942 0 1.8345297311054183e-03
GC_9_943 b_9 NI_9 NS_943 0 1.0514012606221389e-02
GC_9_944 b_9 NI_9 NS_944 0 -1.9642833995147824e-02
GC_9_945 b_9 NI_9 NS_945 0 -1.7746430659650599e-02
GC_9_946 b_9 NI_9 NS_946 0 1.9129850712233349e-02
GC_9_947 b_9 NI_9 NS_947 0 7.6846929972949393e-03
GC_9_948 b_9 NI_9 NS_948 0 -1.4647961343414878e-03
GC_9_949 b_9 NI_9 NS_949 0 -1.5663695356294131e-02
GC_9_950 b_9 NI_9 NS_950 0 -4.7646585392284585e-03
GC_9_951 b_9 NI_9 NS_951 0 8.0859975997433758e-03
GC_9_952 b_9 NI_9 NS_952 0 7.2458392344718070e-03
GC_9_953 b_9 NI_9 NS_953 0 8.1137527442081674e-03
GC_9_954 b_9 NI_9 NS_954 0 -6.0473592427647800e-03
GC_9_955 b_9 NI_9 NS_955 0 -1.3987009841277456e-02
GC_9_956 b_9 NI_9 NS_956 0 4.5767044118306200e-03
GC_9_957 b_9 NI_9 NS_957 0 6.2436878133990837e-03
GC_9_958 b_9 NI_9 NS_958 0 2.3779886766406759e-03
GC_9_959 b_9 NI_9 NS_959 0 -6.3098266680049805e-03
GC_9_960 b_9 NI_9 NS_960 0 -1.1127813894253881e-02
GC_9_961 b_9 NI_9 NS_961 0 2.1503507497208532e-03
GC_9_962 b_9 NI_9 NS_962 0 1.1938066038686362e-02
GC_9_963 b_9 NI_9 NS_963 0 4.2146509118331978e-03
GC_9_964 b_9 NI_9 NS_964 0 -1.1800115880074085e-03
GC_9_965 b_9 NI_9 NS_965 0 -4.9267465127460471e-03
GC_9_966 b_9 NI_9 NS_966 0 1.0434789746039490e-03
GC_9_967 b_9 NI_9 NS_967 0 3.0295918234717590e-03
GC_9_968 b_9 NI_9 NS_968 0 6.8509421433343427e-04
GC_9_969 b_9 NI_9 NS_969 0 -2.2185442028713788e-03
GC_9_970 b_9 NI_9 NS_970 0 4.8987925557770421e-04
GC_9_971 b_9 NI_9 NS_971 0 3.0814366936513802e-03
GC_9_972 b_9 NI_9 NS_972 0 2.2937712263651944e-03
GC_9_973 b_9 NI_9 NS_973 0 -1.5261903156410220e-03
GC_9_974 b_9 NI_9 NS_974 0 -6.8311090771638785e-04
GC_9_975 b_9 NI_9 NS_975 0 1.8943367520300959e-03
GC_9_976 b_9 NI_9 NS_976 0 6.7631629385852903e-04
GC_9_977 b_9 NI_9 NS_977 0 -1.5560125360784798e-03
GC_9_978 b_9 NI_9 NS_978 0 1.2187771813988782e-03
GC_9_979 b_9 NI_9 NS_979 0 3.9927828059971807e-03
GC_9_980 b_9 NI_9 NS_980 0 1.4034832744516481e-03
GC_9_981 b_9 NI_9 NS_981 0 -1.5356518598095947e-03
GC_9_982 b_9 NI_9 NS_982 0 5.9546630884189944e-05
GC_9_983 b_9 NI_9 NS_983 0 2.8410943534162890e-03
GC_9_984 b_9 NI_9 NS_984 0 -6.9178251938510551e-04
GC_9_985 b_9 NI_9 NS_985 0 -1.8626304934044279e-03
GC_9_986 b_9 NI_9 NS_986 0 1.9986019937520113e-03
GC_9_987 b_9 NI_9 NS_987 0 4.9308339550331592e-03
GC_9_988 b_9 NI_9 NS_988 0 -1.7294296437696615e-04
GC_9_989 b_9 NI_9 NS_989 0 -1.6210911037052920e-03
GC_9_990 b_9 NI_9 NS_990 0 9.0628766643394804e-04
GC_9_991 b_9 NI_9 NS_991 0 3.0921542848532458e-03
GC_9_992 b_9 NI_9 NS_992 0 -2.8475023084149451e-03
GC_9_993 b_9 NI_9 NS_993 0 -1.4246678020848173e-03
GC_9_994 b_9 NI_9 NS_994 0 3.1958012338290944e-03
GC_9_995 b_9 NI_9 NS_995 0 3.8550219538652257e-03
GC_9_996 b_9 NI_9 NS_996 0 -2.9522299049287055e-03
GC_9_997 b_9 NI_9 NS_997 0 -2.0071714227067401e-03
GC_9_998 b_9 NI_9 NS_998 0 -4.1861199998799378e-03
GC_9_999 b_9 NI_9 NS_999 0 -3.5103813548552977e-04
GC_9_1000 b_9 NI_9 NS_1000 0 2.2864621989012912e-03
GC_9_1001 b_9 NI_9 NS_1001 0 -1.0763404492469775e-05
GC_9_1002 b_9 NI_9 NS_1002 0 -2.3358512622479606e-05
GC_9_1003 b_9 NI_9 NS_1003 0 8.7769872405550598e-04
GC_9_1004 b_9 NI_9 NS_1004 0 -3.8352110073250028e-03
GC_9_1005 b_9 NI_9 NS_1005 0 3.5234250997916085e-04
GC_9_1006 b_9 NI_9 NS_1006 0 3.3067871907684052e-03
GC_9_1007 b_9 NI_9 NS_1007 0 1.3988574453094251e-03
GC_9_1008 b_9 NI_9 NS_1008 0 -2.3422177521989799e-03
GC_9_1009 b_9 NI_9 NS_1009 0 2.2595473446470238e-03
GC_9_1010 b_9 NI_9 NS_1010 0 3.3689502297269041e-03
GC_9_1011 b_9 NI_9 NS_1011 0 1.1614261634618061e-03
GC_9_1012 b_9 NI_9 NS_1012 0 2.4048209520122726e-03
GC_9_1013 b_9 NI_9 NS_1013 0 -8.2758772881358844e-04
GC_9_1014 b_9 NI_9 NS_1014 0 -1.9684509236774237e-03
GC_9_1015 b_9 NI_9 NS_1015 0 3.9845160819744718e-04
GC_9_1016 b_9 NI_9 NS_1016 0 -2.6910251894529313e-03
GC_9_1017 b_9 NI_9 NS_1017 0 9.7822682465522259e-04
GC_9_1018 b_9 NI_9 NS_1018 0 2.7413561725081704e-03
GC_9_1019 b_9 NI_9 NS_1019 0 1.0427102867671349e-03
GC_9_1020 b_9 NI_9 NS_1020 0 -2.4233095739191863e-03
GC_9_1021 b_9 NI_9 NS_1021 0 -1.0796390318191177e-03
GC_9_1022 b_9 NI_9 NS_1022 0 1.5897876532715682e-03
GC_9_1023 b_9 NI_9 NS_1023 0 -1.0823809464560397e-08
GC_9_1024 b_9 NI_9 NS_1024 0 -2.6612215031517179e-09
GC_9_1025 b_9 NI_9 NS_1025 0 2.3026014584190990e-06
GC_9_1026 b_9 NI_9 NS_1026 0 5.5056631416519076e-07
GC_9_1027 b_9 NI_9 NS_1027 0 1.8435412401579032e-02
GC_9_1028 b_9 NI_9 NS_1028 0 6.7474797529250008e-03
GC_9_1029 b_9 NI_9 NS_1029 0 4.6857917199005810e-07
GC_9_1030 b_9 NI_9 NS_1030 0 1.4597152662160697e-06
GC_9_1031 b_9 NI_9 NS_1031 0 6.0883563693663106e-03
GC_9_1032 b_9 NI_9 NS_1032 0 1.8079697378841103e-03
GC_9_1033 b_9 NI_9 NS_1033 0 -6.0692939311995679e-03
GC_9_1034 b_9 NI_9 NS_1034 0 -6.1755323612633633e-04
GC_9_1035 b_9 NI_9 NS_1035 0 7.3052495337176818e-03
GC_9_1036 b_9 NI_9 NS_1036 0 -1.2868624997723349e-02
GC_9_1037 b_9 NI_9 NS_1037 0 8.4478397845725080e-03
GC_9_1038 b_9 NI_9 NS_1038 0 -2.4318216813365757e-04
GC_9_1039 b_9 NI_9 NS_1039 0 -9.6437745087863420e-03
GC_9_1040 b_9 NI_9 NS_1040 0 2.6145169223877386e-03
GC_9_1041 b_9 NI_9 NS_1041 0 -8.8623538353725419e-03
GC_9_1042 b_9 NI_9 NS_1042 0 -2.4394274563080073e-02
GC_9_1043 b_9 NI_9 NS_1043 0 -8.6173540188209160e-04
GC_9_1044 b_9 NI_9 NS_1044 0 4.1811215342885998e-03
GC_9_1045 b_9 NI_9 NS_1045 0 7.1873632449022673e-03
GC_9_1046 b_9 NI_9 NS_1046 0 -1.0295225277454480e-03
GC_9_1047 b_9 NI_9 NS_1047 0 -2.5161203599690620e-02
GC_9_1048 b_9 NI_9 NS_1048 0 4.8304218498001136e-03
GC_9_1049 b_9 NI_9 NS_1049 0 -1.9677166603242386e-02
GC_9_1050 b_9 NI_9 NS_1050 0 8.9700837900282590e-04
GC_9_1051 b_9 NI_9 NS_1051 0 1.0760342813884747e-02
GC_9_1052 b_9 NI_9 NS_1052 0 -2.7834959874194149e-03
GC_9_1053 b_9 NI_9 NS_1053 0 -4.7877934427124850e-03
GC_9_1054 b_9 NI_9 NS_1054 0 4.5022521267384222e-02
GC_9_1055 b_9 NI_9 NS_1055 0 -1.2656477991338434e-02
GC_9_1056 b_9 NI_9 NS_1056 0 -2.7337493562051683e-04
GC_9_1057 b_9 NI_9 NS_1057 0 1.5916673587996606e-02
GC_9_1058 b_9 NI_9 NS_1058 0 -4.0521710780090049e-03
GC_9_1059 b_9 NI_9 NS_1059 0 3.2201056380365710e-02
GC_9_1060 b_9 NI_9 NS_1060 0 1.8584910760078243e-02
GC_9_1061 b_9 NI_9 NS_1061 0 -1.2597870748215459e-02
GC_9_1062 b_9 NI_9 NS_1062 0 1.6058531755385052e-04
GC_9_1063 b_9 NI_9 NS_1063 0 1.7204454051842139e-02
GC_9_1064 b_9 NI_9 NS_1064 0 -3.5162914624202644e-02
GC_9_1065 b_9 NI_9 NS_1065 0 1.4015912178214728e-02
GC_9_1066 b_9 NI_9 NS_1066 0 4.7859288565677274e-03
GC_9_1067 b_9 NI_9 NS_1067 0 -1.4402608782691693e-02
GC_9_1068 b_9 NI_9 NS_1068 0 2.3858803247397013e-04
GC_9_1069 b_9 NI_9 NS_1069 0 -2.0144316656752162e-02
GC_9_1070 b_9 NI_9 NS_1070 0 -3.0186671502125666e-02
GC_9_1071 b_9 NI_9 NS_1071 0 1.0530823242429047e-02
GC_9_1072 b_9 NI_9 NS_1072 0 3.5935710975885473e-03
GC_9_1073 b_9 NI_9 NS_1073 0 -2.6797802179773046e-02
GC_9_1074 b_9 NI_9 NS_1074 0 1.1150563015180862e-02
GC_9_1075 b_9 NI_9 NS_1075 0 -1.4133808841566165e-02
GC_9_1076 b_9 NI_9 NS_1076 0 -2.5194655416744646e-03
GC_9_1077 b_9 NI_9 NS_1077 0 7.5552555789602177e-03
GC_9_1078 b_9 NI_9 NS_1078 0 1.5923973161430026e-03
GC_9_1079 b_9 NI_9 NS_1079 0 -8.5552848479123606e-04
GC_9_1080 b_9 NI_9 NS_1080 0 2.4403185070971518e-02
GC_9_1081 b_9 NI_9 NS_1081 0 -7.6201582359672311e-03
GC_9_1082 b_9 NI_9 NS_1082 0 2.8214473281528752e-04
GC_9_1083 b_9 NI_9 NS_1083 0 -5.5977007458570319e-04
GC_9_1084 b_9 NI_9 NS_1084 0 -5.5368534776433671e-03
GC_9_1085 b_9 NI_9 NS_1085 0 8.2660198609056726e-03
GC_9_1086 b_9 NI_9 NS_1086 0 7.0201649795975027e-03
GC_9_1087 b_9 NI_9 NS_1087 0 -7.1913673292448043e-04
GC_9_1088 b_9 NI_9 NS_1088 0 1.2092542130593447e-02
GC_9_1089 b_9 NI_9 NS_1089 0 -5.1474202836320161e-03
GC_9_1090 b_9 NI_9 NS_1090 0 -1.3697057642152481e-04
GC_9_1091 b_9 NI_9 NS_1091 0 -1.8303673921581086e-03
GC_9_1092 b_9 NI_9 NS_1092 0 -5.1700312801403209e-03
GC_9_1093 b_9 NI_9 NS_1093 0 9.2878948415415427e-03
GC_9_1094 b_9 NI_9 NS_1094 0 5.4155078209547260e-03
GC_9_1095 b_9 NI_9 NS_1095 0 3.5153192734402971e-03
GC_9_1096 b_9 NI_9 NS_1096 0 1.1689902301887689e-02
GC_9_1097 b_9 NI_9 NS_1097 0 -6.1369968679813036e-03
GC_9_1098 b_9 NI_9 NS_1098 0 1.4286839696451726e-03
GC_9_1099 b_9 NI_9 NS_1099 0 -2.8171450948823585e-03
GC_9_1100 b_9 NI_9 NS_1100 0 -7.3461609234601113e-03
GC_9_1101 b_9 NI_9 NS_1101 0 9.9560514722193474e-03
GC_9_1102 b_9 NI_9 NS_1102 0 3.3690008335945138e-03
GC_9_1103 b_9 NI_9 NS_1103 0 8.1686478330978782e-03
GC_9_1104 b_9 NI_9 NS_1104 0 1.0244265668732743e-02
GC_9_1105 b_9 NI_9 NS_1105 0 -6.9844909552791027e-03
GC_9_1106 b_9 NI_9 NS_1106 0 2.9356666602424995e-03
GC_9_1107 b_9 NI_9 NS_1107 0 -5.6335165515931547e-03
GC_9_1108 b_9 NI_9 NS_1108 0 -8.0963389495466338e-03
GC_9_1109 b_9 NI_9 NS_1109 0 9.8582264347487226e-03
GC_9_1110 b_9 NI_9 NS_1110 0 5.4666337857154745e-04
GC_9_1111 b_9 NI_9 NS_1111 0 -1.0938596974803852e-02
GC_9_1112 b_9 NI_9 NS_1112 0 1.2297963480667482e-02
GC_9_1113 b_9 NI_9 NS_1113 0 9.6448399365143891e-03
GC_9_1114 b_9 NI_9 NS_1114 0 5.0354163388920880e-03
GC_9_1115 b_9 NI_9 NS_1115 0 -1.9866494684974064e-05
GC_9_1116 b_9 NI_9 NS_1116 0 3.1663139722552625e-05
GC_9_1117 b_9 NI_9 NS_1117 0 -7.1316248431642559e-03
GC_9_1118 b_9 NI_9 NS_1118 0 4.4780553837691691e-03
GC_9_1119 b_9 NI_9 NS_1119 0 -7.6761507357491808e-03
GC_9_1120 b_9 NI_9 NS_1120 0 -5.3212201426376714e-03
GC_9_1121 b_9 NI_9 NS_1121 0 9.5161718411133130e-03
GC_9_1122 b_9 NI_9 NS_1122 0 -1.7356724710185214e-03
GC_9_1123 b_9 NI_9 NS_1123 0 1.2474751026288526e-02
GC_9_1124 b_9 NI_9 NS_1124 0 -1.4037761675371708e-03
GC_9_1125 b_9 NI_9 NS_1125 0 -5.0717230645196485e-03
GC_9_1126 b_9 NI_9 NS_1126 0 -2.7497988181118755e-03
GC_9_1127 b_9 NI_9 NS_1127 0 -2.2245921531921942e-03
GC_9_1128 b_9 NI_9 NS_1128 0 6.6015856511003274e-03
GC_9_1129 b_9 NI_9 NS_1129 0 8.9572659788627780e-03
GC_9_1130 b_9 NI_9 NS_1130 0 1.3090365551121915e-04
GC_9_1131 b_9 NI_9 NS_1131 0 1.2487382878024547e-02
GC_9_1132 b_9 NI_9 NS_1132 0 1.7799311417201679e-03
GC_9_1133 b_9 NI_9 NS_1133 0 -5.3780365813402920e-03
GC_9_1134 b_9 NI_9 NS_1134 0 4.1549170169347957e-03
GC_9_1135 b_9 NI_9 NS_1135 0 -1.8499128776165565e-03
GC_9_1136 b_9 NI_9 NS_1136 0 -5.6869431369817505e-03
GC_9_1137 b_9 NI_9 NS_1137 0 2.0796303167458877e-07
GC_9_1138 b_9 NI_9 NS_1138 0 -2.4555623362992996e-07
GC_9_1139 b_9 NI_9 NS_1139 0 -1.1509981861677499e-05
GC_9_1140 b_9 NI_9 NS_1140 0 1.8244024752520902e-05
GC_9_1141 b_9 NI_9 NS_1141 0 7.7517847499608845e-03
GC_9_1142 b_9 NI_9 NS_1142 0 -1.6012309488679694e-03
GC_9_1143 b_9 NI_9 NS_1143 0 -1.2107357777314372e-08
GC_9_1144 b_9 NI_9 NS_1144 0 -8.8419733076257476e-07
GC_9_1145 b_9 NI_9 NS_1145 0 1.0389334678028366e-04
GC_9_1146 b_9 NI_9 NS_1146 0 -5.1165497914145764e-04
GC_9_1147 b_9 NI_9 NS_1147 0 -1.9366722490408849e-03
GC_9_1148 b_9 NI_9 NS_1148 0 -5.9740611531011137e-04
GC_9_1149 b_9 NI_9 NS_1149 0 2.9415496646430423e-03
GC_9_1150 b_9 NI_9 NS_1150 0 2.2646150034270614e-03
GC_9_1151 b_9 NI_9 NS_1151 0 -3.5699560029924934e-03
GC_9_1152 b_9 NI_9 NS_1152 0 -3.0486859049661925e-03
GC_9_1153 b_9 NI_9 NS_1153 0 -1.7071461899151111e-03
GC_9_1154 b_9 NI_9 NS_1154 0 5.8436823019136089e-03
GC_9_1155 b_9 NI_9 NS_1155 0 4.3687526632737190e-03
GC_9_1156 b_9 NI_9 NS_1156 0 -2.4746080186935685e-03
GC_9_1157 b_9 NI_9 NS_1157 0 -1.1051345529904771e-04
GC_9_1158 b_9 NI_9 NS_1158 0 -1.0368748323563517e-04
GC_9_1159 b_9 NI_9 NS_1159 0 -4.4520077614423658e-03
GC_9_1160 b_9 NI_9 NS_1160 0 -9.2458271011419332e-04
GC_9_1161 b_9 NI_9 NS_1161 0 9.1257545990907282e-03
GC_9_1162 b_9 NI_9 NS_1162 0 1.7785323756131934e-02
GC_9_1163 b_9 NI_9 NS_1163 0 -4.0274383895288991e-03
GC_9_1164 b_9 NI_9 NS_1164 0 -1.7847938779752246e-02
GC_9_1165 b_9 NI_9 NS_1165 0 -8.2175426840410473e-03
GC_9_1166 b_9 NI_9 NS_1166 0 4.1736400791746479e-03
GC_9_1167 b_9 NI_9 NS_1167 0 1.7064437340059704e-02
GC_9_1168 b_9 NI_9 NS_1168 0 -4.4006004129423527e-04
GC_9_1169 b_9 NI_9 NS_1169 0 -9.2787957944338081e-03
GC_9_1170 b_9 NI_9 NS_1170 0 -3.2071931228856323e-03
GC_9_1171 b_9 NI_9 NS_1171 0 -1.3712649598662351e-02
GC_9_1172 b_9 NI_9 NS_1172 0 2.2836660703411945e-02
GC_9_1173 b_9 NI_9 NS_1173 0 2.2839352234481268e-02
GC_9_1174 b_9 NI_9 NS_1174 0 -2.2670699964558942e-02
GC_9_1175 b_9 NI_9 NS_1175 0 -9.2392572266465668e-03
GC_9_1176 b_9 NI_9 NS_1176 0 9.0801649156103015e-04
GC_9_1177 b_9 NI_9 NS_1177 0 1.8480444531577048e-02
GC_9_1178 b_9 NI_9 NS_1178 0 6.2433949828413979e-03
GC_9_1179 b_9 NI_9 NS_1179 0 -9.1763265309298108e-03
GC_9_1180 b_9 NI_9 NS_1180 0 -9.4611036353863479e-03
GC_9_1181 b_9 NI_9 NS_1181 0 -9.9741831229017922e-03
GC_9_1182 b_9 NI_9 NS_1182 0 6.3961404491670228e-03
GC_9_1183 b_9 NI_9 NS_1183 0 1.6838378743725058e-02
GC_9_1184 b_9 NI_9 NS_1184 0 -4.8507571343218737e-03
GC_9_1185 b_9 NI_9 NS_1185 0 -7.2149766097677924e-03
GC_9_1186 b_9 NI_9 NS_1186 0 -3.4093170377390426e-03
GC_9_1187 b_9 NI_9 NS_1187 0 6.8284598867639767e-03
GC_9_1188 b_9 NI_9 NS_1188 0 1.3296718008882286e-02
GC_9_1189 b_9 NI_9 NS_1189 0 -1.8198422883994197e-03
GC_9_1190 b_9 NI_9 NS_1190 0 -1.4401884747286533e-02
GC_9_1191 b_9 NI_9 NS_1191 0 -4.9859624292223088e-03
GC_9_1192 b_9 NI_9 NS_1192 0 1.0394192940165706e-03
GC_9_1193 b_9 NI_9 NS_1193 0 6.0026872519326384e-03
GC_9_1194 b_9 NI_9 NS_1194 0 -1.1033379851640990e-03
GC_9_1195 b_9 NI_9 NS_1195 0 -3.4642736715968939e-03
GC_9_1196 b_9 NI_9 NS_1196 0 -1.0877132921070299e-03
GC_9_1197 b_9 NI_9 NS_1197 0 2.7180843228174155e-03
GC_9_1198 b_9 NI_9 NS_1198 0 -5.0793073185805449e-04
GC_9_1199 b_9 NI_9 NS_1199 0 -3.2964042307130261e-03
GC_9_1200 b_9 NI_9 NS_1200 0 -2.8952142993837067e-03
GC_9_1201 b_9 NI_9 NS_1201 0 2.0160582918130536e-03
GC_9_1202 b_9 NI_9 NS_1202 0 7.7561412799204740e-04
GC_9_1203 b_9 NI_9 NS_1203 0 -2.0162391613312517e-03
GC_9_1204 b_9 NI_9 NS_1204 0 -9.6653840622431294e-04
GC_9_1205 b_9 NI_9 NS_1205 0 2.1216791622874426e-03
GC_9_1206 b_9 NI_9 NS_1206 0 -1.4710192928717989e-03
GC_9_1207 b_9 NI_9 NS_1207 0 -4.1846667586618721e-03
GC_9_1208 b_9 NI_9 NS_1208 0 -1.8129789192803303e-03
GC_9_1209 b_9 NI_9 NS_1209 0 2.3699521136933016e-03
GC_9_1210 b_9 NI_9 NS_1210 0 -3.7091804134447908e-04
GC_9_1211 b_9 NI_9 NS_1211 0 -3.0171283246551322e-03
GC_9_1212 b_9 NI_9 NS_1212 0 4.6227809629418378e-04
GC_9_1213 b_9 NI_9 NS_1213 0 2.7066143487271543e-03
GC_9_1214 b_9 NI_9 NS_1214 0 -2.7283529759331462e-03
GC_9_1215 b_9 NI_9 NS_1215 0 -5.0391230855259452e-03
GC_9_1216 b_9 NI_9 NS_1216 0 -1.2777907302011357e-04
GC_9_1217 b_9 NI_9 NS_1217 0 2.4350369276816557e-03
GC_9_1218 b_9 NI_9 NS_1218 0 -2.1722372652507658e-03
GC_9_1219 b_9 NI_9 NS_1219 0 -3.2447335282944079e-03
GC_9_1220 b_9 NI_9 NS_1220 0 2.6004818072959692e-03
GC_9_1221 b_9 NI_9 NS_1221 0 1.7440002919543881e-03
GC_9_1222 b_9 NI_9 NS_1222 0 -4.7506629812875192e-03
GC_9_1223 b_9 NI_9 NS_1223 0 -3.6334526772661170e-03
GC_9_1224 b_9 NI_9 NS_1224 0 2.5968941596441132e-03
GC_9_1225 b_9 NI_9 NS_1225 0 -2.8337529739959791e-03
GC_9_1226 b_9 NI_9 NS_1226 0 3.9869956619983764e-03
GC_9_1227 b_9 NI_9 NS_1227 0 -2.2097510893575136e-04
GC_9_1228 b_9 NI_9 NS_1228 0 -4.2143869040178437e-03
GC_9_1229 b_9 NI_9 NS_1229 0 -9.9004394498567988e-06
GC_9_1230 b_9 NI_9 NS_1230 0 7.5069812221660601e-06
GC_9_1231 b_9 NI_9 NS_1231 0 -1.3536762360025533e-03
GC_9_1232 b_9 NI_9 NS_1232 0 3.3750405193553796e-03
GC_9_1233 b_9 NI_9 NS_1233 0 -9.6980990466844202e-04
GC_9_1234 b_9 NI_9 NS_1234 0 -4.3483855057000051e-03
GC_9_1235 b_9 NI_9 NS_1235 0 -1.0004341440474213e-03
GC_9_1236 b_9 NI_9 NS_1236 0 2.2215368758924290e-03
GC_9_1237 b_9 NI_9 NS_1237 0 -1.6509401654854494e-03
GC_9_1238 b_9 NI_9 NS_1238 0 -4.4091665541816831e-03
GC_9_1239 b_9 NI_9 NS_1239 0 -1.4483893071176224e-03
GC_9_1240 b_9 NI_9 NS_1240 0 -2.4971174640483810e-03
GC_9_1241 b_9 NI_9 NS_1241 0 7.8206336442691274e-04
GC_9_1242 b_9 NI_9 NS_1242 0 2.5934675449261510e-03
GC_9_1243 b_9 NI_9 NS_1243 0 -6.9629910872200248e-04
GC_9_1244 b_9 NI_9 NS_1244 0 2.8791307009008479e-03
GC_9_1245 b_9 NI_9 NS_1245 0 -1.4354331452082450e-03
GC_9_1246 b_9 NI_9 NS_1246 0 -2.7718928615073912e-03
GC_9_1247 b_9 NI_9 NS_1247 0 -1.1678458093008694e-03
GC_9_1248 b_9 NI_9 NS_1248 0 2.6661739013162261e-03
GC_9_1249 b_9 NI_9 NS_1249 0 7.8077011825179591e-04
GC_9_1250 b_9 NI_9 NS_1250 0 -1.8746307413897063e-03
GC_9_1251 b_9 NI_9 NS_1251 0 2.3791496125770761e-08
GC_9_1252 b_9 NI_9 NS_1252 0 -6.0255366166141446e-08
GC_9_1253 b_9 NI_9 NS_1253 0 -9.0379586952769769e-07
GC_9_1254 b_9 NI_9 NS_1254 0 3.2032341124473335e-06
GC_9_1255 b_9 NI_9 NS_1255 0 2.9495679940693912e-03
GC_9_1256 b_9 NI_9 NS_1256 0 -6.1234113326721245e-04
GC_9_1257 b_9 NI_9 NS_1257 0 2.7950027954278982e-08
GC_9_1258 b_9 NI_9 NS_1258 0 -3.1703345463930437e-08
GC_9_1259 b_9 NI_9 NS_1259 0 2.0347235321188236e-04
GC_9_1260 b_9 NI_9 NS_1260 0 1.3799460007516754e-04
GC_9_1261 b_9 NI_9 NS_1261 0 5.6259198180166534e-04
GC_9_1262 b_9 NI_9 NS_1262 0 2.6570831657286224e-04
GC_9_1263 b_9 NI_9 NS_1263 0 3.1064656356366940e-03
GC_9_1264 b_9 NI_9 NS_1264 0 -2.2048908545829193e-03
GC_9_1265 b_9 NI_9 NS_1265 0 -1.5822536260906206e-03
GC_9_1266 b_9 NI_9 NS_1266 0 -2.6870774479138340e-03
GC_9_1267 b_9 NI_9 NS_1267 0 -2.0496561196713978e-03
GC_9_1268 b_9 NI_9 NS_1268 0 -3.7885087020446567e-03
GC_9_1269 b_9 NI_9 NS_1269 0 -4.9745586321529468e-03
GC_9_1270 b_9 NI_9 NS_1270 0 -1.5415288871657277e-03
GC_9_1271 b_9 NI_9 NS_1271 0 2.9290513834002242e-04
GC_9_1272 b_9 NI_9 NS_1272 0 1.9565076845820363e-04
GC_9_1273 b_9 NI_9 NS_1273 0 -2.8663285478989879e-03
GC_9_1274 b_9 NI_9 NS_1274 0 -9.5746354397062384e-04
GC_9_1275 b_9 NI_9 NS_1275 0 -2.2151870465680155e-02
GC_9_1276 b_9 NI_9 NS_1276 0 -1.0226311516934367e-02
GC_9_1277 b_9 NI_9 NS_1277 0 1.1325003956531824e-03
GC_9_1278 b_9 NI_9 NS_1278 0 2.0395318218717522e-02
GC_9_1279 b_9 NI_9 NS_1279 0 -5.8416196342551208e-03
GC_9_1280 b_9 NI_9 NS_1280 0 4.6116300268963248e-03
GC_9_1281 b_9 NI_9 NS_1281 0 5.7171575713024251e-03
GC_9_1282 b_9 NI_9 NS_1282 0 3.4516067884488570e-02
GC_9_1283 b_9 NI_9 NS_1283 0 8.0342764986013875e-03
GC_9_1284 b_9 NI_9 NS_1284 0 2.7930219483789437e-03
GC_9_1285 b_9 NI_9 NS_1285 0 -7.7724143243275588e-03
GC_9_1286 b_9 NI_9 NS_1286 0 2.9556755626563892e-02
GC_9_1287 b_9 NI_9 NS_1287 0 5.0768424387934101e-02
GC_9_1288 b_9 NI_9 NS_1288 0 -2.0072972526211957e-02
GC_9_1289 b_9 NI_9 NS_1289 0 7.9195780552725019e-03
GC_9_1290 b_9 NI_9 NS_1290 0 -1.6364429539933298e-03
GC_9_1291 b_9 NI_9 NS_1291 0 2.9084853638030619e-02
GC_9_1292 b_9 NI_9 NS_1292 0 -2.6464743141271729e-02
GC_9_1293 b_9 NI_9 NS_1293 0 -6.7250699989454136e-03
GC_9_1294 b_9 NI_9 NS_1294 0 -9.8822038532503428e-03
GC_9_1295 b_9 NI_9 NS_1295 0 8.4630804940090607e-03
GC_9_1296 b_9 NI_9 NS_1296 0 -8.0278000547105571e-03
GC_9_1297 b_9 NI_9 NS_1297 0 -1.8994957662684907e-02
GC_9_1298 b_9 NI_9 NS_1298 0 -2.5238416819028910e-02
GC_9_1299 b_9 NI_9 NS_1299 0 -5.4717854415041933e-03
GC_9_1300 b_9 NI_9 NS_1300 0 -2.8547826219760273e-03
GC_9_1301 b_9 NI_9 NS_1301 0 -1.7741075684371159e-02
GC_9_1302 b_9 NI_9 NS_1302 0 -1.3132225692575918e-02
GC_9_1303 b_9 NI_9 NS_1303 0 -4.8177975447712320e-03
GC_9_1304 b_9 NI_9 NS_1304 0 1.2541404139423978e-02
GC_9_1305 b_9 NI_9 NS_1305 0 -3.4590894789614402e-03
GC_9_1306 b_9 NI_9 NS_1306 0 1.5412388388980161e-03
GC_9_1307 b_9 NI_9 NS_1307 0 -7.1864995638827632e-04
GC_9_1308 b_9 NI_9 NS_1308 0 7.0058601089434333e-03
GC_9_1309 b_9 NI_9 NS_1309 0 1.8820413719497166e-03
GC_9_1310 b_9 NI_9 NS_1310 0 8.5748068800394181e-05
GC_9_1311 b_9 NI_9 NS_1311 0 3.1400245499142807e-04
GC_9_1312 b_9 NI_9 NS_1312 0 -1.9467015743245550e-03
GC_9_1313 b_9 NI_9 NS_1313 0 -1.8563355675584421e-03
GC_9_1314 b_9 NI_9 NS_1314 0 -1.6182085847056265e-03
GC_9_1315 b_9 NI_9 NS_1315 0 -2.1290958980289239e-03
GC_9_1316 b_9 NI_9 NS_1316 0 1.6850436216496042e-03
GC_9_1317 b_9 NI_9 NS_1317 0 7.6361045212609076e-04
GC_9_1318 b_9 NI_9 NS_1318 0 1.8527504119130256e-04
GC_9_1319 b_9 NI_9 NS_1319 0 -6.9730374401336093e-04
GC_9_1320 b_9 NI_9 NS_1320 0 -1.6780701358443441e-03
GC_9_1321 b_9 NI_9 NS_1321 0 -2.6815284491109341e-03
GC_9_1322 b_9 NI_9 NS_1322 0 -8.2749108318575502e-04
GC_9_1323 b_9 NI_9 NS_1323 0 -4.9989633057091851e-04
GC_9_1324 b_9 NI_9 NS_1324 0 2.9288644903597816e-03
GC_9_1325 b_9 NI_9 NS_1325 0 1.3533577613275727e-03
GC_9_1326 b_9 NI_9 NS_1326 0 -8.5805582422482862e-04
GC_9_1327 b_9 NI_9 NS_1327 0 -2.4189245083752310e-03
GC_9_1328 b_9 NI_9 NS_1328 0 -2.2676209057864568e-03
GC_9_1329 b_9 NI_9 NS_1329 0 -3.5540455296452483e-03
GC_9_1330 b_9 NI_9 NS_1330 0 7.4852709667471427e-04
GC_9_1331 b_9 NI_9 NS_1331 0 2.4633837046622153e-03
GC_9_1332 b_9 NI_9 NS_1332 0 3.0182802129159452e-03
GC_9_1333 b_9 NI_9 NS_1333 0 9.8455437090501341e-04
GC_9_1334 b_9 NI_9 NS_1334 0 -2.9418099053371517e-03
GC_9_1335 b_9 NI_9 NS_1335 0 -4.7677997600105871e-03
GC_9_1336 b_9 NI_9 NS_1336 0 5.4340110826196837e-05
GC_9_1337 b_9 NI_9 NS_1337 0 -1.7083702474394158e-03
GC_9_1338 b_9 NI_9 NS_1338 0 3.7124268779096200e-03
GC_9_1339 b_9 NI_9 NS_1339 0 -7.6587306598475968e-04
GC_9_1340 b_9 NI_9 NS_1340 0 1.5006759439069592e-03
GC_9_1341 b_9 NI_9 NS_1341 0 3.2213013834260103e-03
GC_9_1342 b_9 NI_9 NS_1342 0 -1.3508681736958974e-03
GC_9_1343 b_9 NI_9 NS_1343 0 -2.9326134613597625e-06
GC_9_1344 b_9 NI_9 NS_1344 0 8.7469996771945133e-06
GC_9_1345 b_9 NI_9 NS_1345 0 -1.8200418131280370e-03
GC_9_1346 b_9 NI_9 NS_1346 0 -2.5277356947917477e-03
GC_9_1347 b_9 NI_9 NS_1347 0 -2.4072528131844251e-03
GC_9_1348 b_9 NI_9 NS_1348 0 2.4886639030400337e-03
GC_9_1349 b_9 NI_9 NS_1349 0 1.0142614019019176e-03
GC_9_1350 b_9 NI_9 NS_1350 0 2.4256823381263743e-03
GC_9_1351 b_9 NI_9 NS_1351 0 8.5775954199840106e-04
GC_9_1352 b_9 NI_9 NS_1352 0 -2.6994832914913267e-03
GC_9_1353 b_9 NI_9 NS_1353 0 -3.0644805767557202e-04
GC_9_1354 b_9 NI_9 NS_1354 0 1.6741356010219937e-03
GC_9_1355 b_9 NI_9 NS_1355 0 -1.7840545176579757e-03
GC_9_1356 b_9 NI_9 NS_1356 0 -3.1181087559361518e-04
GC_9_1357 b_9 NI_9 NS_1357 0 1.4004540025064078e-03
GC_9_1358 b_9 NI_9 NS_1358 0 1.9709614159929439e-03
GC_9_1359 b_9 NI_9 NS_1359 0 1.0449286373672931e-03
GC_9_1360 b_9 NI_9 NS_1360 0 -2.2998046800000805e-03
GC_9_1361 b_9 NI_9 NS_1361 0 -6.9799492357377005e-04
GC_9_1362 b_9 NI_9 NS_1362 0 -1.4668899079096245e-03
GC_9_1363 b_9 NI_9 NS_1363 0 -1.3735490693109877e-03
GC_9_1364 b_9 NI_9 NS_1364 0 -3.1252861795985599e-04
GC_9_1365 b_9 NI_9 NS_1365 0 7.1030495328530861e-09
GC_9_1366 b_9 NI_9 NS_1366 0 -2.4709972806960687e-08
GC_9_1367 b_9 NI_9 NS_1367 0 -4.5275608481998805e-07
GC_9_1368 b_9 NI_9 NS_1368 0 1.6341840534431939e-06
GD_9_1 b_9 NI_9 NA_1 0 -1.8797278172832675e-06
GD_9_2 b_9 NI_9 NA_2 0 5.6280536661590336e-06
GD_9_3 b_9 NI_9 NA_3 0 -5.5537914020317968e-06
GD_9_4 b_9 NI_9 NA_4 0 4.7472069075166415e-07
GD_9_5 b_9 NI_9 NA_5 0 4.5909851974180033e-06
GD_9_6 b_9 NI_9 NA_6 0 1.2379585097852849e-06
GD_9_7 b_9 NI_9 NA_7 0 1.0377145993641142e-04
GD_9_8 b_9 NI_9 NA_8 0 2.6586123964651599e-05
GD_9_9 b_9 NI_9 NA_9 0 -8.6867573911805582e-03
GD_9_10 b_9 NI_9 NA_10 0 -4.2441623974806674e-03
GD_9_11 b_9 NI_9 NA_11 0 1.3006424217651818e-02
GD_9_12 b_9 NI_9 NA_12 0 5.9084240467126682e-04
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 -2.7508893938899258e-05
GC_10_2 b_10 NI_10 NS_2 0 -1.0597481601631146e-08
GC_10_3 b_10 NI_10 NS_3 0 1.0238663393770382e-11
GC_10_4 b_10 NI_10 NS_4 0 -5.9557115759443859e-11
GC_10_5 b_10 NI_10 NS_5 0 -6.3653597462755455e-07
GC_10_6 b_10 NI_10 NS_6 0 -1.0748172610165871e-06
GC_10_7 b_10 NI_10 NS_7 0 -1.4323543785347750e-06
GC_10_8 b_10 NI_10 NS_8 0 2.3248382337241046e-06
GC_10_9 b_10 NI_10 NS_9 0 -3.8131192876609988e-06
GC_10_10 b_10 NI_10 NS_10 0 2.1795952416944330e-06
GC_10_11 b_10 NI_10 NS_11 0 1.9255556240165656e-06
GC_10_12 b_10 NI_10 NS_12 0 -2.3467049885247559e-07
GC_10_13 b_10 NI_10 NS_13 0 1.4104706969632813e-06
GC_10_14 b_10 NI_10 NS_14 0 5.7203904248072498e-06
GC_10_15 b_10 NI_10 NS_15 0 3.7051865945807558e-06
GC_10_16 b_10 NI_10 NS_16 0 3.2538242309460749e-06
GC_10_17 b_10 NI_10 NS_17 0 -1.4742101134044455e-06
GC_10_18 b_10 NI_10 NS_18 0 -9.4918358724248226e-07
GC_10_19 b_10 NI_10 NS_19 0 9.7320233203480378e-07
GC_10_20 b_10 NI_10 NS_20 0 -2.1860365313718368e-06
GC_10_21 b_10 NI_10 NS_21 0 6.4354576589679731e-06
GC_10_22 b_10 NI_10 NS_22 0 8.5306779480363118e-06
GC_10_23 b_10 NI_10 NS_23 0 1.3303187052540580e-06
GC_10_24 b_10 NI_10 NS_24 0 -9.3980189874513159e-07
GC_10_25 b_10 NI_10 NS_25 0 1.0706262246112963e-06
GC_10_26 b_10 NI_10 NS_26 0 -1.9034787007921180e-06
GC_10_27 b_10 NI_10 NS_27 0 1.4528567145120655e-05
GC_10_28 b_10 NI_10 NS_28 0 -4.1922294687513462e-06
GC_10_29 b_10 NI_10 NS_29 0 -2.0124975370554693e-07
GC_10_30 b_10 NI_10 NS_30 0 6.7953948139518564e-07
GC_10_31 b_10 NI_10 NS_31 0 4.9185684200853572e-06
GC_10_32 b_10 NI_10 NS_32 0 -2.1983512390183377e-06
GC_10_33 b_10 NI_10 NS_33 0 -7.4682180848983609e-07
GC_10_34 b_10 NI_10 NS_34 0 -1.4996634517367930e-05
GC_10_35 b_10 NI_10 NS_35 0 -7.6209536310564924e-08
GC_10_36 b_10 NI_10 NS_36 0 9.7376803840110546e-07
GC_10_37 b_10 NI_10 NS_37 0 -7.9309876453926192e-06
GC_10_38 b_10 NI_10 NS_38 0 -8.5785738262438727e-06
GC_10_39 b_10 NI_10 NS_39 0 -6.2161142323342062e-07
GC_10_40 b_10 NI_10 NS_40 0 -2.1586591951480847e-06
GC_10_41 b_10 NI_10 NS_41 0 -8.3548793705322306e-09
GC_10_42 b_10 NI_10 NS_42 0 1.2073831921283967e-06
GC_10_43 b_10 NI_10 NS_43 0 -7.7193083009115523e-06
GC_10_44 b_10 NI_10 NS_44 0 1.9618686729736814e-06
GC_10_45 b_10 NI_10 NS_45 0 2.4499728271273743e-07
GC_10_46 b_10 NI_10 NS_46 0 -1.6819636773941194e-06
GC_10_47 b_10 NI_10 NS_47 0 1.1608837498700348e-06
GC_10_48 b_10 NI_10 NS_48 0 3.0679012932770651e-06
GC_10_49 b_10 NI_10 NS_49 0 -9.7670489376771336e-07
GC_10_50 b_10 NI_10 NS_50 0 2.0311623029336069e-06
GC_10_51 b_10 NI_10 NS_51 0 4.5640486942468979e-07
GC_10_52 b_10 NI_10 NS_52 0 -1.2309756327330380e-06
GC_10_53 b_10 NI_10 NS_53 0 3.2453699145031543e-06
GC_10_54 b_10 NI_10 NS_54 0 -8.8263316145044359e-07
GC_10_55 b_10 NI_10 NS_55 0 -1.6147965006235583e-07
GC_10_56 b_10 NI_10 NS_56 0 5.1317029650990764e-07
GC_10_57 b_10 NI_10 NS_57 0 -8.4629659577497446e-07
GC_10_58 b_10 NI_10 NS_58 0 -4.1983678993160827e-07
GC_10_59 b_10 NI_10 NS_59 0 9.9341481071296947e-07
GC_10_60 b_10 NI_10 NS_60 0 -1.2689975928048251e-06
GC_10_61 b_10 NI_10 NS_61 0 1.4441190330165936e-06
GC_10_62 b_10 NI_10 NS_62 0 -5.7045272122444436e-07
GC_10_63 b_10 NI_10 NS_63 0 -3.4127605821959471e-08
GC_10_64 b_10 NI_10 NS_64 0 9.6990688766001571e-08
GC_10_65 b_10 NI_10 NS_65 0 -5.9769203587798811e-07
GC_10_66 b_10 NI_10 NS_66 0 -3.4060875282201594e-07
GC_10_67 b_10 NI_10 NS_67 0 9.6764720751845541e-07
GC_10_68 b_10 NI_10 NS_68 0 -1.0810513332640344e-06
GC_10_69 b_10 NI_10 NS_69 0 1.3955406610223672e-06
GC_10_70 b_10 NI_10 NS_70 0 -1.2449148205538002e-06
GC_10_71 b_10 NI_10 NS_71 0 1.6144726112836297e-07
GC_10_72 b_10 NI_10 NS_72 0 -4.3249262124936344e-08
GC_10_73 b_10 NI_10 NS_73 0 -4.8924774166157516e-07
GC_10_74 b_10 NI_10 NS_74 0 -5.0361967929717384e-07
GC_10_75 b_10 NI_10 NS_75 0 1.0632933605931252e-06
GC_10_76 b_10 NI_10 NS_76 0 -8.0454656010847581e-07
GC_10_77 b_10 NI_10 NS_77 0 1.2280669013742353e-06
GC_10_78 b_10 NI_10 NS_78 0 -2.1206236695462781e-06
GC_10_79 b_10 NI_10 NS_79 0 4.9661700741507294e-07
GC_10_80 b_10 NI_10 NS_80 0 -2.5356843593468228e-07
GC_10_81 b_10 NI_10 NS_81 0 -2.4768285696471869e-07
GC_10_82 b_10 NI_10 NS_82 0 -9.1984005039562874e-07
GC_10_83 b_10 NI_10 NS_83 0 1.9186405695249642e-06
GC_10_84 b_10 NI_10 NS_84 0 -1.0012898070615084e-06
GC_10_85 b_10 NI_10 NS_85 0 -8.0998127198842194e-06
GC_10_86 b_10 NI_10 NS_86 0 -9.1473015202365743e-07
GC_10_87 b_10 NI_10 NS_87 0 -3.1607425186864268e-07
GC_10_88 b_10 NI_10 NS_88 0 -3.6264956231914102e-06
GC_10_89 b_10 NI_10 NS_89 0 -4.9018343721280301e-08
GC_10_90 b_10 NI_10 NS_90 0 -3.3202875609289374e-08
GC_10_91 b_10 NI_10 NS_91 0 -1.0293941029322123e-07
GC_10_92 b_10 NI_10 NS_92 0 -1.2361446628235974e-06
GC_10_93 b_10 NI_10 NS_93 0 -1.0227326461196870e-06
GC_10_94 b_10 NI_10 NS_94 0 -6.6783059347776406e-07
GC_10_95 b_10 NI_10 NS_95 0 1.4569219292055611e-06
GC_10_96 b_10 NI_10 NS_96 0 -7.6152211950838040e-07
GC_10_97 b_10 NI_10 NS_97 0 1.9436905875234502e-06
GC_10_98 b_10 NI_10 NS_98 0 -1.8722412268954719e-06
GC_10_99 b_10 NI_10 NS_99 0 -2.2230857632009413e-07
GC_10_100 b_10 NI_10 NS_100 0 3.2515823160696578e-07
GC_10_101 b_10 NI_10 NS_101 0 2.1538321541877412e-07
GC_10_102 b_10 NI_10 NS_102 0 5.2991215866141600e-07
GC_10_103 b_10 NI_10 NS_103 0 -1.0774199736020922e-07
GC_10_104 b_10 NI_10 NS_104 0 -2.8383121859725833e-07
GC_10_105 b_10 NI_10 NS_105 0 8.1696518149676524e-09
GC_10_106 b_10 NI_10 NS_106 0 -9.6164615446627034e-08
GC_10_107 b_10 NI_10 NS_107 0 -8.8650248876893230e-08
GC_10_108 b_10 NI_10 NS_108 0 4.2005306428089032e-08
GC_10_109 b_10 NI_10 NS_109 0 -1.2200388749801090e-07
GC_10_110 b_10 NI_10 NS_110 0 -5.3538805826271833e-08
GC_10_111 b_10 NI_10 NS_111 0 6.1367442518211928e-12
GC_10_112 b_10 NI_10 NS_112 0 -1.6270632649026780e-12
GC_10_113 b_10 NI_10 NS_113 0 3.5453380563090943e-10
GC_10_114 b_10 NI_10 NS_114 0 6.9229613174404715e-10
GC_10_115 b_10 NI_10 NS_115 0 1.3439640693240003e-05
GC_10_116 b_10 NI_10 NS_116 0 -5.8811666008385650e-08
GC_10_117 b_10 NI_10 NS_117 0 -1.4973646003055918e-11
GC_10_118 b_10 NI_10 NS_118 0 1.3623458994843434e-10
GC_10_119 b_10 NI_10 NS_119 0 3.6109503686135079e-07
GC_10_120 b_10 NI_10 NS_120 0 -1.7974058858828938e-07
GC_10_121 b_10 NI_10 NS_121 0 2.8426234307402063e-07
GC_10_122 b_10 NI_10 NS_122 0 -3.5218297094117679e-07
GC_10_123 b_10 NI_10 NS_123 0 5.0389364988751635e-07
GC_10_124 b_10 NI_10 NS_124 0 -1.4258624693914526e-06
GC_10_125 b_10 NI_10 NS_125 0 -1.1608911337083200e-06
GC_10_126 b_10 NI_10 NS_126 0 -4.7429562021473418e-07
GC_10_127 b_10 NI_10 NS_127 0 -3.4574784771791459e-07
GC_10_128 b_10 NI_10 NS_128 0 -6.3124048552834442e-07
GC_10_129 b_10 NI_10 NS_129 0 -2.5929911533646223e-06
GC_10_130 b_10 NI_10 NS_130 0 -6.5714139244342719e-07
GC_10_131 b_10 NI_10 NS_131 0 7.1939761724716335e-07
GC_10_132 b_10 NI_10 NS_132 0 3.6304541053016834e-07
GC_10_133 b_10 NI_10 NS_133 0 -7.3971047386472140e-07
GC_10_134 b_10 NI_10 NS_134 0 3.6642637747605424e-07
GC_10_135 b_10 NI_10 NS_135 0 -1.0222414758706251e-06
GC_10_136 b_10 NI_10 NS_136 0 5.8988411479551548e-07
GC_10_137 b_10 NI_10 NS_137 0 -4.1600466528880446e-07
GC_10_138 b_10 NI_10 NS_138 0 2.6264310335134245e-07
GC_10_139 b_10 NI_10 NS_139 0 -8.5727208447419053e-07
GC_10_140 b_10 NI_10 NS_140 0 4.4631299009739902e-07
GC_10_141 b_10 NI_10 NS_141 0 1.5253918567798346e-07
GC_10_142 b_10 NI_10 NS_142 0 1.1341005359320475e-06
GC_10_143 b_10 NI_10 NS_143 0 -5.9583506910494836e-07
GC_10_144 b_10 NI_10 NS_144 0 1.1918705398459169e-07
GC_10_145 b_10 NI_10 NS_145 0 -1.9185659990801744e-06
GC_10_146 b_10 NI_10 NS_146 0 1.2734567750216332e-06
GC_10_147 b_10 NI_10 NS_147 0 2.0855884917555579e-06
GC_10_148 b_10 NI_10 NS_148 0 2.8031336559509748e-07
GC_10_149 b_10 NI_10 NS_149 0 -6.8889830584015935e-07
GC_10_150 b_10 NI_10 NS_150 0 1.8836136207287664e-07
GC_10_151 b_10 NI_10 NS_151 0 9.8343411287414779e-07
GC_10_152 b_10 NI_10 NS_152 0 1.7053682215742242e-06
GC_10_153 b_10 NI_10 NS_153 0 -2.2785250523123510e-07
GC_10_154 b_10 NI_10 NS_154 0 -5.8892787420024620e-07
GC_10_155 b_10 NI_10 NS_155 0 -9.2869872239419507e-07
GC_10_156 b_10 NI_10 NS_156 0 4.1600968569656157e-07
GC_10_157 b_10 NI_10 NS_157 0 1.4319961032232304e-06
GC_10_158 b_10 NI_10 NS_158 0 7.1444776134816752e-07
GC_10_159 b_10 NI_10 NS_159 0 -3.3565454131483826e-07
GC_10_160 b_10 NI_10 NS_160 0 -2.2026679678019241e-07
GC_10_161 b_10 NI_10 NS_161 0 -5.3855050102634444e-08
GC_10_162 b_10 NI_10 NS_162 0 1.4317869082120925e-06
GC_10_163 b_10 NI_10 NS_163 0 4.8359324132777195e-07
GC_10_164 b_10 NI_10 NS_164 0 -7.6448870444620229e-07
GC_10_165 b_10 NI_10 NS_165 0 -3.5361622367917380e-07
GC_10_166 b_10 NI_10 NS_166 0 4.2725039940285871e-08
GC_10_167 b_10 NI_10 NS_167 0 3.2259207545554945e-07
GC_10_168 b_10 NI_10 NS_168 0 3.9012923467491055e-07
GC_10_169 b_10 NI_10 NS_169 0 -1.4407258217473719e-07
GC_10_170 b_10 NI_10 NS_170 0 -1.1227716822679877e-08
GC_10_171 b_10 NI_10 NS_171 0 1.4059231810427961e-07
GC_10_172 b_10 NI_10 NS_172 0 1.2582106804664090e-07
GC_10_173 b_10 NI_10 NS_173 0 -1.9006710291924021e-07
GC_10_174 b_10 NI_10 NS_174 0 -6.9875969405310443e-08
GC_10_175 b_10 NI_10 NS_175 0 3.8836468553831369e-08
GC_10_176 b_10 NI_10 NS_176 0 1.9898312979364533e-07
GC_10_177 b_10 NI_10 NS_177 0 -1.1133969178163624e-07
GC_10_178 b_10 NI_10 NS_178 0 9.3792281107001147e-09
GC_10_179 b_10 NI_10 NS_179 0 4.6150699415331688e-08
GC_10_180 b_10 NI_10 NS_180 0 7.8744471232099304e-09
GC_10_181 b_10 NI_10 NS_181 0 -2.9781816341704256e-07
GC_10_182 b_10 NI_10 NS_182 0 -5.3926574254057845e-08
GC_10_183 b_10 NI_10 NS_183 0 -9.1414102955848027e-08
GC_10_184 b_10 NI_10 NS_184 0 6.3222368843421536e-08
GC_10_185 b_10 NI_10 NS_185 0 -2.3130301351472309e-07
GC_10_186 b_10 NI_10 NS_186 0 7.8668897407888449e-08
GC_10_187 b_10 NI_10 NS_187 0 -1.3284208501394498e-07
GC_10_188 b_10 NI_10 NS_188 0 -6.8245309211401685e-08
GC_10_189 b_10 NI_10 NS_189 0 -4.3126490404563878e-07
GC_10_190 b_10 NI_10 NS_190 0 -5.7483731109076123e-08
GC_10_191 b_10 NI_10 NS_191 0 -4.2237571843699952e-07
GC_10_192 b_10 NI_10 NS_192 0 6.4399124743593131e-08
GC_10_193 b_10 NI_10 NS_193 0 -4.4356288797698890e-07
GC_10_194 b_10 NI_10 NS_194 0 1.4475411635026056e-07
GC_10_195 b_10 NI_10 NS_195 0 -5.1285003200858690e-07
GC_10_196 b_10 NI_10 NS_196 0 1.0392220982010024e-07
GC_10_197 b_10 NI_10 NS_197 0 -9.6728438753322614e-07
GC_10_198 b_10 NI_10 NS_198 0 -1.0044906203774691e-07
GC_10_199 b_10 NI_10 NS_199 0 2.6364145009008402e-06
GC_10_200 b_10 NI_10 NS_200 0 3.0037223311771137e-06
GC_10_201 b_10 NI_10 NS_201 0 -6.1832966087248098e-07
GC_10_202 b_10 NI_10 NS_202 0 1.0424218773090233e-06
GC_10_203 b_10 NI_10 NS_203 0 9.1726162755511159e-09
GC_10_204 b_10 NI_10 NS_204 0 2.5504725300819851e-08
GC_10_205 b_10 NI_10 NS_205 0 -4.7322577839723769e-07
GC_10_206 b_10 NI_10 NS_206 0 8.3082224127054195e-07
GC_10_207 b_10 NI_10 NS_207 0 9.3288647172995513e-09
GC_10_208 b_10 NI_10 NS_208 0 3.8802053610268844e-07
GC_10_209 b_10 NI_10 NS_209 0 -8.7284250858741594e-07
GC_10_210 b_10 NI_10 NS_210 0 -7.3755431755560803e-08
GC_10_211 b_10 NI_10 NS_211 0 -9.8359171058835966e-07
GC_10_212 b_10 NI_10 NS_212 0 -1.8073798650152695e-07
GC_10_213 b_10 NI_10 NS_213 0 1.0888657360597277e-07
GC_10_214 b_10 NI_10 NS_214 0 -1.4767566898149960e-07
GC_10_215 b_10 NI_10 NS_215 0 6.7378677600121364e-08
GC_10_216 b_10 NI_10 NS_216 0 1.3250454687938397e-08
GC_10_217 b_10 NI_10 NS_217 0 -6.9949645642393464e-08
GC_10_218 b_10 NI_10 NS_218 0 1.6113308001781018e-07
GC_10_219 b_10 NI_10 NS_219 0 2.9099319628728294e-08
GC_10_220 b_10 NI_10 NS_220 0 -4.0233237403988016e-08
GC_10_221 b_10 NI_10 NS_221 0 -8.1240467882732254e-08
GC_10_222 b_10 NI_10 NS_222 0 1.6008187902973840e-07
GC_10_223 b_10 NI_10 NS_223 0 5.6406778176825075e-08
GC_10_224 b_10 NI_10 NS_224 0 -1.6261373630679063e-08
GC_10_225 b_10 NI_10 NS_225 0 -1.1764284278228091e-11
GC_10_226 b_10 NI_10 NS_226 0 5.1442945511337749e-12
GC_10_227 b_10 NI_10 NS_227 0 -3.3968994727325316e-10
GC_10_228 b_10 NI_10 NS_228 0 -9.7415206911195679e-10
GC_10_229 b_10 NI_10 NS_229 0 -2.1854824181534118e-05
GC_10_230 b_10 NI_10 NS_230 0 2.4289840867103552e-07
GC_10_231 b_10 NI_10 NS_231 0 1.6216473311092679e-11
GC_10_232 b_10 NI_10 NS_232 0 -4.8482543583374967e-10
GC_10_233 b_10 NI_10 NS_233 0 3.7393828882243125e-07
GC_10_234 b_10 NI_10 NS_234 0 -1.3861922442073096e-06
GC_10_235 b_10 NI_10 NS_235 0 -1.4298858485246249e-07
GC_10_236 b_10 NI_10 NS_236 0 1.1185368133418358e-06
GC_10_237 b_10 NI_10 NS_237 0 -3.5074189516207827e-06
GC_10_238 b_10 NI_10 NS_238 0 -2.2370251912804962e-06
GC_10_239 b_10 NI_10 NS_239 0 -7.4943835210617608e-07
GC_10_240 b_10 NI_10 NS_240 0 -1.1227634732201164e-06
GC_10_241 b_10 NI_10 NS_241 0 -6.8343749381662218e-07
GC_10_242 b_10 NI_10 NS_242 0 2.6595633943878516e-06
GC_10_243 b_10 NI_10 NS_243 0 -5.0813960031553604e-06
GC_10_244 b_10 NI_10 NS_244 0 3.8742887002431590e-06
GC_10_245 b_10 NI_10 NS_245 0 9.5053093124888614e-07
GC_10_246 b_10 NI_10 NS_246 0 -1.5553499561287053e-07
GC_10_247 b_10 NI_10 NS_247 0 -2.6358441499810520e-07
GC_10_248 b_10 NI_10 NS_248 0 -5.2938698712025441e-07
GC_10_249 b_10 NI_10 NS_249 0 -1.4742607443294712e-06
GC_10_250 b_10 NI_10 NS_250 0 1.1166392432907620e-05
GC_10_251 b_10 NI_10 NS_251 0 5.7536166350421955e-06
GC_10_252 b_10 NI_10 NS_252 0 2.9700709611774540e-06
GC_10_253 b_10 NI_10 NS_253 0 7.6103335969304785e-07
GC_10_254 b_10 NI_10 NS_254 0 -4.0059674069265993e-07
GC_10_255 b_10 NI_10 NS_255 0 1.7105182645060764e-05
GC_10_256 b_10 NI_10 NS_256 0 -2.9783341803994562e-07
GC_10_257 b_10 NI_10 NS_257 0 7.0007322269049621e-07
GC_10_258 b_10 NI_10 NS_258 0 1.7703040262907053e-07
GC_10_259 b_10 NI_10 NS_259 0 6.4126693051944232e-06
GC_10_260 b_10 NI_10 NS_260 0 -4.4402795209175741e-07
GC_10_261 b_10 NI_10 NS_261 0 -8.2381542858721524e-07
GC_10_262 b_10 NI_10 NS_262 0 -1.7747640760616073e-05
GC_10_263 b_10 NI_10 NS_263 0 -2.8347507106615259e-07
GC_10_264 b_10 NI_10 NS_264 0 2.3003600300994768e-07
GC_10_265 b_10 NI_10 NS_265 0 -1.0769398775547954e-05
GC_10_266 b_10 NI_10 NS_266 0 -9.4805213900930322e-06
GC_10_267 b_10 NI_10 NS_267 0 -1.3423576161756929e-06
GC_10_268 b_10 NI_10 NS_268 0 -8.1223868676925698e-07
GC_10_269 b_10 NI_10 NS_269 0 -1.6041426447729598e-06
GC_10_270 b_10 NI_10 NS_270 0 4.5694582482007085e-07
GC_10_271 b_10 NI_10 NS_271 0 -9.3337965656378544e-06
GC_10_272 b_10 NI_10 NS_272 0 6.4384875704870836e-06
GC_10_273 b_10 NI_10 NS_273 0 6.7351571978914004e-08
GC_10_274 b_10 NI_10 NS_274 0 -3.9969604228286110e-07
GC_10_275 b_10 NI_10 NS_275 0 -7.1799616247048604e-07
GC_10_276 b_10 NI_10 NS_276 0 7.2325979566752324e-06
GC_10_277 b_10 NI_10 NS_277 0 2.0739496448834925e-06
GC_10_278 b_10 NI_10 NS_278 0 2.4611622249746592e-06
GC_10_279 b_10 NI_10 NS_279 0 6.1968363344327277e-07
GC_10_280 b_10 NI_10 NS_280 0 -2.5247660497586016e-07
GC_10_281 b_10 NI_10 NS_281 0 4.6128204652247434e-06
GC_10_282 b_10 NI_10 NS_282 0 3.3398362773747416e-07
GC_10_283 b_10 NI_10 NS_283 0 1.7628560386958352e-07
GC_10_284 b_10 NI_10 NS_284 0 5.3873458675226089e-07
GC_10_285 b_10 NI_10 NS_285 0 -7.4074132228843031e-07
GC_10_286 b_10 NI_10 NS_286 0 -4.2045448029220341e-08
GC_10_287 b_10 NI_10 NS_287 0 7.4598003455167206e-07
GC_10_288 b_10 NI_10 NS_288 0 -5.2039439009258632e-07
GC_10_289 b_10 NI_10 NS_289 0 1.8298789851079102e-06
GC_10_290 b_10 NI_10 NS_290 0 4.7566089586321300e-07
GC_10_291 b_10 NI_10 NS_291 0 1.7708157027597233e-07
GC_10_292 b_10 NI_10 NS_292 0 4.5205088773319512e-07
GC_10_293 b_10 NI_10 NS_293 0 -4.4618876107424408e-07
GC_10_294 b_10 NI_10 NS_294 0 2.3604808847101294e-07
GC_10_295 b_10 NI_10 NS_295 0 6.4977369682003090e-07
GC_10_296 b_10 NI_10 NS_296 0 -3.4554293652722451e-07
GC_10_297 b_10 NI_10 NS_297 0 1.8733454496046690e-06
GC_10_298 b_10 NI_10 NS_298 0 -2.9392961633038187e-08
GC_10_299 b_10 NI_10 NS_299 0 2.9827021133195238e-07
GC_10_300 b_10 NI_10 NS_300 0 5.0985802864844817e-07
GC_10_301 b_10 NI_10 NS_301 0 -3.1520261921200810e-07
GC_10_302 b_10 NI_10 NS_302 0 4.5596894734557638e-07
GC_10_303 b_10 NI_10 NS_303 0 5.5349888707699758e-07
GC_10_304 b_10 NI_10 NS_304 0 -4.4724726757592287e-08
GC_10_305 b_10 NI_10 NS_305 0 1.9808667318150351e-06
GC_10_306 b_10 NI_10 NS_306 0 -4.0113621314326930e-07
GC_10_307 b_10 NI_10 NS_307 0 4.1702866762858368e-07
GC_10_308 b_10 NI_10 NS_308 0 7.7175836119869562e-07
GC_10_309 b_10 NI_10 NS_309 0 5.0615073961731703e-07
GC_10_310 b_10 NI_10 NS_310 0 7.2776826373128273e-07
GC_10_311 b_10 NI_10 NS_311 0 9.0283372262659960e-07
GC_10_312 b_10 NI_10 NS_312 0 9.8988568606943553e-07
GC_10_313 b_10 NI_10 NS_313 0 1.6386495062545877e-06
GC_10_314 b_10 NI_10 NS_314 0 -9.9921380651401517e-06
GC_10_315 b_10 NI_10 NS_315 0 2.8725442042594931e-06
GC_10_316 b_10 NI_10 NS_316 0 -1.2252067791747313e-06
GC_10_317 b_10 NI_10 NS_317 0 3.1669876095654662e-08
GC_10_318 b_10 NI_10 NS_318 0 -4.6445368419859596e-08
GC_10_319 b_10 NI_10 NS_319 0 1.4054983260902581e-06
GC_10_320 b_10 NI_10 NS_320 0 1.6971625581671121e-07
GC_10_321 b_10 NI_10 NS_321 0 9.7902320027646515e-07
GC_10_322 b_10 NI_10 NS_322 0 -4.9521637227866741e-07
GC_10_323 b_10 NI_10 NS_323 0 6.9358707904684425e-07
GC_10_324 b_10 NI_10 NS_324 0 1.3039617954541945e-06
GC_10_325 b_10 NI_10 NS_325 0 1.3369660341040503e-06
GC_10_326 b_10 NI_10 NS_326 0 1.9875920972081629e-06
GC_10_327 b_10 NI_10 NS_327 0 -9.2425227190845217e-08
GC_10_328 b_10 NI_10 NS_328 0 -2.7737400185972450e-08
GC_10_329 b_10 NI_10 NS_329 0 -5.3471683800798109e-07
GC_10_330 b_10 NI_10 NS_330 0 1.8250408663143228e-07
GC_10_331 b_10 NI_10 NS_331 0 3.1922773690705717e-07
GC_10_332 b_10 NI_10 NS_332 0 -3.6120294788622826e-07
GC_10_333 b_10 NI_10 NS_333 0 1.1467857443846447e-08
GC_10_334 b_10 NI_10 NS_334 0 -6.0659816732823582e-07
GC_10_335 b_10 NI_10 NS_335 0 5.2308726482152674e-08
GC_10_336 b_10 NI_10 NS_336 0 1.0683024044237987e-07
GC_10_337 b_10 NI_10 NS_337 0 2.9594390296720962e-07
GC_10_338 b_10 NI_10 NS_338 0 -1.4212193459180051e-09
GC_10_339 b_10 NI_10 NS_339 0 -2.9859155703170653e-12
GC_10_340 b_10 NI_10 NS_340 0 -1.0058359908351870e-11
GC_10_341 b_10 NI_10 NS_341 0 9.3177973909710418e-10
GC_10_342 b_10 NI_10 NS_342 0 3.3553895759417524e-09
GC_10_343 b_10 NI_10 NS_343 0 4.4177058756412571e-05
GC_10_344 b_10 NI_10 NS_344 0 -2.5097185976971737e-07
GC_10_345 b_10 NI_10 NS_345 0 -1.3616178142802775e-11
GC_10_346 b_10 NI_10 NS_346 0 3.6730833737290534e-10
GC_10_347 b_10 NI_10 NS_347 0 9.4985814116014279e-07
GC_10_348 b_10 NI_10 NS_348 0 -2.0373719148032102e-07
GC_10_349 b_10 NI_10 NS_349 0 1.1052050242776341e-06
GC_10_350 b_10 NI_10 NS_350 0 -6.5604994150677658e-07
GC_10_351 b_10 NI_10 NS_351 0 1.6285500655269714e-06
GC_10_352 b_10 NI_10 NS_352 0 -3.6724994872850312e-06
GC_10_353 b_10 NI_10 NS_353 0 -2.3667651046472988e-06
GC_10_354 b_10 NI_10 NS_354 0 -1.3304689516724547e-06
GC_10_355 b_10 NI_10 NS_355 0 -2.0333762511678727e-07
GC_10_356 b_10 NI_10 NS_356 0 -2.4445405867375502e-06
GC_10_357 b_10 NI_10 NS_357 0 -7.1157294626427683e-06
GC_10_358 b_10 NI_10 NS_358 0 -2.8107549360528674e-06
GC_10_359 b_10 NI_10 NS_359 0 1.7244823302000209e-06
GC_10_360 b_10 NI_10 NS_360 0 1.3116575553700636e-06
GC_10_361 b_10 NI_10 NS_361 0 -1.6513151316776930e-06
GC_10_362 b_10 NI_10 NS_362 0 9.9666903735613134e-07
GC_10_363 b_10 NI_10 NS_363 0 -2.8707126708271034e-06
GC_10_364 b_10 NI_10 NS_364 0 -1.6218902905018721e-06
GC_10_365 b_10 NI_10 NS_365 0 -2.0401147221493395e-06
GC_10_366 b_10 NI_10 NS_366 0 2.9683219015782797e-06
GC_10_367 b_10 NI_10 NS_367 0 -1.1731160575690848e-06
GC_10_368 b_10 NI_10 NS_368 0 1.1051278401406073e-06
GC_10_369 b_10 NI_10 NS_369 0 -2.0978475281227394e-06
GC_10_370 b_10 NI_10 NS_370 0 1.5286379238462809e-06
GC_10_371 b_10 NI_10 NS_371 0 -9.4302721224118188e-07
GC_10_372 b_10 NI_10 NS_372 0 1.4307779985960094e-06
GC_10_373 b_10 NI_10 NS_373 0 -1.4824685735080182e-06
GC_10_374 b_10 NI_10 NS_374 0 1.7943981322486918e-06
GC_10_375 b_10 NI_10 NS_375 0 2.5484689485347362e-07
GC_10_376 b_10 NI_10 NS_376 0 1.3612764232112203e-06
GC_10_377 b_10 NI_10 NS_377 0 -8.4240919624936235e-07
GC_10_378 b_10 NI_10 NS_378 0 1.3600821991339907e-06
GC_10_379 b_10 NI_10 NS_379 0 9.0836750885493792e-07
GC_10_380 b_10 NI_10 NS_380 0 1.8504793646667519e-06
GC_10_381 b_10 NI_10 NS_381 0 -7.6710503249460834e-07
GC_10_382 b_10 NI_10 NS_382 0 5.7087097917879402e-07
GC_10_383 b_10 NI_10 NS_383 0 -8.0356110607436406e-07
GC_10_384 b_10 NI_10 NS_384 0 1.5919272107558748e-06
GC_10_385 b_10 NI_10 NS_385 0 1.2779892185741621e-06
GC_10_386 b_10 NI_10 NS_386 0 5.6822833482548029e-07
GC_10_387 b_10 NI_10 NS_387 0 -6.6680311187522927e-07
GC_10_388 b_10 NI_10 NS_388 0 6.5598677171597432e-07
GC_10_389 b_10 NI_10 NS_389 0 5.3996076731832292e-07
GC_10_390 b_10 NI_10 NS_390 0 1.7896996108890446e-06
GC_10_391 b_10 NI_10 NS_391 0 -2.5639117768020130e-07
GC_10_392 b_10 NI_10 NS_392 0 -3.2550602044478226e-07
GC_10_393 b_10 NI_10 NS_393 0 -4.7492387217527699e-07
GC_10_394 b_10 NI_10 NS_394 0 6.1074272694250184e-07
GC_10_395 b_10 NI_10 NS_395 0 1.1438524523975435e-07
GC_10_396 b_10 NI_10 NS_396 0 5.8913341759661273e-07
GC_10_397 b_10 NI_10 NS_397 0 -3.1820144433433134e-07
GC_10_398 b_10 NI_10 NS_398 0 4.4618023716200336e-07
GC_10_399 b_10 NI_10 NS_399 0 6.3950306596320749e-08
GC_10_400 b_10 NI_10 NS_400 0 2.2647532618326536e-07
GC_10_401 b_10 NI_10 NS_401 0 -6.7253818092280791e-07
GC_10_402 b_10 NI_10 NS_402 0 2.4744292896819104e-07
GC_10_403 b_10 NI_10 NS_403 0 -1.6416019577283530e-07
GC_10_404 b_10 NI_10 NS_404 0 5.7606109555119905e-07
GC_10_405 b_10 NI_10 NS_405 0 -3.0458062962460850e-07
GC_10_406 b_10 NI_10 NS_406 0 2.5969235446821322e-07
GC_10_407 b_10 NI_10 NS_407 0 -9.8766963657604588e-08
GC_10_408 b_10 NI_10 NS_408 0 2.0869421615237375e-07
GC_10_409 b_10 NI_10 NS_409 0 -7.6623270341429134e-07
GC_10_410 b_10 NI_10 NS_410 0 5.3639713138339777e-08
GC_10_411 b_10 NI_10 NS_411 0 -4.8039104289140095e-07
GC_10_412 b_10 NI_10 NS_412 0 4.3217423456070499e-07
GC_10_413 b_10 NI_10 NS_413 0 -5.3152812493496467e-07
GC_10_414 b_10 NI_10 NS_414 0 2.1427236590764409e-07
GC_10_415 b_10 NI_10 NS_415 0 -5.2278837067383255e-07
GC_10_416 b_10 NI_10 NS_416 0 1.4454166646075546e-07
GC_10_417 b_10 NI_10 NS_417 0 -1.0033849103695405e-06
GC_10_418 b_10 NI_10 NS_418 0 -3.4734932437484340e-07
GC_10_419 b_10 NI_10 NS_419 0 -1.4397696731828185e-06
GC_10_420 b_10 NI_10 NS_420 0 5.4836664748643148e-07
GC_10_421 b_10 NI_10 NS_421 0 -1.1943883902071787e-06
GC_10_422 b_10 NI_10 NS_422 0 1.3609843632082551e-07
GC_10_423 b_10 NI_10 NS_423 0 -1.4806566628860723e-06
GC_10_424 b_10 NI_10 NS_424 0 7.7902408153874046e-07
GC_10_425 b_10 NI_10 NS_425 0 -2.2609433586651506e-06
GC_10_426 b_10 NI_10 NS_426 0 -8.4608319743100696e-07
GC_10_427 b_10 NI_10 NS_427 0 5.6638037179555604e-06
GC_10_428 b_10 NI_10 NS_428 0 1.1197138037696441e-05
GC_10_429 b_10 NI_10 NS_429 0 -2.2219655331121259e-06
GC_10_430 b_10 NI_10 NS_430 0 3.0963831015458493e-06
GC_10_431 b_10 NI_10 NS_431 0 1.1649814779462421e-08
GC_10_432 b_10 NI_10 NS_432 0 7.3477924756055766e-08
GC_10_433 b_10 NI_10 NS_433 0 -1.2473677402867223e-06
GC_10_434 b_10 NI_10 NS_434 0 1.6458030544194929e-06
GC_10_435 b_10 NI_10 NS_435 0 -6.3373475137545416e-07
GC_10_436 b_10 NI_10 NS_436 0 1.4520519918223930e-06
GC_10_437 b_10 NI_10 NS_437 0 -1.6479511415355572e-06
GC_10_438 b_10 NI_10 NS_438 0 -1.2214123114007827e-06
GC_10_439 b_10 NI_10 NS_439 0 -3.3894898432851765e-06
GC_10_440 b_10 NI_10 NS_440 0 -1.1083936000238382e-06
GC_10_441 b_10 NI_10 NS_441 0 7.1944918045719482e-09
GC_10_442 b_10 NI_10 NS_442 0 -1.2021669987144030e-07
GC_10_443 b_10 NI_10 NS_443 0 6.2008596995251484e-07
GC_10_444 b_10 NI_10 NS_444 0 -3.6780547767836943e-07
GC_10_445 b_10 NI_10 NS_445 0 -4.6880498169103736e-08
GC_10_446 b_10 NI_10 NS_446 0 3.9700348950169886e-07
GC_10_447 b_10 NI_10 NS_447 0 -5.1636700406534546e-08
GC_10_448 b_10 NI_10 NS_448 0 2.9619666824393344e-08
GC_10_449 b_10 NI_10 NS_449 0 -2.7362372843018544e-07
GC_10_450 b_10 NI_10 NS_450 0 1.7742432585102030e-07
GC_10_451 b_10 NI_10 NS_451 0 -2.2775884096956304e-07
GC_10_452 b_10 NI_10 NS_452 0 -6.5495360630964149e-09
GC_10_453 b_10 NI_10 NS_453 0 -8.0168023506537676e-12
GC_10_454 b_10 NI_10 NS_454 0 -8.1402869043672076e-13
GC_10_455 b_10 NI_10 NS_455 0 -1.1403329611539745e-09
GC_10_456 b_10 NI_10 NS_456 0 -2.4259801080780428e-09
GC_10_457 b_10 NI_10 NS_457 0 -3.2389974502221883e-05
GC_10_458 b_10 NI_10 NS_458 0 2.2145967009130675e-06
GC_10_459 b_10 NI_10 NS_459 0 6.9003316422542671e-11
GC_10_460 b_10 NI_10 NS_460 0 3.0548373837264004e-09
GC_10_461 b_10 NI_10 NS_461 0 -1.7288670868743920e-06
GC_10_462 b_10 NI_10 NS_462 0 -1.8218362019188048e-06
GC_10_463 b_10 NI_10 NS_463 0 -5.3710531896368151e-06
GC_10_464 b_10 NI_10 NS_464 0 2.8657834815324020e-06
GC_10_465 b_10 NI_10 NS_465 0 -1.6530932831995716e-05
GC_10_466 b_10 NI_10 NS_466 0 1.8435247673079520e-05
GC_10_467 b_10 NI_10 NS_467 0 1.5105428472839859e-05
GC_10_468 b_10 NI_10 NS_468 0 9.7996086710662168e-06
GC_10_469 b_10 NI_10 NS_469 0 1.7319499564464938e-05
GC_10_470 b_10 NI_10 NS_470 0 2.2757389030072377e-05
GC_10_471 b_10 NI_10 NS_471 0 2.9272126507735250e-05
GC_10_472 b_10 NI_10 NS_472 0 4.9456665872715460e-06
GC_10_473 b_10 NI_10 NS_473 0 -3.0091164954258030e-06
GC_10_474 b_10 NI_10 NS_474 0 -1.8920538317546962e-06
GC_10_475 b_10 NI_10 NS_475 0 1.6961530529784328e-05
GC_10_476 b_10 NI_10 NS_476 0 -2.2247619820703023e-06
GC_10_477 b_10 NI_10 NS_477 0 1.2893964023962944e-04
GC_10_478 b_10 NI_10 NS_478 0 3.4692029287842780e-05
GC_10_479 b_10 NI_10 NS_479 0 -2.8903411085923844e-05
GC_10_480 b_10 NI_10 NS_480 0 -9.8807188611716554e-05
GC_10_481 b_10 NI_10 NS_481 0 2.4942414461451039e-05
GC_10_482 b_10 NI_10 NS_482 0 -3.1439756800468188e-05
GC_10_483 b_10 NI_10 NS_483 0 -4.1725652482356032e-05
GC_10_484 b_10 NI_10 NS_484 0 -1.6659190411742384e-04
GC_10_485 b_10 NI_10 NS_485 0 -4.1856507250592021e-05
GC_10_486 b_10 NI_10 NS_486 0 -4.9686954907460089e-06
GC_10_487 b_10 NI_10 NS_487 0 2.1526362443299074e-05
GC_10_488 b_10 NI_10 NS_488 0 -1.5189810732891851e-04
GC_10_489 b_10 NI_10 NS_489 0 -2.3067319251690927e-04
GC_10_490 b_10 NI_10 NS_490 0 1.1454500857731533e-04
GC_10_491 b_10 NI_10 NS_491 0 -3.7434335174917871e-05
GC_10_492 b_10 NI_10 NS_492 0 1.4285229464253979e-05
GC_10_493 b_10 NI_10 NS_493 0 -1.3769141305538604e-04
GC_10_494 b_10 NI_10 NS_494 0 1.3059618042209032e-04
GC_10_495 b_10 NI_10 NS_495 0 3.6482050737766318e-05
GC_10_496 b_10 NI_10 NS_496 0 4.1333285293284282e-05
GC_10_497 b_10 NI_10 NS_497 0 -3.8174086623468575e-05
GC_10_498 b_10 NI_10 NS_498 0 4.3297473346981236e-05
GC_10_499 b_10 NI_10 NS_499 0 8.7698359711752057e-05
GC_10_500 b_10 NI_10 NS_500 0 1.1839031238995674e-04
GC_10_501 b_10 NI_10 NS_501 0 2.7360612959487369e-05
GC_10_502 b_10 NI_10 NS_502 0 1.0188100790386358e-05
GC_10_503 b_10 NI_10 NS_503 0 8.7309714542693488e-05
GC_10_504 b_10 NI_10 NS_504 0 6.5588845899845649e-05
GC_10_505 b_10 NI_10 NS_505 0 2.0355360933398170e-05
GC_10_506 b_10 NI_10 NS_506 0 -5.7134031164321949e-05
GC_10_507 b_10 NI_10 NS_507 0 1.6985921912692275e-05
GC_10_508 b_10 NI_10 NS_508 0 -8.8834606061901057e-06
GC_10_509 b_10 NI_10 NS_509 0 8.5005635393730049e-06
GC_10_510 b_10 NI_10 NS_510 0 -3.2939557357715242e-05
GC_10_511 b_10 NI_10 NS_511 0 -8.8537842597458358e-06
GC_10_512 b_10 NI_10 NS_512 0 5.2634498184240111e-07
GC_10_513 b_10 NI_10 NS_513 0 -2.4131095081509925e-06
GC_10_514 b_10 NI_10 NS_514 0 8.5086293659092779e-06
GC_10_515 b_10 NI_10 NS_515 0 1.0220484830656530e-05
GC_10_516 b_10 NI_10 NS_516 0 6.0869799422349938e-06
GC_10_517 b_10 NI_10 NS_517 0 1.2161238350723526e-05
GC_10_518 b_10 NI_10 NS_518 0 -7.8265404236314022e-06
GC_10_519 b_10 NI_10 NS_519 0 -3.4879197426136550e-06
GC_10_520 b_10 NI_10 NS_520 0 -4.4672717138987877e-07
GC_10_521 b_10 NI_10 NS_521 0 2.4880758873233267e-06
GC_10_522 b_10 NI_10 NS_522 0 7.4078970364710457e-06
GC_10_523 b_10 NI_10 NS_523 0 1.3650684610456888e-05
GC_10_524 b_10 NI_10 NS_524 0 2.6358824256900554e-06
GC_10_525 b_10 NI_10 NS_525 0 4.5207281043601576e-06
GC_10_526 b_10 NI_10 NS_526 0 -1.4188660962500318e-05
GC_10_527 b_10 NI_10 NS_527 0 -5.9269895484773369e-06
GC_10_528 b_10 NI_10 NS_528 0 4.2582615316445775e-06
GC_10_529 b_10 NI_10 NS_529 0 1.0309892907974963e-05
GC_10_530 b_10 NI_10 NS_530 0 9.9374583190469039e-06
GC_10_531 b_10 NI_10 NS_531 0 1.7307676827728319e-05
GC_10_532 b_10 NI_10 NS_532 0 -4.2709478737764331e-06
GC_10_533 b_10 NI_10 NS_533 0 -9.2921149939368261e-06
GC_10_534 b_10 NI_10 NS_534 0 -1.5315721932597516e-05
GC_10_535 b_10 NI_10 NS_535 0 -4.0817850412987391e-06
GC_10_536 b_10 NI_10 NS_536 0 1.3516462490615352e-05
GC_10_537 b_10 NI_10 NS_537 0 2.0928880153636002e-05
GC_10_538 b_10 NI_10 NS_538 0 -5.6272479649021733e-07
GC_10_539 b_10 NI_10 NS_539 0 8.8752265282926065e-06
GC_10_540 b_10 NI_10 NS_540 0 -1.7452662792171185e-05
GC_10_541 b_10 NI_10 NS_541 0 2.4046508519929129e-06
GC_10_542 b_10 NI_10 NS_542 0 -1.3697829013681407e-05
GC_10_543 b_10 NI_10 NS_543 0 -1.3815733182847775e-05
GC_10_544 b_10 NI_10 NS_544 0 4.3766471073644000e-06
GC_10_545 b_10 NI_10 NS_545 0 1.5474916554983773e-08
GC_10_546 b_10 NI_10 NS_546 0 -4.2109927868921434e-08
GC_10_547 b_10 NI_10 NS_547 0 8.6210497250404280e-06
GC_10_548 b_10 NI_10 NS_548 0 1.1597864434486722e-05
GC_10_549 b_10 NI_10 NS_549 0 1.0904639560444432e-05
GC_10_550 b_10 NI_10 NS_550 0 -1.1278376488113791e-05
GC_10_551 b_10 NI_10 NS_551 0 -3.7306486876522349e-06
GC_10_552 b_10 NI_10 NS_552 0 -1.0216313648449865e-05
GC_10_553 b_10 NI_10 NS_553 0 -2.2939446048296910e-06
GC_10_554 b_10 NI_10 NS_554 0 1.2865853068045407e-05
GC_10_555 b_10 NI_10 NS_555 0 9.6692486309210434e-07
GC_10_556 b_10 NI_10 NS_556 0 -7.2694842129671858e-06
GC_10_557 b_10 NI_10 NS_557 0 7.5166672040590454e-06
GC_10_558 b_10 NI_10 NS_558 0 1.6932076312693757e-06
GC_10_559 b_10 NI_10 NS_559 0 -6.1012275295067497e-06
GC_10_560 b_10 NI_10 NS_560 0 -8.8953906675978644e-06
GC_10_561 b_10 NI_10 NS_561 0 -4.1215016564640965e-06
GC_10_562 b_10 NI_10 NS_562 0 9.6659699045377215e-06
GC_10_563 b_10 NI_10 NS_563 0 3.3268384836576660e-06
GC_10_564 b_10 NI_10 NS_564 0 6.0367149464996757e-06
GC_10_565 b_10 NI_10 NS_565 0 5.6518830304141353e-06
GC_10_566 b_10 NI_10 NS_566 0 5.1680983173980033e-07
GC_10_567 b_10 NI_10 NS_567 0 6.1804964637194873e-11
GC_10_568 b_10 NI_10 NS_568 0 1.4894763316179579e-10
GC_10_569 b_10 NI_10 NS_569 0 5.9431497211701728e-09
GC_10_570 b_10 NI_10 NS_570 0 -8.3385338908140002e-09
GC_10_571 b_10 NI_10 NS_571 0 -1.1776551461720217e-04
GC_10_572 b_10 NI_10 NS_572 0 -2.1390368515459633e-06
GC_10_573 b_10 NI_10 NS_573 0 -2.5034436131423259e-10
GC_10_574 b_10 NI_10 NS_574 0 2.5994078450878429e-09
GC_10_575 b_10 NI_10 NS_575 0 1.6865026238180974e-06
GC_10_576 b_10 NI_10 NS_576 0 -1.5557519362165553e-06
GC_10_577 b_10 NI_10 NS_577 0 1.0498558843242763e-07
GC_10_578 b_10 NI_10 NS_578 0 -6.3346749929243938e-06
GC_10_579 b_10 NI_10 NS_579 0 -7.5924902663616430e-06
GC_10_580 b_10 NI_10 NS_580 0 2.3113173326033996e-07
GC_10_581 b_10 NI_10 NS_581 0 -1.1742330362450999e-06
GC_10_582 b_10 NI_10 NS_582 0 -4.6213207581394862e-06
GC_10_583 b_10 NI_10 NS_583 0 -1.5831640687897620e-05
GC_10_584 b_10 NI_10 NS_584 0 -1.5727949115492175e-06
GC_10_585 b_10 NI_10 NS_585 0 -6.0025250449227453e-06
GC_10_586 b_10 NI_10 NS_586 0 1.9095125165787802e-05
GC_10_587 b_10 NI_10 NS_587 0 4.6272149776709703e-06
GC_10_588 b_10 NI_10 NS_588 0 -3.0068109908687378e-06
GC_10_589 b_10 NI_10 NS_589 0 -1.4071465114005033e-08
GC_10_590 b_10 NI_10 NS_590 0 -2.6089082315928240e-06
GC_10_591 b_10 NI_10 NS_591 0 -2.5759905823740121e-05
GC_10_592 b_10 NI_10 NS_592 0 2.8490204435505850e-05
GC_10_593 b_10 NI_10 NS_593 0 2.8211388188237114e-05
GC_10_594 b_10 NI_10 NS_594 0 -8.6038970174859051e-06
GC_10_595 b_10 NI_10 NS_595 0 -8.0514515941833058e-06
GC_10_596 b_10 NI_10 NS_596 0 -4.3168390762385454e-06
GC_10_597 b_10 NI_10 NS_597 0 1.2692846224078782e-05
GC_10_598 b_10 NI_10 NS_598 0 2.6907360012001874e-05
GC_10_599 b_10 NI_10 NS_599 0 1.4541619814496883e-06
GC_10_600 b_10 NI_10 NS_600 0 -9.0171640421720176e-06
GC_10_601 b_10 NI_10 NS_601 0 -2.8297055007021552e-05
GC_10_602 b_10 NI_10 NS_602 0 4.7690831571145489e-06
GC_10_603 b_10 NI_10 NS_603 0 4.1340036151944069e-05
GC_10_604 b_10 NI_10 NS_604 0 1.0566874579290607e-05
GC_10_605 b_10 NI_10 NS_605 0 -2.9777178476171994e-06
GC_10_606 b_10 NI_10 NS_606 0 -4.5076722961716897e-06
GC_10_607 b_10 NI_10 NS_607 0 1.2968810375095684e-05
GC_10_608 b_10 NI_10 NS_608 0 1.8946405469852699e-05
GC_10_609 b_10 NI_10 NS_609 0 3.7956313627462358e-06
GC_10_610 b_10 NI_10 NS_610 0 -1.0952540345334997e-05
GC_10_611 b_10 NI_10 NS_611 0 -6.4190507922680981e-06
GC_10_612 b_10 NI_10 NS_612 0 8.3208976578062671e-07
GC_10_613 b_10 NI_10 NS_613 0 1.8890182720098678e-05
GC_10_614 b_10 NI_10 NS_614 0 5.3956718038971199e-06
GC_10_615 b_10 NI_10 NS_615 0 -7.6255020815251924e-08
GC_10_616 b_10 NI_10 NS_616 0 -4.2077104724770865e-06
GC_10_617 b_10 NI_10 NS_617 0 4.9306595611388882e-06
GC_10_618 b_10 NI_10 NS_618 0 1.4263142570829639e-05
GC_10_619 b_10 NI_10 NS_619 0 7.8225222619777397e-06
GC_10_620 b_10 NI_10 NS_620 0 -1.1202028010026539e-05
GC_10_621 b_10 NI_10 NS_621 0 -1.3847719303184284e-06
GC_10_622 b_10 NI_10 NS_622 0 9.2712254971477811e-07
GC_10_623 b_10 NI_10 NS_623 0 1.0915582198909381e-05
GC_10_624 b_10 NI_10 NS_624 0 4.0962626104606264e-06
GC_10_625 b_10 NI_10 NS_625 0 1.7204806914048593e-06
GC_10_626 b_10 NI_10 NS_626 0 -6.4492695062307245e-07
GC_10_627 b_10 NI_10 NS_627 0 5.6901266733296360e-06
GC_10_628 b_10 NI_10 NS_628 0 1.6919134498159918e-06
GC_10_629 b_10 NI_10 NS_629 0 3.4275670794771960e-06
GC_10_630 b_10 NI_10 NS_630 0 2.0300852800046538e-06
GC_10_631 b_10 NI_10 NS_631 0 1.0987681049266041e-05
GC_10_632 b_10 NI_10 NS_632 0 3.7699911387628219e-06
GC_10_633 b_10 NI_10 NS_633 0 4.8689033424170457e-06
GC_10_634 b_10 NI_10 NS_634 0 -9.2939730933963618e-08
GC_10_635 b_10 NI_10 NS_635 0 9.9989118537185802e-06
GC_10_636 b_10 NI_10 NS_636 0 -1.0950577426235229e-06
GC_10_637 b_10 NI_10 NS_637 0 8.2824377005002641e-06
GC_10_638 b_10 NI_10 NS_638 0 2.9417405465178048e-06
GC_10_639 b_10 NI_10 NS_639 0 1.9094674823090674e-05
GC_10_640 b_10 NI_10 NS_640 0 -5.5863941180706701e-06
GC_10_641 b_10 NI_10 NS_641 0 7.2293231682137443e-06
GC_10_642 b_10 NI_10 NS_642 0 -4.0341369126695585e-06
GC_10_643 b_10 NI_10 NS_643 0 1.3781905581504494e-05
GC_10_644 b_10 NI_10 NS_644 0 -1.1917593506685299e-05
GC_10_645 b_10 NI_10 NS_645 0 1.2441236798984121e-05
GC_10_646 b_10 NI_10 NS_646 0 -3.9380664873189161e-06
GC_10_647 b_10 NI_10 NS_647 0 9.3021680213687537e-06
GC_10_648 b_10 NI_10 NS_648 0 -2.6814459397140017e-05
GC_10_649 b_10 NI_10 NS_649 0 2.4411468785506072e-06
GC_10_650 b_10 NI_10 NS_650 0 -1.2372670222207556e-05
GC_10_651 b_10 NI_10 NS_651 0 -8.1267819259083364e-06
GC_10_652 b_10 NI_10 NS_652 0 -1.8722451416533736e-05
GC_10_653 b_10 NI_10 NS_653 0 -4.6961711209198162e-06
GC_10_654 b_10 NI_10 NS_654 0 -1.1981122996537474e-05
GC_10_655 b_10 NI_10 NS_655 0 5.4399751296180106e-05
GC_10_656 b_10 NI_10 NS_656 0 -8.9383199208204804e-05
GC_10_657 b_10 NI_10 NS_657 0 -9.7660123324562107e-06
GC_10_658 b_10 NI_10 NS_658 0 9.8738767200171019e-07
GC_10_659 b_10 NI_10 NS_659 0 3.8976890424328567e-07
GC_10_660 b_10 NI_10 NS_660 0 -1.3364778388710622e-07
GC_10_661 b_10 NI_10 NS_661 0 -2.5756629382340502e-06
GC_10_662 b_10 NI_10 NS_662 0 -2.1120209498830940e-06
GC_10_663 b_10 NI_10 NS_663 0 -4.3189711203575308e-06
GC_10_664 b_10 NI_10 NS_664 0 3.8846841584597188e-07
GC_10_665 b_10 NI_10 NS_665 0 -1.7308660635894613e-05
GC_10_666 b_10 NI_10 NS_666 0 9.7288645157079538e-06
GC_10_667 b_10 NI_10 NS_667 0 -8.8649391894937442e-06
GC_10_668 b_10 NI_10 NS_668 0 3.7519899851562219e-05
GC_10_669 b_10 NI_10 NS_669 0 -7.2572372364732125e-06
GC_10_670 b_10 NI_10 NS_670 0 3.2751347239825551e-07
GC_10_671 b_10 NI_10 NS_671 0 -1.3477623905567284e-05
GC_10_672 b_10 NI_10 NS_672 0 1.9011794892823876e-06
GC_10_673 b_10 NI_10 NS_673 0 -4.6310018894736851e-06
GC_10_674 b_10 NI_10 NS_674 0 -3.4347516693066980e-06
GC_10_675 b_10 NI_10 NS_675 0 -6.4037965310354422e-06
GC_10_676 b_10 NI_10 NS_676 0 1.0107229840919118e-06
GC_10_677 b_10 NI_10 NS_677 0 -3.0174080581711607e-06
GC_10_678 b_10 NI_10 NS_678 0 8.7541100383846798e-07
GC_10_679 b_10 NI_10 NS_679 0 -1.7610332385599502e-06
GC_10_680 b_10 NI_10 NS_680 0 -9.6128228626078696e-07
GC_10_681 b_10 NI_10 NS_681 0 -2.6099340575917180e-10
GC_10_682 b_10 NI_10 NS_682 0 4.2237628183225884e-10
GC_10_683 b_10 NI_10 NS_683 0 2.2553960169049018e-09
GC_10_684 b_10 NI_10 NS_684 0 -2.6817127091618116e-08
GC_10_685 b_10 NI_10 NS_685 0 -2.0263963628982398e-04
GC_10_686 b_10 NI_10 NS_686 0 -3.3244780532495325e-06
GC_10_687 b_10 NI_10 NS_687 0 1.2949489848671545e-09
GC_10_688 b_10 NI_10 NS_688 0 9.6762672090673728e-09
GC_10_689 b_10 NI_10 NS_689 0 -4.1489176135951258e-06
GC_10_690 b_10 NI_10 NS_690 0 6.1899620056422917e-06
GC_10_691 b_10 NI_10 NS_691 0 3.7984415510072006e-06
GC_10_692 b_10 NI_10 NS_692 0 -8.1732064404747184e-06
GC_10_693 b_10 NI_10 NS_693 0 2.1695002639545139e-05
GC_10_694 b_10 NI_10 NS_694 0 -8.8474241196300580e-06
GC_10_695 b_10 NI_10 NS_695 0 -2.1457573908123663e-05
GC_10_696 b_10 NI_10 NS_696 0 -1.1750548194464220e-06
GC_10_697 b_10 NI_10 NS_697 0 -2.9650340654350850e-05
GC_10_698 b_10 NI_10 NS_698 0 -2.8288024542408708e-05
GC_10_699 b_10 NI_10 NS_699 0 -5.5338667599008491e-06
GC_10_700 b_10 NI_10 NS_700 0 1.6528825236645039e-05
GC_10_701 b_10 NI_10 NS_701 0 -2.4253110908661133e-06
GC_10_702 b_10 NI_10 NS_702 0 -7.1416175746950210e-06
GC_10_703 b_10 NI_10 NS_703 0 -2.2543160497000961e-05
GC_10_704 b_10 NI_10 NS_704 0 6.0040521753633361e-06
GC_10_705 b_10 NI_10 NS_705 0 -1.8562633180392696e-04
GC_10_706 b_10 NI_10 NS_706 0 -4.4048585383783577e-05
GC_10_707 b_10 NI_10 NS_707 0 6.2607976114367238e-05
GC_10_708 b_10 NI_10 NS_708 0 1.3739432914795032e-04
GC_10_709 b_10 NI_10 NS_709 0 -3.7276505808107970e-05
GC_10_710 b_10 NI_10 NS_710 0 5.6604129926282646e-05
GC_10_711 b_10 NI_10 NS_711 0 9.5167630553905387e-05
GC_10_712 b_10 NI_10 NS_712 0 2.4608316035922413e-04
GC_10_713 b_10 NI_10 NS_713 0 7.3783611630807289e-05
GC_10_714 b_10 NI_10 NS_714 0 4.9169983124307951e-07
GC_10_715 b_10 NI_10 NS_715 0 -1.5399686000653092e-05
GC_10_716 b_10 NI_10 NS_716 0 2.6123481919894089e-04
GC_10_717 b_10 NI_10 NS_717 0 3.6434226552072057e-04
GC_10_718 b_10 NI_10 NS_718 0 -2.4310562774006210e-04
GC_10_719 b_10 NI_10 NS_719 0 6.5642863025694277e-05
GC_10_720 b_10 NI_10 NS_720 0 -2.8524091572626553e-05
GC_10_721 b_10 NI_10 NS_721 0 2.0802916845815840e-04
GC_10_722 b_10 NI_10 NS_722 0 -2.4138717244711347e-04
GC_10_723 b_10 NI_10 NS_723 0 -7.1282968537476226e-05
GC_10_724 b_10 NI_10 NS_724 0 -7.1463392760900507e-05
GC_10_725 b_10 NI_10 NS_725 0 6.4487018401072246e-05
GC_10_726 b_10 NI_10 NS_726 0 -7.5529274046343847e-05
GC_10_727 b_10 NI_10 NS_727 0 -1.7047212365183209e-04
GC_10_728 b_10 NI_10 NS_728 0 -1.8309631777007365e-04
GC_10_729 b_10 NI_10 NS_729 0 -4.8833094147667620e-05
GC_10_730 b_10 NI_10 NS_730 0 -1.9097917163061292e-05
GC_10_731 b_10 NI_10 NS_731 0 -1.4491742456254365e-04
GC_10_732 b_10 NI_10 NS_732 0 -9.5347160799139039e-05
GC_10_733 b_10 NI_10 NS_733 0 -2.7318506925979338e-05
GC_10_734 b_10 NI_10 NS_734 0 1.0360166417973302e-04
GC_10_735 b_10 NI_10 NS_735 0 -2.7242628494026643e-05
GC_10_736 b_10 NI_10 NS_736 0 1.3907339355548771e-05
GC_10_737 b_10 NI_10 NS_737 0 2.1261971449045688e-06
GC_10_738 b_10 NI_10 NS_738 0 5.0767019133639894e-05
GC_10_739 b_10 NI_10 NS_739 0 1.6811819638257065e-05
GC_10_740 b_10 NI_10 NS_740 0 -5.9722075951259808e-07
GC_10_741 b_10 NI_10 NS_741 0 1.8082649041348037e-06
GC_10_742 b_10 NI_10 NS_742 0 -1.5452703432938696e-05
GC_10_743 b_10 NI_10 NS_743 0 -1.5113318494782255e-05
GC_10_744 b_10 NI_10 NS_744 0 -1.3586604188668553e-05
GC_10_745 b_10 NI_10 NS_745 0 -1.3111591995046604e-05
GC_10_746 b_10 NI_10 NS_746 0 1.2341873844998559e-05
GC_10_747 b_10 NI_10 NS_747 0 7.7827968323684235e-06
GC_10_748 b_10 NI_10 NS_748 0 1.2547800048416064e-06
GC_10_749 b_10 NI_10 NS_749 0 -5.1388190424279550e-06
GC_10_750 b_10 NI_10 NS_750 0 -1.2683796289690612e-05
GC_10_751 b_10 NI_10 NS_751 0 -2.0805173053355698e-05
GC_10_752 b_10 NI_10 NS_752 0 -5.8763644860211728e-06
GC_10_753 b_10 NI_10 NS_753 0 1.0765874701110819e-06
GC_10_754 b_10 NI_10 NS_754 0 2.1822936112556163e-05
GC_10_755 b_10 NI_10 NS_755 0 1.2863935780003859e-05
GC_10_756 b_10 NI_10 NS_756 0 -6.8611685637603265e-06
GC_10_757 b_10 NI_10 NS_757 0 -1.7284419626354100e-05
GC_10_758 b_10 NI_10 NS_758 0 -1.5977690652121488e-05
GC_10_759 b_10 NI_10 NS_759 0 -2.7118726313694003e-05
GC_10_760 b_10 NI_10 NS_760 0 8.8182311606614176e-06
GC_10_761 b_10 NI_10 NS_761 0 2.7088809810657749e-05
GC_10_762 b_10 NI_10 NS_762 0 2.2448437367663997e-05
GC_10_763 b_10 NI_10 NS_763 0 1.0940725251332743e-05
GC_10_764 b_10 NI_10 NS_764 0 -2.1302018937095683e-05
GC_10_765 b_10 NI_10 NS_765 0 -3.0617491319202968e-05
GC_10_766 b_10 NI_10 NS_766 0 3.9079209185197667e-06
GC_10_767 b_10 NI_10 NS_767 0 -9.8041691949897935e-06
GC_10_768 b_10 NI_10 NS_768 0 3.9250448242771024e-05
GC_10_769 b_10 NI_10 NS_769 0 1.9741565775743468e-05
GC_10_770 b_10 NI_10 NS_770 0 -6.8523910249076818e-05
GC_10_771 b_10 NI_10 NS_771 0 4.3396457579440968e-05
GC_10_772 b_10 NI_10 NS_772 0 -1.6864115259784935e-05
GC_10_773 b_10 NI_10 NS_773 0 2.0643883791562192e-07
GC_10_774 b_10 NI_10 NS_774 0 -2.4337034284896838e-07
GC_10_775 b_10 NI_10 NS_775 0 -3.6341780228727793e-06
GC_10_776 b_10 NI_10 NS_776 0 -2.0830491939960720e-05
GC_10_777 b_10 NI_10 NS_777 0 -1.0493729410382638e-05
GC_10_778 b_10 NI_10 NS_778 0 1.6700704299302682e-05
GC_10_779 b_10 NI_10 NS_779 0 9.1927140700557514e-06
GC_10_780 b_10 NI_10 NS_780 0 3.1865113979895401e-05
GC_10_781 b_10 NI_10 NS_781 0 1.4275077678599970e-05
GC_10_782 b_10 NI_10 NS_782 0 -3.0125662154022213e-06
GC_10_783 b_10 NI_10 NS_783 0 -3.9047775616605914e-06
GC_10_784 b_10 NI_10 NS_784 0 1.2499363510117550e-05
GC_10_785 b_10 NI_10 NS_785 0 -1.8573490083046014e-05
GC_10_786 b_10 NI_10 NS_786 0 -3.6270080883277521e-06
GC_10_787 b_10 NI_10 NS_787 0 1.3215675485141635e-05
GC_10_788 b_10 NI_10 NS_788 0 1.3176843427005795e-05
GC_10_789 b_10 NI_10 NS_789 0 7.6359157351265730e-06
GC_10_790 b_10 NI_10 NS_790 0 -2.3019060497659072e-05
GC_10_791 b_10 NI_10 NS_791 0 -3.8460168433091301e-06
GC_10_792 b_10 NI_10 NS_792 0 -1.1722919120261895e-05
GC_10_793 b_10 NI_10 NS_793 0 -8.7362198271700651e-06
GC_10_794 b_10 NI_10 NS_794 0 -2.6278894811769813e-06
GC_10_795 b_10 NI_10 NS_795 0 5.5142464303504647e-10
GC_10_796 b_10 NI_10 NS_796 0 2.9347469013933922e-10
GC_10_797 b_10 NI_10 NS_797 0 4.2109542589220991e-08
GC_10_798 b_10 NI_10 NS_798 0 3.6939224436857854e-08
GC_10_799 b_10 NI_10 NS_799 0 2.8651768438229825e-04
GC_10_800 b_10 NI_10 NS_800 0 -1.4350270448486925e-05
GC_10_801 b_10 NI_10 NS_801 0 -1.2376921224925990e-09
GC_10_802 b_10 NI_10 NS_802 0 -1.9231838034228682e-08
GC_10_803 b_10 NI_10 NS_803 0 2.6656319935377171e-06
GC_10_804 b_10 NI_10 NS_804 0 -3.8233434185388790e-06
GC_10_805 b_10 NI_10 NS_805 0 -1.3224305989273408e-05
GC_10_806 b_10 NI_10 NS_806 0 -5.0206338989427430e-07
GC_10_807 b_10 NI_10 NS_807 0 3.9456084812921974e-05
GC_10_808 b_10 NI_10 NS_808 0 2.7908358420999095e-06
GC_10_809 b_10 NI_10 NS_809 0 -4.1773666439223985e-05
GC_10_810 b_10 NI_10 NS_810 0 -2.3731190971672866e-05
GC_10_811 b_10 NI_10 NS_811 0 1.7633809429442870e-06
GC_10_812 b_10 NI_10 NS_812 0 4.4847668927322557e-05
GC_10_813 b_10 NI_10 NS_813 0 1.4507221252490528e-05
GC_10_814 b_10 NI_10 NS_814 0 -4.8182186918792043e-05
GC_10_815 b_10 NI_10 NS_815 0 1.9346478886634887e-06
GC_10_816 b_10 NI_10 NS_816 0 5.6524855560923454e-06
GC_10_817 b_10 NI_10 NS_817 0 -4.4992649112913179e-05
GC_10_818 b_10 NI_10 NS_818 0 1.5680701338528858e-06
GC_10_819 b_10 NI_10 NS_819 0 1.0311100372429572e-04
GC_10_820 b_10 NI_10 NS_820 0 1.2335725378699738e-04
GC_10_821 b_10 NI_10 NS_821 0 -7.5524315876189873e-05
GC_10_822 b_10 NI_10 NS_822 0 -1.3698768782838329e-04
GC_10_823 b_10 NI_10 NS_823 0 -6.7108091699533799e-05
GC_10_824 b_10 NI_10 NS_824 0 4.9269053939498822e-05
GC_10_825 b_10 NI_10 NS_825 0 1.3517316951942740e-04
GC_10_826 b_10 NI_10 NS_826 0 -2.8539512828524372e-05
GC_10_827 b_10 NI_10 NS_827 0 -8.7330355738415131e-05
GC_10_828 b_10 NI_10 NS_828 0 -1.1763765248760676e-05
GC_10_829 b_10 NI_10 NS_829 0 -9.4644586909568645e-05
GC_10_830 b_10 NI_10 NS_830 0 2.1148789535736063e-04
GC_10_831 b_10 NI_10 NS_831 0 1.6429528244631033e-04
GC_10_832 b_10 NI_10 NS_832 0 -2.1487718437087833e-04
GC_10_833 b_10 NI_10 NS_833 0 -8.1683784350222531e-05
GC_10_834 b_10 NI_10 NS_834 0 1.9188652314575233e-05
GC_10_835 b_10 NI_10 NS_835 0 1.6096945080755861e-04
GC_10_836 b_10 NI_10 NS_836 0 4.2088604071384386e-05
GC_10_837 b_10 NI_10 NS_837 0 -8.8878228113558043e-05
GC_10_838 b_10 NI_10 NS_838 0 -7.1909714175783919e-05
GC_10_839 b_10 NI_10 NS_839 0 -8.4866179898445841e-05
GC_10_840 b_10 NI_10 NS_840 0 6.3595962066375326e-05
GC_10_841 b_10 NI_10 NS_841 0 1.4068739980874366e-04
GC_10_842 b_10 NI_10 NS_842 0 -4.8520533829852498e-05
GC_10_843 b_10 NI_10 NS_843 0 -6.6207336013452642e-05
GC_10_844 b_10 NI_10 NS_844 0 -2.4251182959761381e-05
GC_10_845 b_10 NI_10 NS_845 0 6.1224274376909453e-05
GC_10_846 b_10 NI_10 NS_846 0 1.1375729331985532e-04
GC_10_847 b_10 NI_10 NS_847 0 -2.2917748216958931e-05
GC_10_848 b_10 NI_10 NS_848 0 -1.2153249744517164e-04
GC_10_849 b_10 NI_10 NS_849 0 -4.4313280189284081e-05
GC_10_850 b_10 NI_10 NS_850 0 1.0974879882650974e-05
GC_10_851 b_10 NI_10 NS_851 0 4.7535701858958794e-05
GC_10_852 b_10 NI_10 NS_852 0 -1.0608044856660445e-05
GC_10_853 b_10 NI_10 NS_853 0 -3.2085808510156403e-05
GC_10_854 b_10 NI_10 NS_854 0 -7.6434683715659013e-06
GC_10_855 b_10 NI_10 NS_855 0 2.1333627514217371e-05
GC_10_856 b_10 NI_10 NS_856 0 -4.8747026035539158e-06
GC_10_857 b_10 NI_10 NS_857 0 -3.2213267134371418e-05
GC_10_858 b_10 NI_10 NS_858 0 -2.5250971007912633e-05
GC_10_859 b_10 NI_10 NS_859 0 1.2710451843713451e-05
GC_10_860 b_10 NI_10 NS_860 0 6.1766879515726346e-06
GC_10_861 b_10 NI_10 NS_861 0 -2.0358851534567794e-05
GC_10_862 b_10 NI_10 NS_862 0 -7.7255063887856975e-06
GC_10_863 b_10 NI_10 NS_863 0 1.4086791184870683e-05
GC_10_864 b_10 NI_10 NS_864 0 -1.2504716650363657e-05
GC_10_865 b_10 NI_10 NS_865 0 -4.1281855301042332e-05
GC_10_866 b_10 NI_10 NS_866 0 -1.6953860513389984e-05
GC_10_867 b_10 NI_10 NS_867 0 1.1908060172564644e-05
GC_10_868 b_10 NI_10 NS_868 0 -1.7650834808358253e-06
GC_10_869 b_10 NI_10 NS_869 0 -3.0212165036005371e-05
GC_10_870 b_10 NI_10 NS_870 0 5.5332080102369234e-06
GC_10_871 b_10 NI_10 NS_871 0 1.6333206838547735e-05
GC_10_872 b_10 NI_10 NS_872 0 -2.0848888600911417e-05
GC_10_873 b_10 NI_10 NS_873 0 -4.9845705923767752e-05
GC_10_874 b_10 NI_10 NS_874 0 -1.6671132723826352e-06
GC_10_875 b_10 NI_10 NS_875 0 1.2248920898216945e-05
GC_10_876 b_10 NI_10 NS_876 0 -1.1718134812977420e-05
GC_10_877 b_10 NI_10 NS_877 0 -3.1907776896236733e-05
GC_10_878 b_10 NI_10 NS_878 0 2.5076448373737974e-05
GC_10_879 b_10 NI_10 NS_879 0 1.0836001565423488e-05
GC_10_880 b_10 NI_10 NS_880 0 -3.6497129665666970e-05
GC_10_881 b_10 NI_10 NS_881 0 -3.3854597050089454e-05
GC_10_882 b_10 NI_10 NS_882 0 1.8659942791585278e-05
GC_10_883 b_10 NI_10 NS_883 0 -5.9885035208891419e-05
GC_10_884 b_10 NI_10 NS_884 0 1.2846809764678762e-04
GC_10_885 b_10 NI_10 NS_885 0 -1.4510116856344772e-05
GC_10_886 b_10 NI_10 NS_886 0 -3.3372795603968142e-05
GC_10_887 b_10 NI_10 NS_887 0 -3.8792938731151877e-07
GC_10_888 b_10 NI_10 NS_888 0 3.6143459659618729e-07
GC_10_889 b_10 NI_10 NS_889 0 -1.9684608197340685e-05
GC_10_890 b_10 NI_10 NS_890 0 3.1288239076063724e-05
GC_10_891 b_10 NI_10 NS_891 0 -1.4242871927678666e-05
GC_10_892 b_10 NI_10 NS_892 0 -3.4197769822527202e-05
GC_10_893 b_10 NI_10 NS_893 0 -5.2907344102376377e-06
GC_10_894 b_10 NI_10 NS_894 0 5.5319735019986129e-06
GC_10_895 b_10 NI_10 NS_895 0 -1.9742370929042573e-05
GC_10_896 b_10 NI_10 NS_896 0 -6.5467166602342939e-05
GC_10_897 b_10 NI_10 NS_897 0 -9.2829821007292189e-06
GC_10_898 b_10 NI_10 NS_898 0 -2.0586456629480900e-05
GC_10_899 b_10 NI_10 NS_899 0 1.4777323901268116e-05
GC_10_900 b_10 NI_10 NS_900 0 2.2998758471097569e-05
GC_10_901 b_10 NI_10 NS_901 0 -6.8231217996964186e-06
GC_10_902 b_10 NI_10 NS_902 0 2.7592360454025724e-05
GC_10_903 b_10 NI_10 NS_903 0 -1.1136047017056686e-05
GC_10_904 b_10 NI_10 NS_904 0 -2.1577810516870336e-05
GC_10_905 b_10 NI_10 NS_905 0 -1.1024479589081584e-05
GC_10_906 b_10 NI_10 NS_906 0 2.3799265339339046e-05
GC_10_907 b_10 NI_10 NS_907 0 5.1499622761218124e-06
GC_10_908 b_10 NI_10 NS_908 0 -1.5352080888778858e-05
GC_10_909 b_10 NI_10 NS_909 0 -4.7263520771193302e-10
GC_10_910 b_10 NI_10 NS_910 0 -9.1862443785234280e-10
GC_10_911 b_10 NI_10 NS_911 0 -5.5412150347946333e-08
GC_10_912 b_10 NI_10 NS_912 0 7.6391281608963577e-09
GC_10_913 b_10 NI_10 NS_913 0 1.8435612387900820e-02
GC_10_914 b_10 NI_10 NS_914 0 6.7474792462818879e-03
GC_10_915 b_10 NI_10 NS_915 0 4.6857909521630048e-07
GC_10_916 b_10 NI_10 NS_916 0 1.4597166157385376e-06
GC_10_917 b_10 NI_10 NS_917 0 6.0883382547653603e-03
GC_10_918 b_10 NI_10 NS_918 0 1.8079600753466082e-03
GC_10_919 b_10 NI_10 NS_919 0 -6.0692580951308191e-03
GC_10_920 b_10 NI_10 NS_920 0 -6.1755768633673454e-04
GC_10_921 b_10 NI_10 NS_921 0 7.3052156135983513e-03
GC_10_922 b_10 NI_10 NS_922 0 -1.2868624824463194e-02
GC_10_923 b_10 NI_10 NS_923 0 8.4477683390281333e-03
GC_10_924 b_10 NI_10 NS_924 0 -2.4318274740153429e-04
GC_10_925 b_10 NI_10 NS_925 0 -9.6437905714249154e-03
GC_10_926 b_10 NI_10 NS_926 0 2.6145221996552327e-03
GC_10_927 b_10 NI_10 NS_927 0 -8.8622836153546044e-03
GC_10_928 b_10 NI_10 NS_928 0 -2.4394128248657040e-02
GC_10_929 b_10 NI_10 NS_929 0 -8.6175319273995978e-04
GC_10_930 b_10 NI_10 NS_930 0 4.1810854508503130e-03
GC_10_931 b_10 NI_10 NS_931 0 7.1873283396622235e-03
GC_10_932 b_10 NI_10 NS_932 0 -1.0295239433862347e-03
GC_10_933 b_10 NI_10 NS_933 0 -2.5161229319595312e-02
GC_10_934 b_10 NI_10 NS_934 0 4.8304471822816887e-03
GC_10_935 b_10 NI_10 NS_935 0 -1.9677030912687268e-02
GC_10_936 b_10 NI_10 NS_936 0 8.9707759594789143e-04
GC_10_937 b_10 NI_10 NS_937 0 1.0760310610544478e-02
GC_10_938 b_10 NI_10 NS_938 0 -2.7834508967899494e-03
GC_10_939 b_10 NI_10 NS_939 0 -4.7876006379652071e-03
GC_10_940 b_10 NI_10 NS_940 0 4.5022478041561544e-02
GC_10_941 b_10 NI_10 NS_941 0 -1.2656406134047442e-02
GC_10_942 b_10 NI_10 NS_942 0 -2.7339913069220518e-04
GC_10_943 b_10 NI_10 NS_943 0 1.5916761592030815e-02
GC_10_944 b_10 NI_10 NS_944 0 -4.0520346254961769e-03
GC_10_945 b_10 NI_10 NS_945 0 3.2201025794269068e-02
GC_10_946 b_10 NI_10 NS_946 0 1.8584534075239034e-02
GC_10_947 b_10 NI_10 NS_947 0 -1.2597833765416669e-02
GC_10_948 b_10 NI_10 NS_948 0 1.6053792226193483e-04
GC_10_949 b_10 NI_10 NS_949 0 1.7204328451060624e-02
GC_10_950 b_10 NI_10 NS_950 0 -3.5163060968447429e-02
GC_10_951 b_10 NI_10 NS_951 0 1.4015821086511384e-02
GC_10_952 b_10 NI_10 NS_952 0 4.7859336291068292e-03
GC_10_953 b_10 NI_10 NS_953 0 -1.4402607502130077e-02
GC_10_954 b_10 NI_10 NS_954 0 2.3853428762401867e-04
GC_10_955 b_10 NI_10 NS_955 0 -2.0144450242618937e-02
GC_10_956 b_10 NI_10 NS_956 0 -3.0186581043413187e-02
GC_10_957 b_10 NI_10 NS_957 0 1.0530784410771163e-02
GC_10_958 b_10 NI_10 NS_958 0 3.5935816882730343e-03
GC_10_959 b_10 NI_10 NS_959 0 -2.6797859934872013e-02
GC_10_960 b_10 NI_10 NS_960 0 1.1150595320241624e-02
GC_10_961 b_10 NI_10 NS_961 0 -1.4133756529886309e-02
GC_10_962 b_10 NI_10 NS_962 0 -2.5194134591562012e-03
GC_10_963 b_10 NI_10 NS_963 0 7.5552443433922010e-03
GC_10_964 b_10 NI_10 NS_964 0 1.5924065838335123e-03
GC_10_965 b_10 NI_10 NS_965 0 -8.5551318004766538e-04
GC_10_966 b_10 NI_10 NS_966 0 2.4403181360446780e-02
GC_10_967 b_10 NI_10 NS_967 0 -7.6201522462998397e-03
GC_10_968 b_10 NI_10 NS_968 0 2.8214368606402503e-04
GC_10_969 b_10 NI_10 NS_969 0 -5.5977717561078331e-04
GC_10_970 b_10 NI_10 NS_970 0 -5.5368502880339511e-03
GC_10_971 b_10 NI_10 NS_971 0 8.2660089980678420e-03
GC_10_972 b_10 NI_10 NS_972 0 7.0201620426320437e-03
GC_10_973 b_10 NI_10 NS_973 0 -7.1913804290868368e-04
GC_10_974 b_10 NI_10 NS_974 0 1.2092544993009798e-02
GC_10_975 b_10 NI_10 NS_975 0 -5.1474185382068827e-03
GC_10_976 b_10 NI_10 NS_976 0 -1.3696932930463182e-04
GC_10_977 b_10 NI_10 NS_977 0 -1.8303692749879715e-03
GC_10_978 b_10 NI_10 NS_978 0 -5.1700319873287989e-03
GC_10_979 b_10 NI_10 NS_979 0 9.2878948173655100e-03
GC_10_980 b_10 NI_10 NS_980 0 5.4154992080077220e-03
GC_10_981 b_10 NI_10 NS_981 0 3.5153075179857407e-03
GC_10_982 b_10 NI_10 NS_982 0 1.1689889648684141e-02
GC_10_983 b_10 NI_10 NS_983 0 -6.1370073008033864e-03
GC_10_984 b_10 NI_10 NS_984 0 1.4286793877627947e-03
GC_10_985 b_10 NI_10 NS_985 0 -2.8171633788654903e-03
GC_10_986 b_10 NI_10 NS_986 0 -7.3461618660298949e-03
GC_10_987 b_10 NI_10 NS_987 0 9.9560406663700401e-03
GC_10_988 b_10 NI_10 NS_988 0 3.3689907072541746e-03
GC_10_989 b_10 NI_10 NS_989 0 8.1686220156131605e-03
GC_10_990 b_10 NI_10 NS_990 0 1.0244275070614890e-02
GC_10_991 b_10 NI_10 NS_991 0 -6.9845048311159598e-03
GC_10_992 b_10 NI_10 NS_992 0 2.9356663461760752e-03
GC_10_993 b_10 NI_10 NS_993 0 -5.6335386548206773e-03
GC_10_994 b_10 NI_10 NS_994 0 -8.0963294470990498e-03
GC_10_995 b_10 NI_10 NS_995 0 9.8581972345700188e-03
GC_10_996 b_10 NI_10 NS_996 0 5.4665539307218326e-04
GC_10_997 b_10 NI_10 NS_997 0 -1.0938520808792545e-02
GC_10_998 b_10 NI_10 NS_998 0 1.2298023816752254e-02
GC_10_999 b_10 NI_10 NS_999 0 9.6448262780441472e-03
GC_10_1000 b_10 NI_10 NS_1000 0 5.0354583750261634e-03
GC_10_1001 b_10 NI_10 NS_1001 0 -1.9866265838165424e-05
GC_10_1002 b_10 NI_10 NS_1002 0 3.1663472790160285e-05
GC_10_1003 b_10 NI_10 NS_1003 0 -7.1316359428667854e-03
GC_10_1004 b_10 NI_10 NS_1004 0 4.4780705489146375e-03
GC_10_1005 b_10 NI_10 NS_1005 0 -7.6761534021381958e-03
GC_10_1006 b_10 NI_10 NS_1006 0 -5.3212035142945965e-03
GC_10_1007 b_10 NI_10 NS_1007 0 9.5161505677169352e-03
GC_10_1008 b_10 NI_10 NS_1008 0 -1.7356766760073161e-03
GC_10_1009 b_10 NI_10 NS_1009 0 1.2474723125596766e-02
GC_10_1010 b_10 NI_10 NS_1010 0 -1.4037693413163968e-03
GC_10_1011 b_10 NI_10 NS_1011 0 -5.0717230701993951e-03
GC_10_1012 b_10 NI_10 NS_1012 0 -2.7497986747740929e-03
GC_10_1013 b_10 NI_10 NS_1013 0 -2.2245920941412122e-03
GC_10_1014 b_10 NI_10 NS_1014 0 6.6015817866906957e-03
GC_10_1015 b_10 NI_10 NS_1015 0 8.9572644668998846e-03
GC_10_1016 b_10 NI_10 NS_1016 0 1.3090554101629067e-04
GC_10_1017 b_10 NI_10 NS_1017 0 1.2487384426645529e-02
GC_10_1018 b_10 NI_10 NS_1018 0 1.7799335453745899e-03
GC_10_1019 b_10 NI_10 NS_1019 0 -5.3780370241361380e-03
GC_10_1020 b_10 NI_10 NS_1020 0 4.1549178222469937e-03
GC_10_1021 b_10 NI_10 NS_1021 0 -1.8499134658876957e-03
GC_10_1022 b_10 NI_10 NS_1022 0 -5.6869425728524187e-03
GC_10_1023 b_10 NI_10 NS_1023 0 2.0796297442000640e-07
GC_10_1024 b_10 NI_10 NS_1024 0 -2.4555621120735843e-07
GC_10_1025 b_10 NI_10 NS_1025 0 -1.1509978778505771e-05
GC_10_1026 b_10 NI_10 NS_1026 0 1.8244020940655961e-05
GC_10_1027 b_10 NI_10 NS_1027 0 -1.4190176474220327e-02
GC_10_1028 b_10 NI_10 NS_1028 0 1.3879312341883953e-03
GC_10_1029 b_10 NI_10 NS_1029 0 -2.6214184849950144e-07
GC_10_1030 b_10 NI_10 NS_1030 0 -3.7469278865742377e-06
GC_10_1031 b_10 NI_10 NS_1031 0 -2.9950674534530582e-04
GC_10_1032 b_10 NI_10 NS_1032 0 4.7112893106071937e-04
GC_10_1033 b_10 NI_10 NS_1033 0 1.2936046057264467e-03
GC_10_1034 b_10 NI_10 NS_1034 0 5.6342157087486489e-04
GC_10_1035 b_10 NI_10 NS_1035 0 -2.7928160469022955e-03
GC_10_1036 b_10 NI_10 NS_1036 0 -7.1086069176997703e-04
GC_10_1037 b_10 NI_10 NS_1037 0 3.5977253048651960e-03
GC_10_1038 b_10 NI_10 NS_1038 0 2.5454524034536625e-03
GC_10_1039 b_10 NI_10 NS_1039 0 1.1770634223598891e-03
GC_10_1040 b_10 NI_10 NS_1040 0 -4.1367913016189242e-03
GC_10_1041 b_10 NI_10 NS_1041 0 -1.5549027037888023e-03
GC_10_1042 b_10 NI_10 NS_1042 0 2.7530000456524855e-03
GC_10_1043 b_10 NI_10 NS_1043 0 -3.5992331282733571e-04
GC_10_1044 b_10 NI_10 NS_1044 0 -2.1737589242752325e-04
GC_10_1045 b_10 NI_10 NS_1045 0 4.0014065019011681e-03
GC_10_1046 b_10 NI_10 NS_1046 0 2.5737097308923726e-04
GC_10_1047 b_10 NI_10 NS_1047 0 -7.3983847206900953e-03
GC_10_1048 b_10 NI_10 NS_1048 0 -1.3542082509393908e-02
GC_10_1049 b_10 NI_10 NS_1049 0 4.4843114449712078e-03
GC_10_1050 b_10 NI_10 NS_1050 0 1.3402112655176941e-02
GC_10_1051 b_10 NI_10 NS_1051 0 6.7170369768755501e-03
GC_10_1052 b_10 NI_10 NS_1052 0 -4.0292270424359782e-03
GC_10_1053 b_10 NI_10 NS_1053 0 -1.3321389325134499e-02
GC_10_1054 b_10 NI_10 NS_1054 0 6.8614134659406424e-04
GC_10_1055 b_10 NI_10 NS_1055 0 7.8581326391374585e-03
GC_10_1056 b_10 NI_10 NS_1056 0 1.8345297311059361e-03
GC_10_1057 b_10 NI_10 NS_1057 0 1.0514012606219340e-02
GC_10_1058 b_10 NI_10 NS_1058 0 -1.9642833995147563e-02
GC_10_1059 b_10 NI_10 NS_1059 0 -1.7746430659648205e-02
GC_10_1060 b_10 NI_10 NS_1060 0 1.9129850712236548e-02
GC_10_1061 b_10 NI_10 NS_1061 0 7.6846929972949757e-03
GC_10_1062 b_10 NI_10 NS_1062 0 -1.4647961343409329e-03
GC_10_1063 b_10 NI_10 NS_1063 0 -1.5663695356293233e-02
GC_10_1064 b_10 NI_10 NS_1064 0 -4.7646585392253594e-03
GC_10_1065 b_10 NI_10 NS_1065 0 8.0859975997443455e-03
GC_10_1066 b_10 NI_10 NS_1066 0 7.2458392344718781e-03
GC_10_1067 b_10 NI_10 NS_1067 0 8.1137527442078691e-03
GC_10_1068 b_10 NI_10 NS_1068 0 -6.0473592427638199e-03
GC_10_1069 b_10 NI_10 NS_1069 0 -1.3987009841274784e-02
GC_10_1070 b_10 NI_10 NS_1070 0 4.5767044118322671e-03
GC_10_1071 b_10 NI_10 NS_1071 0 6.2436878133995790e-03
GC_10_1072 b_10 NI_10 NS_1072 0 2.3779886766409743e-03
GC_10_1073 b_10 NI_10 NS_1073 0 -6.3098266680039197e-03
GC_10_1074 b_10 NI_10 NS_1074 0 -1.1127813894251493e-02
GC_10_1075 b_10 NI_10 NS_1075 0 2.1503507497223641e-03
GC_10_1076 b_10 NI_10 NS_1076 0 1.1938066038685687e-02
GC_10_1077 b_10 NI_10 NS_1077 0 4.2146509118333739e-03
GC_10_1078 b_10 NI_10 NS_1078 0 -1.1800115880068387e-03
GC_10_1079 b_10 NI_10 NS_1079 0 -4.9267465127444563e-03
GC_10_1080 b_10 NI_10 NS_1080 0 1.0434789746052628e-03
GC_10_1081 b_10 NI_10 NS_1081 0 3.0295918234723943e-03
GC_10_1082 b_10 NI_10 NS_1082 0 6.8509421433378328e-04
GC_10_1083 b_10 NI_10 NS_1083 0 -2.2185442028706368e-03
GC_10_1084 b_10 NI_10 NS_1084 0 4.8987925557821747e-04
GC_10_1085 b_10 NI_10 NS_1085 0 3.0814366936518360e-03
GC_10_1086 b_10 NI_10 NS_1086 0 2.2937712263661645e-03
GC_10_1087 b_10 NI_10 NS_1087 0 -1.5261903156397979e-03
GC_10_1088 b_10 NI_10 NS_1088 0 -6.8311090771520889e-04
GC_10_1089 b_10 NI_10 NS_1089 0 1.8943367520306814e-03
GC_10_1090 b_10 NI_10 NS_1090 0 6.7631629385907536e-04
GC_10_1091 b_10 NI_10 NS_1091 0 -1.5560125360775550e-03
GC_10_1092 b_10 NI_10 NS_1092 0 1.2187771813996424e-03
GC_10_1093 b_10 NI_10 NS_1093 0 3.9927828059973100e-03
GC_10_1094 b_10 NI_10 NS_1094 0 1.4034832744531302e-03
GC_10_1095 b_10 NI_10 NS_1095 0 -1.5356518598079699e-03
GC_10_1096 b_10 NI_10 NS_1096 0 5.9546630886372070e-05
GC_10_1097 b_10 NI_10 NS_1097 0 2.8410943534169404e-03
GC_10_1098 b_10 NI_10 NS_1098 0 -6.9178251938379883e-04
GC_10_1099 b_10 NI_10 NS_1099 0 -1.8626304934026411e-03
GC_10_1100 b_10 NI_10 NS_1100 0 1.9986019937544021e-03
GC_10_1101 b_10 NI_10 NS_1101 0 4.9308339550326223e-03
GC_10_1102 b_10 NI_10 NS_1102 0 -1.7294296437359708e-04
GC_10_1103 b_10 NI_10 NS_1103 0 -1.6210911036999205e-03
GC_10_1104 b_10 NI_10 NS_1104 0 9.0628766643911709e-04
GC_10_1105 b_10 NI_10 NS_1105 0 3.0921542848554710e-03
GC_10_1106 b_10 NI_10 NS_1106 0 -2.8475023084105675e-03
GC_10_1107 b_10 NI_10 NS_1107 0 -1.4246678020761543e-03
GC_10_1108 b_10 NI_10 NS_1108 0 3.1958012338328770e-03
GC_10_1109 b_10 NI_10 NS_1109 0 3.8550219538698600e-03
GC_10_1110 b_10 NI_10 NS_1110 0 -2.9522299049154670e-03
GC_10_1111 b_10 NI_10 NS_1111 0 -2.0071714227440779e-03
GC_10_1112 b_10 NI_10 NS_1112 0 -4.1861199999256834e-03
GC_10_1113 b_10 NI_10 NS_1113 0 -3.5103813546213676e-04
GC_10_1114 b_10 NI_10 NS_1114 0 2.2864621988934347e-03
GC_10_1115 b_10 NI_10 NS_1115 0 -1.0763404492238676e-05
GC_10_1116 b_10 NI_10 NS_1116 0 -2.3358512623060993e-05
GC_10_1117 b_10 NI_10 NS_1117 0 8.7769872406692089e-04
GC_10_1118 b_10 NI_10 NS_1118 0 -3.8352110073319014e-03
GC_10_1119 b_10 NI_10 NS_1119 0 3.5234250998337233e-04
GC_10_1120 b_10 NI_10 NS_1120 0 3.3067871907586396e-03
GC_10_1121 b_10 NI_10 NS_1121 0 1.3988574453202541e-03
GC_10_1122 b_10 NI_10 NS_1122 0 -2.3422177521932562e-03
GC_10_1123 b_10 NI_10 NS_1123 0 2.2595473446642656e-03
GC_10_1124 b_10 NI_10 NS_1124 0 3.3689502297281015e-03
GC_10_1125 b_10 NI_10 NS_1125 0 1.1614261634610734e-03
GC_10_1126 b_10 NI_10 NS_1126 0 2.4048209520131343e-03
GC_10_1127 b_10 NI_10 NS_1127 0 -8.2758772881499833e-04
GC_10_1128 b_10 NI_10 NS_1128 0 -1.9684509236745596e-03
GC_10_1129 b_10 NI_10 NS_1129 0 3.9845160819691142e-04
GC_10_1130 b_10 NI_10 NS_1130 0 -2.6910251894535276e-03
GC_10_1131 b_10 NI_10 NS_1131 0 9.7822682465456513e-04
GC_10_1132 b_10 NI_10 NS_1132 0 2.7413561725082268e-03
GC_10_1133 b_10 NI_10 NS_1133 0 1.0427102867670752e-03
GC_10_1134 b_10 NI_10 NS_1134 0 -2.4233095739193480e-03
GC_10_1135 b_10 NI_10 NS_1135 0 -1.0796390318190917e-03
GC_10_1136 b_10 NI_10 NS_1136 0 1.5897876532714650e-03
GC_10_1137 b_10 NI_10 NS_1137 0 -1.0823809464565049e-08
GC_10_1138 b_10 NI_10 NS_1138 0 -2.6612215031558517e-09
GC_10_1139 b_10 NI_10 NS_1139 0 2.3026014584191993e-06
GC_10_1140 b_10 NI_10 NS_1140 0 5.5056631416549071e-07
GC_10_1141 b_10 NI_10 NS_1141 0 2.9495811742531273e-03
GC_10_1142 b_10 NI_10 NS_1142 0 -6.1234115645140367e-04
GC_10_1143 b_10 NI_10 NS_1143 0 2.7950026892218843e-08
GC_10_1144 b_10 NI_10 NS_1144 0 -3.1703309089459317e-08
GC_10_1145 b_10 NI_10 NS_1145 0 2.0347268045948325e-04
GC_10_1146 b_10 NI_10 NS_1146 0 1.3799475864180493e-04
GC_10_1147 b_10 NI_10 NS_1147 0 5.6259278798346417e-04
GC_10_1148 b_10 NI_10 NS_1148 0 2.6570821007289828e-04
GC_10_1149 b_10 NI_10 NS_1149 0 3.1064663771861300e-03
GC_10_1150 b_10 NI_10 NS_1150 0 -2.2048923437347451e-03
GC_10_1151 b_10 NI_10 NS_1151 0 -1.5822544766565816e-03
GC_10_1152 b_10 NI_10 NS_1152 0 -2.6870781070182548e-03
GC_10_1153 b_10 NI_10 NS_1153 0 -2.0496561640580930e-03
GC_10_1154 b_10 NI_10 NS_1154 0 -3.7885098604893363e-03
GC_10_1155 b_10 NI_10 NS_1155 0 -4.9745616994666866e-03
GC_10_1156 b_10 NI_10 NS_1156 0 -1.5415300131158059e-03
GC_10_1157 b_10 NI_10 NS_1157 0 2.9290591200195544e-04
GC_10_1158 b_10 NI_10 NS_1158 0 1.9565149288311562e-04
GC_10_1159 b_10 NI_10 NS_1159 0 -2.8663291160091497e-03
GC_10_1160 b_10 NI_10 NS_1160 0 -9.5746315550123470e-04
GC_10_1161 b_10 NI_10 NS_1161 0 -2.2151872817684864e-02
GC_10_1162 b_10 NI_10 NS_1162 0 -1.0226311643604316e-02
GC_10_1163 b_10 NI_10 NS_1163 0 1.1325012384533458e-03
GC_10_1164 b_10 NI_10 NS_1164 0 2.0395319979965042e-02
GC_10_1165 b_10 NI_10 NS_1165 0 -5.8416198939845506e-03
GC_10_1166 b_10 NI_10 NS_1166 0 4.6116305228382131e-03
GC_10_1167 b_10 NI_10 NS_1167 0 5.7171588901381767e-03
GC_10_1168 b_10 NI_10 NS_1168 0 3.4516068684395697e-02
GC_10_1169 b_10 NI_10 NS_1169 0 8.0342767433485198e-03
GC_10_1170 b_10 NI_10 NS_1170 0 2.7930216040076544e-03
GC_10_1171 b_10 NI_10 NS_1171 0 -7.7724132588519561e-03
GC_10_1172 b_10 NI_10 NS_1172 0 2.9556755330065354e-02
GC_10_1173 b_10 NI_10 NS_1173 0 5.0768422614382636e-02
GC_10_1174 b_10 NI_10 NS_1174 0 -2.0072973638957270e-02
GC_10_1175 b_10 NI_10 NS_1175 0 7.9195777574569935e-03
GC_10_1176 b_10 NI_10 NS_1176 0 -1.6364431161031603e-03
GC_10_1177 b_10 NI_10 NS_1177 0 2.9084851984565549e-02
GC_10_1178 b_10 NI_10 NS_1178 0 -2.6464742845081272e-02
GC_10_1179 b_10 NI_10 NS_1179 0 -6.7250699733901994e-03
GC_10_1180 b_10 NI_10 NS_1180 0 -9.8822034204616126e-03
GC_10_1181 b_10 NI_10 NS_1181 0 8.4630802992075559e-03
GC_10_1182 b_10 NI_10 NS_1182 0 -8.0277999869234305e-03
GC_10_1183 b_10 NI_10 NS_1183 0 -1.8994958082058745e-02
GC_10_1184 b_10 NI_10 NS_1184 0 -2.5238416401572646e-02
GC_10_1185 b_10 NI_10 NS_1185 0 -5.4717856762337824e-03
GC_10_1186 b_10 NI_10 NS_1186 0 -2.8547826260396044e-03
GC_10_1187 b_10 NI_10 NS_1187 0 -1.7741076974559841e-02
GC_10_1188 b_10 NI_10 NS_1188 0 -1.3132225703051047e-02
GC_10_1189 b_10 NI_10 NS_1189 0 -4.8177974099876345e-03
GC_10_1190 b_10 NI_10 NS_1190 0 1.2541405033607783e-02
GC_10_1191 b_10 NI_10 NS_1191 0 -3.4590897686922421e-03
GC_10_1192 b_10 NI_10 NS_1192 0 1.5412389401679772e-03
GC_10_1193 b_10 NI_10 NS_1193 0 -7.1865040470905526e-04
GC_10_1194 b_10 NI_10 NS_1194 0 7.0058608634819665e-03
GC_10_1195 b_10 NI_10 NS_1195 0 1.8820413105141956e-03
GC_10_1196 b_10 NI_10 NS_1196 0 8.5748332613687725e-05
GC_10_1197 b_10 NI_10 NS_1197 0 3.1400233418790052e-04
GC_10_1198 b_10 NI_10 NS_1198 0 -1.9467013334576585e-03
GC_10_1199 b_10 NI_10 NS_1199 0 -1.8563359968445899e-03
GC_10_1200 b_10 NI_10 NS_1200 0 -1.6182084461863887e-03
GC_10_1201 b_10 NI_10 NS_1201 0 -2.1290963464937352e-03
GC_10_1202 b_10 NI_10 NS_1202 0 1.6850444056223900e-03
GC_10_1203 b_10 NI_10 NS_1203 0 7.6361045253130135e-04
GC_10_1204 b_10 NI_10 NS_1204 0 1.8527551194215308e-04
GC_10_1205 b_10 NI_10 NS_1205 0 -6.9730355788848349e-04
GC_10_1206 b_10 NI_10 NS_1206 0 -1.6780696732776939e-03
GC_10_1207 b_10 NI_10 NS_1207 0 -2.6815284286397347e-03
GC_10_1208 b_10 NI_10 NS_1208 0 -8.2749066456769011e-04
GC_10_1209 b_10 NI_10 NS_1209 0 -4.9989599398789729e-04
GC_10_1210 b_10 NI_10 NS_1210 0 2.9288646880063539e-03
GC_10_1211 b_10 NI_10 NS_1211 0 1.3533577628722939e-03
GC_10_1212 b_10 NI_10 NS_1212 0 -8.5805585573830556e-04
GC_10_1213 b_10 NI_10 NS_1213 0 -2.4189246512610952e-03
GC_10_1214 b_10 NI_10 NS_1214 0 -2.2676208469955303e-03
GC_10_1215 b_10 NI_10 NS_1215 0 -3.5540457750803177e-03
GC_10_1216 b_10 NI_10 NS_1216 0 7.4852698690677788e-04
GC_10_1217 b_10 NI_10 NS_1217 0 2.4633831864147048e-03
GC_10_1218 b_10 NI_10 NS_1218 0 3.0182806570870310e-03
GC_10_1219 b_10 NI_10 NS_1219 0 9.8455404187781231e-04
GC_10_1220 b_10 NI_10 NS_1220 0 -2.9418095402951269e-03
GC_10_1221 b_10 NI_10 NS_1221 0 -4.7677995762038534e-03
GC_10_1222 b_10 NI_10 NS_1222 0 5.4340723728901622e-05
GC_10_1223 b_10 NI_10 NS_1223 0 -1.7083701070289704e-03
GC_10_1224 b_10 NI_10 NS_1224 0 3.7124272466180033e-03
GC_10_1225 b_10 NI_10 NS_1225 0 -7.6587239284450282e-04
GC_10_1226 b_10 NI_10 NS_1226 0 1.5006822167187904e-03
GC_10_1227 b_10 NI_10 NS_1227 0 3.2213016471490754e-03
GC_10_1228 b_10 NI_10 NS_1228 0 -1.3508686361711482e-03
GC_10_1229 b_10 NI_10 NS_1229 0 -2.9326244145418727e-06
GC_10_1230 b_10 NI_10 NS_1230 0 8.7469676315159365e-06
GC_10_1231 b_10 NI_10 NS_1231 0 -1.8200423201619083e-03
GC_10_1232 b_10 NI_10 NS_1232 0 -2.5277362755914425e-03
GC_10_1233 b_10 NI_10 NS_1233 0 -2.4072536483496806e-03
GC_10_1234 b_10 NI_10 NS_1234 0 2.4886640637733133e-03
GC_10_1235 b_10 NI_10 NS_1235 0 1.0142609867773501e-03
GC_10_1236 b_10 NI_10 NS_1236 0 2.4256812370204088e-03
GC_10_1237 b_10 NI_10 NS_1237 0 8.5775821240963472e-04
GC_10_1238 b_10 NI_10 NS_1238 0 -2.6994845899480785e-03
GC_10_1239 b_10 NI_10 NS_1239 0 -3.0644790150903631e-04
GC_10_1240 b_10 NI_10 NS_1240 0 1.6741355472200657e-03
GC_10_1241 b_10 NI_10 NS_1241 0 -1.7840541426726918e-03
GC_10_1242 b_10 NI_10 NS_1242 0 -3.1181108409156390e-04
GC_10_1243 b_10 NI_10 NS_1243 0 1.4004540369821888e-03
GC_10_1244 b_10 NI_10 NS_1244 0 1.9709615356371655e-03
GC_10_1245 b_10 NI_10 NS_1245 0 1.0449287331449361e-03
GC_10_1246 b_10 NI_10 NS_1246 0 -2.2998046401287316e-03
GC_10_1247 b_10 NI_10 NS_1247 0 -6.9799493589196328e-04
GC_10_1248 b_10 NI_10 NS_1248 0 -1.4668898763355238e-03
GC_10_1249 b_10 NI_10 NS_1249 0 -1.3735490954940638e-03
GC_10_1250 b_10 NI_10 NS_1250 0 -3.1252859547377290e-04
GC_10_1251 b_10 NI_10 NS_1251 0 7.1030487328272083e-09
GC_10_1252 b_10 NI_10 NS_1252 0 -2.4709966348712714e-08
GC_10_1253 b_10 NI_10 NS_1253 0 -4.5275596766090129e-07
GC_10_1254 b_10 NI_10 NS_1254 0 1.6341837978301841e-06
GC_10_1255 b_10 NI_10 NS_1255 0 7.7624118558382582e-03
GC_10_1256 b_10 NI_10 NS_1256 0 -1.6012430130799111e-03
GC_10_1257 b_10 NI_10 NS_1257 0 -1.2108955808884595e-08
GC_10_1258 b_10 NI_10 NS_1258 0 -8.8417701864810631e-07
GC_10_1259 b_10 NI_10 NS_1259 0 1.0417949015734674e-04
GC_10_1260 b_10 NI_10 NS_1260 0 -5.1169960681443009e-04
GC_10_1261 b_10 NI_10 NS_1261 0 -1.9362876174674781e-03
GC_10_1262 b_10 NI_10 NS_1262 0 -5.9765058655085912e-04
GC_10_1263 b_10 NI_10 NS_1263 0 2.9418170709409521e-03
GC_10_1264 b_10 NI_10 NS_1264 0 2.2635987277035800e-03
GC_10_1265 b_10 NI_10 NS_1265 0 -3.5704321000968845e-03
GC_10_1266 b_10 NI_10 NS_1266 0 -3.0490699932925348e-03
GC_10_1267 b_10 NI_10 NS_1267 0 -1.7073690282817197e-03
GC_10_1268 b_10 NI_10 NS_1268 0 5.8427804732026434e-03
GC_10_1269 b_10 NI_10 NS_1269 0 4.3666880349392465e-03
GC_10_1270 b_10 NI_10 NS_1270 0 -2.4751072749372950e-03
GC_10_1271 b_10 NI_10 NS_1271 0 -1.1000736114668372e-04
GC_10_1272 b_10 NI_10 NS_1272 0 -1.0334111022581018e-04
GC_10_1273 b_10 NI_10 NS_1273 0 -4.4523080010265394e-03
GC_10_1274 b_10 NI_10 NS_1274 0 -9.2440216644957781e-04
GC_10_1275 b_10 NI_10 NS_1275 0 9.1241451991947286e-03
GC_10_1276 b_10 NI_10 NS_1276 0 1.7784743700107655e-02
GC_10_1277 b_10 NI_10 NS_1277 0 -4.0272952724853513e-03
GC_10_1278 b_10 NI_10 NS_1278 0 -1.7846764115834898e-02
GC_10_1279 b_10 NI_10 NS_1279 0 -8.2177715159456339e-03
GC_10_1280 b_10 NI_10 NS_1280 0 4.1736031904648580e-03
GC_10_1281 b_10 NI_10 NS_1281 0 1.7063488480834652e-02
GC_10_1282 b_10 NI_10 NS_1282 0 -4.3909755959806916e-04
GC_10_1283 b_10 NI_10 NS_1283 0 -9.2787149378705698e-03
GC_10_1284 b_10 NI_10 NS_1284 0 -3.2069945232172932e-03
GC_10_1285 b_10 NI_10 NS_1285 0 -1.3713354902277505e-02
GC_10_1286 b_10 NI_10 NS_1286 0 2.2836241728451129e-02
GC_10_1287 b_10 NI_10 NS_1287 0 2.2839545856672493e-02
GC_10_1288 b_10 NI_10 NS_1288 0 -2.2669178990011935e-02
GC_10_1289 b_10 NI_10 NS_1289 0 -9.2392853390804754e-03
GC_10_1290 b_10 NI_10 NS_1290 0 9.0811412226233547e-04
GC_10_1291 b_10 NI_10 NS_1291 0 1.8480129598970878e-02
GC_10_1292 b_10 NI_10 NS_1292 0 6.2442194291569145e-03
GC_10_1293 b_10 NI_10 NS_1293 0 -9.1760825917089842e-03
GC_10_1294 b_10 NI_10 NS_1294 0 -9.4609771756993481e-03
GC_10_1295 b_10 NI_10 NS_1295 0 -9.9743257214595770e-03
GC_10_1296 b_10 NI_10 NS_1296 0 6.3961893660862976e-03
GC_10_1297 b_10 NI_10 NS_1297 0 1.6838478148080139e-02
GC_10_1298 b_10 NI_10 NS_1298 0 -4.8501226537065291e-03
GC_10_1299 b_10 NI_10 NS_1299 0 -7.2149234000147451e-03
GC_10_1300 b_10 NI_10 NS_1300 0 -3.4092345264253401e-03
GC_10_1301 b_10 NI_10 NS_1301 0 6.8281951752810410e-03
GC_10_1302 b_10 NI_10 NS_1302 0 1.3297050871185209e-02
GC_10_1303 b_10 NI_10 NS_1303 0 -1.8195853055223126e-03
GC_10_1304 b_10 NI_10 NS_1304 0 -1.4401718425428797e-02
GC_10_1305 b_10 NI_10 NS_1305 0 -4.9860075666278234e-03
GC_10_1306 b_10 NI_10 NS_1306 0 1.0394632537667442e-03
GC_10_1307 b_10 NI_10 NS_1307 0 6.0026082178580636e-03
GC_10_1308 b_10 NI_10 NS_1308 0 -1.1030577012290056e-03
GC_10_1309 b_10 NI_10 NS_1309 0 -3.4642738155391023e-03
GC_10_1310 b_10 NI_10 NS_1310 0 -1.0876296808350686e-03
GC_10_1311 b_10 NI_10 NS_1311 0 2.7180506512249842e-03
GC_10_1312 b_10 NI_10 NS_1312 0 -5.0782197071479694e-04
GC_10_1313 b_10 NI_10 NS_1313 0 -3.2964875840286382e-03
GC_10_1314 b_10 NI_10 NS_1314 0 -2.8951322147139822e-03
GC_10_1315 b_10 NI_10 NS_1315 0 2.0159599130026603e-03
GC_10_1316 b_10 NI_10 NS_1316 0 7.7577878023798519e-04
GC_10_1317 b_10 NI_10 NS_1317 0 -2.0162769558034269e-03
GC_10_1318 b_10 NI_10 NS_1318 0 -9.6646490666639669e-04
GC_10_1319 b_10 NI_10 NS_1319 0 2.1216204026185837e-03
GC_10_1320 b_10 NI_10 NS_1320 0 -1.4709119213605578e-03
GC_10_1321 b_10 NI_10 NS_1321 0 -4.1847966358709273e-03
GC_10_1322 b_10 NI_10 NS_1322 0 -1.8129451333208349e-03
GC_10_1323 b_10 NI_10 NS_1323 0 2.3697775066020910e-03
GC_10_1324 b_10 NI_10 NS_1324 0 -3.7075616305296623e-04
GC_10_1325 b_10 NI_10 NS_1325 0 -3.0172236709727763e-03
GC_10_1326 b_10 NI_10 NS_1326 0 4.6233814230720006e-04
GC_10_1327 b_10 NI_10 NS_1327 0 2.7064424611681730e-03
GC_10_1328 b_10 NI_10 NS_1328 0 -2.7282228980239995e-03
GC_10_1329 b_10 NI_10 NS_1329 0 -5.0393302507005869e-03
GC_10_1330 b_10 NI_10 NS_1330 0 -1.2782932411566273e-04
GC_10_1331 b_10 NI_10 NS_1331 0 2.4346766646885809e-03
GC_10_1332 b_10 NI_10 NS_1332 0 -2.1719792852930380e-03
GC_10_1333 b_10 NI_10 NS_1333 0 -3.2449817597156689e-03
GC_10_1334 b_10 NI_10 NS_1334 0 2.6005317677844932e-03
GC_10_1335 b_10 NI_10 NS_1335 0 1.7436666478569435e-03
GC_10_1336 b_10 NI_10 NS_1336 0 -4.7503531473250043e-03
GC_10_1337 b_10 NI_10 NS_1337 0 -3.6339988945856641e-03
GC_10_1338 b_10 NI_10 NS_1338 0 2.5967287839337694e-03
GC_10_1339 b_10 NI_10 NS_1339 0 -2.8319048140421645e-03
GC_10_1340 b_10 NI_10 NS_1340 0 3.9895731634650442e-03
GC_10_1341 b_10 NI_10 NS_1341 0 -2.2141478368044025e-04
GC_10_1342 b_10 NI_10 NS_1342 0 -4.2135113287555120e-03
GC_10_1343 b_10 NI_10 NS_1343 0 -9.8957945628013259e-06
GC_10_1344 b_10 NI_10 NS_1344 0 7.5258087897587903e-06
GC_10_1345 b_10 NI_10 NS_1345 0 -1.3539535487032362e-03
GC_10_1346 b_10 NI_10 NS_1346 0 3.3754883304646017e-03
GC_10_1347 b_10 NI_10 NS_1347 0 -9.6985119084811746e-04
GC_10_1348 b_10 NI_10 NS_1348 0 -4.3479509979951385e-03
GC_10_1349 b_10 NI_10 NS_1349 0 -1.0009112717441013e-03
GC_10_1350 b_10 NI_10 NS_1350 0 2.2213051273753492e-03
GC_10_1351 b_10 NI_10 NS_1351 0 -1.6517283917427648e-03
GC_10_1352 b_10 NI_10 NS_1352 0 -4.4093139762067324e-03
GC_10_1353 b_10 NI_10 NS_1353 0 -1.4483159798036028e-03
GC_10_1354 b_10 NI_10 NS_1354 0 -2.4971456887776704e-03
GC_10_1355 b_10 NI_10 NS_1355 0 7.8219595711522742e-04
GC_10_1356 b_10 NI_10 NS_1356 0 2.5933469659666342e-03
GC_10_1357 b_10 NI_10 NS_1357 0 -6.9628533778962618e-04
GC_10_1358 b_10 NI_10 NS_1358 0 2.8792042523863299e-03
GC_10_1359 b_10 NI_10 NS_1359 0 -1.4353705247931842e-03
GC_10_1360 b_10 NI_10 NS_1360 0 -2.7718613469606048e-03
GC_10_1361 b_10 NI_10 NS_1361 0 -1.1678495830825645e-03
GC_10_1362 b_10 NI_10 NS_1362 0 2.6661995998535910e-03
GC_10_1363 b_10 NI_10 NS_1363 0 7.8075940709442947e-04
GC_10_1364 b_10 NI_10 NS_1364 0 -1.8746154576252442e-03
GC_10_1365 b_10 NI_10 NS_1365 0 2.3789744546651722e-08
GC_10_1366 b_10 NI_10 NS_1366 0 -6.0253429559730513e-08
GC_10_1367 b_10 NI_10 NS_1367 0 -9.0373524595306165e-07
GC_10_1368 b_10 NI_10 NS_1368 0 3.2031377343762641e-06
GD_10_1 b_10 NI_10 NA_1 0 5.6280346764792760e-06
GD_10_2 b_10 NI_10 NA_2 0 -1.8680220013075213e-06
GD_10_3 b_10 NI_10 NA_3 0 4.7457956852591431e-07
GD_10_4 b_10 NI_10 NA_4 0 -5.5534207809670377e-06
GD_10_5 b_10 NI_10 NA_5 0 1.2382044181522569e-06
GD_10_6 b_10 NI_10 NA_6 0 4.8704198361389570e-06
GD_10_7 b_10 NI_10 NA_7 0 2.6580138883612736e-05
GD_10_8 b_10 NI_10 NA_8 0 1.0377477843714573e-04
GD_10_9 b_10 NI_10 NA_9 0 -4.2441668755691490e-03
GD_10_10 b_10 NI_10 NA_10 0 -8.6867573911805149e-03
GD_10_11 b_10 NI_10 NA_11 0 5.9084121393460738e-04
GD_10_12 b_10 NI_10 NA_12 0 1.3004900789018288e-02
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 5.5755236666141958e-06
GC_11_2 b_11 NI_11 NS_2 0 -6.0660004250714066e-08
GC_11_3 b_11 NI_11 NS_3 0 -3.1618489752449203e-11
GC_11_4 b_11 NI_11 NS_4 0 4.1807631323172803e-10
GC_11_5 b_11 NI_11 NS_5 0 8.6995339194311467e-08
GC_11_6 b_11 NI_11 NS_6 0 -7.3605823320682992e-08
GC_11_7 b_11 NI_11 NS_7 0 3.8660601318163010e-09
GC_11_8 b_11 NI_11 NS_8 0 8.3840027522250360e-08
GC_11_9 b_11 NI_11 NS_9 0 6.3124920217853004e-07
GC_11_10 b_11 NI_11 NS_10 0 -8.3236115365640159e-07
GC_11_11 b_11 NI_11 NS_11 0 -9.1896949991296092e-07
GC_11_12 b_11 NI_11 NS_12 0 7.4767398205034276e-08
GC_11_13 b_11 NI_11 NS_13 0 5.4102904789133648e-07
GC_11_14 b_11 NI_11 NS_14 0 4.6009314449325679e-08
GC_11_15 b_11 NI_11 NS_15 0 -1.3827631087527056e-06
GC_11_16 b_11 NI_11 NS_16 0 -9.7963480835588509e-07
GC_11_17 b_11 NI_11 NS_17 0 3.0638171743443738e-07
GC_11_18 b_11 NI_11 NS_18 0 2.0537906257599618e-07
GC_11_19 b_11 NI_11 NS_19 0 -5.6258819251759194e-07
GC_11_20 b_11 NI_11 NS_20 0 7.1028206322094044e-07
GC_11_21 b_11 NI_11 NS_21 0 1.9977094806604460e-06
GC_11_22 b_11 NI_11 NS_22 0 -6.2823241848958011e-07
GC_11_23 b_11 NI_11 NS_23 0 -2.6418324854900423e-06
GC_11_24 b_11 NI_11 NS_24 0 3.8227289346353810e-07
GC_11_25 b_11 NI_11 NS_25 0 4.1279235555666214e-08
GC_11_26 b_11 NI_11 NS_26 0 1.4294009862038351e-06
GC_11_27 b_11 NI_11 NS_27 0 2.3354979947511601e-07
GC_11_28 b_11 NI_11 NS_28 0 -1.8328019763605085e-06
GC_11_29 b_11 NI_11 NS_29 0 -8.6530551514861955e-07
GC_11_30 b_11 NI_11 NS_30 0 1.3761334376667921e-06
GC_11_31 b_11 NI_11 NS_31 0 2.2852343485517291e-06
GC_11_32 b_11 NI_11 NS_32 0 2.9655735293204102e-06
GC_11_33 b_11 NI_11 NS_33 0 -2.0507621167849545e-06
GC_11_34 b_11 NI_11 NS_34 0 -3.4924530935456853e-06
GC_11_35 b_11 NI_11 NS_35 0 -2.8718750781547062e-07
GC_11_36 b_11 NI_11 NS_36 0 1.5382141390845420e-06
GC_11_37 b_11 NI_11 NS_37 0 1.7081593407363720e-06
GC_11_38 b_11 NI_11 NS_38 0 -1.8793185945067098e-06
GC_11_39 b_11 NI_11 NS_39 0 -1.6427720404991461e-06
GC_11_40 b_11 NI_11 NS_40 0 1.0311044607325779e-06
GC_11_41 b_11 NI_11 NS_41 0 4.2910642968010851e-07
GC_11_42 b_11 NI_11 NS_42 0 1.8543444486597642e-06
GC_11_43 b_11 NI_11 NS_43 0 2.5925851909270456e-07
GC_11_44 b_11 NI_11 NS_44 0 -2.2599443668814207e-06
GC_11_45 b_11 NI_11 NS_45 0 -7.4200630585986862e-07
GC_11_46 b_11 NI_11 NS_46 0 9.6144879355062762e-07
GC_11_47 b_11 NI_11 NS_47 0 2.0833940943737946e-06
GC_11_48 b_11 NI_11 NS_48 0 -1.8914137986180384e-08
GC_11_49 b_11 NI_11 NS_49 0 -1.8132847794760759e-06
GC_11_50 b_11 NI_11 NS_50 0 -3.2980288223464446e-07
GC_11_51 b_11 NI_11 NS_51 0 -9.5351397519391526e-08
GC_11_52 b_11 NI_11 NS_52 0 7.6456718315705571e-07
GC_11_53 b_11 NI_11 NS_53 0 2.1964047094442798e-07
GC_11_54 b_11 NI_11 NS_54 0 -5.5288916743159263e-07
GC_11_55 b_11 NI_11 NS_55 0 -2.4027541354216717e-07
GC_11_56 b_11 NI_11 NS_56 0 4.2924000391220568e-07
GC_11_57 b_11 NI_11 NS_57 0 1.0687575450697487e-07
GC_11_58 b_11 NI_11 NS_58 0 -2.2411989275836596e-07
GC_11_59 b_11 NI_11 NS_59 0 -4.5513574740349919e-07
GC_11_60 b_11 NI_11 NS_60 0 3.0524960920782961e-07
GC_11_61 b_11 NI_11 NS_61 0 2.0652137026861765e-07
GC_11_62 b_11 NI_11 NS_62 0 1.6753684212852121e-08
GC_11_63 b_11 NI_11 NS_63 0 -1.4742331963584045e-07
GC_11_64 b_11 NI_11 NS_64 0 1.9350230652539337e-07
GC_11_65 b_11 NI_11 NS_65 0 2.4903153443082525e-08
GC_11_66 b_11 NI_11 NS_66 0 -1.4137794883297758e-07
GC_11_67 b_11 NI_11 NS_67 0 -3.4514289280496584e-07
GC_11_68 b_11 NI_11 NS_68 0 2.7931881165258628e-07
GC_11_69 b_11 NI_11 NS_69 0 1.1043781787671364e-07
GC_11_70 b_11 NI_11 NS_70 0 -2.3194401318501036e-08
GC_11_71 b_11 NI_11 NS_71 0 -1.1145130132379048e-07
GC_11_72 b_11 NI_11 NS_72 0 2.2574263131585403e-07
GC_11_73 b_11 NI_11 NS_73 0 -1.8935033865007169e-08
GC_11_74 b_11 NI_11 NS_74 0 -1.6882348365593798e-07
GC_11_75 b_11 NI_11 NS_75 0 -2.8639914622843239e-07
GC_11_76 b_11 NI_11 NS_76 0 1.8674281449061859e-07
GC_11_77 b_11 NI_11 NS_77 0 -1.1162243171570951e-07
GC_11_78 b_11 NI_11 NS_78 0 -5.9977771353852103e-08
GC_11_79 b_11 NI_11 NS_79 0 -1.7478653594344419e-07
GC_11_80 b_11 NI_11 NS_80 0 2.0344673648025456e-07
GC_11_81 b_11 NI_11 NS_81 0 -2.9228577563658386e-07
GC_11_82 b_11 NI_11 NS_82 0 -3.9974371571890977e-08
GC_11_83 b_11 NI_11 NS_83 0 -4.9673877236028460e-07
GC_11_84 b_11 NI_11 NS_84 0 5.7782713366873832e-08
GC_11_85 b_11 NI_11 NS_85 0 2.7716620970686399e-06
GC_11_86 b_11 NI_11 NS_86 0 4.3274910284927486e-07
GC_11_87 b_11 NI_11 NS_87 0 -3.2405411759649701e-07
GC_11_88 b_11 NI_11 NS_88 0 6.7628408041162407e-07
GC_11_89 b_11 NI_11 NS_89 0 1.2397621043474626e-08
GC_11_90 b_11 NI_11 NS_90 0 1.2810073349475503e-08
GC_11_91 b_11 NI_11 NS_91 0 -6.7252784729564591e-09
GC_11_92 b_11 NI_11 NS_92 0 4.6490261709748042e-07
GC_11_93 b_11 NI_11 NS_93 0 -1.2602623324804433e-07
GC_11_94 b_11 NI_11 NS_94 0 2.6648530367178724e-07
GC_11_95 b_11 NI_11 NS_95 0 -4.8106096751822948e-07
GC_11_96 b_11 NI_11 NS_96 0 9.8571716156935796e-08
GC_11_97 b_11 NI_11 NS_97 0 -9.4580716854553927e-07
GC_11_98 b_11 NI_11 NS_98 0 4.8604612082697954e-07
GC_11_99 b_11 NI_11 NS_99 0 -1.8710926592817507e-07
GC_11_100 b_11 NI_11 NS_100 0 -7.9276776252217464e-08
GC_11_101 b_11 NI_11 NS_101 0 1.6398871949711904e-08
GC_11_102 b_11 NI_11 NS_102 0 -1.4792141897853921e-07
GC_11_103 b_11 NI_11 NS_103 0 8.6143299412193223e-08
GC_11_104 b_11 NI_11 NS_104 0 1.0231044803711723e-07
GC_11_105 b_11 NI_11 NS_105 0 -1.1792080781972772e-07
GC_11_106 b_11 NI_11 NS_106 0 -1.5795712522898897e-07
GC_11_107 b_11 NI_11 NS_107 0 -7.0287862343113647e-08
GC_11_108 b_11 NI_11 NS_108 0 8.1119501789227969e-08
GC_11_109 b_11 NI_11 NS_109 0 -4.4653819236226497e-10
GC_11_110 b_11 NI_11 NS_110 0 -3.7628552539837902e-08
GC_11_111 b_11 NI_11 NS_111 0 -8.0395437914484086e-12
GC_11_112 b_11 NI_11 NS_112 0 7.1577823988983396e-12
GC_11_113 b_11 NI_11 NS_113 0 9.6678245989145203e-10
GC_11_114 b_11 NI_11 NS_114 0 -3.3560587245374733e-10
GC_11_115 b_11 NI_11 NS_115 0 -1.2624809307115051e-05
GC_11_116 b_11 NI_11 NS_116 0 1.6614662640935741e-08
GC_11_117 b_11 NI_11 NS_117 0 2.1156928083993149e-11
GC_11_118 b_11 NI_11 NS_118 0 -3.0722865469899574e-10
GC_11_119 b_11 NI_11 NS_119 0 -3.4980953676618041e-07
GC_11_120 b_11 NI_11 NS_120 0 -9.9927141669836975e-07
GC_11_121 b_11 NI_11 NS_121 0 -9.3440256998009971e-07
GC_11_122 b_11 NI_11 NS_122 0 1.7812972225185147e-06
GC_11_123 b_11 NI_11 NS_123 0 -3.3145737109136827e-06
GC_11_124 b_11 NI_11 NS_124 0 8.1232076302461920e-07
GC_11_125 b_11 NI_11 NS_125 0 9.4647105633553833e-07
GC_11_126 b_11 NI_11 NS_126 0 -2.3710044844775857e-07
GC_11_127 b_11 NI_11 NS_127 0 5.4136939106297060e-07
GC_11_128 b_11 NI_11 NS_128 0 4.5112155285682987e-06
GC_11_129 b_11 NI_11 NS_129 0 1.6155090724882848e-06
GC_11_130 b_11 NI_11 NS_130 0 3.0375513412667175e-06
GC_11_131 b_11 NI_11 NS_131 0 -8.7083860710227516e-07
GC_11_132 b_11 NI_11 NS_132 0 -5.9646444503774751e-07
GC_11_133 b_11 NI_11 NS_133 0 4.7061613839263935e-07
GC_11_134 b_11 NI_11 NS_134 0 -1.1586865293525802e-06
GC_11_135 b_11 NI_11 NS_135 0 2.8699786071425417e-06
GC_11_136 b_11 NI_11 NS_136 0 1.0313963508282344e-05
GC_11_137 b_11 NI_11 NS_137 0 4.5228652676375217e-06
GC_11_138 b_11 NI_11 NS_138 0 -7.5298326708627592e-07
GC_11_139 b_11 NI_11 NS_139 0 1.6523558573381327e-06
GC_11_140 b_11 NI_11 NS_140 0 -4.2608453978673586e-07
GC_11_141 b_11 NI_11 NS_141 0 1.6706030169471077e-05
GC_11_142 b_11 NI_11 NS_142 0 -4.4199344819947536e-06
GC_11_143 b_11 NI_11 NS_143 0 2.2368658800246875e-07
GC_11_144 b_11 NI_11 NS_144 0 -1.0416416292728954e-06
GC_11_145 b_11 NI_11 NS_145 0 9.3469258329669422e-06
GC_11_146 b_11 NI_11 NS_146 0 -7.0992745182520472e-07
GC_11_147 b_11 NI_11 NS_147 0 -5.5727596587626390e-06
GC_11_148 b_11 NI_11 NS_148 0 -1.9751248004374708e-05
GC_11_149 b_11 NI_11 NS_149 0 -6.0103023454437466e-07
GC_11_150 b_11 NI_11 NS_150 0 -8.9964460750712303e-07
GC_11_151 b_11 NI_11 NS_151 0 -1.1428657685274264e-05
GC_11_152 b_11 NI_11 NS_152 0 -1.0988294924499851e-05
GC_11_153 b_11 NI_11 NS_153 0 -2.2555833689012247e-06
GC_11_154 b_11 NI_11 NS_154 0 2.5926756429101487e-07
GC_11_155 b_11 NI_11 NS_155 0 -1.9214224334732414e-06
GC_11_156 b_11 NI_11 NS_156 0 -7.8273490281394828e-07
GC_11_157 b_11 NI_11 NS_157 0 -9.6694391284153966e-06
GC_11_158 b_11 NI_11 NS_158 0 5.8238596867244867e-06
GC_11_159 b_11 NI_11 NS_159 0 -3.0070390226804888e-07
GC_11_160 b_11 NI_11 NS_160 0 1.6096110101283435e-07
GC_11_161 b_11 NI_11 NS_161 0 -1.6035952413652707e-06
GC_11_162 b_11 NI_11 NS_162 0 5.7948445508251016e-06
GC_11_163 b_11 NI_11 NS_163 0 2.0456012303100733e-06
GC_11_164 b_11 NI_11 NS_164 0 1.9760432784622389e-06
GC_11_165 b_11 NI_11 NS_165 0 6.0757109983679242e-07
GC_11_166 b_11 NI_11 NS_166 0 -8.9292213599713589e-08
GC_11_167 b_11 NI_11 NS_167 0 3.3238986525765459e-06
GC_11_168 b_11 NI_11 NS_168 0 -4.3020983083018192e-07
GC_11_169 b_11 NI_11 NS_169 0 -5.1720178575616883e-08
GC_11_170 b_11 NI_11 NS_170 0 3.3332486727726133e-08
GC_11_171 b_11 NI_11 NS_171 0 -8.0692562509312688e-07
GC_11_172 b_11 NI_11 NS_172 0 -2.3783621105866186e-07
GC_11_173 b_11 NI_11 NS_173 0 3.8089999386972390e-07
GC_11_174 b_11 NI_11 NS_174 0 -5.1763484438157882e-07
GC_11_175 b_11 NI_11 NS_175 0 1.1838643063863073e-06
GC_11_176 b_11 NI_11 NS_176 0 -3.2905320343163989e-08
GC_11_177 b_11 NI_11 NS_177 0 2.3909301389773830e-08
GC_11_178 b_11 NI_11 NS_178 0 4.9140113678944839e-08
GC_11_179 b_11 NI_11 NS_179 0 -5.6752129035539005e-07
GC_11_180 b_11 NI_11 NS_180 0 -5.4511752949739278e-08
GC_11_181 b_11 NI_11 NS_181 0 4.9423811223595759e-07
GC_11_182 b_11 NI_11 NS_182 0 -5.0922567426342014e-07
GC_11_183 b_11 NI_11 NS_183 0 1.1633700202406792e-06
GC_11_184 b_11 NI_11 NS_184 0 -6.8915236953313537e-07
GC_11_185 b_11 NI_11 NS_185 0 5.6879120469692410e-08
GC_11_186 b_11 NI_11 NS_186 0 -7.6274718122722824e-12
GC_11_187 b_11 NI_11 NS_187 0 -5.7572912950039112e-07
GC_11_188 b_11 NI_11 NS_188 0 -6.5420403244152713e-08
GC_11_189 b_11 NI_11 NS_189 0 6.3198127009596859e-07
GC_11_190 b_11 NI_11 NS_190 0 -5.0017472133900703e-07
GC_11_191 b_11 NI_11 NS_191 0 8.4908883072695976e-07
GC_11_192 b_11 NI_11 NS_192 0 -1.3993597598688759e-06
GC_11_193 b_11 NI_11 NS_193 0 1.0851631658914172e-07
GC_11_194 b_11 NI_11 NS_194 0 -6.0235217519219857e-08
GC_11_195 b_11 NI_11 NS_195 0 -3.9931014177459837e-07
GC_11_196 b_11 NI_11 NS_196 0 -2.0521059208802435e-07
GC_11_197 b_11 NI_11 NS_197 0 1.1352424758494213e-06
GC_11_198 b_11 NI_11 NS_198 0 -8.8090144564375791e-07
GC_11_199 b_11 NI_11 NS_199 0 -4.1524178458292170e-06
GC_11_200 b_11 NI_11 NS_200 0 6.0076205822858946e-07
GC_11_201 b_11 NI_11 NS_201 0 -5.6337357053751464e-07
GC_11_202 b_11 NI_11 NS_202 0 -1.9350600144600659e-06
GC_11_203 b_11 NI_11 NS_203 0 -2.9192734685673568e-08
GC_11_204 b_11 NI_11 NS_204 0 -9.6996378506101586e-09
GC_11_205 b_11 NI_11 NS_205 0 -3.5869181568187895e-07
GC_11_206 b_11 NI_11 NS_206 0 -2.9247742836783107e-07
GC_11_207 b_11 NI_11 NS_207 0 -4.7717814161115129e-07
GC_11_208 b_11 NI_11 NS_208 0 -1.7395804033882855e-07
GC_11_209 b_11 NI_11 NS_209 0 8.5945770614713840e-07
GC_11_210 b_11 NI_11 NS_210 0 -7.5659643131171687e-07
GC_11_211 b_11 NI_11 NS_211 0 6.0934832601820242e-07
GC_11_212 b_11 NI_11 NS_212 0 -1.0778276645711785e-06
GC_11_213 b_11 NI_11 NS_213 0 9.0828652496316249e-08
GC_11_214 b_11 NI_11 NS_214 0 1.4506981264193302e-07
GC_11_215 b_11 NI_11 NS_215 0 1.5780166300889988e-07
GC_11_216 b_11 NI_11 NS_216 0 4.4524675035644386e-07
GC_11_217 b_11 NI_11 NS_217 0 2.3130719170550260e-08
GC_11_218 b_11 NI_11 NS_218 0 -1.6507917224643207e-07
GC_11_219 b_11 NI_11 NS_219 0 -3.7596932109660995e-08
GC_11_220 b_11 NI_11 NS_220 0 -1.2378315342334743e-07
GC_11_221 b_11 NI_11 NS_221 0 -8.6474435815201701e-08
GC_11_222 b_11 NI_11 NS_222 0 1.2324392508960156e-07
GC_11_223 b_11 NI_11 NS_223 0 -9.0131162962698241e-09
GC_11_224 b_11 NI_11 NS_224 0 -3.7918655735831909e-09
GC_11_225 b_11 NI_11 NS_225 0 2.2957005692125217e-12
GC_11_226 b_11 NI_11 NS_226 0 -3.3975213846155314e-12
GC_11_227 b_11 NI_11 NS_227 0 -7.3117549347338839e-10
GC_11_228 b_11 NI_11 NS_228 0 -8.2653557722608890e-11
GC_11_229 b_11 NI_11 NS_229 0 1.3351809288195114e-05
GC_11_230 b_11 NI_11 NS_230 0 -5.9008750923864211e-08
GC_11_231 b_11 NI_11 NS_231 0 -1.4919045099925479e-11
GC_11_232 b_11 NI_11 NS_232 0 1.3565936058984920e-10
GC_11_233 b_11 NI_11 NS_233 0 3.5691508694796307e-07
GC_11_234 b_11 NI_11 NS_234 0 -1.8036855785474590e-07
GC_11_235 b_11 NI_11 NS_235 0 2.7982053503420791e-07
GC_11_236 b_11 NI_11 NS_236 0 -3.4839665083453148e-07
GC_11_237 b_11 NI_11 NS_237 0 4.9688859194333686e-07
GC_11_238 b_11 NI_11 NS_238 0 -1.4211337628594796e-06
GC_11_239 b_11 NI_11 NS_239 0 -1.1580122978420691e-06
GC_11_240 b_11 NI_11 NS_240 0 -4.6157863595205710e-07
GC_11_241 b_11 NI_11 NS_241 0 -3.3852691545884133e-07
GC_11_242 b_11 NI_11 NS_242 0 -6.2315324588818936e-07
GC_11_243 b_11 NI_11 NS_243 0 -2.5799929714316297e-06
GC_11_244 b_11 NI_11 NS_244 0 -6.4781522436897912e-07
GC_11_245 b_11 NI_11 NS_245 0 7.1553442867100396e-07
GC_11_246 b_11 NI_11 NS_246 0 3.5782581913668396e-07
GC_11_247 b_11 NI_11 NS_247 0 -7.3448892007739897e-07
GC_11_248 b_11 NI_11 NS_248 0 3.7214420332345964e-07
GC_11_249 b_11 NI_11 NS_249 0 -9.8995946753587378e-07
GC_11_250 b_11 NI_11 NS_250 0 5.8052909844835030e-07
GC_11_251 b_11 NI_11 NS_251 0 -4.3434610103860359e-07
GC_11_252 b_11 NI_11 NS_252 0 2.6522545080181336e-07
GC_11_253 b_11 NI_11 NS_253 0 -8.4585927842600358e-07
GC_11_254 b_11 NI_11 NS_254 0 4.5732483789770261e-07
GC_11_255 b_11 NI_11 NS_255 0 1.5918319116360643e-07
GC_11_256 b_11 NI_11 NS_256 0 1.1045473228641425e-06
GC_11_257 b_11 NI_11 NS_257 0 -5.9724299603774906e-07
GC_11_258 b_11 NI_11 NS_258 0 1.3109632901594172e-07
GC_11_259 b_11 NI_11 NS_259 0 -1.8767397174429001e-06
GC_11_260 b_11 NI_11 NS_260 0 1.2955869096619141e-06
GC_11_261 b_11 NI_11 NS_261 0 2.0522690066996279e-06
GC_11_262 b_11 NI_11 NS_262 0 2.3513020289895809e-07
GC_11_263 b_11 NI_11 NS_263 0 -6.8553510359534961e-07
GC_11_264 b_11 NI_11 NS_264 0 2.0088554450894459e-07
GC_11_265 b_11 NI_11 NS_265 0 9.9851450651825409e-07
GC_11_266 b_11 NI_11 NS_266 0 1.6701841790290672e-06
GC_11_267 b_11 NI_11 NS_267 0 -2.4331624331578343e-07
GC_11_268 b_11 NI_11 NS_268 0 -5.7760829602983208e-07
GC_11_269 b_11 NI_11 NS_269 0 -9.1795090917066364e-07
GC_11_270 b_11 NI_11 NS_270 0 4.3082211091808717e-07
GC_11_271 b_11 NI_11 NS_271 0 1.4279737860394248e-06
GC_11_272 b_11 NI_11 NS_272 0 6.8214168898893333e-07
GC_11_273 b_11 NI_11 NS_273 0 -3.4147110124355281e-07
GC_11_274 b_11 NI_11 NS_274 0 -2.1170572833683183e-07
GC_11_275 b_11 NI_11 NS_275 0 -2.9973032421819261e-08
GC_11_276 b_11 NI_11 NS_276 0 1.4218684235262772e-06
GC_11_277 b_11 NI_11 NS_277 0 4.6149646692223300e-07
GC_11_278 b_11 NI_11 NS_278 0 -7.6771761030964285e-07
GC_11_279 b_11 NI_11 NS_279 0 -3.5264144432294186e-07
GC_11_280 b_11 NI_11 NS_280 0 4.8843601983341796e-08
GC_11_281 b_11 NI_11 NS_281 0 3.2445647290774525e-07
GC_11_282 b_11 NI_11 NS_282 0 3.7912989590733076e-07
GC_11_283 b_11 NI_11 NS_283 0 -1.4602248050188876e-07
GC_11_284 b_11 NI_11 NS_284 0 -8.6160914645058870e-09
GC_11_285 b_11 NI_11 NS_285 0 1.4120907853612055e-07
GC_11_286 b_11 NI_11 NS_286 0 1.2124342576912799e-07
GC_11_287 b_11 NI_11 NS_287 0 -1.9293193938516225e-07
GC_11_288 b_11 NI_11 NS_288 0 -6.8413909402798505e-08
GC_11_289 b_11 NI_11 NS_289 0 4.0854757841072955e-08
GC_11_290 b_11 NI_11 NS_290 0 1.9500430984673773e-07
GC_11_291 b_11 NI_11 NS_291 0 -1.1264869659048661e-07
GC_11_292 b_11 NI_11 NS_292 0 1.0076507602258905e-08
GC_11_293 b_11 NI_11 NS_293 0 4.5458878612895846e-08
GC_11_294 b_11 NI_11 NS_294 0 4.5514996226706029e-09
GC_11_295 b_11 NI_11 NS_295 0 -2.9963279919047614e-07
GC_11_296 b_11 NI_11 NS_296 0 -5.1511631288802537e-08
GC_11_297 b_11 NI_11 NS_297 0 -9.0274574510775435e-08
GC_11_298 b_11 NI_11 NS_298 0 6.0418075826641529e-08
GC_11_299 b_11 NI_11 NS_299 0 -2.3104816358488882e-07
GC_11_300 b_11 NI_11 NS_300 0 8.0694666168598535e-08
GC_11_301 b_11 NI_11 NS_301 0 -1.3259201454851455e-07
GC_11_302 b_11 NI_11 NS_302 0 -7.1016408018328023e-08
GC_11_303 b_11 NI_11 NS_303 0 -4.3085747419434909e-07
GC_11_304 b_11 NI_11 NS_304 0 -5.3628272140111442e-08
GC_11_305 b_11 NI_11 NS_305 0 -4.1936641858199375e-07
GC_11_306 b_11 NI_11 NS_306 0 6.1406870809296802e-08
GC_11_307 b_11 NI_11 NS_307 0 -4.4043839319192315e-07
GC_11_308 b_11 NI_11 NS_308 0 1.4691505936524078e-07
GC_11_309 b_11 NI_11 NS_309 0 -5.1097781673547644e-07
GC_11_310 b_11 NI_11 NS_310 0 9.9964491320560746e-08
GC_11_311 b_11 NI_11 NS_311 0 -9.6170605065650153e-07
GC_11_312 b_11 NI_11 NS_312 0 -9.6202559803950012e-08
GC_11_313 b_11 NI_11 NS_313 0 2.6182503860444805e-06
GC_11_314 b_11 NI_11 NS_314 0 2.9793849856569535e-06
GC_11_315 b_11 NI_11 NS_315 0 -6.1475114699314173e-07
GC_11_316 b_11 NI_11 NS_316 0 1.0339424523968106e-06
GC_11_317 b_11 NI_11 NS_317 0 9.1584998372080205e-09
GC_11_318 b_11 NI_11 NS_318 0 2.5337450515882057e-08
GC_11_319 b_11 NI_11 NS_319 0 -4.6874934250373500e-07
GC_11_320 b_11 NI_11 NS_320 0 8.2782641463831221e-07
GC_11_321 b_11 NI_11 NS_321 0 8.6792753414864640e-09
GC_11_322 b_11 NI_11 NS_322 0 3.8300019463063100e-07
GC_11_323 b_11 NI_11 NS_323 0 -8.6727475550593379e-07
GC_11_324 b_11 NI_11 NS_324 0 -7.0681872986867138e-08
GC_11_325 b_11 NI_11 NS_325 0 -9.7701451821693728e-07
GC_11_326 b_11 NI_11 NS_326 0 -1.7981804627726955e-07
GC_11_327 b_11 NI_11 NS_327 0 1.0738479246823597e-07
GC_11_328 b_11 NI_11 NS_328 0 -1.4754523679006921e-07
GC_11_329 b_11 NI_11 NS_329 0 6.6801840462151122e-08
GC_11_330 b_11 NI_11 NS_330 0 1.4718289185617590e-08
GC_11_331 b_11 NI_11 NS_331 0 -6.9818607200401221e-08
GC_11_332 b_11 NI_11 NS_332 0 1.6103509354122330e-07
GC_11_333 b_11 NI_11 NS_333 0 2.7786822844396172e-08
GC_11_334 b_11 NI_11 NS_334 0 -4.0821778534128821e-08
GC_11_335 b_11 NI_11 NS_335 0 -8.1243018206344208e-08
GC_11_336 b_11 NI_11 NS_336 0 1.6047197847309771e-07
GC_11_337 b_11 NI_11 NS_337 0 5.6556666141436279e-08
GC_11_338 b_11 NI_11 NS_338 0 -1.6778174566831400e-08
GC_11_339 b_11 NI_11 NS_339 0 -1.1804137311831385e-11
GC_11_340 b_11 NI_11 NS_340 0 5.2790194428412893e-12
GC_11_341 b_11 NI_11 NS_341 0 -3.4095489306712524e-10
GC_11_342 b_11 NI_11 NS_342 0 -9.7317210036866128e-10
GC_11_343 b_11 NI_11 NS_343 0 -2.7457116274305798e-05
GC_11_344 b_11 NI_11 NS_344 0 -1.0861416416346822e-08
GC_11_345 b_11 NI_11 NS_345 0 1.0271925129146228e-11
GC_11_346 b_11 NI_11 NS_346 0 -5.9963123483584810e-11
GC_11_347 b_11 NI_11 NS_347 0 -6.3441258445568957e-07
GC_11_348 b_11 NI_11 NS_348 0 -1.0701455391168440e-06
GC_11_349 b_11 NI_11 NS_349 0 -1.4351360125686452e-06
GC_11_350 b_11 NI_11 NS_350 0 2.3180833529912637e-06
GC_11_351 b_11 NI_11 NS_351 0 -3.8038674493693708e-06
GC_11_352 b_11 NI_11 NS_352 0 2.1755711742175594e-06
GC_11_353 b_11 NI_11 NS_353 0 1.9264451993277429e-06
GC_11_354 b_11 NI_11 NS_354 0 -2.2569193427501215e-07
GC_11_355 b_11 NI_11 NS_355 0 1.3997842057547016e-06
GC_11_356 b_11 NI_11 NS_356 0 5.7146518307279389e-06
GC_11_357 b_11 NI_11 NS_357 0 3.7149801521801161e-06
GC_11_358 b_11 NI_11 NS_358 0 3.2450679883401650e-06
GC_11_359 b_11 NI_11 NS_359 0 -1.4756060915753978e-06
GC_11_360 b_11 NI_11 NS_360 0 -9.4893529057189424e-07
GC_11_361 b_11 NI_11 NS_361 0 9.7598883137450343e-07
GC_11_362 b_11 NI_11 NS_362 0 -2.1769791970228486e-06
GC_11_363 b_11 NI_11 NS_363 0 6.4144573498058141e-06
GC_11_364 b_11 NI_11 NS_364 0 8.5314123664066499e-06
GC_11_365 b_11 NI_11 NS_365 0 1.3418230687535474e-06
GC_11_366 b_11 NI_11 NS_366 0 -9.5630628324226146e-07
GC_11_367 b_11 NI_11 NS_367 0 1.0785518765111698e-06
GC_11_368 b_11 NI_11 NS_368 0 -1.8906349462416897e-06
GC_11_369 b_11 NI_11 NS_369 0 1.4514949316372176e-05
GC_11_370 b_11 NI_11 NS_370 0 -4.1896481878040817e-06
GC_11_371 b_11 NI_11 NS_371 0 -2.0072622124420180e-07
GC_11_372 b_11 NI_11 NS_372 0 6.6359791822390559e-07
GC_11_373 b_11 NI_11 NS_373 0 4.9434744734746733e-06
GC_11_374 b_11 NI_11 NS_374 0 -2.1797934858154105e-06
GC_11_375 b_11 NI_11 NS_375 0 -7.7232618610028279e-07
GC_11_376 b_11 NI_11 NS_376 0 -1.5002610725189169e-05
GC_11_377 b_11 NI_11 NS_377 0 -7.8145956055893735e-08
GC_11_378 b_11 NI_11 NS_378 0 9.5809137869342357e-07
GC_11_379 b_11 NI_11 NS_379 0 -7.9221109285856375e-06
GC_11_380 b_11 NI_11 NS_380 0 -8.5843025198563364e-06
GC_11_381 b_11 NI_11 NS_381 0 -6.3256806868088361e-07
GC_11_382 b_11 NI_11 NS_382 0 -2.1422065998015091e-06
GC_11_383 b_11 NI_11 NS_383 0 -1.4555361633508426e-08
GC_11_384 b_11 NI_11 NS_384 0 1.1898562729845837e-06
GC_11_385 b_11 NI_11 NS_385 0 -7.7141173569142266e-06
GC_11_386 b_11 NI_11 NS_386 0 1.9653003255010448e-06
GC_11_387 b_11 NI_11 NS_387 0 2.3902057324950742e-07
GC_11_388 b_11 NI_11 NS_388 0 -1.6696994368076353e-06
GC_11_389 b_11 NI_11 NS_389 0 1.1429281058409575e-06
GC_11_390 b_11 NI_11 NS_390 0 3.0633288695732583e-06
GC_11_391 b_11 NI_11 NS_391 0 -9.6195459732978996e-07
GC_11_392 b_11 NI_11 NS_392 0 2.0271933705429169e-06
GC_11_393 b_11 NI_11 NS_393 0 4.5489649353217938e-07
GC_11_394 b_11 NI_11 NS_394 0 -1.2226883853941834e-06
GC_11_395 b_11 NI_11 NS_395 0 3.2356524353846653e-06
GC_11_396 b_11 NI_11 NS_396 0 -8.8238270585750551e-07
GC_11_397 b_11 NI_11 NS_397 0 -1.6005582729865135e-07
GC_11_398 b_11 NI_11 NS_398 0 5.0797765355727397e-07
GC_11_399 b_11 NI_11 NS_399 0 -8.4404696556218667e-07
GC_11_400 b_11 NI_11 NS_400 0 -4.1915992582540232e-07
GC_11_401 b_11 NI_11 NS_401 0 9.8705196739470441e-07
GC_11_402 b_11 NI_11 NS_402 0 -1.2634866134121166e-06
GC_11_403 b_11 NI_11 NS_403 0 1.4385529744577145e-06
GC_11_404 b_11 NI_11 NS_404 0 -5.6892309258109349e-07
GC_11_405 b_11 NI_11 NS_405 0 -3.3371916568801030e-08
GC_11_406 b_11 NI_11 NS_406 0 9.4899307520356583e-08
GC_11_407 b_11 NI_11 NS_407 0 -5.9608804315541099e-07
GC_11_408 b_11 NI_11 NS_408 0 -3.3988440066187845e-07
GC_11_409 b_11 NI_11 NS_409 0 9.6297819100606869e-07
GC_11_410 b_11 NI_11 NS_410 0 -1.0755606753992298e-06
GC_11_411 b_11 NI_11 NS_411 0 1.3913853505751093e-06
GC_11_412 b_11 NI_11 NS_412 0 -1.2415313471417361e-06
GC_11_413 b_11 NI_11 NS_413 0 1.6086493386951408e-07
GC_11_414 b_11 NI_11 NS_414 0 -4.5335273310913402e-08
GC_11_415 b_11 NI_11 NS_415 0 -4.8805854462887644e-07
GC_11_416 b_11 NI_11 NS_416 0 -5.0217695011910963e-07
GC_11_417 b_11 NI_11 NS_417 0 1.0601453818744863e-06
GC_11_418 b_11 NI_11 NS_418 0 -7.9957814936655465e-07
GC_11_419 b_11 NI_11 NS_419 0 1.2253752362460668e-06
GC_11_420 b_11 NI_11 NS_420 0 -2.1157360846420026e-06
GC_11_421 b_11 NI_11 NS_421 0 4.9451561060864110e-07
GC_11_422 b_11 NI_11 NS_422 0 -2.5501377388401963e-07
GC_11_423 b_11 NI_11 NS_423 0 -2.4640820247002772e-07
GC_11_424 b_11 NI_11 NS_424 0 -9.1750578611834430e-07
GC_11_425 b_11 NI_11 NS_425 0 1.9158047560070014e-06
GC_11_426 b_11 NI_11 NS_426 0 -9.9682471519435097e-07
GC_11_427 b_11 NI_11 NS_427 0 -8.0875005185356590e-06
GC_11_428 b_11 NI_11 NS_428 0 -9.1348565999229453e-07
GC_11_429 b_11 NI_11 NS_429 0 -3.1590611067453786e-07
GC_11_430 b_11 NI_11 NS_430 0 -3.6199056703646797e-06
GC_11_431 b_11 NI_11 NS_431 0 -4.8932270967711575e-08
GC_11_432 b_11 NI_11 NS_432 0 -3.3150813834730535e-08
GC_11_433 b_11 NI_11 NS_433 0 -1.0395727516854505e-07
GC_11_434 b_11 NI_11 NS_434 0 -1.2351416381125989e-06
GC_11_435 b_11 NI_11 NS_435 0 -1.0202864668351254e-06
GC_11_436 b_11 NI_11 NS_436 0 -6.6669686235342572e-07
GC_11_437 b_11 NI_11 NS_437 0 1.4550409845361842e-06
GC_11_438 b_11 NI_11 NS_438 0 -7.5894383497289286e-07
GC_11_439 b_11 NI_11 NS_439 0 1.9403533740223758e-06
GC_11_440 b_11 NI_11 NS_440 0 -1.8687465682841088e-06
GC_11_441 b_11 NI_11 NS_441 0 -2.2166695062197889e-07
GC_11_442 b_11 NI_11 NS_442 0 3.2466584366792171e-07
GC_11_443 b_11 NI_11 NS_443 0 2.1427805783732442e-07
GC_11_444 b_11 NI_11 NS_444 0 5.2885356731864283e-07
GC_11_445 b_11 NI_11 NS_445 0 -1.0742387794989876e-07
GC_11_446 b_11 NI_11 NS_446 0 -2.8271652230465506e-07
GC_11_447 b_11 NI_11 NS_447 0 7.8976027316850654e-09
GC_11_448 b_11 NI_11 NS_448 0 -9.5824314712196048e-08
GC_11_449 b_11 NI_11 NS_449 0 -8.8821447176799961e-08
GC_11_450 b_11 NI_11 NS_450 0 4.1483529025969118e-08
GC_11_451 b_11 NI_11 NS_451 0 -1.2204416056890153e-07
GC_11_452 b_11 NI_11 NS_452 0 -5.3450871590051749e-08
GC_11_453 b_11 NI_11 NS_453 0 6.1484538762158726e-12
GC_11_454 b_11 NI_11 NS_454 0 -1.7070422884008581e-12
GC_11_455 b_11 NI_11 NS_455 0 3.5216720149104188e-10
GC_11_456 b_11 NI_11 NS_456 0 6.9300699950415924e-10
GC_11_457 b_11 NI_11 NS_457 0 8.4580444223879178e-05
GC_11_458 b_11 NI_11 NS_458 0 1.9045626105667682e-07
GC_11_459 b_11 NI_11 NS_459 0 2.0155274496148803e-11
GC_11_460 b_11 NI_11 NS_460 0 -9.4458295807957883e-10
GC_11_461 b_11 NI_11 NS_461 0 8.8329947726713279e-07
GC_11_462 b_11 NI_11 NS_462 0 5.7933425880103152e-08
GC_11_463 b_11 NI_11 NS_463 0 1.1602010077557045e-06
GC_11_464 b_11 NI_11 NS_464 0 6.9968105261025649e-08
GC_11_465 b_11 NI_11 NS_465 0 3.3628862048474323e-06
GC_11_466 b_11 NI_11 NS_466 0 -3.2258608605592207e-06
GC_11_467 b_11 NI_11 NS_467 0 -2.0855280312256105e-06
GC_11_468 b_11 NI_11 NS_468 0 -1.7319080763419381e-06
GC_11_469 b_11 NI_11 NS_469 0 1.9313031097616848e-06
GC_11_470 b_11 NI_11 NS_470 0 -2.2094016347459393e-06
GC_11_471 b_11 NI_11 NS_471 0 -5.8922110604462330e-06
GC_11_472 b_11 NI_11 NS_472 0 -7.1422706064320229e-06
GC_11_473 b_11 NI_11 NS_473 0 9.4972535928061161e-07
GC_11_474 b_11 NI_11 NS_474 0 2.2263820796417764e-06
GC_11_475 b_11 NI_11 NS_475 0 -2.2764210873014525e-06
GC_11_476 b_11 NI_11 NS_476 0 8.0098703003545140e-07
GC_11_477 b_11 NI_11 NS_477 0 5.8207644674714172e-07
GC_11_478 b_11 NI_11 NS_478 0 -4.8941597637291085e-06
GC_11_479 b_11 NI_11 NS_479 0 -6.4023894383029666e-06
GC_11_480 b_11 NI_11 NS_480 0 2.7555984854984618e-06
GC_11_481 b_11 NI_11 NS_481 0 -1.0155998316542175e-06
GC_11_482 b_11 NI_11 NS_482 0 1.6581852477160933e-06
GC_11_483 b_11 NI_11 NS_483 0 -3.3720580846898163e-06
GC_11_484 b_11 NI_11 NS_484 0 -2.5292967797300869e-06
GC_11_485 b_11 NI_11 NS_485 0 -2.2047549298747554e-06
GC_11_486 b_11 NI_11 NS_486 0 2.3621389568241038e-06
GC_11_487 b_11 NI_11 NS_487 0 1.5152440479194506e-06
GC_11_488 b_11 NI_11 NS_488 0 2.6088613388854030e-06
GC_11_489 b_11 NI_11 NS_489 0 -5.1183461052463439e-06
GC_11_490 b_11 NI_11 NS_490 0 -2.0383785607321994e-06
GC_11_491 b_11 NI_11 NS_491 0 -1.4940206057811735e-06
GC_11_492 b_11 NI_11 NS_492 0 2.2226897803345989e-06
GC_11_493 b_11 NI_11 NS_493 0 -4.8359641797109115e-08
GC_11_494 b_11 NI_11 NS_494 0 -1.0715150338090601e-06
GC_11_495 b_11 NI_11 NS_495 0 -2.7776174817228212e-06
GC_11_496 b_11 NI_11 NS_496 0 1.7676086722363852e-06
GC_11_497 b_11 NI_11 NS_497 0 -7.8765239373512284e-07
GC_11_498 b_11 NI_11 NS_498 0 2.3415814041636951e-06
GC_11_499 b_11 NI_11 NS_499 0 -1.0034713210210130e-06
GC_11_500 b_11 NI_11 NS_500 0 -1.3434469544755512e-06
GC_11_501 b_11 NI_11 NS_501 0 -1.8384294998337534e-06
GC_11_502 b_11 NI_11 NS_502 0 1.3364981930409243e-06
GC_11_503 b_11 NI_11 NS_503 0 5.5164880955705404e-07
GC_11_504 b_11 NI_11 NS_504 0 1.6482318250341835e-07
GC_11_505 b_11 NI_11 NS_505 0 -2.9422070809255354e-06
GC_11_506 b_11 NI_11 NS_506 0 3.7599796260834070e-07
GC_11_507 b_11 NI_11 NS_507 0 -9.6502852166146697e-07
GC_11_508 b_11 NI_11 NS_508 0 7.1171507970713853e-07
GC_11_509 b_11 NI_11 NS_509 0 -1.9725522363563264e-06
GC_11_510 b_11 NI_11 NS_510 0 -7.9508491540134712e-07
GC_11_511 b_11 NI_11 NS_511 0 -1.4687384186706020e-06
GC_11_512 b_11 NI_11 NS_512 0 6.2098843424795178e-07
GC_11_513 b_11 NI_11 NS_513 0 -1.1171724357837201e-06
GC_11_514 b_11 NI_11 NS_514 0 -3.9225835013168238e-07
GC_11_515 b_11 NI_11 NS_515 0 -2.4594675070046001e-06
GC_11_516 b_11 NI_11 NS_516 0 -6.3473558757363386e-07
GC_11_517 b_11 NI_11 NS_517 0 -3.0280709149246042e-06
GC_11_518 b_11 NI_11 NS_518 0 -3.1143930841390479e-07
GC_11_519 b_11 NI_11 NS_519 0 -2.1722198011863700e-06
GC_11_520 b_11 NI_11 NS_520 0 3.1818641840297836e-07
GC_11_521 b_11 NI_11 NS_521 0 -2.7406254636243139e-06
GC_11_522 b_11 NI_11 NS_522 0 3.0317817816327682e-07
GC_11_523 b_11 NI_11 NS_523 0 -4.2061080180847485e-06
GC_11_524 b_11 NI_11 NS_524 0 -7.3435620226901688e-07
GC_11_525 b_11 NI_11 NS_525 0 -5.6819242708197152e-06
GC_11_526 b_11 NI_11 NS_526 0 2.2499642522214055e-06
GC_11_527 b_11 NI_11 NS_527 0 -3.1747527620975799e-06
GC_11_528 b_11 NI_11 NS_528 0 1.8635246952527558e-06
GC_11_529 b_11 NI_11 NS_529 0 -4.1153814370569324e-06
GC_11_530 b_11 NI_11 NS_530 0 3.2994552957701525e-06
GC_11_531 b_11 NI_11 NS_531 0 -5.6740252534126332e-06
GC_11_532 b_11 NI_11 NS_532 0 1.3489955797872204e-06
GC_11_533 b_11 NI_11 NS_533 0 -3.5119894705847739e-06
GC_11_534 b_11 NI_11 NS_534 0 8.2346882899706213e-06
GC_11_535 b_11 NI_11 NS_535 0 -2.3076938386385822e-06
GC_11_536 b_11 NI_11 NS_536 0 4.5638149156953067e-06
GC_11_537 b_11 NI_11 NS_537 0 1.1261130714072121e-06
GC_11_538 b_11 NI_11 NS_538 0 5.4139213433355775e-06
GC_11_539 b_11 NI_11 NS_539 0 -1.8428020065489739e-06
GC_11_540 b_11 NI_11 NS_540 0 3.4530151107922822e-06
GC_11_541 b_11 NI_11 NS_541 0 -7.0172848715939272e-06
GC_11_542 b_11 NI_11 NS_542 0 3.7168282265697131e-05
GC_11_543 b_11 NI_11 NS_543 0 6.9494316448313509e-07
GC_11_544 b_11 NI_11 NS_544 0 2.6509038508028006e-06
GC_11_545 b_11 NI_11 NS_545 0 -8.4712154291533521e-08
GC_11_546 b_11 NI_11 NS_546 0 1.1840329431228899e-07
GC_11_547 b_11 NI_11 NS_547 0 -7.2440198324294493e-07
GC_11_548 b_11 NI_11 NS_548 0 3.4149225486108697e-06
GC_11_549 b_11 NI_11 NS_549 0 6.7713243778266922e-07
GC_11_550 b_11 NI_11 NS_550 0 8.6106598554714661e-07
GC_11_551 b_11 NI_11 NS_551 0 2.2825495040750223e-06
GC_11_552 b_11 NI_11 NS_552 0 -3.1366057486517447e-06
GC_11_553 b_11 NI_11 NS_553 0 -1.5483050919445345e-06
GC_11_554 b_11 NI_11 NS_554 0 -1.1843703893156053e-05
GC_11_555 b_11 NI_11 NS_555 0 2.0447490035509154e-06
GC_11_556 b_11 NI_11 NS_556 0 -7.3740383286643397e-07
GC_11_557 b_11 NI_11 NS_557 0 4.5135000508968605e-06
GC_11_558 b_11 NI_11 NS_558 0 -4.0110367010178724e-07
GC_11_559 b_11 NI_11 NS_559 0 1.2442190688948713e-06
GC_11_560 b_11 NI_11 NS_560 0 1.9853481328671771e-06
GC_11_561 b_11 NI_11 NS_561 0 1.7411980671585392e-06
GC_11_562 b_11 NI_11 NS_562 0 -7.6164713208814375e-07
GC_11_563 b_11 NI_11 NS_563 0 5.8319426172573245e-07
GC_11_564 b_11 NI_11 NS_564 0 5.1104633954696583e-07
GC_11_565 b_11 NI_11 NS_565 0 6.5669153833478978e-07
GC_11_566 b_11 NI_11 NS_566 0 -7.6193902185868505e-08
GC_11_567 b_11 NI_11 NS_567 0 2.2925820252429275e-11
GC_11_568 b_11 NI_11 NS_568 0 -9.3367295004400399e-11
GC_11_569 b_11 NI_11 NS_569 0 -1.8302754337372487e-09
GC_11_570 b_11 NI_11 NS_570 0 4.0623346478956023e-09
GC_11_571 b_11 NI_11 NS_571 0 -6.3086683869682209e-05
GC_11_572 b_11 NI_11 NS_572 0 3.1407861644456421e-07
GC_11_573 b_11 NI_11 NS_573 0 1.6213783984299794e-11
GC_11_574 b_11 NI_11 NS_574 0 -9.0526371008467824e-11
GC_11_575 b_11 NI_11 NS_575 0 -1.1178117688183584e-06
GC_11_576 b_11 NI_11 NS_576 0 -1.7847514932852855e-06
GC_11_577 b_11 NI_11 NS_577 0 -1.9986034286070562e-06
GC_11_578 b_11 NI_11 NS_578 0 1.9870799516978829e-06
GC_11_579 b_11 NI_11 NS_579 0 -9.6875215984189863e-06
GC_11_580 b_11 NI_11 NS_580 0 6.6934231309478623e-07
GC_11_581 b_11 NI_11 NS_581 0 -2.3280748123349641e-07
GC_11_582 b_11 NI_11 NS_582 0 3.4992284186455021e-06
GC_11_583 b_11 NI_11 NS_583 0 -2.1124292791001670e-06
GC_11_584 b_11 NI_11 NS_584 0 1.1812011421232556e-05
GC_11_585 b_11 NI_11 NS_585 0 6.7540260318347113e-06
GC_11_586 b_11 NI_11 NS_586 0 1.2474521970903150e-05
GC_11_587 b_11 NI_11 NS_587 0 -1.9954535313637184e-06
GC_11_588 b_11 NI_11 NS_588 0 -2.3039262604070079e-06
GC_11_589 b_11 NI_11 NS_589 0 1.6659032589243336e-06
GC_11_590 b_11 NI_11 NS_590 0 9.5797578680143739e-07
GC_11_591 b_11 NI_11 NS_591 0 7.5629425686997020e-06
GC_11_592 b_11 NI_11 NS_592 0 3.8828223145173483e-05
GC_11_593 b_11 NI_11 NS_593 0 2.3010293943395847e-05
GC_11_594 b_11 NI_11 NS_594 0 -1.1868418147204981e-05
GC_11_595 b_11 NI_11 NS_595 0 8.3672992794143778e-06
GC_11_596 b_11 NI_11 NS_596 0 1.6445433310500279e-06
GC_11_597 b_11 NI_11 NS_597 0 4.8509113307476302e-05
GC_11_598 b_11 NI_11 NS_598 0 -2.5181071657765159e-05
GC_11_599 b_11 NI_11 NS_599 0 -8.8536770958468418e-07
GC_11_600 b_11 NI_11 NS_600 0 -7.8651568708001922e-06
GC_11_601 b_11 NI_11 NS_601 0 3.4167775442414077e-05
GC_11_602 b_11 NI_11 NS_602 0 -7.8499518819513066e-06
GC_11_603 b_11 NI_11 NS_603 0 -3.8183058309379491e-05
GC_11_604 b_11 NI_11 NS_604 0 -5.2548377571092351e-05
GC_11_605 b_11 NI_11 NS_605 0 -4.5027056411737533e-06
GC_11_606 b_11 NI_11 NS_606 0 -4.3379495753987538e-06
GC_11_607 b_11 NI_11 NS_607 0 -3.9815357297173128e-05
GC_11_608 b_11 NI_11 NS_608 0 -2.0116799697586378e-05
GC_11_609 b_11 NI_11 NS_609 0 -4.8511662055573176e-06
GC_11_610 b_11 NI_11 NS_610 0 6.2282653960587718e-06
GC_11_611 b_11 NI_11 NS_611 0 -8.5210924052821246e-06
GC_11_612 b_11 NI_11 NS_612 0 -4.5734610210173262e-07
GC_11_613 b_11 NI_11 NS_613 0 -1.5552800923999749e-05
GC_11_614 b_11 NI_11 NS_614 0 2.4319405066934624e-05
GC_11_615 b_11 NI_11 NS_615 0 1.1127392626597661e-06
GC_11_616 b_11 NI_11 NS_616 0 2.3765185500278477e-06
GC_11_617 b_11 NI_11 NS_617 0 3.2444559116654848e-06
GC_11_618 b_11 NI_11 NS_618 0 1.8514020574786194e-05
GC_11_619 b_11 NI_11 NS_619 0 7.5499006387489316e-06
GC_11_620 b_11 NI_11 NS_620 0 -1.4049663834718512e-06
GC_11_621 b_11 NI_11 NS_621 0 2.9997389478206481e-06
GC_11_622 b_11 NI_11 NS_622 0 -5.0735572303566729e-07
GC_11_623 b_11 NI_11 NS_623 0 7.6482559978961723e-06
GC_11_624 b_11 NI_11 NS_624 0 -4.5383939791329968e-06
GC_11_625 b_11 NI_11 NS_625 0 -8.6323797573449399e-07
GC_11_626 b_11 NI_11 NS_626 0 -4.4782454596052580e-07
GC_11_627 b_11 NI_11 NS_627 0 -1.7220281997726822e-06
GC_11_628 b_11 NI_11 NS_628 0 1.8650796350269996e-07
GC_11_629 b_11 NI_11 NS_629 0 1.6124747321701393e-06
GC_11_630 b_11 NI_11 NS_630 0 -2.3831634763138513e-08
GC_11_631 b_11 NI_11 NS_631 0 3.7027762597270841e-06
GC_11_632 b_11 NI_11 NS_632 0 -9.2679544867830183e-07
GC_11_633 b_11 NI_11 NS_633 0 -8.7846709291032456e-08
GC_11_634 b_11 NI_11 NS_634 0 -3.4244766562819230e-07
GC_11_635 b_11 NI_11 NS_635 0 -5.7040323478614785e-07
GC_11_636 b_11 NI_11 NS_636 0 5.1106396608040938e-07
GC_11_637 b_11 NI_11 NS_637 0 2.4651899982570030e-06
GC_11_638 b_11 NI_11 NS_638 0 1.0968737282728920e-07
GC_11_639 b_11 NI_11 NS_639 0 3.4039022124554938e-06
GC_11_640 b_11 NI_11 NS_640 0 -2.8600680635866036e-06
GC_11_641 b_11 NI_11 NS_641 0 -2.6935566574374985e-07
GC_11_642 b_11 NI_11 NS_642 0 -4.9653654659598325e-08
GC_11_643 b_11 NI_11 NS_643 0 7.1909533001190973e-07
GC_11_644 b_11 NI_11 NS_644 0 1.0039442969558248e-06
GC_11_645 b_11 NI_11 NS_645 0 3.5525134673748668e-06
GC_11_646 b_11 NI_11 NS_646 0 3.5545284883164120e-08
GC_11_647 b_11 NI_11 NS_647 0 2.4198816383953975e-06
GC_11_648 b_11 NI_11 NS_648 0 -4.6562321120814863e-06
GC_11_649 b_11 NI_11 NS_649 0 4.5356122457631713e-07
GC_11_650 b_11 NI_11 NS_650 0 1.1318779847402097e-06
GC_11_651 b_11 NI_11 NS_651 0 3.6738640502719682e-06
GC_11_652 b_11 NI_11 NS_652 0 -6.8877932822912533e-07
GC_11_653 b_11 NI_11 NS_653 0 5.6188352233486683e-06
GC_11_654 b_11 NI_11 NS_654 0 -9.6836418328652552e-07
GC_11_655 b_11 NI_11 NS_655 0 -1.6176046078432396e-05
GC_11_656 b_11 NI_11 NS_656 0 -1.0667592246453710e-05
GC_11_657 b_11 NI_11 NS_657 0 9.4793381353664641e-07
GC_11_658 b_11 NI_11 NS_658 0 -7.4950695056465363e-06
GC_11_659 b_11 NI_11 NS_659 0 -6.7190847624418021e-08
GC_11_660 b_11 NI_11 NS_660 0 -1.4892254481570223e-07
GC_11_661 b_11 NI_11 NS_661 0 1.8092922886064027e-06
GC_11_662 b_11 NI_11 NS_662 0 -1.8934246859680776e-06
GC_11_663 b_11 NI_11 NS_663 0 5.4099511390168843e-07
GC_11_664 b_11 NI_11 NS_664 0 -3.3989100143044172e-06
GC_11_665 b_11 NI_11 NS_665 0 3.4155741078635617e-06
GC_11_666 b_11 NI_11 NS_666 0 -1.3122436946519261e-06
GC_11_667 b_11 NI_11 NS_667 0 4.5903000778627845e-06
GC_11_668 b_11 NI_11 NS_668 0 -7.9885899116713642e-07
GC_11_669 b_11 NI_11 NS_669 0 -1.9723770389684806e-07
GC_11_670 b_11 NI_11 NS_670 0 -2.0613810491344983e-07
GC_11_671 b_11 NI_11 NS_671 0 7.0253899739999072e-07
GC_11_672 b_11 NI_11 NS_672 0 1.4071793610437722e-06
GC_11_673 b_11 NI_11 NS_673 0 -7.0005281001599812e-07
GC_11_674 b_11 NI_11 NS_674 0 -1.4722238274682817e-06
GC_11_675 b_11 NI_11 NS_675 0 -6.2852517976928968e-07
GC_11_676 b_11 NI_11 NS_676 0 8.2374772720113704e-07
GC_11_677 b_11 NI_11 NS_677 0 2.2513785359008874e-07
GC_11_678 b_11 NI_11 NS_678 0 6.5418603541886232e-07
GC_11_679 b_11 NI_11 NS_679 0 6.0606475511975824e-07
GC_11_680 b_11 NI_11 NS_680 0 2.1063112244758158e-08
GC_11_681 b_11 NI_11 NS_681 0 1.3943978147208569e-11
GC_11_682 b_11 NI_11 NS_682 0 5.4830595139577640e-13
GC_11_683 b_11 NI_11 NS_683 0 4.3772452088799673e-10
GC_11_684 b_11 NI_11 NS_684 0 1.6923729878328266e-09
GC_11_685 b_11 NI_11 NS_685 0 -1.1277210786203245e-04
GC_11_686 b_11 NI_11 NS_686 0 -2.1518464769279575e-06
GC_11_687 b_11 NI_11 NS_687 0 -2.4613965129134436e-10
GC_11_688 b_11 NI_11 NS_688 0 2.5681351049888242e-09
GC_11_689 b_11 NI_11 NS_689 0 1.7816033662098149e-06
GC_11_690 b_11 NI_11 NS_690 0 -1.5815621155464114e-06
GC_11_691 b_11 NI_11 NS_691 0 2.3533689977139154e-07
GC_11_692 b_11 NI_11 NS_692 0 -6.4013237316979109e-06
GC_11_693 b_11 NI_11 NS_693 0 -7.4872988338856100e-06
GC_11_694 b_11 NI_11 NS_694 0 -2.0463982632243115e-07
GC_11_695 b_11 NI_11 NS_695 0 -1.3991988953532271e-06
GC_11_696 b_11 NI_11 NS_696 0 -4.6879150808647445e-06
GC_11_697 b_11 NI_11 NS_697 0 -1.5829941785818928e-05
GC_11_698 b_11 NI_11 NS_698 0 -1.8864567648885549e-06
GC_11_699 b_11 NI_11 NS_699 0 -6.8244339792956212e-06
GC_11_700 b_11 NI_11 NS_700 0 1.8864266834729853e-05
GC_11_701 b_11 NI_11 NS_701 0 4.8188265900013667e-06
GC_11_702 b_11 NI_11 NS_702 0 -2.8796975653713559e-06
GC_11_703 b_11 NI_11 NS_703 0 -1.3563214707975785e-07
GC_11_704 b_11 NI_11 NS_704 0 -2.4716414218674549e-06
GC_11_705 b_11 NI_11 NS_705 0 -2.6117097797787346e-05
GC_11_706 b_11 NI_11 NS_706 0 2.8150832302653728e-05
GC_11_707 b_11 NI_11 NS_707 0 2.8021136251792301e-05
GC_11_708 b_11 NI_11 NS_708 0 -8.1067138956420475e-06
GC_11_709 b_11 NI_11 NS_709 0 -8.0870808233292159e-06
GC_11_710 b_11 NI_11 NS_710 0 -4.2194541638888881e-06
GC_11_711 b_11 NI_11 NS_711 0 1.2345315585526195e-05
GC_11_712 b_11 NI_11 NS_712 0 2.7049491977171819e-05
GC_11_713 b_11 NI_11 NS_713 0 1.4325014334520080e-06
GC_11_714 b_11 NI_11 NS_714 0 -8.8303088946745078e-06
GC_11_715 b_11 NI_11 NS_715 0 -2.8319562997335517e-05
GC_11_716 b_11 NI_11 NS_716 0 4.8085423274449224e-06
GC_11_717 b_11 NI_11 NS_717 0 4.1184590117051691e-05
GC_11_718 b_11 NI_11 NS_718 0 1.0835845468590339e-05
GC_11_719 b_11 NI_11 NS_719 0 -3.0015681934964476e-06
GC_11_720 b_11 NI_11 NS_720 0 -4.3670101538050487e-06
GC_11_721 b_11 NI_11 NS_721 0 1.2955898676300235e-05
GC_11_722 b_11 NI_11 NS_722 0 1.9080714764958941e-05
GC_11_723 b_11 NI_11 NS_723 0 3.7635944130425238e-06
GC_11_724 b_11 NI_11 NS_724 0 -1.0833681891382544e-05
GC_11_725 b_11 NI_11 NS_725 0 -6.4466353103392831e-06
GC_11_726 b_11 NI_11 NS_726 0 9.6349173042500093e-07
GC_11_727 b_11 NI_11 NS_727 0 1.8926188284032420e-05
GC_11_728 b_11 NI_11 NS_728 0 5.4714303780027754e-06
GC_11_729 b_11 NI_11 NS_729 0 -1.1342490437568887e-07
GC_11_730 b_11 NI_11 NS_730 0 -4.1223382561935413e-06
GC_11_731 b_11 NI_11 NS_731 0 4.9483400785335101e-06
GC_11_732 b_11 NI_11 NS_732 0 1.4379800960982239e-05
GC_11_733 b_11 NI_11 NS_733 0 7.7968519537862621e-06
GC_11_734 b_11 NI_11 NS_734 0 -1.1164421057361544e-05
GC_11_735 b_11 NI_11 NS_735 0 -1.4154740088833200e-06
GC_11_736 b_11 NI_11 NS_736 0 9.8362929926054339e-07
GC_11_737 b_11 NI_11 NS_737 0 1.0884949593993562e-05
GC_11_738 b_11 NI_11 NS_738 0 4.1621733737805311e-06
GC_11_739 b_11 NI_11 NS_739 0 1.6970822798690003e-06
GC_11_740 b_11 NI_11 NS_740 0 -5.9090565832352541e-07
GC_11_741 b_11 NI_11 NS_741 0 5.6760840611175015e-06
GC_11_742 b_11 NI_11 NS_742 0 1.7180061137786339e-06
GC_11_743 b_11 NI_11 NS_743 0 3.3604893739545593e-06
GC_11_744 b_11 NI_11 NS_744 0 2.0717605506848228e-06
GC_11_745 b_11 NI_11 NS_745 0 1.0946296489747717e-05
GC_11_746 b_11 NI_11 NS_746 0 3.8300823165481868e-06
GC_11_747 b_11 NI_11 NS_747 0 4.8385991607017169e-06
GC_11_748 b_11 NI_11 NS_748 0 -5.2549180698228284e-08
GC_11_749 b_11 NI_11 NS_749 0 9.9675844446766836e-06
GC_11_750 b_11 NI_11 NS_750 0 -1.0598260062023872e-06
GC_11_751 b_11 NI_11 NS_751 0 8.2081792685010753e-06
GC_11_752 b_11 NI_11 NS_752 0 2.9740306469603556e-06
GC_11_753 b_11 NI_11 NS_753 0 1.9026488785986705e-05
GC_11_754 b_11 NI_11 NS_754 0 -5.5233826128892799e-06
GC_11_755 b_11 NI_11 NS_755 0 7.1917044921243087e-06
GC_11_756 b_11 NI_11 NS_756 0 -3.9943585022325621e-06
GC_11_757 b_11 NI_11 NS_757 0 1.3712813691243259e-05
GC_11_758 b_11 NI_11 NS_758 0 -1.1879978878053086e-05
GC_11_759 b_11 NI_11 NS_759 0 1.2365923391439787e-05
GC_11_760 b_11 NI_11 NS_760 0 -3.9393633422189438e-06
GC_11_761 b_11 NI_11 NS_761 0 9.1636805321919920e-06
GC_11_762 b_11 NI_11 NS_762 0 -2.6747062579591323e-05
GC_11_763 b_11 NI_11 NS_763 0 2.3618350542030239e-06
GC_11_764 b_11 NI_11 NS_764 0 -1.2358488737114878e-05
GC_11_765 b_11 NI_11 NS_765 0 -8.2831497475932082e-06
GC_11_766 b_11 NI_11 NS_766 0 -1.8645470334922066e-05
GC_11_767 b_11 NI_11 NS_767 0 -4.8702696217547839e-06
GC_11_768 b_11 NI_11 NS_768 0 -1.2077489879306745e-05
GC_11_769 b_11 NI_11 NS_769 0 5.4674645295482846e-05
GC_11_770 b_11 NI_11 NS_770 0 -8.8166253369074388e-05
GC_11_771 b_11 NI_11 NS_771 0 -1.0018835464702479e-05
GC_11_772 b_11 NI_11 NS_772 0 1.2701497229550513e-06
GC_11_773 b_11 NI_11 NS_773 0 3.8983284796819513e-07
GC_11_774 b_11 NI_11 NS_774 0 -1.2677284199467955e-07
GC_11_775 b_11 NI_11 NS_775 0 -2.7052832156928818e-06
GC_11_776 b_11 NI_11 NS_776 0 -1.9795977785539399e-06
GC_11_777 b_11 NI_11 NS_777 0 -4.4027975598772235e-06
GC_11_778 b_11 NI_11 NS_778 0 5.4784844523691559e-07
GC_11_779 b_11 NI_11 NS_779 0 -1.7423550302082378e-05
GC_11_780 b_11 NI_11 NS_780 0 9.5920517951428180e-06
GC_11_781 b_11 NI_11 NS_781 0 -9.1285281268714924e-06
GC_11_782 b_11 NI_11 NS_782 0 3.7355110740785198e-05
GC_11_783 b_11 NI_11 NS_783 0 -7.2451100075424161e-06
GC_11_784 b_11 NI_11 NS_784 0 3.3527604454305460e-07
GC_11_785 b_11 NI_11 NS_785 0 -1.3395935272804419e-05
GC_11_786 b_11 NI_11 NS_786 0 1.8751236121959655e-06
GC_11_787 b_11 NI_11 NS_787 0 -4.6442422014426192e-06
GC_11_788 b_11 NI_11 NS_788 0 -3.3978550327239070e-06
GC_11_789 b_11 NI_11 NS_789 0 -6.4046490466764472e-06
GC_11_790 b_11 NI_11 NS_790 0 1.0361834594963778e-06
GC_11_791 b_11 NI_11 NS_791 0 -3.0540566103477308e-06
GC_11_792 b_11 NI_11 NS_792 0 8.8642143154041784e-07
GC_11_793 b_11 NI_11 NS_793 0 -1.7952292063618197e-06
GC_11_794 b_11 NI_11 NS_794 0 -9.3643238317164582e-07
GC_11_795 b_11 NI_11 NS_795 0 -2.6050211534336509e-10
GC_11_796 b_11 NI_11 NS_796 0 4.2261540855450003e-10
GC_11_797 b_11 NI_11 NS_797 0 2.3349518572001670e-09
GC_11_798 b_11 NI_11 NS_798 0 -2.6679272653033660e-08
GC_11_799 b_11 NI_11 NS_799 0 -3.7757926301782143e-05
GC_11_800 b_11 NI_11 NS_800 0 2.2260818924540788e-06
GC_11_801 b_11 NI_11 NS_801 0 6.0497519034676064e-11
GC_11_802 b_11 NI_11 NS_802 0 3.0748149740279912e-09
GC_11_803 b_11 NI_11 NS_803 0 -1.9314697237325641e-06
GC_11_804 b_11 NI_11 NS_804 0 -1.7211201004480580e-06
GC_11_805 b_11 NI_11 NS_805 0 -5.6037063146461473e-06
GC_11_806 b_11 NI_11 NS_806 0 2.9249829424147494e-06
GC_11_807 b_11 NI_11 NS_807 0 -1.6662619245859438e-05
GC_11_808 b_11 NI_11 NS_808 0 1.9136408509925351e-05
GC_11_809 b_11 NI_11 NS_809 0 1.5401444989273528e-05
GC_11_810 b_11 NI_11 NS_810 0 1.0211362852644530e-05
GC_11_811 b_11 NI_11 NS_811 0 1.7356961749479004e-05
GC_11_812 b_11 NI_11 NS_812 0 2.3278420772984116e-05
GC_11_813 b_11 NI_11 NS_813 0 3.0898150773782620e-05
GC_11_814 b_11 NI_11 NS_814 0 5.3461970324299734e-06
GC_11_815 b_11 NI_11 NS_815 0 -3.3856238138808187e-06
GC_11_816 b_11 NI_11 NS_816 0 -2.1458381472888381e-06
GC_11_817 b_11 NI_11 NS_817 0 1.7190879971579605e-05
GC_11_818 b_11 NI_11 NS_818 0 -2.2223157343882964e-06
GC_11_819 b_11 NI_11 NS_819 0 1.2979334904903513e-04
GC_11_820 b_11 NI_11 NS_820 0 3.5245900906440898e-05
GC_11_821 b_11 NI_11 NS_821 0 -2.8532249493516027e-05
GC_11_822 b_11 NI_11 NS_822 0 -9.9831824368078724e-05
GC_11_823 b_11 NI_11 NS_823 0 2.5236662429538445e-05
GC_11_824 b_11 NI_11 NS_824 0 -3.1266673826410022e-05
GC_11_825 b_11 NI_11 NS_825 0 -4.0929314097212900e-05
GC_11_826 b_11 NI_11 NS_826 0 -1.6750258977753216e-04
GC_11_827 b_11 NI_11 NS_827 0 -4.1821230098493446e-05
GC_11_828 b_11 NI_11 NS_828 0 -5.3848026548872113e-06
GC_11_829 b_11 NI_11 NS_829 0 2.2549798698928803e-05
GC_11_830 b_11 NI_11 NS_830 0 -1.5151993988982721e-04
GC_11_831 b_11 NI_11 NS_831 0 -2.3148578994629709e-04
GC_11_832 b_11 NI_11 NS_832 0 1.1299682855767654e-04
GC_11_833 b_11 NI_11 NS_833 0 -3.7411184224793296e-05
GC_11_834 b_11 NI_11 NS_834 0 1.3952070456709377e-05
GC_11_835 b_11 NI_11 NS_835 0 -1.3781868631210014e-04
GC_11_836 b_11 NI_11 NS_836 0 1.2973370401669137e-04
GC_11_837 b_11 NI_11 NS_837 0 3.6131599536200630e-05
GC_11_838 b_11 NI_11 NS_838 0 4.1461238625778583e-05
GC_11_839 b_11 NI_11 NS_839 0 -3.8173653947803063e-05
GC_11_840 b_11 NI_11 NS_840 0 4.2970718353182850e-05
GC_11_841 b_11 NI_11 NS_841 0 8.7353506371169403e-05
GC_11_842 b_11 NI_11 NS_842 0 1.1821522000521526e-04
GC_11_843 b_11 NI_11 NS_843 0 2.7244714405443371e-05
GC_11_844 b_11 NI_11 NS_844 0 1.0262298035725672e-05
GC_11_845 b_11 NI_11 NS_845 0 8.7157828294067902e-05
GC_11_846 b_11 NI_11 NS_846 0 6.5380837168884008e-05
GC_11_847 b_11 NI_11 NS_847 0 2.0401053684571904e-05
GC_11_848 b_11 NI_11 NS_848 0 -5.7168349314372884e-05
GC_11_849 b_11 NI_11 NS_849 0 1.7001785515744761e-05
GC_11_850 b_11 NI_11 NS_850 0 -8.8439359491393649e-06
GC_11_851 b_11 NI_11 NS_851 0 8.4707981187111964e-06
GC_11_852 b_11 NI_11 NS_852 0 -3.3126354418953930e-05
GC_11_853 b_11 NI_11 NS_853 0 -8.8428225692262233e-06
GC_11_854 b_11 NI_11 NS_854 0 4.1504017798523653e-07
GC_11_855 b_11 NI_11 NS_855 0 -2.4023060465208659e-06
GC_11_856 b_11 NI_11 NS_856 0 8.4362063642728738e-06
GC_11_857 b_11 NI_11 NS_857 0 1.0207724315508014e-05
GC_11_858 b_11 NI_11 NS_858 0 6.0581933411192760e-06
GC_11_859 b_11 NI_11 NS_859 0 1.2154854488613014e-05
GC_11_860 b_11 NI_11 NS_860 0 -7.9359481714647789e-06
GC_11_861 b_11 NI_11 NS_861 0 -3.4649634450698435e-06
GC_11_862 b_11 NI_11 NS_862 0 -5.2259415046011141e-07
GC_11_863 b_11 NI_11 NS_863 0 2.5131894265998390e-06
GC_11_864 b_11 NI_11 NS_864 0 7.3270595727917945e-06
GC_11_865 b_11 NI_11 NS_865 0 1.3691622834761276e-05
GC_11_866 b_11 NI_11 NS_866 0 2.6181495018310290e-06
GC_11_867 b_11 NI_11 NS_867 0 4.5508845158866018e-06
GC_11_868 b_11 NI_11 NS_868 0 -1.4312595760624794e-05
GC_11_869 b_11 NI_11 NS_869 0 -5.8920262715116212e-06
GC_11_870 b_11 NI_11 NS_870 0 4.1741001584516349e-06
GC_11_871 b_11 NI_11 NS_871 0 1.0370342810987565e-05
GC_11_872 b_11 NI_11 NS_872 0 9.8155121109596108e-06
GC_11_873 b_11 NI_11 NS_873 0 1.7399291424255534e-05
GC_11_874 b_11 NI_11 NS_874 0 -4.2746525173037201e-06
GC_11_875 b_11 NI_11 NS_875 0 -9.2261099086653355e-06
GC_11_876 b_11 NI_11 NS_876 0 -1.5489849364519141e-05
GC_11_877 b_11 NI_11 NS_877 0 -4.0027571103055507e-06
GC_11_878 b_11 NI_11 NS_878 0 1.3420111671351486e-05
GC_11_879 b_11 NI_11 NS_879 0 2.1008719680714694e-05
GC_11_880 b_11 NI_11 NS_880 0 -7.6339067689859759e-07
GC_11_881 b_11 NI_11 NS_881 0 9.1217865036373384e-06
GC_11_882 b_11 NI_11 NS_882 0 -1.7455397327771109e-05
GC_11_883 b_11 NI_11 NS_883 0 1.4586631433466695e-06
GC_11_884 b_11 NI_11 NS_884 0 -1.4427274352068245e-05
GC_11_885 b_11 NI_11 NS_885 0 -1.3809208253672856e-05
GC_11_886 b_11 NI_11 NS_886 0 3.9887202257562670e-06
GC_11_887 b_11 NI_11 NS_887 0 9.7959541015655244e-09
GC_11_888 b_11 NI_11 NS_888 0 -4.8131127625566654e-08
GC_11_889 b_11 NI_11 NS_889 0 8.6297977547125970e-06
GC_11_890 b_11 NI_11 NS_890 0 1.1373551527385569e-05
GC_11_891 b_11 NI_11 NS_891 0 1.0873479499508927e-05
GC_11_892 b_11 NI_11 NS_892 0 -1.1464240745494702e-05
GC_11_893 b_11 NI_11 NS_893 0 -3.5306961052499688e-06
GC_11_894 b_11 NI_11 NS_894 0 -1.0164963675336544e-05
GC_11_895 b_11 NI_11 NS_895 0 -2.0125069595705539e-06
GC_11_896 b_11 NI_11 NS_896 0 1.2870399607916829e-05
GC_11_897 b_11 NI_11 NS_897 0 9.7605828278171986e-07
GC_11_898 b_11 NI_11 NS_898 0 -7.2620172971093457e-06
GC_11_899 b_11 NI_11 NS_899 0 7.4715757645550915e-06
GC_11_900 b_11 NI_11 NS_900 0 1.7440633904989828e-06
GC_11_901 b_11 NI_11 NS_901 0 -6.1165745399360316e-06
GC_11_902 b_11 NI_11 NS_902 0 -8.8986358089421235e-06
GC_11_903 b_11 NI_11 NS_903 0 -4.1366737079388532e-06
GC_11_904 b_11 NI_11 NS_904 0 9.6569026238196345e-06
GC_11_905 b_11 NI_11 NS_905 0 3.3152442958467304e-06
GC_11_906 b_11 NI_11 NS_906 0 6.0578134918479475e-06
GC_11_907 b_11 NI_11 NS_907 0 5.7049730471468685e-06
GC_11_908 b_11 NI_11 NS_908 0 5.2025363723990840e-07
GC_11_909 b_11 NI_11 NS_909 0 5.9120283220308041e-11
GC_11_910 b_11 NI_11 NS_910 0 1.4784841056498898e-10
GC_11_911 b_11 NI_11 NS_911 0 5.9030599493105053e-09
GC_11_912 b_11 NI_11 NS_912 0 -8.4601872172234582e-09
GC_11_913 b_11 NI_11 NS_913 0 7.7624118557887119e-03
GC_11_914 b_11 NI_11 NS_914 0 -1.6012430130798107e-03
GC_11_915 b_11 NI_11 NS_915 0 -1.2108955808903303e-08
GC_11_916 b_11 NI_11 NS_916 0 -8.8417701864832760e-07
GC_11_917 b_11 NI_11 NS_917 0 1.0417949015757194e-04
GC_11_918 b_11 NI_11 NS_918 0 -5.1169960681450024e-04
GC_11_919 b_11 NI_11 NS_919 0 -1.9362876174670964e-03
GC_11_920 b_11 NI_11 NS_920 0 -5.9765058655115186e-04
GC_11_921 b_11 NI_11 NS_921 0 2.9418170709411273e-03
GC_11_922 b_11 NI_11 NS_922 0 2.2635987277022491e-03
GC_11_923 b_11 NI_11 NS_923 0 -3.5704321000976950e-03
GC_11_924 b_11 NI_11 NS_924 0 -3.0490699932929385e-03
GC_11_925 b_11 NI_11 NS_925 0 -1.7073690282823429e-03
GC_11_926 b_11 NI_11 NS_926 0 5.8427804732014456e-03
GC_11_927 b_11 NI_11 NS_927 0 4.3666880349356842e-03
GC_11_928 b_11 NI_11 NS_928 0 -2.4751072749372850e-03
GC_11_929 b_11 NI_11 NS_929 0 -1.1000736114569339e-04
GC_11_930 b_11 NI_11 NS_930 0 -1.0334111022543572e-04
GC_11_931 b_11 NI_11 NS_931 0 -4.4523080010270364e-03
GC_11_932 b_11 NI_11 NS_932 0 -9.2440216644904460e-04
GC_11_933 b_11 NI_11 NS_933 0 9.1241451991915315e-03
GC_11_934 b_11 NI_11 NS_934 0 1.7784743700107700e-02
GC_11_935 b_11 NI_11 NS_935 0 -4.0272952724844727e-03
GC_11_936 b_11 NI_11 NS_936 0 -1.7846764115832709e-02
GC_11_937 b_11 NI_11 NS_937 0 -8.2177715159461699e-03
GC_11_938 b_11 NI_11 NS_938 0 4.1736031904651850e-03
GC_11_939 b_11 NI_11 NS_939 0 1.7063488480833732e-02
GC_11_940 b_11 NI_11 NS_940 0 -4.3909755959498521e-04
GC_11_941 b_11 NI_11 NS_941 0 -9.2787149378702020e-03
GC_11_942 b_11 NI_11 NS_942 0 -3.2069945232167333e-03
GC_11_943 b_11 NI_11 NS_943 0 -1.3713354902279840e-02
GC_11_944 b_11 NI_11 NS_944 0 2.2836241728451612e-02
GC_11_945 b_11 NI_11 NS_945 0 2.2839545856675605e-02
GC_11_946 b_11 NI_11 NS_946 0 -2.2669178990008618e-02
GC_11_947 b_11 NI_11 NS_947 0 -9.2392853390803487e-03
GC_11_948 b_11 NI_11 NS_948 0 9.0811412226296506e-04
GC_11_949 b_11 NI_11 NS_949 0 1.8480129598972734e-02
GC_11_950 b_11 NI_11 NS_950 0 6.2442194291600110e-03
GC_11_951 b_11 NI_11 NS_951 0 -9.1760825917079590e-03
GC_11_952 b_11 NI_11 NS_952 0 -9.4609771756995857e-03
GC_11_953 b_11 NI_11 NS_953 0 -9.9743257214594799e-03
GC_11_954 b_11 NI_11 NS_954 0 6.3961893660873593e-03
GC_11_955 b_11 NI_11 NS_955 0 1.6838478148083223e-02
GC_11_956 b_11 NI_11 NS_956 0 -4.8501226537060165e-03
GC_11_957 b_11 NI_11 NS_957 0 -7.2149234000141614e-03
GC_11_958 b_11 NI_11 NS_958 0 -3.4092345264253084e-03
GC_11_959 b_11 NI_11 NS_959 0 6.8281951752828607e-03
GC_11_960 b_11 NI_11 NS_960 0 1.3297050871186541e-02
GC_11_961 b_11 NI_11 NS_961 0 -1.8195853055215537e-03
GC_11_962 b_11 NI_11 NS_962 0 -1.4401718425429944e-02
GC_11_963 b_11 NI_11 NS_963 0 -4.9860075666274938e-03
GC_11_964 b_11 NI_11 NS_964 0 1.0394632537669935e-03
GC_11_965 b_11 NI_11 NS_965 0 6.0026082178593421e-03
GC_11_966 b_11 NI_11 NS_966 0 -1.1030577012288558e-03
GC_11_967 b_11 NI_11 NS_967 0 -3.4642738155387172e-03
GC_11_968 b_11 NI_11 NS_968 0 -1.0876296808350985e-03
GC_11_969 b_11 NI_11 NS_969 0 2.7180506512254040e-03
GC_11_970 b_11 NI_11 NS_970 0 -5.0782197071475379e-04
GC_11_971 b_11 NI_11 NS_971 0 -3.2964875840283334e-03
GC_11_972 b_11 NI_11 NS_972 0 -2.8951322147136769e-03
GC_11_973 b_11 NI_11 NS_973 0 2.0159599130031951e-03
GC_11_974 b_11 NI_11 NS_974 0 7.7577878023835122e-04
GC_11_975 b_11 NI_11 NS_975 0 -2.0162769558032213e-03
GC_11_976 b_11 NI_11 NS_976 0 -9.6646490666619654e-04
GC_11_977 b_11 NI_11 NS_977 0 2.1216204026188652e-03
GC_11_978 b_11 NI_11 NS_978 0 -1.4709119213601866e-03
GC_11_979 b_11 NI_11 NS_979 0 -4.1847966358711441e-03
GC_11_980 b_11 NI_11 NS_980 0 -1.8129451333201436e-03
GC_11_981 b_11 NI_11 NS_981 0 2.3697775066024761e-03
GC_11_982 b_11 NI_11 NS_982 0 -3.7075616305148179e-04
GC_11_983 b_11 NI_11 NS_983 0 -3.0172236709726909e-03
GC_11_984 b_11 NI_11 NS_984 0 4.6233814230811664e-04
GC_11_985 b_11 NI_11 NS_985 0 2.7064424611687784e-03
GC_11_986 b_11 NI_11 NS_986 0 -2.7282228980221512e-03
GC_11_987 b_11 NI_11 NS_987 0 -5.0393302507016347e-03
GC_11_988 b_11 NI_11 NS_988 0 -1.2782932411362481e-04
GC_11_989 b_11 NI_11 NS_989 0 2.4346766646909414e-03
GC_11_990 b_11 NI_11 NS_990 0 -2.1719792852885242e-03
GC_11_991 b_11 NI_11 NS_991 0 -3.2449817597152877e-03
GC_11_992 b_11 NI_11 NS_992 0 2.6005317677879267e-03
GC_11_993 b_11 NI_11 NS_993 0 1.7436666478618768e-03
GC_11_994 b_11 NI_11 NS_994 0 -4.7503531473200846e-03
GC_11_995 b_11 NI_11 NS_995 0 -3.6339988945863189e-03
GC_11_996 b_11 NI_11 NS_996 0 2.5967287839450126e-03
GC_11_997 b_11 NI_11 NS_997 0 -2.8319048140698407e-03
GC_11_998 b_11 NI_11 NS_998 0 3.9895731634161588e-03
GC_11_999 b_11 NI_11 NS_999 0 -2.2141478365981122e-04
GC_11_1000 b_11 NI_11 NS_1000 0 -4.2135113287542552e-03
GC_11_1001 b_11 NI_11 NS_1001 0 -9.8957945623950686e-06
GC_11_1002 b_11 NI_11 NS_1002 0 7.5258087893796660e-06
GC_11_1003 b_11 NI_11 NS_1003 0 -1.3539535486911832e-03
GC_11_1004 b_11 NI_11 NS_1004 0 3.3754883304623340e-03
GC_11_1005 b_11 NI_11 NS_1005 0 -9.6985119084135854e-04
GC_11_1006 b_11 NI_11 NS_1006 0 -4.3479509980028520e-03
GC_11_1007 b_11 NI_11 NS_1007 0 -1.0009112717346330e-03
GC_11_1008 b_11 NI_11 NS_1008 0 2.2213051273832054e-03
GC_11_1009 b_11 NI_11 NS_1009 0 -1.6517283917261037e-03
GC_11_1010 b_11 NI_11 NS_1010 0 -4.4093139762028787e-03
GC_11_1011 b_11 NI_11 NS_1011 0 -1.4483159798043181e-03
GC_11_1012 b_11 NI_11 NS_1012 0 -2.4971456887770138e-03
GC_11_1013 b_11 NI_11 NS_1013 0 7.8219595711366942e-04
GC_11_1014 b_11 NI_11 NS_1014 0 2.5933469659691253e-03
GC_11_1015 b_11 NI_11 NS_1015 0 -6.9628533778992650e-04
GC_11_1016 b_11 NI_11 NS_1016 0 2.8792042523857276e-03
GC_11_1017 b_11 NI_11 NS_1017 0 -1.4353705247937556e-03
GC_11_1018 b_11 NI_11 NS_1018 0 -2.7718613469607501e-03
GC_11_1019 b_11 NI_11 NS_1019 0 -1.1678495830825517e-03
GC_11_1020 b_11 NI_11 NS_1020 0 2.6661995998534045e-03
GC_11_1021 b_11 NI_11 NS_1021 0 7.8075940709451891e-04
GC_11_1022 b_11 NI_11 NS_1022 0 -1.8746154576253610e-03
GC_11_1023 b_11 NI_11 NS_1023 0 2.3789744546657182e-08
GC_11_1024 b_11 NI_11 NS_1024 0 -6.0253429559747520e-08
GC_11_1025 b_11 NI_11 NS_1025 0 -9.0373524595352942e-07
GC_11_1026 b_11 NI_11 NS_1026 0 3.2031377343772348e-06
GC_11_1027 b_11 NI_11 NS_1027 0 2.9495688897880549e-03
GC_11_1028 b_11 NI_11 NS_1028 0 -6.1234114299872004e-04
GC_11_1029 b_11 NI_11 NS_1029 0 2.7950027461630188e-08
GC_11_1030 b_11 NI_11 NS_1030 0 -3.1703326955533772e-08
GC_11_1031 b_11 NI_11 NS_1031 0 2.0347235583961215e-04
GC_11_1032 b_11 NI_11 NS_1032 0 1.3799460333053254e-04
GC_11_1033 b_11 NI_11 NS_1033 0 5.6259198714739462e-04
GC_11_1034 b_11 NI_11 NS_1034 0 2.6570831983870627e-04
GC_11_1035 b_11 NI_11 NS_1035 0 3.1064656501059319e-03
GC_11_1036 b_11 NI_11 NS_1036 0 -2.2048908558380933e-03
GC_11_1037 b_11 NI_11 NS_1037 0 -1.5822536236692868e-03
GC_11_1038 b_11 NI_11 NS_1038 0 -2.6870774555434974e-03
GC_11_1039 b_11 NI_11 NS_1039 0 -2.0496561115956697e-03
GC_11_1040 b_11 NI_11 NS_1040 0 -3.7885087032059417e-03
GC_11_1041 b_11 NI_11 NS_1041 0 -4.9745586090373878e-03
GC_11_1042 b_11 NI_11 NS_1042 0 -1.5415288989221938e-03
GC_11_1043 b_11 NI_11 NS_1043 0 2.9290513156797140e-04
GC_11_1044 b_11 NI_11 NS_1044 0 1.9565076647451985e-04
GC_11_1045 b_11 NI_11 NS_1045 0 -2.8663285430045884e-03
GC_11_1046 b_11 NI_11 NS_1046 0 -9.5746355550839393e-04
GC_11_1047 b_11 NI_11 NS_1047 0 -2.2151870424099298e-02
GC_11_1048 b_11 NI_11 NS_1048 0 -1.0226311566058353e-02
GC_11_1049 b_11 NI_11 NS_1049 0 1.1325003492652806e-03
GC_11_1050 b_11 NI_11 NS_1050 0 2.0395318206839867e-02
GC_11_1051 b_11 NI_11 NS_1051 0 -5.8416196347151851e-03
GC_11_1052 b_11 NI_11 NS_1052 0 4.6116300148141918e-03
GC_11_1053 b_11 NI_11 NS_1053 0 5.7171575312122136e-03
GC_11_1054 b_11 NI_11 NS_1054 0 3.4516067845661892e-02
GC_11_1055 b_11 NI_11 NS_1055 0 8.0342764878597855e-03
GC_11_1056 b_11 NI_11 NS_1056 0 2.7930219494437972e-03
GC_11_1057 b_11 NI_11 NS_1057 0 -7.7724143150378873e-03
GC_11_1058 b_11 NI_11 NS_1058 0 2.9556755592449521e-02
GC_11_1059 b_11 NI_11 NS_1059 0 5.0768424324015404e-02
GC_11_1060 b_11 NI_11 NS_1060 0 -2.0072972509441133e-02
GC_11_1061 b_11 NI_11 NS_1061 0 7.9195780475259780e-03
GC_11_1062 b_11 NI_11 NS_1062 0 -1.6364429566542843e-03
GC_11_1063 b_11 NI_11 NS_1063 0 2.9084853593921076e-02
GC_11_1064 b_11 NI_11 NS_1064 0 -2.6464743146716811e-02
GC_11_1065 b_11 NI_11 NS_1065 0 -6.7250700047082838e-03
GC_11_1066 b_11 NI_11 NS_1066 0 -9.8822038426658963e-03
GC_11_1067 b_11 NI_11 NS_1067 0 8.4630804861070604e-03
GC_11_1068 b_11 NI_11 NS_1068 0 -8.0278000634926416e-03
GC_11_1069 b_11 NI_11 NS_1069 0 -1.8994957697072844e-02
GC_11_1070 b_11 NI_11 NS_1070 0 -2.5238416803829797e-02
GC_11_1071 b_11 NI_11 NS_1071 0 -5.4717854479283583e-03
GC_11_1072 b_11 NI_11 NS_1072 0 -2.8547826196595695e-03
GC_11_1073 b_11 NI_11 NS_1073 0 -1.7741075714951728e-02
GC_11_1074 b_11 NI_11 NS_1074 0 -1.3132225703460614e-02
GC_11_1075 b_11 NI_11 NS_1075 0 -4.8177975522807337e-03
GC_11_1076 b_11 NI_11 NS_1076 0 1.2541404159100567e-02
GC_11_1077 b_11 NI_11 NS_1077 0 -3.4590894860970500e-03
GC_11_1078 b_11 NI_11 NS_1078 0 1.5412388346450210e-03
GC_11_1079 b_11 NI_11 NS_1079 0 -7.1864998745200734e-04
GC_11_1080 b_11 NI_11 NS_1080 0 7.0058601123304046e-03
GC_11_1081 b_11 NI_11 NS_1081 0 1.8820413603393414e-03
GC_11_1082 b_11 NI_11 NS_1082 0 8.5748073651130801e-05
GC_11_1083 b_11 NI_11 NS_1083 0 3.1400244222160609e-04
GC_11_1084 b_11 NI_11 NS_1084 0 -1.9467015672588891e-03
GC_11_1085 b_11 NI_11 NS_1085 0 -1.8563355820308892e-03
GC_11_1086 b_11 NI_11 NS_1086 0 -1.6182085843550256e-03
GC_11_1087 b_11 NI_11 NS_1087 0 -2.1290959190495063e-03
GC_11_1088 b_11 NI_11 NS_1088 0 1.6850436298704388e-03
GC_11_1089 b_11 NI_11 NS_1089 0 7.6361044220855608e-04
GC_11_1090 b_11 NI_11 NS_1090 0 1.8527504704870620e-04
GC_11_1091 b_11 NI_11 NS_1091 0 -6.9730375377938562e-04
GC_11_1092 b_11 NI_11 NS_1092 0 -1.6780701256937950e-03
GC_11_1093 b_11 NI_11 NS_1093 0 -2.6815284605536459e-03
GC_11_1094 b_11 NI_11 NS_1094 0 -8.2749108293081214e-04
GC_11_1095 b_11 NI_11 NS_1095 0 -4.9989634712239387e-04
GC_11_1096 b_11 NI_11 NS_1096 0 2.9288644974138152e-03
GC_11_1097 b_11 NI_11 NS_1097 0 1.3533577525682077e-03
GC_11_1098 b_11 NI_11 NS_1098 0 -8.5805582310373083e-04
GC_11_1099 b_11 NI_11 NS_1099 0 -2.4189245251177559e-03
GC_11_1100 b_11 NI_11 NS_1100 0 -2.2676209007467321e-03
GC_11_1101 b_11 NI_11 NS_1101 0 -3.5540455455156249e-03
GC_11_1102 b_11 NI_11 NS_1102 0 7.4852709191338329e-04
GC_11_1103 b_11 NI_11 NS_1103 0 2.4633836864989605e-03
GC_11_1104 b_11 NI_11 NS_1104 0 3.0182802279719451e-03
GC_11_1105 b_11 NI_11 NS_1105 0 9.8455436592599231e-04
GC_11_1106 b_11 NI_11 NS_1106 0 -2.9418099057198777e-03
GC_11_1107 b_11 NI_11 NS_1107 0 -4.7677997716361834e-03
GC_11_1108 b_11 NI_11 NS_1108 0 5.4340106908619244e-05
GC_11_1109 b_11 NI_11 NS_1109 0 -1.7083702421896248e-03
GC_11_1110 b_11 NI_11 NS_1110 0 3.7124268513342882e-03
GC_11_1111 b_11 NI_11 NS_1111 0 -7.6587333777938587e-04
GC_11_1112 b_11 NI_11 NS_1112 0 1.5006762460863762e-03
GC_11_1113 b_11 NI_11 NS_1113 0 3.2213013307031174e-03
GC_11_1114 b_11 NI_11 NS_1114 0 -1.3508681933053289e-03
GC_11_1115 b_11 NI_11 NS_1115 0 -2.9326147319160507e-06
GC_11_1116 b_11 NI_11 NS_1116 0 8.7469999201409861e-06
GC_11_1117 b_11 NI_11 NS_1117 0 -1.8200418480663822e-03
GC_11_1118 b_11 NI_11 NS_1118 0 -2.5277357131666071e-03
GC_11_1119 b_11 NI_11 NS_1119 0 -2.4072528515181068e-03
GC_11_1120 b_11 NI_11 NS_1120 0 2.4886639017697746e-03
GC_11_1121 b_11 NI_11 NS_1121 0 1.0142614252845108e-03
GC_11_1122 b_11 NI_11 NS_1122 0 2.4256822809683048e-03
GC_11_1123 b_11 NI_11 NS_1123 0 8.5775954933653062e-04
GC_11_1124 b_11 NI_11 NS_1124 0 -2.6994833951142386e-03
GC_11_1125 b_11 NI_11 NS_1125 0 -3.0644805107856430e-04
GC_11_1126 b_11 NI_11 NS_1126 0 1.6741356131013108e-03
GC_11_1127 b_11 NI_11 NS_1127 0 -1.7840544963941686e-03
GC_11_1128 b_11 NI_11 NS_1128 0 -3.1181085817973044e-04
GC_11_1129 b_11 NI_11 NS_1129 0 1.4004539851165234e-03
GC_11_1130 b_11 NI_11 NS_1130 0 1.9709614214838472e-03
GC_11_1131 b_11 NI_11 NS_1131 0 1.0449286310742108e-03
GC_11_1132 b_11 NI_11 NS_1132 0 -2.2998046594622113e-03
GC_11_1133 b_11 NI_11 NS_1133 0 -6.9799493710965025e-04
GC_11_1134 b_11 NI_11 NS_1134 0 -1.4668899050094522e-03
GC_11_1135 b_11 NI_11 NS_1135 0 -1.3735490844138513e-03
GC_11_1136 b_11 NI_11 NS_1136 0 -3.1252861358753171e-04
GC_11_1137 b_11 NI_11 NS_1137 0 7.1030485756397359e-09
GC_11_1138 b_11 NI_11 NS_1138 0 -2.4709970475652812e-08
GC_11_1139 b_11 NI_11 NS_1139 0 -4.5275603084989712e-07
GC_11_1140 b_11 NI_11 NS_1140 0 1.6341839314124877e-06
GC_11_1141 b_11 NI_11 NS_1141 0 -1.3077626181950885e-02
GC_11_1142 b_11 NI_11 NS_1142 0 1.3851822870423515e-03
GC_11_1143 b_11 NI_11 NS_1143 0 -2.6206484157238706e-07
GC_11_1144 b_11 NI_11 NS_1144 0 -3.7495559724260546e-06
GC_11_1145 b_11 NI_11 NS_1145 0 -2.7819372045824914e-04
GC_11_1146 b_11 NI_11 NS_1146 0 4.6297784968867738e-04
GC_11_1147 b_11 NI_11 NS_1147 0 1.3195321554402711e-03
GC_11_1148 b_11 NI_11 NS_1148 0 5.4935775116451394e-04
GC_11_1149 b_11 NI_11 NS_1149 0 -2.7628705965086300e-03
GC_11_1150 b_11 NI_11 NS_1150 0 -8.1703054050131401e-04
GC_11_1151 b_11 NI_11 NS_1151 0 3.5326192481361838e-03
GC_11_1152 b_11 NI_11 NS_1152 0 2.5338002367322602e-03
GC_11_1153 b_11 NI_11 NS_1153 0 1.1824232660161524e-03
GC_11_1154 b_11 NI_11 NS_1154 0 -4.1997922523624035e-03
GC_11_1155 b_11 NI_11 NS_1155 0 -1.7498503089831820e-03
GC_11_1156 b_11 NI_11 NS_1156 0 2.6968800977728710e-03
GC_11_1157 b_11 NI_11 NS_1157 0 -3.1387333304585592e-04
GC_11_1158 b_11 NI_11 NS_1158 0 -1.8984121393569484e-04
GC_11_1159 b_11 NI_11 NS_1159 0 3.9674889269260601e-03
GC_11_1160 b_11 NI_11 NS_1160 0 2.9857839207260379e-04
GC_11_1161 b_11 NI_11 NS_1161 0 -7.4413975684285176e-03
GC_11_1162 b_11 NI_11 NS_1162 0 -1.3618339017549776e-02
GC_11_1163 b_11 NI_11 NS_1163 0 4.4052505494701875e-03
GC_11_1164 b_11 NI_11 NS_1164 0 1.3511458829104445e-02
GC_11_1165 b_11 NI_11 NS_1165 0 6.7110109769434583e-03
GC_11_1166 b_11 NI_11 NS_1166 0 -3.9862631677579554e-03
GC_11_1167 b_11 NI_11 NS_1167 0 -1.3390055117710379e-02
GC_11_1168 b_11 NI_11 NS_1168 0 6.9024316026117466e-04
GC_11_1169 b_11 NI_11 NS_1169 0 7.8426044093509173e-03
GC_11_1170 b_11 NI_11 NS_1170 0 1.8947671797552503e-03
GC_11_1171 b_11 NI_11 NS_1171 0 1.0544112092795136e-02
GC_11_1172 b_11 NI_11 NS_1172 0 -1.9595447135794183e-02
GC_11_1173 b_11 NI_11 NS_1173 0 -1.7809609065537191e-02
GC_11_1174 b_11 NI_11 NS_1174 0 1.9141982245256314e-02
GC_11_1175 b_11 NI_11 NS_1175 0 7.6787750431322700e-03
GC_11_1176 b_11 NI_11 NS_1176 0 -1.4142909528423082e-03
GC_11_1177 b_11 NI_11 NS_1177 0 -1.5647914336480228e-02
GC_11_1178 b_11 NI_11 NS_1178 0 -4.7614896901247107e-03
GC_11_1179 b_11 NI_11 NS_1179 0 8.0618573016896389e-03
GC_11_1180 b_11 NI_11 NS_1180 0 7.2869891809915341e-03
GC_11_1181 b_11 NI_11 NS_1181 0 8.1170047185718189e-03
GC_11_1182 b_11 NI_11 NS_1182 0 -5.9990832035982430e-03
GC_11_1183 b_11 NI_11 NS_1183 0 -1.3980586997120653e-02
GC_11_1184 b_11 NI_11 NS_1184 0 4.5682719333453607e-03
GC_11_1185 b_11 NI_11 NS_1185 0 6.2307820113007249e-03
GC_11_1186 b_11 NI_11 NS_1186 0 2.4081612519185531e-03
GC_11_1187 b_11 NI_11 NS_1187 0 -6.2859264355150614e-03
GC_11_1188 b_11 NI_11 NS_1188 0 -1.1107051557285624e-02
GC_11_1189 b_11 NI_11 NS_1189 0 2.1280730573089665e-03
GC_11_1190 b_11 NI_11 NS_1190 0 1.1947397205329082e-02
GC_11_1191 b_11 NI_11 NS_1191 0 4.2092178851988581e-03
GC_11_1192 b_11 NI_11 NS_1192 0 -1.1609522005070299e-03
GC_11_1193 b_11 NI_11 NS_1193 0 -4.9313045763678494e-03
GC_11_1194 b_11 NI_11 NS_1194 0 1.0532438103220839e-03
GC_11_1195 b_11 NI_11 NS_1195 0 3.0238807200197327e-03
GC_11_1196 b_11 NI_11 NS_1196 0 6.9985711643237374e-04
GC_11_1197 b_11 NI_11 NS_1197 0 -2.2205262517192834e-03
GC_11_1198 b_11 NI_11 NS_1198 0 4.9428581137972601e-04
GC_11_1199 b_11 NI_11 NS_1199 0 3.0655102801236587e-03
GC_11_1200 b_11 NI_11 NS_1200 0 2.3037302634439836e-03
GC_11_1201 b_11 NI_11 NS_1201 0 -1.5339091967097984e-03
GC_11_1202 b_11 NI_11 NS_1202 0 -6.6977447033582458e-04
GC_11_1203 b_11 NI_11 NS_1203 0 1.8873378600738927e-03
GC_11_1204 b_11 NI_11 NS_1204 0 6.8441649659159443e-04
GC_11_1205 b_11 NI_11 NS_1205 0 -1.5620993801149304e-03
GC_11_1206 b_11 NI_11 NS_1206 0 1.2263492645297222e-03
GC_11_1207 b_11 NI_11 NS_1207 0 3.9751893811776967e-03
GC_11_1208 b_11 NI_11 NS_1208 0 1.4060884820820531e-03
GC_11_1209 b_11 NI_11 NS_1209 0 -1.5528106206009961e-03
GC_11_1210 b_11 NI_11 NS_1210 0 7.4661566659931457e-05
GC_11_1211 b_11 NI_11 NS_1211 0 2.8290380091206152e-03
GC_11_1212 b_11 NI_11 NS_1212 0 -6.8616923824458013e-04
GC_11_1213 b_11 NI_11 NS_1213 0 -1.8781833910554364e-03
GC_11_1214 b_11 NI_11 NS_1214 0 2.0100728806594689e-03
GC_11_1215 b_11 NI_11 NS_1215 0 4.9079320153824473e-03
GC_11_1216 b_11 NI_11 NS_1216 0 -1.8215321236843656e-04
GC_11_1217 b_11 NI_11 NS_1217 0 -1.6564588825827961e-03
GC_11_1218 b_11 NI_11 NS_1218 0 9.3019323073935596e-04
GC_11_1219 b_11 NI_11 NS_1219 0 3.0643003907121565e-03
GC_11_1220 b_11 NI_11 NS_1220 0 -2.8465101716213131e-03
GC_11_1221 b_11 NI_11 NS_1221 0 -1.4568553769444580e-03
GC_11_1222 b_11 NI_11 NS_1222 0 3.2233613952251808e-03
GC_11_1223 b_11 NI_11 NS_1223 0 3.8009920814151246e-03
GC_11_1224 b_11 NI_11 NS_1224 0 -2.9784186698552191e-03
GC_11_1225 b_11 NI_11 NS_1225 0 -1.8786582710828927e-03
GC_11_1226 b_11 NI_11 NS_1226 0 -3.8879556392316869e-03
GC_11_1227 b_11 NI_11 NS_1227 0 -4.0379406914628393e-04
GC_11_1228 b_11 NI_11 NS_1228 0 2.3675280190566341e-03
GC_11_1229 b_11 NI_11 NS_1229 0 -1.0556590125632033e-05
GC_11_1230 b_11 NI_11 NS_1230 0 -2.1452520938685761e-05
GC_11_1231 b_11 NI_11 NS_1231 0 8.4230055209683378e-04
GC_11_1232 b_11 NI_11 NS_1232 0 -3.7965136864239009e-03
GC_11_1233 b_11 NI_11 NS_1233 0 3.4279644062311132e-04
GC_11_1234 b_11 NI_11 NS_1234 0 3.3487743163436554e-03
GC_11_1235 b_11 NI_11 NS_1235 0 1.3577034085074490e-03
GC_11_1236 b_11 NI_11 NS_1236 0 -2.3752403677718267e-03
GC_11_1237 b_11 NI_11 NS_1237 0 2.1858930129685485e-03
GC_11_1238 b_11 NI_11 NS_1238 0 3.3360532781765888e-03
GC_11_1239 b_11 NI_11 NS_1239 0 1.1689674476250656e-03
GC_11_1240 b_11 NI_11 NS_1240 0 2.4033191298493536e-03
GC_11_1241 b_11 NI_11 NS_1241 0 -8.1092511614918867e-04
GC_11_1242 b_11 NI_11 NS_1242 0 -1.9781530790467612e-03
GC_11_1243 b_11 NI_11 NS_1243 0 3.9749601063585933e-04
GC_11_1244 b_11 NI_11 NS_1244 0 -2.6833654762312108e-03
GC_11_1245 b_11 NI_11 NS_1245 0 9.8234543226962475e-04
GC_11_1246 b_11 NI_11 NS_1246 0 2.7459675674614795e-03
GC_11_1247 b_11 NI_11 NS_1247 0 1.0390538027585377e-03
GC_11_1248 b_11 NI_11 NS_1248 0 -2.4207682785439043e-03
GC_11_1249 b_11 NI_11 NS_1249 0 -1.0837509675524512e-03
GC_11_1250 b_11 NI_11 NS_1250 0 1.5920956231316975e-03
GC_11_1251 b_11 NI_11 NS_1251 0 -1.1067035140379793e-08
GC_11_1252 b_11 NI_11 NS_1252 0 -2.8126814937096164e-09
GC_11_1253 b_11 NI_11 NS_1253 0 2.2672981072121503e-06
GC_11_1254 b_11 NI_11 NS_1254 0 5.3151740922522633e-07
GC_11_1255 b_11 NI_11 NS_1255 0 1.8226558401297190e-02
GC_11_1256 b_11 NI_11 NS_1256 0 6.7518773451198215e-03
GC_11_1257 b_11 NI_11 NS_1257 0 4.8241140797484367e-07
GC_11_1258 b_11 NI_11 NS_1258 0 1.4304303894833612e-06
GC_11_1259 b_11 NI_11 NS_1259 0 6.0825153122807882e-03
GC_11_1260 b_11 NI_11 NS_1260 0 1.8254957225330652e-03
GC_11_1261 b_11 NI_11 NS_1261 0 -6.0662904926585045e-03
GC_11_1262 b_11 NI_11 NS_1262 0 -6.4127966387047077e-04
GC_11_1263 b_11 NI_11 NS_1263 0 7.3353747880288249e-03
GC_11_1264 b_11 NI_11 NS_1264 0 -1.2858474181208107e-02
GC_11_1265 b_11 NI_11 NS_1265 0 8.4354447291468421e-03
GC_11_1266 b_11 NI_11 NS_1266 0 -2.1170041271973390e-04
GC_11_1267 b_11 NI_11 NS_1267 0 -9.6680461703341821e-03
GC_11_1268 b_11 NI_11 NS_1268 0 2.5853122431647967e-03
GC_11_1269 b_11 NI_11 NS_1269 0 -8.8082179864397911e-03
GC_11_1270 b_11 NI_11 NS_1270 0 -2.4395000016513874e-02
GC_11_1271 b_11 NI_11 NS_1271 0 -8.6843598488188392e-04
GC_11_1272 b_11 NI_11 NS_1272 0 4.1759356243908797e-03
GC_11_1273 b_11 NI_11 NS_1273 0 7.1854221032982323e-03
GC_11_1274 b_11 NI_11 NS_1274 0 -9.9748569418021439e-04
GC_11_1275 b_11 NI_11 NS_1275 0 -2.5220085129980668e-02
GC_11_1276 b_11 NI_11 NS_1276 0 4.8140848744996434e-03
GC_11_1277 b_11 NI_11 NS_1277 0 -1.9618495641927663e-02
GC_11_1278 b_11 NI_11 NS_1278 0 8.5380894792422973e-04
GC_11_1279 b_11 NI_11 NS_1279 0 1.0773060773795574e-02
GC_11_1280 b_11 NI_11 NS_1280 0 -2.7350673782021002e-03
GC_11_1281 b_11 NI_11 NS_1281 0 -4.8271290233661886e-03
GC_11_1282 b_11 NI_11 NS_1282 0 4.5019621963325394e-02
GC_11_1283 b_11 NI_11 NS_1283 0 -1.2641866883878727e-02
GC_11_1284 b_11 NI_11 NS_1284 0 -3.2181979212595347e-04
GC_11_1285 b_11 NI_11 NS_1285 0 1.5975197581399155e-02
GC_11_1286 b_11 NI_11 NS_1286 0 -3.9759623685589329e-03
GC_11_1287 b_11 NI_11 NS_1287 0 3.2145941912160102e-02
GC_11_1288 b_11 NI_11 NS_1288 0 1.8555419449381796e-02
GC_11_1289 b_11 NI_11 NS_1289 0 -1.2594989808622498e-02
GC_11_1290 b_11 NI_11 NS_1290 0 1.1571471500205085e-04
GC_11_1291 b_11 NI_11 NS_1291 0 1.7251913665928761e-02
GC_11_1292 b_11 NI_11 NS_1292 0 -3.5175767581701212e-02
GC_11_1293 b_11 NI_11 NS_1293 0 1.3984048379077270e-02
GC_11_1294 b_11 NI_11 NS_1294 0 4.8235533570249144e-03
GC_11_1295 b_11 NI_11 NS_1295 0 -1.4410969266873453e-02
GC_11_1296 b_11 NI_11 NS_1296 0 1.9247495865411387e-04
GC_11_1297 b_11 NI_11 NS_1297 0 -2.0124126275040229e-02
GC_11_1298 b_11 NI_11 NS_1298 0 -3.0196846984724343e-02
GC_11_1299 b_11 NI_11 NS_1299 0 1.0516061918837586e-02
GC_11_1300 b_11 NI_11 NS_1300 0 3.6210539818726881e-03
GC_11_1301 b_11 NI_11 NS_1301 0 -2.6839350445827293e-02
GC_11_1302 b_11 NI_11 NS_1302 0 1.1127553613557604e-02
GC_11_1303 b_11 NI_11 NS_1303 0 -1.4106800383209906e-02
GC_11_1304 b_11 NI_11 NS_1304 0 -2.5292621507084462e-03
GC_11_1305 b_11 NI_11 NS_1305 0 7.5511305299930612e-03
GC_11_1306 b_11 NI_11 NS_1306 0 1.6110865726161215e-03
GC_11_1307 b_11 NI_11 NS_1307 0 -8.7781419241282719e-04
GC_11_1308 b_11 NI_11 NS_1308 0 2.4406549452682433e-02
GC_11_1309 b_11 NI_11 NS_1309 0 -7.6159445781354531e-03
GC_11_1310 b_11 NI_11 NS_1310 0 2.7283454542378612e-04
GC_11_1311 b_11 NI_11 NS_1311 0 -5.5397169072155623e-04
GC_11_1312 b_11 NI_11 NS_1312 0 -5.5347197021903844e-03
GC_11_1313 b_11 NI_11 NS_1313 0 8.2549158338449790e-03
GC_11_1314 b_11 NI_11 NS_1314 0 7.0292097422187403e-03
GC_11_1315 b_11 NI_11 NS_1315 0 -7.2657245690646187e-04
GC_11_1316 b_11 NI_11 NS_1316 0 1.2096327849002482e-02
GC_11_1317 b_11 NI_11 NS_1317 0 -5.1449872370469786e-03
GC_11_1318 b_11 NI_11 NS_1318 0 -1.3732679561072187e-04
GC_11_1319 b_11 NI_11 NS_1319 0 -1.8277731745325332e-03
GC_11_1320 b_11 NI_11 NS_1320 0 -5.1663196047603121e-03
GC_11_1321 b_11 NI_11 NS_1321 0 9.2805746883016117e-03
GC_11_1322 b_11 NI_11 NS_1322 0 5.4202571546288787e-03
GC_11_1323 b_11 NI_11 NS_1323 0 3.5140269664283310e-03
GC_11_1324 b_11 NI_11 NS_1324 0 1.1697048665664149e-02
GC_11_1325 b_11 NI_11 NS_1325 0 -6.1352117495547384e-03
GC_11_1326 b_11 NI_11 NS_1326 0 1.4323536018075889e-03
GC_11_1327 b_11 NI_11 NS_1327 0 -2.8179114132830256e-03
GC_11_1328 b_11 NI_11 NS_1328 0 -7.3385865112807237e-03
GC_11_1329 b_11 NI_11 NS_1329 0 9.9490953820989721e-03
GC_11_1330 b_11 NI_11 NS_1330 0 3.3702689893436045e-03
GC_11_1331 b_11 NI_11 NS_1331 0 8.1728141361503068e-03
GC_11_1332 b_11 NI_11 NS_1332 0 1.0256566116436645e-02
GC_11_1333 b_11 NI_11 NS_1333 0 -6.9843294494699639e-03
GC_11_1334 b_11 NI_11 NS_1334 0 2.9456481549008325e-03
GC_11_1335 b_11 NI_11 NS_1335 0 -5.6338028865628616e-03
GC_11_1336 b_11 NI_11 NS_1336 0 -8.0802574913391989e-03
GC_11_1337 b_11 NI_11 NS_1337 0 9.8429423872190922e-03
GC_11_1338 b_11 NI_11 NS_1338 0 5.5983489821727860e-04
GC_11_1339 b_11 NI_11 NS_1339 0 -1.0787139007492863e-02
GC_11_1340 b_11 NI_11 NS_1340 0 1.2188746257468656e-02
GC_11_1341 b_11 NI_11 NS_1341 0 9.6751304237299440e-03
GC_11_1342 b_11 NI_11 NS_1342 0 5.0628524765796903e-03
GC_11_1343 b_11 NI_11 NS_1343 0 -1.9007150021624534e-05
GC_11_1344 b_11 NI_11 NS_1344 0 3.1757118551863463e-05
GC_11_1345 b_11 NI_11 NS_1345 0 -7.1154983497078647e-03
GC_11_1346 b_11 NI_11 NS_1346 0 4.4968633763016689e-03
GC_11_1347 b_11 NI_11 NS_1347 0 -7.6588015262057541e-03
GC_11_1348 b_11 NI_11 NS_1348 0 -5.3140585001085917e-03
GC_11_1349 b_11 NI_11 NS_1349 0 9.4988888941623766e-03
GC_11_1350 b_11 NI_11 NS_1350 0 -1.7110127975792590e-03
GC_11_1351 b_11 NI_11 NS_1351 0 1.2462819698046393e-02
GC_11_1352 b_11 NI_11 NS_1352 0 -1.3552953196774280e-03
GC_11_1353 b_11 NI_11 NS_1353 0 -5.0734355575875389e-03
GC_11_1354 b_11 NI_11 NS_1354 0 -2.7550310988677519e-03
GC_11_1355 b_11 NI_11 NS_1355 0 -2.2334790621585114e-03
GC_11_1356 b_11 NI_11 NS_1356 0 6.5927069523012329e-03
GC_11_1357 b_11 NI_11 NS_1357 0 8.9637858333551507e-03
GC_11_1358 b_11 NI_11 NS_1358 0 1.2891576707251744e-04
GC_11_1359 b_11 NI_11 NS_1359 0 1.2489969491654530e-02
GC_11_1360 b_11 NI_11 NS_1360 0 1.7707492273427885e-03
GC_11_1361 b_11 NI_11 NS_1361 0 -5.3740565164713972e-03
GC_11_1362 b_11 NI_11 NS_1362 0 4.1561446469687022e-03
GC_11_1363 b_11 NI_11 NS_1363 0 -1.8426485698956646e-03
GC_11_1364 b_11 NI_11 NS_1364 0 -5.6872682784694407e-03
GC_11_1365 b_11 NI_11 NS_1365 0 2.0880735207101956e-07
GC_11_1366 b_11 NI_11 NS_1366 0 -2.4392496418157611e-07
GC_11_1367 b_11 NI_11 NS_1367 0 -1.1440672520200850e-05
GC_11_1368 b_11 NI_11 NS_1368 0 1.8294492803427793e-05
GD_11_1 b_11 NI_11 NA_1 0 -6.4862660429223661e-07
GD_11_2 b_11 NI_11 NA_2 0 3.5859774240729921e-06
GD_11_3 b_11 NI_11 NA_3 0 -1.8573497842381583e-06
GD_11_4 b_11 NI_11 NA_4 0 5.6258474695865988e-06
GD_11_5 b_11 NI_11 NA_5 0 -6.7028356362235435e-06
GD_11_6 b_11 NI_11 NA_6 0 1.0203937741638903e-05
GD_11_7 b_11 NI_11 NA_7 0 4.1424654069122602e-06
GD_11_8 b_11 NI_11 NA_8 0 2.4546235260497769e-06
GD_11_9 b_11 NI_11 NA_9 0 1.3004900789018385e-02
GD_11_10 b_11 NI_11 NA_10 0 5.9084237279017227e-04
GD_11_11 b_11 NI_11 NA_11 0 -8.8592637656549431e-03
GD_11_12 b_11 NI_11 NA_12 0 -4.2259745752110259e-03
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -1.2624340515034760e-05
GC_12_2 b_12 NI_12 NS_2 0 1.6605298164753227e-08
GC_12_3 b_12 NI_12 NS_3 0 2.1156744655284066e-11
GC_12_4 b_12 NI_12 NS_4 0 -3.0722497214500394e-10
GC_12_5 b_12 NI_12 NS_5 0 -3.4970559251814183e-07
GC_12_6 b_12 NI_12 NS_6 0 -9.9914998952592473e-07
GC_12_7 b_12 NI_12 NS_7 0 -9.3464152611640296e-07
GC_12_8 b_12 NI_12 NS_8 0 1.7814213161160438e-06
GC_12_9 b_12 NI_12 NS_9 0 -3.3141591559097762e-06
GC_12_10 b_12 NI_12 NS_10 0 8.1245933087178972e-07
GC_12_11 b_12 NI_12 NS_11 0 9.4712163415693670e-07
GC_12_12 b_12 NI_12 NS_12 0 -2.3716147598292826e-07
GC_12_13 b_12 NI_12 NS_13 0 5.4159331040102278e-07
GC_12_14 b_12 NI_12 NS_14 0 4.5114370859113298e-06
GC_12_15 b_12 NI_12 NS_15 0 1.6161413147413057e-06
GC_12_16 b_12 NI_12 NS_16 0 3.0361310842891111e-06
GC_12_17 b_12 NI_12 NS_17 0 -8.7112003293702495e-07
GC_12_18 b_12 NI_12 NS_18 0 -5.9629327801701094e-07
GC_12_19 b_12 NI_12 NS_19 0 4.7104111891186193e-07
GC_12_20 b_12 NI_12 NS_20 0 -1.1590526278300133e-06
GC_12_21 b_12 NI_12 NS_21 0 2.8710438724336843e-06
GC_12_22 b_12 NI_12 NS_22 0 1.0312478226154637e-05
GC_12_23 b_12 NI_12 NS_23 0 4.5202360662808911e-06
GC_12_24 b_12 NI_12 NS_24 0 -7.5372083274458585e-07
GC_12_25 b_12 NI_12 NS_25 0 1.6526199944217339e-06
GC_12_26 b_12 NI_12 NS_26 0 -4.2690992482837990e-07
GC_12_27 b_12 NI_12 NS_27 0 1.6702708176962984e-05
GC_12_28 b_12 NI_12 NS_28 0 -4.4193887237214928e-06
GC_12_29 b_12 NI_12 NS_29 0 2.2260080325251955e-07
GC_12_30 b_12 NI_12 NS_30 0 -1.0410954221381860e-06
GC_12_31 b_12 NI_12 NS_31 0 9.3453502361590692e-06
GC_12_32 b_12 NI_12 NS_32 0 -7.1208014985314854e-07
GC_12_33 b_12 NI_12 NS_33 0 -5.5720409880366869e-06
GC_12_34 b_12 NI_12 NS_34 0 -1.9745304730738119e-05
GC_12_35 b_12 NI_12 NS_35 0 -6.0170130319256210e-07
GC_12_36 b_12 NI_12 NS_36 0 -8.9886625381265841e-07
GC_12_37 b_12 NI_12 NS_37 0 -1.1426761427643588e-05
GC_12_38 b_12 NI_12 NS_38 0 -1.0985921469464177e-05
GC_12_39 b_12 NI_12 NS_39 0 -2.2538842410777954e-06
GC_12_40 b_12 NI_12 NS_40 0 2.5922622444926245e-07
GC_12_41 b_12 NI_12 NS_41 0 -1.9214958712212896e-06
GC_12_42 b_12 NI_12 NS_42 0 -7.8162590226550682e-07
GC_12_43 b_12 NI_12 NS_43 0 -9.6669570049279494e-06
GC_12_44 b_12 NI_12 NS_44 0 5.8218582463314292e-06
GC_12_45 b_12 NI_12 NS_45 0 -2.9986996297857565e-07
GC_12_46 b_12 NI_12 NS_46 0 1.6066143391827670e-07
GC_12_47 b_12 NI_12 NS_47 0 -1.6024803967812621e-06
GC_12_48 b_12 NI_12 NS_48 0 5.7938341105299180e-06
GC_12_49 b_12 NI_12 NS_49 0 2.0440931139334887e-06
GC_12_50 b_12 NI_12 NS_50 0 1.9749667856009079e-06
GC_12_51 b_12 NI_12 NS_51 0 6.0777009188761986e-07
GC_12_52 b_12 NI_12 NS_52 0 -8.9639263698381167e-08
GC_12_53 b_12 NI_12 NS_53 0 3.3231646491471137e-06
GC_12_54 b_12 NI_12 NS_54 0 -4.3001152157148866e-07
GC_12_55 b_12 NI_12 NS_55 0 -5.2000556646678111e-08
GC_12_56 b_12 NI_12 NS_56 0 3.3451710249961541e-08
GC_12_57 b_12 NI_12 NS_57 0 -8.0680171053655832e-07
GC_12_58 b_12 NI_12 NS_58 0 -2.3790065592334585e-07
GC_12_59 b_12 NI_12 NS_59 0 3.8123046276251326e-07
GC_12_60 b_12 NI_12 NS_60 0 -5.1760902101189238e-07
GC_12_61 b_12 NI_12 NS_61 0 1.1837454510122792e-06
GC_12_62 b_12 NI_12 NS_62 0 -3.2959258987373482e-08
GC_12_63 b_12 NI_12 NS_63 0 2.3780673196600600e-08
GC_12_64 b_12 NI_12 NS_64 0 4.9143002011366758e-08
GC_12_65 b_12 NI_12 NS_65 0 -5.6742679910438302e-07
GC_12_66 b_12 NI_12 NS_66 0 -5.4636882874839765e-08
GC_12_67 b_12 NI_12 NS_67 0 4.9448371152764963e-07
GC_12_68 b_12 NI_12 NS_68 0 -5.0932303950330165e-07
GC_12_69 b_12 NI_12 NS_69 0 1.1632167981662096e-06
GC_12_70 b_12 NI_12 NS_70 0 -6.8919840760112292e-07
GC_12_71 b_12 NI_12 NS_71 0 5.6825116871929705e-08
GC_12_72 b_12 NI_12 NS_72 0 3.5514385144880148e-11
GC_12_73 b_12 NI_12 NS_73 0 -5.7560497138160219e-07
GC_12_74 b_12 NI_12 NS_74 0 -6.5638144749678529e-08
GC_12_75 b_12 NI_12 NS_75 0 6.3212351580200766e-07
GC_12_76 b_12 NI_12 NS_76 0 -5.0035596231341207e-07
GC_12_77 b_12 NI_12 NS_77 0 8.4892138387681240e-07
GC_12_78 b_12 NI_12 NS_78 0 -1.3993923777121608e-06
GC_12_79 b_12 NI_12 NS_79 0 1.0856894176998518e-07
GC_12_80 b_12 NI_12 NS_80 0 -6.0252879171408315e-08
GC_12_81 b_12 NI_12 NS_81 0 -3.9935318736630618e-07
GC_12_82 b_12 NI_12 NS_82 0 -2.0554230569360452e-07
GC_12_83 b_12 NI_12 NS_83 0 1.1352911656178605e-06
GC_12_84 b_12 NI_12 NS_84 0 -8.8116538504994555e-07
GC_12_85 b_12 NI_12 NS_85 0 -4.1532476552210630e-06
GC_12_86 b_12 NI_12 NS_86 0 6.0162328407520717e-07
GC_12_87 b_12 NI_12 NS_87 0 -5.6369200513792926e-07
GC_12_88 b_12 NI_12 NS_88 0 -1.9351435846743098e-06
GC_12_89 b_12 NI_12 NS_89 0 -2.9200099305289900e-08
GC_12_90 b_12 NI_12 NS_90 0 -9.6976909657027651e-09
GC_12_91 b_12 NI_12 NS_91 0 -3.5883311761571637e-07
GC_12_92 b_12 NI_12 NS_92 0 -2.9257646436666423e-07
GC_12_93 b_12 NI_12 NS_93 0 -4.7734141564159216e-07
GC_12_94 b_12 NI_12 NS_94 0 -1.7399214149755265e-07
GC_12_95 b_12 NI_12 NS_95 0 8.5953338110574397e-07
GC_12_96 b_12 NI_12 NS_96 0 -7.5679188976681852e-07
GC_12_97 b_12 NI_12 NS_97 0 6.0934547863968378e-07
GC_12_98 b_12 NI_12 NS_98 0 -1.0781605902458984e-06
GC_12_99 b_12 NI_12 NS_99 0 9.0838948526275156e-08
GC_12_100 b_12 NI_12 NS_100 0 1.4512005826595624e-07
GC_12_101 b_12 NI_12 NS_101 0 1.5784606592809249e-07
GC_12_102 b_12 NI_12 NS_102 0 4.4529247489669853e-07
GC_12_103 b_12 NI_12 NS_103 0 2.3088526749001930e-08
GC_12_104 b_12 NI_12 NS_104 0 -1.6503980625855481e-07
GC_12_105 b_12 NI_12 NS_105 0 -3.7569230298299491e-08
GC_12_106 b_12 NI_12 NS_106 0 -1.2372686405968820e-07
GC_12_107 b_12 NI_12 NS_107 0 -8.6481660731132930e-08
GC_12_108 b_12 NI_12 NS_108 0 1.2325181425473164e-07
GC_12_109 b_12 NI_12 NS_109 0 -9.0264068330166675e-09
GC_12_110 b_12 NI_12 NS_110 0 -3.7855603820812815e-09
GC_12_111 b_12 NI_12 NS_111 0 2.2964572971866422e-12
GC_12_112 b_12 NI_12 NS_112 0 -3.3973157977027348e-12
GC_12_113 b_12 NI_12 NS_113 0 -7.3122987357502343e-10
GC_12_114 b_12 NI_12 NS_114 0 -8.2733841589519198e-11
GC_12_115 b_12 NI_12 NS_115 0 5.5770342646746362e-06
GC_12_116 b_12 NI_12 NS_116 0 -6.0661734556460391e-08
GC_12_117 b_12 NI_12 NS_117 0 -3.1618805112495728e-11
GC_12_118 b_12 NI_12 NS_118 0 4.1808080763510930e-10
GC_12_119 b_12 NI_12 NS_119 0 8.7028954262963440e-08
GC_12_120 b_12 NI_12 NS_120 0 -7.3629545499673162e-08
GC_12_121 b_12 NI_12 NS_121 0 3.8985572758694229e-09
GC_12_122 b_12 NI_12 NS_122 0 8.3796080511404351e-08
GC_12_123 b_12 NI_12 NS_123 0 6.3125380168506290e-07
GC_12_124 b_12 NI_12 NS_124 0 -8.3251282170956119e-07
GC_12_125 b_12 NI_12 NS_125 0 -9.1906435300967819e-07
GC_12_126 b_12 NI_12 NS_126 0 7.4744325045922499e-08
GC_12_127 b_12 NI_12 NS_127 0 5.4098498782682534e-07
GC_12_128 b_12 NI_12 NS_128 0 4.5916100138418416e-08
GC_12_129 b_12 NI_12 NS_129 0 -1.3830487463507988e-06
GC_12_130 b_12 NI_12 NS_130 0 -9.7965333021299006e-07
GC_12_131 b_12 NI_12 NS_131 0 3.0645726639518803e-07
GC_12_132 b_12 NI_12 NS_132 0 2.0540829609486133e-07
GC_12_133 b_12 NI_12 NS_133 0 -5.6263414137143580e-07
GC_12_134 b_12 NI_12 NS_134 0 7.1032651137303631e-07
GC_12_135 b_12 NI_12 NS_135 0 1.9975475748894595e-06
GC_12_136 b_12 NI_12 NS_136 0 -6.2826569637596251e-07
GC_12_137 b_12 NI_12 NS_137 0 -2.6418464478543042e-06
GC_12_138 b_12 NI_12 NS_138 0 3.8240853745332423e-07
GC_12_139 b_12 NI_12 NS_139 0 4.1242826955290817e-08
GC_12_140 b_12 NI_12 NS_140 0 1.4294319730479508e-06
GC_12_141 b_12 NI_12 NS_141 0 2.3346789663249041e-07
GC_12_142 b_12 NI_12 NS_142 0 -1.8326923177113972e-06
GC_12_143 b_12 NI_12 NS_143 0 -8.6531549618839780e-07
GC_12_144 b_12 NI_12 NS_144 0 1.3761787968677958e-06
GC_12_145 b_12 NI_12 NS_145 0 2.2851556894171110e-06
GC_12_146 b_12 NI_12 NS_146 0 2.9656044273633323e-06
GC_12_147 b_12 NI_12 NS_147 0 -2.0507151065540329e-06
GC_12_148 b_12 NI_12 NS_148 0 -3.4923364218270941e-06
GC_12_149 b_12 NI_12 NS_149 0 -2.8720393074610754e-07
GC_12_150 b_12 NI_12 NS_150 0 1.5382510849442903e-06
GC_12_151 b_12 NI_12 NS_151 0 1.7081737437118549e-06
GC_12_152 b_12 NI_12 NS_152 0 -1.8792221789353494e-06
GC_12_153 b_12 NI_12 NS_153 0 -1.6427702913770572e-06
GC_12_154 b_12 NI_12 NS_154 0 1.0311220770718560e-06
GC_12_155 b_12 NI_12 NS_155 0 4.2908073203536260e-07
GC_12_156 b_12 NI_12 NS_156 0 1.8543841373604474e-06
GC_12_157 b_12 NI_12 NS_157 0 2.5930376139251309e-07
GC_12_158 b_12 NI_12 NS_158 0 -2.2598885631856182e-06
GC_12_159 b_12 NI_12 NS_159 0 -7.4201414524560124e-07
GC_12_160 b_12 NI_12 NS_160 0 9.6146795983993518e-07
GC_12_161 b_12 NI_12 NS_161 0 2.0833922011960684e-06
GC_12_162 b_12 NI_12 NS_162 0 -1.8848659027160382e-08
GC_12_163 b_12 NI_12 NS_163 0 -1.8132678507282323e-06
GC_12_164 b_12 NI_12 NS_164 0 -3.2980078004817465e-07
GC_12_165 b_12 NI_12 NS_165 0 -9.5362760898797733e-08
GC_12_166 b_12 NI_12 NS_166 0 7.6458383141278367e-07
GC_12_167 b_12 NI_12 NS_167 0 2.1964067508762576e-07
GC_12_168 b_12 NI_12 NS_168 0 -5.5285387155829359e-07
GC_12_169 b_12 NI_12 NS_169 0 -2.4027916160821678e-07
GC_12_170 b_12 NI_12 NS_170 0 4.2925626705979780e-07
GC_12_171 b_12 NI_12 NS_171 0 1.0687535507745125e-07
GC_12_172 b_12 NI_12 NS_172 0 -2.2410620308940182e-07
GC_12_173 b_12 NI_12 NS_173 0 -4.5515335762647922e-07
GC_12_174 b_12 NI_12 NS_174 0 3.0526536441941567e-07
GC_12_175 b_12 NI_12 NS_175 0 2.0651311582650302e-07
GC_12_176 b_12 NI_12 NS_176 0 1.6780378384431621e-08
GC_12_177 b_12 NI_12 NS_177 0 -1.4742975916443225e-07
GC_12_178 b_12 NI_12 NS_178 0 1.9351604268094015e-07
GC_12_179 b_12 NI_12 NS_179 0 2.4897560900003375e-08
GC_12_180 b_12 NI_12 NS_180 0 -1.4136264098152233e-07
GC_12_181 b_12 NI_12 NS_181 0 -3.4516553777056247e-07
GC_12_182 b_12 NI_12 NS_182 0 2.7933059014359064e-07
GC_12_183 b_12 NI_12 NS_183 0 1.1041860926222167e-07
GC_12_184 b_12 NI_12 NS_184 0 -2.3166479027627731e-08
GC_12_185 b_12 NI_12 NS_185 0 -1.1146410092974311e-07
GC_12_186 b_12 NI_12 NS_186 0 2.2575709532411602e-07
GC_12_187 b_12 NI_12 NS_187 0 -1.8955184182405841e-08
GC_12_188 b_12 NI_12 NS_188 0 -1.6880172231994002e-07
GC_12_189 b_12 NI_12 NS_189 0 -2.8643062544148802e-07
GC_12_190 b_12 NI_12 NS_190 0 1.8674647712019689e-07
GC_12_191 b_12 NI_12 NS_191 0 -1.1166099415636608e-07
GC_12_192 b_12 NI_12 NS_192 0 -5.9934081059626595e-08
GC_12_193 b_12 NI_12 NS_193 0 -1.7481563849002855e-07
GC_12_194 b_12 NI_12 NS_194 0 2.0346172165963460e-07
GC_12_195 b_12 NI_12 NS_195 0 -2.9232268591847585e-07
GC_12_196 b_12 NI_12 NS_196 0 -3.9929793974533433e-08
GC_12_197 b_12 NI_12 NS_197 0 -4.9681199415775654e-07
GC_12_198 b_12 NI_12 NS_198 0 5.7772281396125621e-08
GC_12_199 b_12 NI_12 NS_199 0 2.7719570972637322e-06
GC_12_200 b_12 NI_12 NS_200 0 4.3304157303459167e-07
GC_12_201 b_12 NI_12 NS_201 0 -3.2409769149246616e-07
GC_12_202 b_12 NI_12 NS_202 0 6.7640652839991354e-07
GC_12_203 b_12 NI_12 NS_203 0 1.2398647155442557e-08
GC_12_204 b_12 NI_12 NS_204 0 1.2812489382938916e-08
GC_12_205 b_12 NI_12 NS_205 0 -6.7517231619751840e-09
GC_12_206 b_12 NI_12 NS_206 0 4.6496662538076238e-07
GC_12_207 b_12 NI_12 NS_207 0 -1.2602595866251918e-07
GC_12_208 b_12 NI_12 NS_208 0 2.6654224812818203e-07
GC_12_209 b_12 NI_12 NS_209 0 -4.8112937803454633e-07
GC_12_210 b_12 NI_12 NS_210 0 9.8550192576070880e-08
GC_12_211 b_12 NI_12 NS_211 0 -9.4591668290226211e-07
GC_12_212 b_12 NI_12 NS_212 0 4.8604669943459734e-07
GC_12_213 b_12 NI_12 NS_213 0 -1.8710254072709219e-07
GC_12_214 b_12 NI_12 NS_214 0 -7.9281385729734727e-08
GC_12_215 b_12 NI_12 NS_215 0 1.6412000956131669e-08
GC_12_216 b_12 NI_12 NS_216 0 -1.4793966732245660e-07
GC_12_217 b_12 NI_12 NS_217 0 8.6145546689325196e-08
GC_12_218 b_12 NI_12 NS_218 0 1.0231854932295099e-07
GC_12_219 b_12 NI_12 NS_219 0 -1.1791426263486852e-07
GC_12_220 b_12 NI_12 NS_220 0 -1.5795358369642100e-07
GC_12_221 b_12 NI_12 NS_221 0 -7.0288347847308830e-08
GC_12_222 b_12 NI_12 NS_222 0 8.1122611351489169e-08
GC_12_223 b_12 NI_12 NS_223 0 -4.4819706485192683e-10
GC_12_224 b_12 NI_12 NS_224 0 -3.7626835524543887e-08
GC_12_225 b_12 NI_12 NS_225 0 -8.0398873433896169e-12
GC_12_226 b_12 NI_12 NS_226 0 7.1578767894626875e-12
GC_12_227 b_12 NI_12 NS_227 0 9.6679467793816081e-10
GC_12_228 b_12 NI_12 NS_228 0 -3.3562036291267884e-10
GC_12_229 b_12 NI_12 NS_229 0 -2.7457198081352710e-05
GC_12_230 b_12 NI_12 NS_230 0 -1.0861269286693789e-08
GC_12_231 b_12 NI_12 NS_231 0 1.0272026304243843e-11
GC_12_232 b_12 NI_12 NS_232 0 -5.9964124873790826e-11
GC_12_233 b_12 NI_12 NS_233 0 -6.3440465848442807e-07
GC_12_234 b_12 NI_12 NS_234 0 -1.0701543154576423e-06
GC_12_235 b_12 NI_12 NS_235 0 -1.4351547579762262e-06
GC_12_236 b_12 NI_12 NS_236 0 2.3181029086755251e-06
GC_12_237 b_12 NI_12 NS_237 0 -3.8038702802996590e-06
GC_12_238 b_12 NI_12 NS_238 0 2.1755687328721488e-06
GC_12_239 b_12 NI_12 NS_239 0 1.9264787935302682e-06
GC_12_240 b_12 NI_12 NS_240 0 -2.2570782726326129e-07
GC_12_241 b_12 NI_12 NS_241 0 1.3997899620215362e-06
GC_12_242 b_12 NI_12 NS_242 0 5.7146733655811099e-06
GC_12_243 b_12 NI_12 NS_243 0 3.7149822073220796e-06
GC_12_244 b_12 NI_12 NS_244 0 3.2450366902692029e-06
GC_12_245 b_12 NI_12 NS_245 0 -1.4756134333568631e-06
GC_12_246 b_12 NI_12 NS_246 0 -9.4893577282280419e-07
GC_12_247 b_12 NI_12 NS_247 0 9.7600553356673144e-07
GC_12_248 b_12 NI_12 NS_248 0 -2.1770032464572028e-06
GC_12_249 b_12 NI_12 NS_249 0 6.4144780968236094e-06
GC_12_250 b_12 NI_12 NS_250 0 8.5313670815811913e-06
GC_12_251 b_12 NI_12 NS_251 0 1.3417320719968775e-06
GC_12_252 b_12 NI_12 NS_252 0 -9.5629790505220177e-07
GC_12_253 b_12 NI_12 NS_253 0 1.0785529915449994e-06
GC_12_254 b_12 NI_12 NS_254 0 -1.8906605506822056e-06
GC_12_255 b_12 NI_12 NS_255 0 1.4514874708048406e-05
GC_12_256 b_12 NI_12 NS_256 0 -4.1895944442332062e-06
GC_12_257 b_12 NI_12 NS_257 0 -2.0074935887909947e-07
GC_12_258 b_12 NI_12 NS_258 0 6.6361946137055432e-07
GC_12_259 b_12 NI_12 NS_259 0 4.9434222377041487e-06
GC_12_260 b_12 NI_12 NS_260 0 -2.1798298619719179e-06
GC_12_261 b_12 NI_12 NS_261 0 -7.7226308983758603e-07
GC_12_262 b_12 NI_12 NS_262 0 -1.5002469863078683e-05
GC_12_263 b_12 NI_12 NS_263 0 -7.8155801195303544e-08
GC_12_264 b_12 NI_12 NS_264 0 9.5811193829899488e-07
GC_12_265 b_12 NI_12 NS_265 0 -7.9220438157255751e-06
GC_12_266 b_12 NI_12 NS_266 0 -8.5842508912402321e-06
GC_12_267 b_12 NI_12 NS_267 0 -6.3253050837645003e-07
GC_12_268 b_12 NI_12 NS_268 0 -2.1422153111262797e-06
GC_12_269 b_12 NI_12 NS_269 0 -1.4549580911885479e-08
GC_12_270 b_12 NI_12 NS_270 0 1.1898787980369554e-06
GC_12_271 b_12 NI_12 NS_271 0 -7.7140594608565480e-06
GC_12_272 b_12 NI_12 NS_272 0 1.9652464508959753e-06
GC_12_273 b_12 NI_12 NS_273 0 2.3903649755308694e-07
GC_12_274 b_12 NI_12 NS_274 0 -1.6697063855202155e-06
GC_12_275 b_12 NI_12 NS_275 0 1.1429579149110565e-06
GC_12_276 b_12 NI_12 NS_276 0 3.0633038754050632e-06
GC_12_277 b_12 NI_12 NS_277 0 -9.6198427684319757e-07
GC_12_278 b_12 NI_12 NS_278 0 2.0271675349649848e-06
GC_12_279 b_12 NI_12 NS_279 0 4.5490131075044643e-07
GC_12_280 b_12 NI_12 NS_280 0 -1.2226950262642844e-06
GC_12_281 b_12 NI_12 NS_281 0 3.2356395948179478e-06
GC_12_282 b_12 NI_12 NS_282 0 -8.8238653313751630e-07
GC_12_283 b_12 NI_12 NS_283 0 -1.6006117773004264e-07
GC_12_284 b_12 NI_12 NS_284 0 5.0797766348978020e-07
GC_12_285 b_12 NI_12 NS_285 0 -8.4404473403598021e-07
GC_12_286 b_12 NI_12 NS_286 0 -4.1916218693652144e-07
GC_12_287 b_12 NI_12 NS_287 0 9.8705772653589023e-07
GC_12_288 b_12 NI_12 NS_288 0 -1.2634882933042166e-06
GC_12_289 b_12 NI_12 NS_289 0 1.4385478890026995e-06
GC_12_290 b_12 NI_12 NS_290 0 -5.6892752092285399e-07
GC_12_291 b_12 NI_12 NS_291 0 -3.3376530327779547e-08
GC_12_292 b_12 NI_12 NS_292 0 9.4899058573473301e-08
GC_12_293 b_12 NI_12 NS_293 0 -5.9608886847789584e-07
GC_12_294 b_12 NI_12 NS_294 0 -3.3988395664657937e-07
GC_12_295 b_12 NI_12 NS_295 0 9.6297947506862885e-07
GC_12_296 b_12 NI_12 NS_296 0 -1.0755592897191044e-06
GC_12_297 b_12 NI_12 NS_297 0 1.3913839776651086e-06
GC_12_298 b_12 NI_12 NS_298 0 -1.2415262747624892e-06
GC_12_299 b_12 NI_12 NS_299 0 1.6086496094433045e-07
GC_12_300 b_12 NI_12 NS_300 0 -4.5331700612490420e-08
GC_12_301 b_12 NI_12 NS_301 0 -4.8805319197381161e-07
GC_12_302 b_12 NI_12 NS_302 0 -5.0217527997926838e-07
GC_12_303 b_12 NI_12 NS_303 0 1.0601485229327623e-06
GC_12_304 b_12 NI_12 NS_304 0 -7.9957387247443440e-07
GC_12_305 b_12 NI_12 NS_305 0 1.2253856203039733e-06
GC_12_306 b_12 NI_12 NS_306 0 -2.1157312410361120e-06
GC_12_307 b_12 NI_12 NS_307 0 4.9452382328579030e-07
GC_12_308 b_12 NI_12 NS_308 0 -2.5500927009654916e-07
GC_12_309 b_12 NI_12 NS_309 0 -2.4639470318427703e-07
GC_12_310 b_12 NI_12 NS_310 0 -9.1751538413044107e-07
GC_12_311 b_12 NI_12 NS_311 0 1.9158197793311291e-06
GC_12_312 b_12 NI_12 NS_312 0 -9.9682461721228231e-07
GC_12_313 b_12 NI_12 NS_313 0 -8.0875222479123087e-06
GC_12_314 b_12 NI_12 NS_314 0 -9.1353127569708977e-07
GC_12_315 b_12 NI_12 NS_315 0 -3.1590337162050994e-07
GC_12_316 b_12 NI_12 NS_316 0 -3.6199255928385935e-06
GC_12_317 b_12 NI_12 NS_317 0 -4.8932606870547487e-08
GC_12_318 b_12 NI_12 NS_318 0 -3.3151000630122027e-08
GC_12_319 b_12 NI_12 NS_319 0 -1.0395690363734654e-07
GC_12_320 b_12 NI_12 NS_320 0 -1.2351493642510593e-06
GC_12_321 b_12 NI_12 NS_321 0 -1.0202892156738405e-06
GC_12_322 b_12 NI_12 NS_322 0 -6.6670133956182011e-07
GC_12_323 b_12 NI_12 NS_323 0 1.4550429510970709e-06
GC_12_324 b_12 NI_12 NS_324 0 -7.5893722247604287e-07
GC_12_325 b_12 NI_12 NS_325 0 1.9403669323438399e-06
GC_12_326 b_12 NI_12 NS_326 0 -1.8687373273549339e-06
GC_12_327 b_12 NI_12 NS_327 0 -2.2166860393825838e-07
GC_12_328 b_12 NI_12 NS_328 0 3.2466693800172733e-07
GC_12_329 b_12 NI_12 NS_329 0 2.1427531647984712e-07
GC_12_330 b_12 NI_12 NS_330 0 5.2885628425311394e-07
GC_12_331 b_12 NI_12 NS_331 0 -1.0742536344145290e-07
GC_12_332 b_12 NI_12 NS_332 0 -2.8271670388044420e-07
GC_12_333 b_12 NI_12 NS_333 0 7.8974202095665451e-09
GC_12_334 b_12 NI_12 NS_334 0 -9.5823355717609504e-08
GC_12_335 b_12 NI_12 NS_335 0 -8.8821323035092991e-08
GC_12_336 b_12 NI_12 NS_336 0 4.1483554343504027e-08
GC_12_337 b_12 NI_12 NS_337 0 -1.2204396709347823e-07
GC_12_338 b_12 NI_12 NS_338 0 -5.3450952266581933e-08
GC_12_339 b_12 NI_12 NS_339 0 6.1485578174179177e-12
GC_12_340 b_12 NI_12 NS_340 0 -1.7070652305939210e-12
GC_12_341 b_12 NI_12 NS_341 0 3.5216382834262060e-10
GC_12_342 b_12 NI_12 NS_342 0 6.9300824301121442e-10
GC_12_343 b_12 NI_12 NS_343 0 1.3355932951297539e-05
GC_12_344 b_12 NI_12 NS_344 0 -5.8997603119928608e-08
GC_12_345 b_12 NI_12 NS_345 0 -1.4899440183364424e-11
GC_12_346 b_12 NI_12 NS_346 0 1.3547819599370960e-10
GC_12_347 b_12 NI_12 NS_347 0 3.5636794409702870e-07
GC_12_348 b_12 NI_12 NS_348 0 -1.8177453337286710e-07
GC_12_349 b_12 NI_12 NS_349 0 2.7825893835895665e-07
GC_12_350 b_12 NI_12 NS_350 0 -3.4971823743689429e-07
GC_12_351 b_12 NI_12 NS_351 0 4.9250094039030385e-07
GC_12_352 b_12 NI_12 NS_352 0 -1.4213854673073219e-06
GC_12_353 b_12 NI_12 NS_353 0 -1.1592228397382233e-06
GC_12_354 b_12 NI_12 NS_354 0 -4.5897566855666529e-07
GC_12_355 b_12 NI_12 NS_355 0 -3.4112968388928967e-07
GC_12_356 b_12 NI_12 NS_356 0 -6.2118976506788748e-07
GC_12_357 b_12 NI_12 NS_357 0 -2.5796968392297985e-06
GC_12_358 b_12 NI_12 NS_358 0 -6.4054865770412626e-07
GC_12_359 b_12 NI_12 NS_359 0 7.1614973479565585e-07
GC_12_360 b_12 NI_12 NS_360 0 3.5572604135347639e-07
GC_12_361 b_12 NI_12 NS_361 0 -7.3376231007674419e-07
GC_12_362 b_12 NI_12 NS_362 0 3.7327424674723680e-07
GC_12_363 b_12 NI_12 NS_363 0 -9.8858907516469266e-07
GC_12_364 b_12 NI_12 NS_364 0 5.8562359543093700e-07
GC_12_365 b_12 NI_12 NS_365 0 -4.3258674469238149e-07
GC_12_366 b_12 NI_12 NS_366 0 2.6363663053606762e-07
GC_12_367 b_12 NI_12 NS_367 0 -8.4568603282038302e-07
GC_12_368 b_12 NI_12 NS_368 0 4.5886023131142242e-07
GC_12_369 b_12 NI_12 NS_369 0 1.6312867697947954e-07
GC_12_370 b_12 NI_12 NS_370 0 1.1048464340039689e-06
GC_12_371 b_12 NI_12 NS_371 0 -5.9745446629731512e-07
GC_12_372 b_12 NI_12 NS_372 0 1.3142481604168005e-07
GC_12_373 b_12 NI_12 NS_373 0 -1.8757719338098584e-06
GC_12_374 b_12 NI_12 NS_374 0 1.2999559433293131e-06
GC_12_375 b_12 NI_12 NS_375 0 2.0548077283299167e-06
GC_12_376 b_12 NI_12 NS_376 0 2.3036205632832794e-07
GC_12_377 b_12 NI_12 NS_377 0 -6.8567143777723086e-07
GC_12_378 b_12 NI_12 NS_378 0 2.0176516663253602e-07
GC_12_379 b_12 NI_12 NS_379 0 1.0020785347404325e-06
GC_12_380 b_12 NI_12 NS_380 0 1.6689080705406472e-06
GC_12_381 b_12 NI_12 NS_381 0 -2.4458558880739803e-07
GC_12_382 b_12 NI_12 NS_382 0 -5.7788280239181339e-07
GC_12_383 b_12 NI_12 NS_383 0 -9.1772848967104885e-07
GC_12_384 b_12 NI_12 NS_384 0 4.3231176340661655e-07
GC_12_385 b_12 NI_12 NS_385 0 1.4296285643215004e-06
GC_12_386 b_12 NI_12 NS_386 0 6.7975838223097577e-07
GC_12_387 b_12 NI_12 NS_387 0 -3.4205148895973859e-07
GC_12_388 b_12 NI_12 NS_388 0 -2.1142717522805926e-07
GC_12_389 b_12 NI_12 NS_389 0 -2.7750216653542332e-08
GC_12_390 b_12 NI_12 NS_390 0 1.4222469024175978e-06
GC_12_391 b_12 NI_12 NS_391 0 4.6031330471391123e-07
GC_12_392 b_12 NI_12 NS_392 0 -7.6889121334016489e-07
GC_12_393 b_12 NI_12 NS_393 0 -3.5271748865367967e-07
GC_12_394 b_12 NI_12 NS_394 0 4.9305992416818345e-08
GC_12_395 b_12 NI_12 NS_395 0 3.2510590237404916e-07
GC_12_396 b_12 NI_12 NS_396 0 3.7853232709312218e-07
GC_12_397 b_12 NI_12 NS_397 0 -1.4616429442199842e-07
GC_12_398 b_12 NI_12 NS_398 0 -8.4907376064080893e-09
GC_12_399 b_12 NI_12 NS_399 0 1.4143252893827973e-07
GC_12_400 b_12 NI_12 NS_400 0 1.2099137535792413e-07
GC_12_401 b_12 NI_12 NS_401 0 -1.9313704513766834e-07
GC_12_402 b_12 NI_12 NS_402 0 -6.8313805867983678e-08
GC_12_403 b_12 NI_12 NS_403 0 4.1149263993140064e-08
GC_12_404 b_12 NI_12 NS_404 0 1.9490952823555560e-07
GC_12_405 b_12 NI_12 NS_405 0 -1.1272482511266778e-07
GC_12_406 b_12 NI_12 NS_406 0 1.0158086664314896e-08
GC_12_407 b_12 NI_12 NS_407 0 4.5539216151541987e-08
GC_12_408 b_12 NI_12 NS_408 0 4.4122094186739165e-09
GC_12_409 b_12 NI_12 NS_409 0 -2.9983391388662794e-07
GC_12_410 b_12 NI_12 NS_410 0 -5.1244849392697095e-08
GC_12_411 b_12 NI_12 NS_411 0 -9.0041916524272147e-08
GC_12_412 b_12 NI_12 NS_412 0 6.0468622408778248e-08
GC_12_413 b_12 NI_12 NS_413 0 -2.3102772772423203e-07
GC_12_414 b_12 NI_12 NS_414 0 8.0940792457824097e-08
GC_12_415 b_12 NI_12 NS_415 0 -1.3243199276390781e-07
GC_12_416 b_12 NI_12 NS_416 0 -7.1040742428343156e-08
GC_12_417 b_12 NI_12 NS_417 0 -4.3092860568759395e-07
GC_12_418 b_12 NI_12 NS_418 0 -5.3209975320041420e-08
GC_12_419 b_12 NI_12 NS_419 0 -4.1895507229298425e-07
GC_12_420 b_12 NI_12 NS_420 0 6.1480320889421376e-08
GC_12_421 b_12 NI_12 NS_421 0 -4.4023024600414184e-07
GC_12_422 b_12 NI_12 NS_422 0 1.4721695792263812e-07
GC_12_423 b_12 NI_12 NS_423 0 -5.1067992362793639e-07
GC_12_424 b_12 NI_12 NS_424 0 9.9879999148486955e-08
GC_12_425 b_12 NI_12 NS_425 0 -9.6150424491954613e-07
GC_12_426 b_12 NI_12 NS_426 0 -9.5716738355108106e-08
GC_12_427 b_12 NI_12 NS_427 0 2.6176284267641073e-06
GC_12_428 b_12 NI_12 NS_428 0 2.9785681077440293e-06
GC_12_429 b_12 NI_12 NS_429 0 -6.1418778371126820e-07
GC_12_430 b_12 NI_12 NS_430 0 1.0336830830980190e-06
GC_12_431 b_12 NI_12 NS_431 0 9.1644702004310847e-09
GC_12_432 b_12 NI_12 NS_432 0 2.5329135803755147e-08
GC_12_433 b_12 NI_12 NS_433 0 -4.6836667282558428e-07
GC_12_434 b_12 NI_12 NS_434 0 8.2780390087802599e-07
GC_12_435 b_12 NI_12 NS_435 0 8.8696783218351241e-09
GC_12_436 b_12 NI_12 NS_436 0 3.8273376762664301e-07
GC_12_437 b_12 NI_12 NS_437 0 -8.6693343470313429e-07
GC_12_438 b_12 NI_12 NS_438 0 -7.0542592551397525e-08
GC_12_439 b_12 NI_12 NS_439 0 -9.7666785407555319e-07
GC_12_440 b_12 NI_12 NS_440 0 -1.7992974993671840e-07
GC_12_441 b_12 NI_12 NS_441 0 1.0735189369959265e-07
GC_12_442 b_12 NI_12 NS_442 0 -1.4754510294506310e-07
GC_12_443 b_12 NI_12 NS_443 0 6.6793613444896520e-08
GC_12_444 b_12 NI_12 NS_444 0 1.4683528477022127e-08
GC_12_445 b_12 NI_12 NS_445 0 -6.9788123400704909e-08
GC_12_446 b_12 NI_12 NS_446 0 1.6094618600718488e-07
GC_12_447 b_12 NI_12 NS_447 0 2.7671224900691884e-08
GC_12_448 b_12 NI_12 NS_448 0 -4.0810011337466634e-08
GC_12_449 b_12 NI_12 NS_449 0 -8.1264163059353863e-08
GC_12_450 b_12 NI_12 NS_450 0 1.6048705050084314e-07
GC_12_451 b_12 NI_12 NS_451 0 5.6542066765028338e-08
GC_12_452 b_12 NI_12 NS_452 0 -1.6756766345953555e-08
GC_12_453 b_12 NI_12 NS_453 0 -1.1794865080653339e-11
GC_12_454 b_12 NI_12 NS_454 0 5.2725137581141396e-12
GC_12_455 b_12 NI_12 NS_455 0 -3.4161810509075794e-10
GC_12_456 b_12 NI_12 NS_456 0 -9.7247779193747477e-10
GC_12_457 b_12 NI_12 NS_457 0 -6.3151479646485242e-05
GC_12_458 b_12 NI_12 NS_458 0 3.1403616382992635e-07
GC_12_459 b_12 NI_12 NS_459 0 1.6220140324436376e-11
GC_12_460 b_12 NI_12 NS_460 0 -9.0649099428488083e-11
GC_12_461 b_12 NI_12 NS_461 0 -1.1289889059201628e-06
GC_12_462 b_12 NI_12 NS_462 0 -1.7888659896650046e-06
GC_12_463 b_12 NI_12 NS_463 0 -1.9838392392693765e-06
GC_12_464 b_12 NI_12 NS_464 0 1.9933847812559950e-06
GC_12_465 b_12 NI_12 NS_465 0 -9.6952313748635819e-06
GC_12_466 b_12 NI_12 NS_466 0 6.8014506380044873e-07
GC_12_467 b_12 NI_12 NS_467 0 -2.5333408623516261e-07
GC_12_468 b_12 NI_12 NS_468 0 3.4894147993865549e-06
GC_12_469 b_12 NI_12 NS_469 0 -2.1026830732386800e-06
GC_12_470 b_12 NI_12 NS_470 0 1.1808595870521234e-05
GC_12_471 b_12 NI_12 NS_471 0 6.7560362819043677e-06
GC_12_472 b_12 NI_12 NS_472 0 1.2503595821363610e-05
GC_12_473 b_12 NI_12 NS_473 0 -1.9973655972299836e-06
GC_12_474 b_12 NI_12 NS_474 0 -2.3069635378795347e-06
GC_12_475 b_12 NI_12 NS_475 0 1.6477115548275695e-06
GC_12_476 b_12 NI_12 NS_476 0 9.5582678205058669e-07
GC_12_477 b_12 NI_12 NS_477 0 7.5392955146103758e-06
GC_12_478 b_12 NI_12 NS_478 0 3.8837522360603382e-05
GC_12_479 b_12 NI_12 NS_479 0 2.3057223750268232e-05
GC_12_480 b_12 NI_12 NS_480 0 -1.1826467579353454e-05
GC_12_481 b_12 NI_12 NS_481 0 8.3538354343182921e-06
GC_12_482 b_12 NI_12 NS_482 0 1.6579965590560142e-06
GC_12_483 b_12 NI_12 NS_483 0 4.8581026502507160e-05
GC_12_484 b_12 NI_12 NS_484 0 -2.5173284138716395e-05
GC_12_485 b_12 NI_12 NS_485 0 -8.6231591195469729e-07
GC_12_486 b_12 NI_12 NS_486 0 -7.8674971074423522e-06
GC_12_487 b_12 NI_12 NS_487 0 3.4181897428830383e-05
GC_12_488 b_12 NI_12 NS_488 0 -7.8071060267114346e-06
GC_12_489 b_12 NI_12 NS_489 0 -3.8154375935252743e-05
GC_12_490 b_12 NI_12 NS_490 0 -5.2649699442514802e-05
GC_12_491 b_12 NI_12 NS_491 0 -4.4897622047404384e-06
GC_12_492 b_12 NI_12 NS_492 0 -4.3444025142607852e-06
GC_12_493 b_12 NI_12 NS_493 0 -3.9819364804270504e-05
GC_12_494 b_12 NI_12 NS_494 0 -2.0163480356375424e-05
GC_12_495 b_12 NI_12 NS_495 0 -4.8690175145382353e-06
GC_12_496 b_12 NI_12 NS_496 0 6.2179216110498622e-06
GC_12_497 b_12 NI_12 NS_497 0 -8.5133364547763216e-06
GC_12_498 b_12 NI_12 NS_498 0 -4.6696241647340785e-07
GC_12_499 b_12 NI_12 NS_499 0 -1.5584987737204824e-05
GC_12_500 b_12 NI_12 NS_500 0 2.4311328781433761e-05
GC_12_501 b_12 NI_12 NS_501 0 1.1061841449537231e-06
GC_12_502 b_12 NI_12 NS_502 0 2.3729737500130170e-06
GC_12_503 b_12 NI_12 NS_503 0 3.2346306877891416e-06
GC_12_504 b_12 NI_12 NS_504 0 1.8506898201813049e-05
GC_12_505 b_12 NI_12 NS_505 0 7.5468321069855793e-06
GC_12_506 b_12 NI_12 NS_506 0 -1.3939235359379944e-06
GC_12_507 b_12 NI_12 NS_507 0 2.9977264752081403e-06
GC_12_508 b_12 NI_12 NS_508 0 -5.0827961847063177e-07
GC_12_509 b_12 NI_12 NS_509 0 7.6492580152603606e-06
GC_12_510 b_12 NI_12 NS_510 0 -4.5387674753971326e-06
GC_12_511 b_12 NI_12 NS_511 0 -8.6278316576892777e-07
GC_12_512 b_12 NI_12 NS_512 0 -4.4779084119082921e-07
GC_12_513 b_12 NI_12 NS_513 0 -1.7230525683939194e-06
GC_12_514 b_12 NI_12 NS_514 0 1.8501990210604801e-07
GC_12_515 b_12 NI_12 NS_515 0 1.6122471780300807e-06
GC_12_516 b_12 NI_12 NS_516 0 -2.6583966987180045e-08
GC_12_517 b_12 NI_12 NS_517 0 3.7023977399018655e-06
GC_12_518 b_12 NI_12 NS_518 0 -9.2832662431562225e-07
GC_12_519 b_12 NI_12 NS_519 0 -8.7821831349275399e-08
GC_12_520 b_12 NI_12 NS_520 0 -3.4286794452128796e-07
GC_12_521 b_12 NI_12 NS_521 0 -5.7131990930226513e-07
GC_12_522 b_12 NI_12 NS_522 0 5.0950898621794342e-07
GC_12_523 b_12 NI_12 NS_523 0 2.4653241194160510e-06
GC_12_524 b_12 NI_12 NS_524 0 1.0743342348455854e-07
GC_12_525 b_12 NI_12 NS_525 0 3.4040158769199476e-06
GC_12_526 b_12 NI_12 NS_526 0 -2.8619461730287980e-06
GC_12_527 b_12 NI_12 NS_527 0 -2.6885138282885733e-07
GC_12_528 b_12 NI_12 NS_528 0 -5.0646602669568013e-08
GC_12_529 b_12 NI_12 NS_529 0 7.1805269310822919e-07
GC_12_530 b_12 NI_12 NS_530 0 1.0014726005936638e-06
GC_12_531 b_12 NI_12 NS_531 0 3.5530359088682934e-06
GC_12_532 b_12 NI_12 NS_532 0 3.3902885580506720e-08
GC_12_533 b_12 NI_12 NS_533 0 2.4205289882146560e-06
GC_12_534 b_12 NI_12 NS_534 0 -4.6592135654399254e-06
GC_12_535 b_12 NI_12 NS_535 0 4.5470749692424026e-07
GC_12_536 b_12 NI_12 NS_536 0 1.1297783182219890e-06
GC_12_537 b_12 NI_12 NS_537 0 3.6719812719131452e-06
GC_12_538 b_12 NI_12 NS_538 0 -6.9207920111322125e-07
GC_12_539 b_12 NI_12 NS_539 0 5.6214540005587947e-06
GC_12_540 b_12 NI_12 NS_540 0 -9.7041075987921387e-07
GC_12_541 b_12 NI_12 NS_541 0 -1.6193981823440883e-05
GC_12_542 b_12 NI_12 NS_542 0 -1.0663748956979456e-05
GC_12_543 b_12 NI_12 NS_543 0 9.4555423720488743e-07
GC_12_544 b_12 NI_12 NS_544 0 -7.5011978029700735e-06
GC_12_545 b_12 NI_12 NS_545 0 -6.7320592401156869e-08
GC_12_546 b_12 NI_12 NS_546 0 -1.4895715851987488e-07
GC_12_547 b_12 NI_12 NS_547 0 1.8076709327555556e-06
GC_12_548 b_12 NI_12 NS_548 0 -1.8968909943718328e-06
GC_12_549 b_12 NI_12 NS_549 0 5.3801649926901576e-07
GC_12_550 b_12 NI_12 NS_550 0 -3.4001984930779956e-06
GC_12_551 b_12 NI_12 NS_551 0 3.4182948497476351e-06
GC_12_552 b_12 NI_12 NS_552 0 -1.3139430598827681e-06
GC_12_553 b_12 NI_12 NS_553 0 4.5934173820076145e-06
GC_12_554 b_12 NI_12 NS_554 0 -8.0351596303825614e-07
GC_12_555 b_12 NI_12 NS_555 0 -1.9741210290143374e-07
GC_12_556 b_12 NI_12 NS_556 0 -2.0545975835566192e-07
GC_12_557 b_12 NI_12 NS_557 0 7.0278285328316060e-07
GC_12_558 b_12 NI_12 NS_558 0 1.4079554507146564e-06
GC_12_559 b_12 NI_12 NS_559 0 -7.0034213540927483e-07
GC_12_560 b_12 NI_12 NS_560 0 -1.4717285215786495e-06
GC_12_561 b_12 NI_12 NS_561 0 -6.2802182597474681e-07
GC_12_562 b_12 NI_12 NS_562 0 8.2383983778095754e-07
GC_12_563 b_12 NI_12 NS_563 0 2.2514746926033982e-07
GC_12_564 b_12 NI_12 NS_564 0 6.5403179905314915e-07
GC_12_565 b_12 NI_12 NS_565 0 6.0595900880915221e-07
GC_12_566 b_12 NI_12 NS_566 0 2.0968576679176088e-08
GC_12_567 b_12 NI_12 NS_567 0 1.3952627010071900e-11
GC_12_568 b_12 NI_12 NS_568 0 5.3746510608447324e-13
GC_12_569 b_12 NI_12 NS_569 0 4.3669365533288495e-10
GC_12_570 b_12 NI_12 NS_570 0 1.6922310274372240e-09
GC_12_571 b_12 NI_12 NS_571 0 8.4593926149263395e-05
GC_12_572 b_12 NI_12 NS_572 0 1.9043596353364018e-07
GC_12_573 b_12 NI_12 NS_573 0 2.0152905601473299e-11
GC_12_574 b_12 NI_12 NS_574 0 -9.4454546245986934e-10
GC_12_575 b_12 NI_12 NS_575 0 8.8362780196969830e-07
GC_12_576 b_12 NI_12 NS_576 0 5.7800597995559662e-08
GC_12_577 b_12 NI_12 NS_577 0 1.1605036451708183e-06
GC_12_578 b_12 NI_12 NS_578 0 6.9649753209708969e-08
GC_12_579 b_12 NI_12 NS_579 0 3.3633120180077879e-06
GC_12_580 b_12 NI_12 NS_580 0 -3.2270900773418764e-06
GC_12_581 b_12 NI_12 NS_581 0 -2.0864348552077136e-06
GC_12_582 b_12 NI_12 NS_582 0 -1.7323698066641211e-06
GC_12_583 b_12 NI_12 NS_583 0 1.9309980643002236e-06
GC_12_584 b_12 NI_12 NS_584 0 -2.2101003139660085e-06
GC_12_585 b_12 NI_12 NS_585 0 -5.8945401559641371e-06
GC_12_586 b_12 NI_12 NS_586 0 -7.1428800561098910e-06
GC_12_587 b_12 NI_12 NS_587 0 9.5034331326945719e-07
GC_12_588 b_12 NI_12 NS_588 0 2.2267365536703217e-06
GC_12_589 b_12 NI_12 NS_589 0 -2.2769834510150930e-06
GC_12_590 b_12 NI_12 NS_590 0 8.0128623192042992e-07
GC_12_591 b_12 NI_12 NS_591 0 5.8088974582295178e-07
GC_12_592 b_12 NI_12 NS_592 0 -4.8941795462781290e-06
GC_12_593 b_12 NI_12 NS_593 0 -6.4026883180881599e-06
GC_12_594 b_12 NI_12 NS_594 0 2.7563305568173496e-06
GC_12_595 b_12 NI_12 NS_595 0 -1.0161048031291296e-06
GC_12_596 b_12 NI_12 NS_596 0 1.6584682219969056e-06
GC_12_597 b_12 NI_12 NS_597 0 -3.3725639422014795e-06
GC_12_598 b_12 NI_12 NS_598 0 -2.5283982785544891e-06
GC_12_599 b_12 NI_12 NS_599 0 -2.2050139890520611e-06
GC_12_600 b_12 NI_12 NS_600 0 2.3624368125054332e-06
GC_12_601 b_12 NI_12 NS_601 0 1.5143149240673696e-06
GC_12_602 b_12 NI_12 NS_602 0 2.6092781502856626e-06
GC_12_603 b_12 NI_12 NS_603 0 -5.1177174707864313e-06
GC_12_604 b_12 NI_12 NS_604 0 -2.0375227433062257e-06
GC_12_605 b_12 NI_12 NS_605 0 -1.4942735811510266e-06
GC_12_606 b_12 NI_12 NS_606 0 2.2229727093621779e-06
GC_12_607 b_12 NI_12 NS_607 0 -4.8186663483279778e-08
GC_12_608 b_12 NI_12 NS_608 0 -1.0705799300334927e-06
GC_12_609 b_12 NI_12 NS_609 0 -2.7776411432456651e-06
GC_12_610 b_12 NI_12 NS_610 0 1.7676654693058952e-06
GC_12_611 b_12 NI_12 NS_611 0 -7.8794272070624831e-07
GC_12_612 b_12 NI_12 NS_612 0 2.3418923612723254e-06
GC_12_613 b_12 NI_12 NS_613 0 -1.0030640163524916e-06
GC_12_614 b_12 NI_12 NS_614 0 -1.3429445376043120e-06
GC_12_615 b_12 NI_12 NS_615 0 -1.8385160115766452e-06
GC_12_616 b_12 NI_12 NS_616 0 1.3366200610854477e-06
GC_12_617 b_12 NI_12 NS_617 0 5.5156984335514135e-07
GC_12_618 b_12 NI_12 NS_618 0 1.6537106679486785e-07
GC_12_619 b_12 NI_12 NS_619 0 -2.9420515402751224e-06
GC_12_620 b_12 NI_12 NS_620 0 3.7600493235065579e-07
GC_12_621 b_12 NI_12 NS_621 0 -9.6513324024708731e-07
GC_12_622 b_12 NI_12 NS_622 0 7.1182582612754483e-07
GC_12_623 b_12 NI_12 NS_623 0 -1.9725834936859443e-06
GC_12_624 b_12 NI_12 NS_624 0 -7.9480746050119919e-07
GC_12_625 b_12 NI_12 NS_625 0 -1.4687825946320634e-06
GC_12_626 b_12 NI_12 NS_626 0 6.2110231123426506e-07
GC_12_627 b_12 NI_12 NS_627 0 -1.1171947598872279e-06
GC_12_628 b_12 NI_12 NS_628 0 -3.9215272633646945e-07
GC_12_629 b_12 NI_12 NS_629 0 -2.4596159063533229e-06
GC_12_630 b_12 NI_12 NS_630 0 -6.3464683244308905e-07
GC_12_631 b_12 NI_12 NS_631 0 -3.0281902254575681e-06
GC_12_632 b_12 NI_12 NS_632 0 -3.1125355329886161e-07
GC_12_633 b_12 NI_12 NS_633 0 -2.1722946400843213e-06
GC_12_634 b_12 NI_12 NS_634 0 3.1827835621035728e-07
GC_12_635 b_12 NI_12 NS_635 0 -2.7407137864623458e-06
GC_12_636 b_12 NI_12 NS_636 0 3.0329398634317531e-07
GC_12_637 b_12 NI_12 NS_637 0 -4.2063160127156936e-06
GC_12_638 b_12 NI_12 NS_638 0 -7.3431026777850807e-07
GC_12_639 b_12 NI_12 NS_639 0 -5.6821673966488860e-06
GC_12_640 b_12 NI_12 NS_640 0 2.2501737066034747e-06
GC_12_641 b_12 NI_12 NS_641 0 -3.1748893419764495e-06
GC_12_642 b_12 NI_12 NS_642 0 1.8636235047452636e-06
GC_12_643 b_12 NI_12 NS_643 0 -4.1156134480057832e-06
GC_12_644 b_12 NI_12 NS_644 0 3.2996228125180558e-06
GC_12_645 b_12 NI_12 NS_645 0 -5.6743075122437924e-06
GC_12_646 b_12 NI_12 NS_646 0 1.3489559168758944e-06
GC_12_647 b_12 NI_12 NS_647 0 -3.5124559272365930e-06
GC_12_648 b_12 NI_12 NS_648 0 8.2350279372963412e-06
GC_12_649 b_12 NI_12 NS_649 0 -2.3080091890229257e-06
GC_12_650 b_12 NI_12 NS_650 0 4.5638944761088940e-06
GC_12_651 b_12 NI_12 NS_651 0 1.1256609112857333e-06
GC_12_652 b_12 NI_12 NS_652 0 5.4143278284707061e-06
GC_12_653 b_12 NI_12 NS_653 0 -1.8435295947777901e-06
GC_12_654 b_12 NI_12 NS_654 0 3.4528269249336065e-06
GC_12_655 b_12 NI_12 NS_655 0 -7.0146452210771115e-06
GC_12_656 b_12 NI_12 NS_656 0 3.7171362690419331e-05
GC_12_657 b_12 NI_12 NS_657 0 6.9438991290122009e-07
GC_12_658 b_12 NI_12 NS_658 0 2.6520866469384482e-06
GC_12_659 b_12 NI_12 NS_659 0 -8.4705172943896649e-08
GC_12_660 b_12 NI_12 NS_660 0 1.1842641879097560e-07
GC_12_661 b_12 NI_12 NS_661 0 -7.2474238089818423e-07
GC_12_662 b_12 NI_12 NS_662 0 3.4155276433231246e-06
GC_12_663 b_12 NI_12 NS_663 0 6.7707655039384947e-07
GC_12_664 b_12 NI_12 NS_664 0 8.6166721693074725e-07
GC_12_665 b_12 NI_12 NS_665 0 2.2818964634523432e-06
GC_12_666 b_12 NI_12 NS_666 0 -3.1368152206912394e-06
GC_12_667 b_12 NI_12 NS_667 0 -1.5493205702460330e-06
GC_12_668 b_12 NI_12 NS_668 0 -1.1843768285299898e-05
GC_12_669 b_12 NI_12 NS_669 0 2.0448386827847780e-06
GC_12_670 b_12 NI_12 NS_670 0 -7.3745640320620696e-07
GC_12_671 b_12 NI_12 NS_671 0 4.5136862882755118e-06
GC_12_672 b_12 NI_12 NS_672 0 -4.0126034440111585e-07
GC_12_673 b_12 NI_12 NS_673 0 1.2442635413716775e-06
GC_12_674 b_12 NI_12 NS_674 0 1.9854521151302685e-06
GC_12_675 b_12 NI_12 NS_675 0 1.7412903996991407e-06
GC_12_676 b_12 NI_12 NS_676 0 -7.6164130640138304e-07
GC_12_677 b_12 NI_12 NS_677 0 5.8319850657314544e-07
GC_12_678 b_12 NI_12 NS_678 0 5.1106040757488562e-07
GC_12_679 b_12 NI_12 NS_679 0 6.5667020224133441e-07
GC_12_680 b_12 NI_12 NS_680 0 -7.6188648604995071e-08
GC_12_681 b_12 NI_12 NS_681 0 2.2923144842456599e-11
GC_12_682 b_12 NI_12 NS_682 0 -9.3363899753944687e-11
GC_12_683 b_12 NI_12 NS_683 0 -1.8301886268116168e-09
GC_12_684 b_12 NI_12 NS_684 0 4.0621509345822190e-09
GC_12_685 b_12 NI_12 NS_685 0 -3.7756381926466130e-05
GC_12_686 b_12 NI_12 NS_686 0 2.2260817727649823e-06
GC_12_687 b_12 NI_12 NS_687 0 6.0497156285814965e-11
GC_12_688 b_12 NI_12 NS_688 0 3.0748225040605811e-09
GC_12_689 b_12 NI_12 NS_689 0 -1.9312551528564528e-06
GC_12_690 b_12 NI_12 NS_690 0 -1.7210842911264364e-06
GC_12_691 b_12 NI_12 NS_691 0 -5.6039609666275821e-06
GC_12_692 b_12 NI_12 NS_692 0 2.9249078517585408e-06
GC_12_693 b_12 NI_12 NS_693 0 -1.6662521232538384e-05
GC_12_694 b_12 NI_12 NS_694 0 1.9136217848583669e-05
GC_12_695 b_12 NI_12 NS_695 0 1.5401878387688226e-05
GC_12_696 b_12 NI_12 NS_696 0 1.0211465239430676e-05
GC_12_697 b_12 NI_12 NS_697 0 1.7356895254832501e-05
GC_12_698 b_12 NI_12 NS_698 0 2.3278503558763436e-05
GC_12_699 b_12 NI_12 NS_699 0 3.0897972692973332e-05
GC_12_700 b_12 NI_12 NS_700 0 5.3455367719961628e-06
GC_12_701 b_12 NI_12 NS_701 0 -3.3855537530674235e-06
GC_12_702 b_12 NI_12 NS_702 0 -2.1457428434071354e-06
GC_12_703 b_12 NI_12 NS_703 0 1.7191268256229552e-05
GC_12_704 b_12 NI_12 NS_704 0 -2.2223448031406201e-06
GC_12_705 b_12 NI_12 NS_705 0 1.2979418727964378e-04
GC_12_706 b_12 NI_12 NS_706 0 3.5245570894507617e-05
GC_12_707 b_12 NI_12 NS_707 0 -2.8533571420483203e-05
GC_12_708 b_12 NI_12 NS_708 0 -9.9832754249268581e-05
GC_12_709 b_12 NI_12 NS_709 0 2.5236941729685763e-05
GC_12_710 b_12 NI_12 NS_710 0 -3.1267147316634176e-05
GC_12_711 b_12 NI_12 NS_711 0 -4.0931247562640653e-05
GC_12_712 b_12 NI_12 NS_712 0 -1.6750292475162435e-04
GC_12_713 b_12 NI_12 NS_713 0 -4.1821890331728534e-05
GC_12_714 b_12 NI_12 NS_714 0 -5.3846148808632730e-06
GC_12_715 b_12 NI_12 NS_715 0 2.2549187450343845e-05
GC_12_716 b_12 NI_12 NS_716 0 -1.5152140313729704e-04
GC_12_717 b_12 NI_12 NS_717 0 -2.3148654672580082e-04
GC_12_718 b_12 NI_12 NS_718 0 1.1299996471385613e-04
GC_12_719 b_12 NI_12 NS_719 0 -3.7411586670333995e-05
GC_12_720 b_12 NI_12 NS_720 0 1.3952382995249238e-05
GC_12_721 b_12 NI_12 NS_721 0 -1.3781859310212557e-04
GC_12_722 b_12 NI_12 NS_722 0 1.2973528123262984e-04
GC_12_723 b_12 NI_12 NS_723 0 3.6132291565477571e-05
GC_12_724 b_12 NI_12 NS_724 0 4.1461476250144669e-05
GC_12_725 b_12 NI_12 NS_725 0 -3.8173870822222744e-05
GC_12_726 b_12 NI_12 NS_726 0 4.2971183739088891e-05
GC_12_727 b_12 NI_12 NS_727 0 8.7354666024668485e-05
GC_12_728 b_12 NI_12 NS_728 0 1.1821531665952493e-04
GC_12_729 b_12 NI_12 NS_729 0 2.7245014869661550e-05
GC_12_730 b_12 NI_12 NS_730 0 1.0262327903278377e-05
GC_12_731 b_12 NI_12 NS_731 0 8.7158314556992170e-05
GC_12_732 b_12 NI_12 NS_732 0 6.5380981031831130e-05
GC_12_733 b_12 NI_12 NS_733 0 2.0400946713469735e-05
GC_12_734 b_12 NI_12 NS_734 0 -5.7168782988975833e-05
GC_12_735 b_12 NI_12 NS_735 0 1.7001878586987111e-05
GC_12_736 b_12 NI_12 NS_736 0 -8.8439679836310878e-06
GC_12_737 b_12 NI_12 NS_737 0 8.4707440687939225e-06
GC_12_738 b_12 NI_12 NS_738 0 -3.3126328093523921e-05
GC_12_739 b_12 NI_12 NS_739 0 -8.8428608762457518e-06
GC_12_740 b_12 NI_12 NS_740 0 4.1505705308858399e-07
GC_12_741 b_12 NI_12 NS_741 0 -2.4022633064500374e-06
GC_12_742 b_12 NI_12 NS_742 0 8.4362258472699224e-06
GC_12_743 b_12 NI_12 NS_743 0 1.0207782701035645e-05
GC_12_744 b_12 NI_12 NS_744 0 6.0582482293486297e-06
GC_12_745 b_12 NI_12 NS_745 0 1.2154867527890102e-05
GC_12_746 b_12 NI_12 NS_746 0 -7.9359225048967089e-06
GC_12_747 b_12 NI_12 NS_747 0 -3.4649723845851143e-06
GC_12_748 b_12 NI_12 NS_748 0 -5.2258255008075030e-07
GC_12_749 b_12 NI_12 NS_749 0 2.5132143750461816e-06
GC_12_750 b_12 NI_12 NS_750 0 7.3270763045030073e-06
GC_12_751 b_12 NI_12 NS_751 0 1.3691635557920648e-05
GC_12_752 b_12 NI_12 NS_752 0 2.6181804793722225e-06
GC_12_753 b_12 NI_12 NS_753 0 4.5508800268634291e-06
GC_12_754 b_12 NI_12 NS_754 0 -1.4312549477996423e-05
GC_12_755 b_12 NI_12 NS_755 0 -5.8920342605727627e-06
GC_12_756 b_12 NI_12 NS_756 0 4.1741258445272523e-06
GC_12_757 b_12 NI_12 NS_757 0 1.0370348903885745e-05
GC_12_758 b_12 NI_12 NS_758 0 9.8155496420341911e-06
GC_12_759 b_12 NI_12 NS_759 0 1.7399256529806333e-05
GC_12_760 b_12 NI_12 NS_760 0 -4.2746286268861718e-06
GC_12_761 b_12 NI_12 NS_761 0 -9.2261162511230191e-06
GC_12_762 b_12 NI_12 NS_762 0 -1.5489746007534268e-05
GC_12_763 b_12 NI_12 NS_763 0 -4.0027782098349653e-06
GC_12_764 b_12 NI_12 NS_764 0 1.3420162887745478e-05
GC_12_765 b_12 NI_12 NS_765 0 2.1008728828449225e-05
GC_12_766 b_12 NI_12 NS_766 0 -7.6329813357895238e-07
GC_12_767 b_12 NI_12 NS_767 0 9.1216872121788214e-06
GC_12_768 b_12 NI_12 NS_768 0 -1.7455310087237491e-05
GC_12_769 b_12 NI_12 NS_769 0 1.4592622215686221e-06
GC_12_770 b_12 NI_12 NS_770 0 -1.4427431571657638e-05
GC_12_771 b_12 NI_12 NS_771 0 -1.3809069230371411e-05
GC_12_772 b_12 NI_12 NS_772 0 3.9888923101473341e-06
GC_12_773 b_12 NI_12 NS_773 0 9.7995432137085831e-09
GC_12_774 b_12 NI_12 NS_774 0 -4.8130472162365125e-08
GC_12_775 b_12 NI_12 NS_775 0 8.6298552215683204e-06
GC_12_776 b_12 NI_12 NS_776 0 1.1373630205874293e-05
GC_12_777 b_12 NI_12 NS_777 0 1.0873523404844628e-05
GC_12_778 b_12 NI_12 NS_778 0 -1.1464205027921602e-05
GC_12_779 b_12 NI_12 NS_779 0 -3.5307993787517500e-06
GC_12_780 b_12 NI_12 NS_780 0 -1.0164881907944783e-05
GC_12_781 b_12 NI_12 NS_781 0 -2.0125620160468493e-06
GC_12_782 b_12 NI_12 NS_782 0 1.2870555605653747e-05
GC_12_783 b_12 NI_12 NS_783 0 9.7604679238933993e-07
GC_12_784 b_12 NI_12 NS_784 0 -7.2620465698303252e-06
GC_12_785 b_12 NI_12 NS_785 0 7.4715654283397044e-06
GC_12_786 b_12 NI_12 NS_786 0 1.7440195079031979e-06
GC_12_787 b_12 NI_12 NS_787 0 -6.1165635161320866e-06
GC_12_788 b_12 NI_12 NS_788 0 -8.8986429009226738e-06
GC_12_789 b_12 NI_12 NS_789 0 -4.1366749985392227e-06
GC_12_790 b_12 NI_12 NS_790 0 9.6568903882806738e-06
GC_12_791 b_12 NI_12 NS_791 0 3.3152499122646773e-06
GC_12_792 b_12 NI_12 NS_792 0 6.0578125670489723e-06
GC_12_793 b_12 NI_12 NS_793 0 5.7049766382441451e-06
GC_12_794 b_12 NI_12 NS_794 0 5.2024814563254172e-07
GC_12_795 b_12 NI_12 NS_795 0 5.9119937131346918e-11
GC_12_796 b_12 NI_12 NS_796 0 1.4784980651341332e-10
GC_12_797 b_12 NI_12 NS_797 0 5.9030980686065757e-09
GC_12_798 b_12 NI_12 NS_798 0 -8.4602307977119755e-09
GC_12_799 b_12 NI_12 NS_799 0 -1.1163639956902446e-04
GC_12_800 b_12 NI_12 NS_800 0 -2.1529158443370188e-06
GC_12_801 b_12 NI_12 NS_801 0 -2.4619850691498288e-10
GC_12_802 b_12 NI_12 NS_802 0 2.5690930378426494e-09
GC_12_803 b_12 NI_12 NS_803 0 1.8039278094274890e-06
GC_12_804 b_12 NI_12 NS_804 0 -1.6072975390178547e-06
GC_12_805 b_12 NI_12 NS_805 0 2.5854821322440738e-07
GC_12_806 b_12 NI_12 NS_806 0 -6.4503863632617060e-06
GC_12_807 b_12 NI_12 NS_807 0 -7.5446339054391656e-06
GC_12_808 b_12 NI_12 NS_808 0 -3.1551865989703316e-07
GC_12_809 b_12 NI_12 NS_809 0 -1.4480433164999897e-06
GC_12_810 b_12 NI_12 NS_810 0 -4.6837952212256389e-06
GC_12_811 b_12 NI_12 NS_811 0 -1.5899387288290652e-05
GC_12_812 b_12 NI_12 NS_812 0 -1.9736059299108864e-06
GC_12_813 b_12 NI_12 NS_813 0 -7.0460530110226972e-06
GC_12_814 b_12 NI_12 NS_814 0 1.8943204714084397e-05
GC_12_815 b_12 NI_12 NS_815 0 4.8825936284962925e-06
GC_12_816 b_12 NI_12 NS_816 0 -2.8766000285347546e-06
GC_12_817 b_12 NI_12 NS_817 0 -1.3982138614898641e-07
GC_12_818 b_12 NI_12 NS_818 0 -2.4404302188285432e-06
GC_12_819 b_12 NI_12 NS_819 0 -2.6317281677602781e-05
GC_12_820 b_12 NI_12 NS_820 0 2.8135822450975784e-05
GC_12_821 b_12 NI_12 NS_821 0 2.8104646088880103e-05
GC_12_822 b_12 NI_12 NS_822 0 -7.9688312860341651e-06
GC_12_823 b_12 NI_12 NS_823 0 -8.0936118314964572e-06
GC_12_824 b_12 NI_12 NS_824 0 -4.2239602905232557e-06
GC_12_825 b_12 NI_12 NS_825 0 1.2266611890990659e-05
GC_12_826 b_12 NI_12 NS_826 0 2.7177893305785217e-05
GC_12_827 b_12 NI_12 NS_827 0 1.4632392613682324e-06
GC_12_828 b_12 NI_12 NS_828 0 -8.8115824074875114e-06
GC_12_829 b_12 NI_12 NS_829 0 -2.8379259765416538e-05
GC_12_830 b_12 NI_12 NS_830 0 4.7636963102827415e-06
GC_12_831 b_12 NI_12 NS_831 0 4.1223376017897051e-05
GC_12_832 b_12 NI_12 NS_832 0 1.0997307186005501e-05
GC_12_833 b_12 NI_12 NS_833 0 -2.9904642862790358e-06
GC_12_834 b_12 NI_12 NS_834 0 -4.3573147748178563e-06
GC_12_835 b_12 NI_12 NS_835 0 1.2935785848030450e-05
GC_12_836 b_12 NI_12 NS_836 0 1.9156001319982458e-05
GC_12_837 b_12 NI_12 NS_837 0 3.7957746011730851e-06
GC_12_838 b_12 NI_12 NS_838 0 -1.0819255573967233e-05
GC_12_839 b_12 NI_12 NS_839 0 -6.4497759600160374e-06
GC_12_840 b_12 NI_12 NS_840 0 9.6990791576127238e-07
GC_12_841 b_12 NI_12 NS_841 0 1.8939860741293300e-05
GC_12_842 b_12 NI_12 NS_842 0 5.5256305510178568e-06
GC_12_843 b_12 NI_12 NS_843 0 -1.0369487720202447e-07
GC_12_844 b_12 NI_12 NS_844 0 -4.1120694563082956e-06
GC_12_845 b_12 NI_12 NS_845 0 4.9329507761176971e-06
GC_12_846 b_12 NI_12 NS_846 0 1.4409307475536643e-05
GC_12_847 b_12 NI_12 NS_847 0 7.8206607745771561e-06
GC_12_848 b_12 NI_12 NS_848 0 -1.1148679773977570e-05
GC_12_849 b_12 NI_12 NS_849 0 -1.4169787380321721e-06
GC_12_850 b_12 NI_12 NS_850 0 9.8983547756725509e-07
GC_12_851 b_12 NI_12 NS_851 0 1.0881123917797364e-05
GC_12_852 b_12 NI_12 NS_852 0 4.1883217093672803e-06
GC_12_853 b_12 NI_12 NS_853 0 1.6989713567469147e-06
GC_12_854 b_12 NI_12 NS_854 0 -5.8201956701050483e-07
GC_12_855 b_12 NI_12 NS_855 0 5.6739379398359018e-06
GC_12_856 b_12 NI_12 NS_856 0 1.7280444088302890e-06
GC_12_857 b_12 NI_12 NS_857 0 3.3535643637889036e-06
GC_12_858 b_12 NI_12 NS_858 0 2.0815596861234222e-06
GC_12_859 b_12 NI_12 NS_859 0 1.0938037528366697e-05
GC_12_860 b_12 NI_12 NS_860 0 3.8462784458899466e-06
GC_12_861 b_12 NI_12 NS_861 0 4.8353426129201777e-06
GC_12_862 b_12 NI_12 NS_862 0 -4.4521259886180949e-08
GC_12_863 b_12 NI_12 NS_863 0 9.9616050540157620e-06
GC_12_864 b_12 NI_12 NS_864 0 -1.0482432472255300e-06
GC_12_865 b_12 NI_12 NS_865 0 8.1946746222199797e-06
GC_12_866 b_12 NI_12 NS_866 0 2.9799205730145754e-06
GC_12_867 b_12 NI_12 NS_867 0 1.9009426587687409e-05
GC_12_868 b_12 NI_12 NS_868 0 -5.5028969399128096e-06
GC_12_869 b_12 NI_12 NS_869 0 7.1831606099636413e-06
GC_12_870 b_12 NI_12 NS_870 0 -3.9855818619096081e-06
GC_12_871 b_12 NI_12 NS_871 0 1.3697382318393967e-05
GC_12_872 b_12 NI_12 NS_872 0 -1.1862008955010945e-05
GC_12_873 b_12 NI_12 NS_873 0 1.2345387857721778e-05
GC_12_874 b_12 NI_12 NS_874 0 -3.9388169194214806e-06
GC_12_875 b_12 NI_12 NS_875 0 9.1353073663964032e-06
GC_12_876 b_12 NI_12 NS_876 0 -2.6714433636524114e-05
GC_12_877 b_12 NI_12 NS_877 0 2.3416332402385855e-06
GC_12_878 b_12 NI_12 NS_878 0 -1.2350035931808488e-05
GC_12_879 b_12 NI_12 NS_879 0 -8.3090395478994854e-06
GC_12_880 b_12 NI_12 NS_880 0 -1.8612842117988349e-05
GC_12_881 b_12 NI_12 NS_881 0 -4.9202384588984253e-06
GC_12_882 b_12 NI_12 NS_882 0 -1.2088815641521426e-05
GC_12_883 b_12 NI_12 NS_883 0 5.4869188421914613e-05
GC_12_884 b_12 NI_12 NS_884 0 -8.7931495102408312e-05
GC_12_885 b_12 NI_12 NS_885 0 -1.0053081392043435e-05
GC_12_886 b_12 NI_12 NS_886 0 1.3554290769003837e-06
GC_12_887 b_12 NI_12 NS_887 0 3.9049610860830325e-07
GC_12_888 b_12 NI_12 NS_888 0 -1.2503197228092230e-07
GC_12_889 b_12 NI_12 NS_889 0 -2.7269125758406371e-06
GC_12_890 b_12 NI_12 NS_890 0 -1.9374888782726351e-06
GC_12_891 b_12 NI_12 NS_891 0 -4.4052554126708421e-06
GC_12_892 b_12 NI_12 NS_892 0 5.8881526725845959e-07
GC_12_893 b_12 NI_12 NS_893 0 -1.7470998450749979e-05
GC_12_894 b_12 NI_12 NS_894 0 9.5706311282159067e-06
GC_12_895 b_12 NI_12 NS_895 0 -9.2073298612844986e-06
GC_12_896 b_12 NI_12 NS_896 0 3.7347453602385911e-05
GC_12_897 b_12 NI_12 NS_897 0 -7.2389890523814598e-06
GC_12_898 b_12 NI_12 NS_898 0 3.3305381361767945e-07
GC_12_899 b_12 NI_12 NS_899 0 -1.3385051586372787e-05
GC_12_900 b_12 NI_12 NS_900 0 1.8624028953697874e-06
GC_12_901 b_12 NI_12 NS_901 0 -4.6430381925861289e-06
GC_12_902 b_12 NI_12 NS_902 0 -3.3916906441230176e-06
GC_12_903 b_12 NI_12 NS_903 0 -6.3994045210883496e-06
GC_12_904 b_12 NI_12 NS_904 0 1.0401448644932981e-06
GC_12_905 b_12 NI_12 NS_905 0 -3.0542884836509914e-06
GC_12_906 b_12 NI_12 NS_906 0 8.8891069345259925e-07
GC_12_907 b_12 NI_12 NS_907 0 -1.7965416764847646e-06
GC_12_908 b_12 NI_12 NS_908 0 -9.3478378023655773e-07
GC_12_909 b_12 NI_12 NS_909 0 -2.6064291861265451e-10
GC_12_910 b_12 NI_12 NS_910 0 4.2284173671267930e-10
GC_12_911 b_12 NI_12 NS_911 0 2.3336442882807486e-09
GC_12_912 b_12 NI_12 NS_912 0 -2.6682895333200740e-08
GC_12_913 b_12 NI_12 NS_913 0 2.9495811923537503e-03
GC_12_914 b_12 NI_12 NS_914 0 -6.1234115659838733e-04
GC_12_915 b_12 NI_12 NS_915 0 2.7950026882784402e-08
GC_12_916 b_12 NI_12 NS_916 0 -3.1703308810825566e-08
GC_12_917 b_12 NI_12 NS_917 0 2.0347267665788766e-04
GC_12_918 b_12 NI_12 NS_918 0 1.3799476263531450e-04
GC_12_919 b_12 NI_12 NS_919 0 5.6259278931877776e-04
GC_12_920 b_12 NI_12 NS_920 0 2.6570822064798239e-04
GC_12_921 b_12 NI_12 NS_921 0 3.1064663995017498e-03
GC_12_922 b_12 NI_12 NS_922 0 -2.2048923377993046e-03
GC_12_923 b_12 NI_12 NS_923 0 -1.5822544729057781e-03
GC_12_924 b_12 NI_12 NS_924 0 -2.6870781195163086e-03
GC_12_925 b_12 NI_12 NS_925 0 -2.0496561562222395e-03
GC_12_926 b_12 NI_12 NS_926 0 -3.7885098699826916e-03
GC_12_927 b_12 NI_12 NS_927 0 -4.9745617115417714e-03
GC_12_928 b_12 NI_12 NS_928 0 -1.5415300338808607e-03
GC_12_929 b_12 NI_12 NS_929 0 2.9290591387105765e-04
GC_12_930 b_12 NI_12 NS_930 0 1.9565149964029271e-04
GC_12_931 b_12 NI_12 NS_931 0 -2.8663291194968620e-03
GC_12_932 b_12 NI_12 NS_932 0 -9.5746315591239452e-04
GC_12_933 b_12 NI_12 NS_933 0 -2.2151872823810342e-02
GC_12_934 b_12 NI_12 NS_934 0 -1.0226311652202039e-02
GC_12_935 b_12 NI_12 NS_935 0 1.1325012348957109e-03
GC_12_936 b_12 NI_12 NS_936 0 2.0395319985909609e-02
GC_12_937 b_12 NI_12 NS_937 0 -5.8416198952844101e-03
GC_12_938 b_12 NI_12 NS_938 0 4.6116305224392935e-03
GC_12_939 b_12 NI_12 NS_939 0 5.7171588852187212e-03
GC_12_940 b_12 NI_12 NS_940 0 3.4516068686460233e-02
GC_12_941 b_12 NI_12 NS_941 0 8.0342767432026105e-03
GC_12_942 b_12 NI_12 NS_942 0 2.7930216049210652e-03
GC_12_943 b_12 NI_12 NS_943 0 -7.7724132610304912e-03
GC_12_944 b_12 NI_12 NS_944 0 2.9556755329158468e-02
GC_12_945 b_12 NI_12 NS_945 0 5.0768422614967855e-02
GC_12_946 b_12 NI_12 NS_946 0 -2.0072973634987768e-02
GC_12_947 b_12 NI_12 NS_947 0 7.9195777573987172e-03
GC_12_948 b_12 NI_12 NS_948 0 -1.6364431156656145e-03
GC_12_949 b_12 NI_12 NS_949 0 2.9084851985046272e-02
GC_12_950 b_12 NI_12 NS_950 0 -2.6464742843239800e-02
GC_12_951 b_12 NI_12 NS_951 0 -6.7250699728445820e-03
GC_12_952 b_12 NI_12 NS_952 0 -9.8822034205078412e-03
GC_12_953 b_12 NI_12 NS_953 0 8.4630802992458967e-03
GC_12_954 b_12 NI_12 NS_954 0 -8.0277999864013534e-03
GC_12_955 b_12 NI_12 NS_955 0 -1.8994958080501462e-02
GC_12_956 b_12 NI_12 NS_956 0 -2.5238416401433643e-02
GC_12_957 b_12 NI_12 NS_957 0 -5.4717856759026956e-03
GC_12_958 b_12 NI_12 NS_958 0 -2.8547826260518659e-03
GC_12_959 b_12 NI_12 NS_959 0 -1.7741076973119479e-02
GC_12_960 b_12 NI_12 NS_960 0 -1.3132225702361526e-02
GC_12_961 b_12 NI_12 NS_961 0 -4.8177974095531375e-03
GC_12_962 b_12 NI_12 NS_962 0 1.2541405032616580e-02
GC_12_963 b_12 NI_12 NS_963 0 -3.4590897682977135e-03
GC_12_964 b_12 NI_12 NS_964 0 1.5412389403709550e-03
GC_12_965 b_12 NI_12 NS_965 0 -7.1865040307237684e-04
GC_12_966 b_12 NI_12 NS_966 0 7.0058608632081959e-03
GC_12_967 b_12 NI_12 NS_967 0 1.8820413111284692e-03
GC_12_968 b_12 NI_12 NS_968 0 8.5748332402728843e-05
GC_12_969 b_12 NI_12 NS_969 0 3.1400233506648391e-04
GC_12_970 b_12 NI_12 NS_970 0 -1.9467013336808764e-03
GC_12_971 b_12 NI_12 NS_971 0 -1.8563359956212089e-03
GC_12_972 b_12 NI_12 NS_972 0 -1.6182084458853004e-03
GC_12_973 b_12 NI_12 NS_973 0 -2.1290963442455913e-03
GC_12_974 b_12 NI_12 NS_974 0 1.6850444052401595e-03
GC_12_975 b_12 NI_12 NS_975 0 7.6361045378036958e-04
GC_12_976 b_12 NI_12 NS_976 0 1.8527551166551114e-04
GC_12_977 b_12 NI_12 NS_977 0 -6.9730355587067818e-04
GC_12_978 b_12 NI_12 NS_978 0 -1.6780696740443422e-03
GC_12_979 b_12 NI_12 NS_979 0 -2.6815284254526951e-03
GC_12_980 b_12 NI_12 NS_980 0 -8.2749066372070986e-04
GC_12_981 b_12 NI_12 NS_981 0 -4.9989598792736208e-04
GC_12_982 b_12 NI_12 NS_982 0 2.9288646850935069e-03
GC_12_983 b_12 NI_12 NS_983 0 1.3533577668197651e-03
GC_12_984 b_12 NI_12 NS_984 0 -8.5805585761030421e-04
GC_12_985 b_12 NI_12 NS_985 0 -2.4189246450171541e-03
GC_12_986 b_12 NI_12 NS_986 0 -2.2676208543534783e-03
GC_12_987 b_12 NI_12 NS_987 0 -3.5540457637606737e-03
GC_12_988 b_12 NI_12 NS_988 0 7.4852698048109346e-04
GC_12_989 b_12 NI_12 NS_989 0 2.4633831805098857e-03
GC_12_990 b_12 NI_12 NS_990 0 3.0182806332560239e-03
GC_12_991 b_12 NI_12 NS_991 0 9.8455403748817978e-04
GC_12_992 b_12 NI_12 NS_992 0 -2.9418095517291603e-03
GC_12_993 b_12 NI_12 NS_993 0 -4.7677995915481408e-03
GC_12_994 b_12 NI_12 NS_994 0 5.4340716195029563e-05
GC_12_995 b_12 NI_12 NS_995 0 -1.7083701125203245e-03
GC_12_996 b_12 NI_12 NS_996 0 3.7124272306012156e-03
GC_12_997 b_12 NI_12 NS_997 0 -7.6587238473877178e-04
GC_12_998 b_12 NI_12 NS_998 0 1.5006822641626277e-03
GC_12_999 b_12 NI_12 NS_999 0 3.2213016220089701e-03
GC_12_1000 b_12 NI_12 NS_1000 0 -1.3508686296772930e-03
GC_12_1001 b_12 NI_12 NS_1001 0 -2.9326246015476770e-06
GC_12_1002 b_12 NI_12 NS_1002 0 8.7469681182399162e-06
GC_12_1003 b_12 NI_12 NS_1003 0 -1.8200423308688235e-03
GC_12_1004 b_12 NI_12 NS_1004 0 -2.5277362718432702e-03
GC_12_1005 b_12 NI_12 NS_1005 0 -2.4072536539359278e-03
GC_12_1006 b_12 NI_12 NS_1006 0 2.4886640702112216e-03
GC_12_1007 b_12 NI_12 NS_1007 0 1.0142609812203104e-03
GC_12_1008 b_12 NI_12 NS_1008 0 2.4256812294375782e-03
GC_12_1009 b_12 NI_12 NS_1009 0 8.5775820128619075e-04
GC_12_1010 b_12 NI_12 NS_1010 0 -2.6994845972613747e-03
GC_12_1011 b_12 NI_12 NS_1011 0 -3.0644790052722354e-04
GC_12_1012 b_12 NI_12 NS_1012 0 1.6741355470716673e-03
GC_12_1013 b_12 NI_12 NS_1013 0 -1.7840541403943862e-03
GC_12_1014 b_12 NI_12 NS_1014 0 -3.1181108525964879e-04
GC_12_1015 b_12 NI_12 NS_1015 0 1.4004540369615714e-03
GC_12_1016 b_12 NI_12 NS_1016 0 1.9709615364841082e-03
GC_12_1017 b_12 NI_12 NS_1017 0 1.0449287337610698e-03
GC_12_1018 b_12 NI_12 NS_1018 0 -2.2998046396501296e-03
GC_12_1019 b_12 NI_12 NS_1019 0 -6.9799493598442762e-04
GC_12_1020 b_12 NI_12 NS_1020 0 -1.4668898760807985e-03
GC_12_1021 b_12 NI_12 NS_1021 0 -1.3735490956513384e-03
GC_12_1022 b_12 NI_12 NS_1022 0 -3.1252859531712319e-04
GC_12_1023 b_12 NI_12 NS_1023 0 7.1030487116399009e-09
GC_12_1024 b_12 NI_12 NS_1024 0 -2.4709966318857688e-08
GC_12_1025 b_12 NI_12 NS_1025 0 -4.5275596677154549e-07
GC_12_1026 b_12 NI_12 NS_1026 0 1.6341837962880834e-06
GC_12_1027 b_12 NI_12 NS_1027 0 7.7517847499170159e-03
GC_12_1028 b_12 NI_12 NS_1028 0 -1.6012309488680962e-03
GC_12_1029 b_12 NI_12 NS_1029 0 -1.2107357777372096e-08
GC_12_1030 b_12 NI_12 NS_1030 0 -8.8419733076225256e-07
GC_12_1031 b_12 NI_12 NS_1031 0 1.0389334678062627e-04
GC_12_1032 b_12 NI_12 NS_1032 0 -5.1165497914171124e-04
GC_12_1033 b_12 NI_12 NS_1033 0 -1.9366722490404861e-03
GC_12_1034 b_12 NI_12 NS_1034 0 -5.9740611531078726e-04
GC_12_1035 b_12 NI_12 NS_1035 0 2.9415496646425054e-03
GC_12_1036 b_12 NI_12 NS_1036 0 2.2646150034249767e-03
GC_12_1037 b_12 NI_12 NS_1037 0 -3.5699560029939215e-03
GC_12_1038 b_12 NI_12 NS_1038 0 -3.0486859049663247e-03
GC_12_1039 b_12 NI_12 NS_1039 0 -1.7071461899168785e-03
GC_12_1040 b_12 NI_12 NS_1040 0 5.8436823019121995e-03
GC_12_1041 b_12 NI_12 NS_1041 0 4.3687526632687481e-03
GC_12_1042 b_12 NI_12 NS_1042 0 -2.4746080186911204e-03
GC_12_1043 b_12 NI_12 NS_1043 0 -1.1051345529748483e-04
GC_12_1044 b_12 NI_12 NS_1044 0 -1.0368748323576710e-04
GC_12_1045 b_12 NI_12 NS_1045 0 -4.4520077614426962e-03
GC_12_1046 b_12 NI_12 NS_1046 0 -9.2458271011306489e-04
GC_12_1047 b_12 NI_12 NS_1047 0 9.1257545990865822e-03
GC_12_1048 b_12 NI_12 NS_1048 0 1.7785323756134501e-02
GC_12_1049 b_12 NI_12 NS_1049 0 -4.0274383895260472e-03
GC_12_1050 b_12 NI_12 NS_1050 0 -1.7847938779750171e-02
GC_12_1051 b_12 NI_12 NS_1051 0 -8.2175426840414220e-03
GC_12_1052 b_12 NI_12 NS_1052 0 4.1736400791754745e-03
GC_12_1053 b_12 NI_12 NS_1053 0 1.7064437340061158e-02
GC_12_1054 b_12 NI_12 NS_1054 0 -4.4006004129026351e-04
GC_12_1055 b_12 NI_12 NS_1055 0 -9.2787957944330327e-03
GC_12_1056 b_12 NI_12 NS_1056 0 -3.2071931228853856e-03
GC_12_1057 b_12 NI_12 NS_1057 0 -1.3712649598663747e-02
GC_12_1058 b_12 NI_12 NS_1058 0 2.2836660703413933e-02
GC_12_1059 b_12 NI_12 NS_1059 0 2.2839352234485612e-02
GC_12_1060 b_12 NI_12 NS_1060 0 -2.2670699964558446e-02
GC_12_1061 b_12 NI_12 NS_1061 0 -9.2392572266461817e-03
GC_12_1062 b_12 NI_12 NS_1062 0 9.0801649156133394e-04
GC_12_1063 b_12 NI_12 NS_1063 0 1.8480444531579071e-02
GC_12_1064 b_12 NI_12 NS_1064 0 6.2433949828427978e-03
GC_12_1065 b_12 NI_12 NS_1065 0 -9.1763265309292540e-03
GC_12_1066 b_12 NI_12 NS_1066 0 -9.4611036353866654e-03
GC_12_1067 b_12 NI_12 NS_1067 0 -9.9741831229017731e-03
GC_12_1068 b_12 NI_12 NS_1068 0 6.3961404491676768e-03
GC_12_1069 b_12 NI_12 NS_1069 0 1.6838378743727202e-02
GC_12_1070 b_12 NI_12 NS_1070 0 -4.8507571343212380e-03
GC_12_1071 b_12 NI_12 NS_1071 0 -7.2149766097673847e-03
GC_12_1072 b_12 NI_12 NS_1072 0 -3.4093170377388717e-03
GC_12_1073 b_12 NI_12 NS_1073 0 6.8284598867650887e-03
GC_12_1074 b_12 NI_12 NS_1074 0 1.3296718008884172e-02
GC_12_1075 b_12 NI_12 NS_1075 0 -1.8198422883981729e-03
GC_12_1076 b_12 NI_12 NS_1076 0 -1.4401884747287253e-02
GC_12_1077 b_12 NI_12 NS_1077 0 -4.9859624292220989e-03
GC_12_1078 b_12 NI_12 NS_1078 0 1.0394192940170717e-03
GC_12_1079 b_12 NI_12 NS_1079 0 6.0026872519342465e-03
GC_12_1080 b_12 NI_12 NS_1080 0 -1.1033379851630248e-03
GC_12_1081 b_12 NI_12 NS_1081 0 -3.4642736715962620e-03
GC_12_1082 b_12 NI_12 NS_1082 0 -1.0877132921067421e-03
GC_12_1083 b_12 NI_12 NS_1083 0 2.7180843228181684e-03
GC_12_1084 b_12 NI_12 NS_1084 0 -5.0793073185757961e-04
GC_12_1085 b_12 NI_12 NS_1085 0 -3.2964042307125105e-03
GC_12_1086 b_12 NI_12 NS_1086 0 -2.8952142993826703e-03
GC_12_1087 b_12 NI_12 NS_1087 0 2.0160582918145454e-03
GC_12_1088 b_12 NI_12 NS_1088 0 7.7561412799337750e-04
GC_12_1089 b_12 NI_12 NS_1089 0 -2.0162391613304334e-03
GC_12_1090 b_12 NI_12 NS_1090 0 -9.6653840622365960e-04
GC_12_1091 b_12 NI_12 NS_1091 0 2.1216791622888586e-03
GC_12_1092 b_12 NI_12 NS_1092 0 -1.4710192928709600e-03
GC_12_1093 b_12 NI_12 NS_1093 0 -4.1846667586610238e-03
GC_12_1094 b_12 NI_12 NS_1094 0 -1.8129789192783327e-03
GC_12_1095 b_12 NI_12 NS_1095 0 2.3699521136967103e-03
GC_12_1096 b_12 NI_12 NS_1096 0 -3.7091804134262553e-04
GC_12_1097 b_12 NI_12 NS_1097 0 -3.0171283246533732e-03
GC_12_1098 b_12 NI_12 NS_1098 0 4.6227809629516509e-04
GC_12_1099 b_12 NI_12 NS_1099 0 2.7066143487306546e-03
GC_12_1100 b_12 NI_12 NS_1100 0 -2.7283529759322355e-03
GC_12_1101 b_12 NI_12 NS_1101 0 -5.0391230855239780e-03
GC_12_1102 b_12 NI_12 NS_1102 0 -1.2777907301728678e-04
GC_12_1103 b_12 NI_12 NS_1103 0 2.4350369276882520e-03
GC_12_1104 b_12 NI_12 NS_1104 0 -2.1722372652505104e-03
GC_12_1105 b_12 NI_12 NS_1105 0 -3.2447335282912138e-03
GC_12_1106 b_12 NI_12 NS_1106 0 2.6004818072975023e-03
GC_12_1107 b_12 NI_12 NS_1107 0 1.7440002919609180e-03
GC_12_1108 b_12 NI_12 NS_1108 0 -4.7506629812880483e-03
GC_12_1109 b_12 NI_12 NS_1109 0 -3.6334526772605338e-03
GC_12_1110 b_12 NI_12 NS_1110 0 2.5968941596526359e-03
GC_12_1111 b_12 NI_12 NS_1111 0 -2.8337529740661100e-03
GC_12_1112 b_12 NI_12 NS_1112 0 3.9869956619756628e-03
GC_12_1113 b_12 NI_12 NS_1113 0 -2.2097510891847568e-04
GC_12_1114 b_12 NI_12 NS_1114 0 -4.2143869040275625e-03
GC_12_1115 b_12 NI_12 NS_1115 0 -9.9004394496546137e-06
GC_12_1116 b_12 NI_12 NS_1116 0 7.5069812216699512e-06
GC_12_1117 b_12 NI_12 NS_1117 0 -1.3536762359922386e-03
GC_12_1118 b_12 NI_12 NS_1118 0 3.3750405193467914e-03
GC_12_1119 b_12 NI_12 NS_1119 0 -9.6980990466620704e-04
GC_12_1120 b_12 NI_12 NS_1120 0 -4.3483855057119842e-03
GC_12_1121 b_12 NI_12 NS_1121 0 -1.0004341440310088e-03
GC_12_1122 b_12 NI_12 NS_1122 0 2.2215368758935518e-03
GC_12_1123 b_12 NI_12 NS_1123 0 -1.6509401654640809e-03
GC_12_1124 b_12 NI_12 NS_1124 0 -4.4091665541923213e-03
GC_12_1125 b_12 NI_12 NS_1125 0 -1.4483893071172741e-03
GC_12_1126 b_12 NI_12 NS_1126 0 -2.4971174640467746e-03
GC_12_1127 b_12 NI_12 NS_1127 0 7.8206336442820132e-04
GC_12_1128 b_12 NI_12 NS_1128 0 2.5934675449305398e-03
GC_12_1129 b_12 NI_12 NS_1129 0 -6.9629910872305936e-04
GC_12_1130 b_12 NI_12 NS_1130 0 2.8791307009012439e-03
GC_12_1131 b_12 NI_12 NS_1131 0 -1.4354331452083717e-03
GC_12_1132 b_12 NI_12 NS_1132 0 -2.7718928615064744e-03
GC_12_1133 b_12 NI_12 NS_1133 0 -1.1678458093011066e-03
GC_12_1134 b_12 NI_12 NS_1134 0 2.6661739013163592e-03
GC_12_1135 b_12 NI_12 NS_1135 0 7.8077011825160422e-04
GC_12_1136 b_12 NI_12 NS_1136 0 -1.8746307413896343e-03
GC_12_1137 b_12 NI_12 NS_1137 0 2.3791496125744685e-08
GC_12_1138 b_12 NI_12 NS_1138 0 -6.0255366166095534e-08
GC_12_1139 b_12 NI_12 NS_1139 0 -9.0379586952661370e-07
GC_12_1140 b_12 NI_12 NS_1140 0 3.2032341124455259e-06
GC_12_1141 b_12 NI_12 NS_1141 0 1.8226639093394684e-02
GC_12_1142 b_12 NI_12 NS_1142 0 6.7518776709956860e-03
GC_12_1143 b_12 NI_12 NS_1143 0 4.8241143035689224e-07
GC_12_1144 b_12 NI_12 NS_1144 0 1.4304300339185533e-06
GC_12_1145 b_12 NI_12 NS_1145 0 6.0825405603485419e-03
GC_12_1146 b_12 NI_12 NS_1146 0 1.8255053945468356e-03
GC_12_1147 b_12 NI_12 NS_1147 0 -6.0663181448941395e-03
GC_12_1148 b_12 NI_12 NS_1148 0 -6.4128061695591120e-04
GC_12_1149 b_12 NI_12 NS_1149 0 7.3354121902149830e-03
GC_12_1150 b_12 NI_12 NS_1150 0 -1.2858493899287247e-02
GC_12_1151 b_12 NI_12 NS_1151 0 8.4355047267817528e-03
GC_12_1152 b_12 NI_12 NS_1152 0 -2.1170237010923596e-04
GC_12_1153 b_12 NI_12 NS_1153 0 -9.6680399981822849e-03
GC_12_1154 b_12 NI_12 NS_1154 0 2.5853163610514290e-03
GC_12_1155 b_12 NI_12 NS_1155 0 -8.8082205211286891e-03
GC_12_1156 b_12 NI_12 NS_1156 0 -2.4395146957781177e-02
GC_12_1157 b_12 NI_12 NS_1157 0 -8.6844452878820507e-04
GC_12_1158 b_12 NI_12 NS_1158 0 4.1759611871123583e-03
GC_12_1159 b_12 NI_12 NS_1159 0 7.1854566561496561e-03
GC_12_1160 b_12 NI_12 NS_1160 0 -9.9750534028919058e-04
GC_12_1161 b_12 NI_12 NS_1161 0 -2.5220033152065183e-02
GC_12_1162 b_12 NI_12 NS_1162 0 4.8139715760926426e-03
GC_12_1163 b_12 NI_12 NS_1163 0 -1.9618700342314742e-02
GC_12_1164 b_12 NI_12 NS_1164 0 8.5375016577444974e-04
GC_12_1165 b_12 NI_12 NS_1165 0 1.0773083089171369e-02
GC_12_1166 b_12 NI_12 NS_1166 0 -2.7351328266457869e-03
GC_12_1167 b_12 NI_12 NS_1167 0 -4.8274331748894110e-03
GC_12_1168 b_12 NI_12 NS_1168 0 4.5019657860878526e-02
GC_12_1169 b_12 NI_12 NS_1169 0 -1.2641951741045121e-02
GC_12_1170 b_12 NI_12 NS_1170 0 -3.2177142892545000e-04
GC_12_1171 b_12 NI_12 NS_1171 0 1.5975052597574597e-02
GC_12_1172 b_12 NI_12 NS_1172 0 -3.9761180146722459e-03
GC_12_1173 b_12 NI_12 NS_1173 0 3.2145985308246819e-02
GC_12_1174 b_12 NI_12 NS_1174 0 1.8555887119905006e-02
GC_12_1175 b_12 NI_12 NS_1175 0 -1.2595033819510692e-02
GC_12_1176 b_12 NI_12 NS_1176 0 1.1576674860419586e-04
GC_12_1177 b_12 NI_12 NS_1177 0 1.7252012112863979e-02
GC_12_1178 b_12 NI_12 NS_1178 0 -3.5175566351817462e-02
GC_12_1179 b_12 NI_12 NS_1179 0 1.3984153722119754e-02
GC_12_1180 b_12 NI_12 NS_1180 0 4.8235598624010853e-03
GC_12_1181 b_12 NI_12 NS_1181 0 -1.4410981988279451e-02
GC_12_1182 b_12 NI_12 NS_1182 0 1.9254056886641588e-04
GC_12_1183 b_12 NI_12 NS_1183 0 -2.0123965939243461e-02
GC_12_1184 b_12 NI_12 NS_1184 0 -3.0196899562290620e-02
GC_12_1185 b_12 NI_12 NS_1185 0 1.0516107326877347e-02
GC_12_1186 b_12 NI_12 NS_1186 0 3.6210484291599528e-03
GC_12_1187 b_12 NI_12 NS_1187 0 -2.6839278492696038e-02
GC_12_1188 b_12 NI_12 NS_1188 0 1.1127542052905087e-02
GC_12_1189 b_12 NI_12 NS_1189 0 -1.4106844356102309e-02
GC_12_1190 b_12 NI_12 NS_1190 0 -2.5293245626218609e-03
GC_12_1191 b_12 NI_12 NS_1191 0 7.5511418333626982e-03
GC_12_1192 b_12 NI_12 NS_1192 0 1.6110774945834250e-03
GC_12_1193 b_12 NI_12 NS_1193 0 -8.7782701212020119e-04
GC_12_1194 b_12 NI_12 NS_1194 0 2.4406558785406349e-02
GC_12_1195 b_12 NI_12 NS_1195 0 -7.6159479844090496e-03
GC_12_1196 b_12 NI_12 NS_1196 0 2.7283646786539165e-04
GC_12_1197 b_12 NI_12 NS_1197 0 -5.5396264048151707e-04
GC_12_1198 b_12 NI_12 NS_1198 0 -5.5347231376909212e-03
GC_12_1199 b_12 NI_12 NS_1199 0 8.2549283975567392e-03
GC_12_1200 b_12 NI_12 NS_1200 0 7.0292117623693973e-03
GC_12_1201 b_12 NI_12 NS_1201 0 -7.2657101415801034e-04
GC_12_1202 b_12 NI_12 NS_1202 0 1.2096321415939807e-02
GC_12_1203 b_12 NI_12 NS_1203 0 -5.1449891401495092e-03
GC_12_1204 b_12 NI_12 NS_1204 0 -1.3733042392405142e-04
GC_12_1205 b_12 NI_12 NS_1205 0 -1.8277729450042253e-03
GC_12_1206 b_12 NI_12 NS_1206 0 -5.1663248385474788e-03
GC_12_1207 b_12 NI_12 NS_1207 0 9.2805749594231345e-03
GC_12_1208 b_12 NI_12 NS_1208 0 5.4202516905103304e-03
GC_12_1209 b_12 NI_12 NS_1209 0 3.5140132276833143e-03
GC_12_1210 b_12 NI_12 NS_1210 0 1.1697043619558700e-02
GC_12_1211 b_12 NI_12 NS_1211 0 -6.1352206029401755e-03
GC_12_1212 b_12 NI_12 NS_1212 0 1.4323530175782008e-03
GC_12_1213 b_12 NI_12 NS_1213 0 -2.8179237740261665e-03
GC_12_1214 b_12 NI_12 NS_1214 0 -7.3385782251106143e-03
GC_12_1215 b_12 NI_12 NS_1215 0 9.9490799174609245e-03
GC_12_1216 b_12 NI_12 NS_1216 0 3.3702684406488243e-03
GC_12_1217 b_12 NI_12 NS_1217 0 8.1727927555613599e-03
GC_12_1218 b_12 NI_12 NS_1218 0 1.0256589319640713e-02
GC_12_1219 b_12 NI_12 NS_1219 0 -6.9843490439527658e-03
GC_12_1220 b_12 NI_12 NS_1220 0 2.9456637906114637e-03
GC_12_1221 b_12 NI_12 NS_1221 0 -5.6338007845899377e-03
GC_12_1222 b_12 NI_12 NS_1222 0 -8.0802091203552931e-03
GC_12_1223 b_12 NI_12 NS_1223 0 9.8429116438253847e-03
GC_12_1224 b_12 NI_12 NS_1224 0 5.5987730382862119e-04
GC_12_1225 b_12 NI_12 NS_1225 0 -1.0787123152828785e-02
GC_12_1226 b_12 NI_12 NS_1226 0 1.2188567634707274e-02
GC_12_1227 b_12 NI_12 NS_1227 0 9.6751942866318188e-03
GC_12_1228 b_12 NI_12 NS_1228 0 5.0629076871176780e-03
GC_12_1229 b_12 NI_12 NS_1229 0 -1.9005129407479682e-05
GC_12_1230 b_12 NI_12 NS_1230 0 3.1757335584331043e-05
GC_12_1231 b_12 NI_12 NS_1231 0 -7.1154533732795486e-03
GC_12_1232 b_12 NI_12 NS_1232 0 4.4968905233308794e-03
GC_12_1233 b_12 NI_12 NS_1233 0 -7.6587589856546090e-03
GC_12_1234 b_12 NI_12 NS_1234 0 -5.3140671940495729e-03
GC_12_1235 b_12 NI_12 NS_1235 0 9.4989054768590906e-03
GC_12_1236 b_12 NI_12 NS_1236 0 -1.7109725485480957e-03
GC_12_1237 b_12 NI_12 NS_1237 0 1.2462859244544862e-02
GC_12_1238 b_12 NI_12 NS_1238 0 -1.3552597453282678e-03
GC_12_1239 b_12 NI_12 NS_1239 0 -5.0734387070050877e-03
GC_12_1240 b_12 NI_12 NS_1240 0 -2.7550314333347997e-03
GC_12_1241 b_12 NI_12 NS_1241 0 -2.2334869277598484e-03
GC_12_1242 b_12 NI_12 NS_1242 0 6.5927094573896014e-03
GC_12_1243 b_12 NI_12 NS_1243 0 8.9637862457898048e-03
GC_12_1244 b_12 NI_12 NS_1244 0 1.2891302023389909e-04
GC_12_1245 b_12 NI_12 NS_1245 0 1.2489967417731057e-02
GC_12_1246 b_12 NI_12 NS_1246 0 1.7707475547818529e-03
GC_12_1247 b_12 NI_12 NS_1247 0 -5.3740562519027984e-03
GC_12_1248 b_12 NI_12 NS_1248 0 4.1561440449526844e-03
GC_12_1249 b_12 NI_12 NS_1249 0 -1.8426481627097577e-03
GC_12_1250 b_12 NI_12 NS_1250 0 -5.6872687344525904e-03
GC_12_1251 b_12 NI_12 NS_1251 0 2.0880737894526377e-07
GC_12_1252 b_12 NI_12 NS_1252 0 -2.4392505773762896e-07
GC_12_1253 b_12 NI_12 NS_1253 0 -1.1440672652985343e-05
GC_12_1254 b_12 NI_12 NS_1254 0 1.8294494930963459e-05
GC_12_1255 b_12 NI_12 NS_1255 0 -1.3077626181952854e-02
GC_12_1256 b_12 NI_12 NS_1256 0 1.3851822870424048e-03
GC_12_1257 b_12 NI_12 NS_1257 0 -2.6206484157238340e-07
GC_12_1258 b_12 NI_12 NS_1258 0 -3.7495559724260936e-06
GC_12_1259 b_12 NI_12 NS_1259 0 -2.7819372045823895e-04
GC_12_1260 b_12 NI_12 NS_1260 0 4.6297784968865710e-04
GC_12_1261 b_12 NI_12 NS_1261 0 1.3195321554402561e-03
GC_12_1262 b_12 NI_12 NS_1262 0 5.4935775116447621e-04
GC_12_1263 b_12 NI_12 NS_1263 0 -2.7628705965086590e-03
GC_12_1264 b_12 NI_12 NS_1264 0 -8.1703054050138513e-04
GC_12_1265 b_12 NI_12 NS_1265 0 3.5326192481360827e-03
GC_12_1266 b_12 NI_12 NS_1266 0 2.5338002367322971e-03
GC_12_1267 b_12 NI_12 NS_1267 0 1.1824232660161515e-03
GC_12_1268 b_12 NI_12 NS_1268 0 -4.1997922523623775e-03
GC_12_1269 b_12 NI_12 NS_1269 0 -1.7498503089834598e-03
GC_12_1270 b_12 NI_12 NS_1270 0 2.6968800977730367e-03
GC_12_1271 b_12 NI_12 NS_1271 0 -3.1387333304569377e-04
GC_12_1272 b_12 NI_12 NS_1272 0 -1.8984121393572973e-04
GC_12_1273 b_12 NI_12 NS_1273 0 3.9674889269261139e-03
GC_12_1274 b_12 NI_12 NS_1274 0 2.9857839207264353e-04
GC_12_1275 b_12 NI_12 NS_1275 0 -7.4413975684283658e-03
GC_12_1276 b_12 NI_12 NS_1276 0 -1.3618339017549618e-02
GC_12_1277 b_12 NI_12 NS_1277 0 4.4052505494702032e-03
GC_12_1278 b_12 NI_12 NS_1278 0 1.3511458829104268e-02
GC_12_1279 b_12 NI_12 NS_1279 0 6.7110109769435052e-03
GC_12_1280 b_12 NI_12 NS_1280 0 -3.9862631677580074e-03
GC_12_1281 b_12 NI_12 NS_1281 0 -1.3390055117710622e-02
GC_12_1282 b_12 NI_12 NS_1282 0 6.9024316026100564e-04
GC_12_1283 b_12 NI_12 NS_1283 0 7.8426044093508635e-03
GC_12_1284 b_12 NI_12 NS_1284 0 1.8947671797552837e-03
GC_12_1285 b_12 NI_12 NS_1285 0 1.0544112092794908e-02
GC_12_1286 b_12 NI_12 NS_1286 0 -1.9595447135794454e-02
GC_12_1287 b_12 NI_12 NS_1287 0 -1.7809609065537284e-02
GC_12_1288 b_12 NI_12 NS_1288 0 1.9141982245256914e-02
GC_12_1289 b_12 NI_12 NS_1289 0 7.6787750431322301e-03
GC_12_1290 b_12 NI_12 NS_1290 0 -1.4142909528422200e-03
GC_12_1291 b_12 NI_12 NS_1291 0 -1.5647914336480159e-02
GC_12_1292 b_12 NI_12 NS_1292 0 -4.7614896901242943e-03
GC_12_1293 b_12 NI_12 NS_1293 0 8.0618573016897534e-03
GC_12_1294 b_12 NI_12 NS_1294 0 7.2869891809915488e-03
GC_12_1295 b_12 NI_12 NS_1295 0 8.1170047185717825e-03
GC_12_1296 b_12 NI_12 NS_1296 0 -5.9990832035981233e-03
GC_12_1297 b_12 NI_12 NS_1297 0 -1.3980586997120310e-02
GC_12_1298 b_12 NI_12 NS_1298 0 4.5682719333455584e-03
GC_12_1299 b_12 NI_12 NS_1299 0 6.2307820113008013e-03
GC_12_1300 b_12 NI_12 NS_1300 0 2.4081612519185852e-03
GC_12_1301 b_12 NI_12 NS_1301 0 -6.2859264355147959e-03
GC_12_1302 b_12 NI_12 NS_1302 0 -1.1107051557285348e-02
GC_12_1303 b_12 NI_12 NS_1303 0 2.1280730573091239e-03
GC_12_1304 b_12 NI_12 NS_1304 0 1.1947397205328898e-02
GC_12_1305 b_12 NI_12 NS_1305 0 4.2092178851989275e-03
GC_12_1306 b_12 NI_12 NS_1306 0 -1.1609522005069772e-03
GC_12_1307 b_12 NI_12 NS_1307 0 -4.9313045763675562e-03
GC_12_1308 b_12 NI_12 NS_1308 0 1.0532438103220748e-03
GC_12_1309 b_12 NI_12 NS_1309 0 3.0238807200198212e-03
GC_12_1310 b_12 NI_12 NS_1310 0 6.9985711643234534e-04
GC_12_1311 b_12 NI_12 NS_1311 0 -2.2205262517191529e-03
GC_12_1312 b_12 NI_12 NS_1312 0 4.9428581137969500e-04
GC_12_1313 b_12 NI_12 NS_1313 0 3.0655102801238135e-03
GC_12_1314 b_12 NI_12 NS_1314 0 2.3037302634440079e-03
GC_12_1315 b_12 NI_12 NS_1315 0 -1.5339091967095620e-03
GC_12_1316 b_12 NI_12 NS_1316 0 -6.6977447033590210e-04
GC_12_1317 b_12 NI_12 NS_1317 0 1.8873378600740025e-03
GC_12_1318 b_12 NI_12 NS_1318 0 6.8441649659154455e-04
GC_12_1319 b_12 NI_12 NS_1319 0 -1.5620993801147751e-03
GC_12_1320 b_12 NI_12 NS_1320 0 1.2263492645296385e-03
GC_12_1321 b_12 NI_12 NS_1321 0 3.9751893811779595e-03
GC_12_1322 b_12 NI_12 NS_1322 0 1.4060884820821051e-03
GC_12_1323 b_12 NI_12 NS_1323 0 -1.5528106206005340e-03
GC_12_1324 b_12 NI_12 NS_1324 0 7.4661566659642788e-05
GC_12_1325 b_12 NI_12 NS_1325 0 2.8290380091208853e-03
GC_12_1326 b_12 NI_12 NS_1326 0 -6.8616923824479188e-04
GC_12_1327 b_12 NI_12 NS_1327 0 -1.8781833910551673e-03
GC_12_1328 b_12 NI_12 NS_1328 0 2.0100728806588782e-03
GC_12_1329 b_12 NI_12 NS_1329 0 4.9079320153830076e-03
GC_12_1330 b_12 NI_12 NS_1330 0 -1.8215321236888759e-04
GC_12_1331 b_12 NI_12 NS_1331 0 -1.6564588825831404e-03
GC_12_1332 b_12 NI_12 NS_1332 0 9.3019323073804548e-04
GC_12_1333 b_12 NI_12 NS_1333 0 3.0643003907121183e-03
GC_12_1334 b_12 NI_12 NS_1334 0 -2.8465101716221132e-03
GC_12_1335 b_12 NI_12 NS_1335 0 -1.4568553769455520e-03
GC_12_1336 b_12 NI_12 NS_1336 0 3.2233613952241500e-03
GC_12_1337 b_12 NI_12 NS_1337 0 3.8009920814148918e-03
GC_12_1338 b_12 NI_12 NS_1338 0 -2.9784186698577327e-03
GC_12_1339 b_12 NI_12 NS_1339 0 -1.8786582710673409e-03
GC_12_1340 b_12 NI_12 NS_1340 0 -3.8879556392330218e-03
GC_12_1341 b_12 NI_12 NS_1341 0 -4.0379406915098704e-04
GC_12_1342 b_12 NI_12 NS_1342 0 2.3675280190575466e-03
GC_12_1343 b_12 NI_12 NS_1343 0 -1.0556590125709999e-05
GC_12_1344 b_12 NI_12 NS_1344 0 -2.1452520938551326e-05
GC_12_1345 b_12 NI_12 NS_1345 0 8.4230055209436484e-04
GC_12_1346 b_12 NI_12 NS_1346 0 -3.7965136864219198e-03
GC_12_1347 b_12 NI_12 NS_1347 0 3.4279644062293107e-04
GC_12_1348 b_12 NI_12 NS_1348 0 3.3487743163464201e-03
GC_12_1349 b_12 NI_12 NS_1349 0 1.3577034085038484e-03
GC_12_1350 b_12 NI_12 NS_1350 0 -2.3752403677709598e-03
GC_12_1351 b_12 NI_12 NS_1351 0 2.1858930129649312e-03
GC_12_1352 b_12 NI_12 NS_1352 0 3.3360532781805713e-03
GC_12_1353 b_12 NI_12 NS_1353 0 1.1689674476248132e-03
GC_12_1354 b_12 NI_12 NS_1354 0 2.4033191298490552e-03
GC_12_1355 b_12 NI_12 NS_1355 0 -8.1092511614991227e-04
GC_12_1356 b_12 NI_12 NS_1356 0 -1.9781530790475318e-03
GC_12_1357 b_12 NI_12 NS_1357 0 3.9749601063605563e-04
GC_12_1358 b_12 NI_12 NS_1358 0 -2.6833654762314328e-03
GC_12_1359 b_12 NI_12 NS_1359 0 9.8234543226954820e-04
GC_12_1360 b_12 NI_12 NS_1360 0 2.7459675674612323e-03
GC_12_1361 b_12 NI_12 NS_1361 0 1.0390538027586018e-03
GC_12_1362 b_12 NI_12 NS_1362 0 -2.4207682785439702e-03
GC_12_1363 b_12 NI_12 NS_1363 0 -1.0837509675523838e-03
GC_12_1364 b_12 NI_12 NS_1364 0 1.5920956231316587e-03
GC_12_1365 b_12 NI_12 NS_1365 0 -1.1067035140367136e-08
GC_12_1366 b_12 NI_12 NS_1366 0 -2.8126814937226801e-09
GC_12_1367 b_12 NI_12 NS_1367 0 2.2672981072117259e-06
GC_12_1368 b_12 NI_12 NS_1368 0 5.3151740922586129e-07
GD_12_1 b_12 NI_12 NA_1 0 3.5860948117629041e-06
GD_12_2 b_12 NI_12 NA_2 0 -6.4899001493163231e-07
GD_12_3 b_12 NI_12 NA_3 0 5.6258472267656250e-06
GD_12_4 b_12 NI_12 NA_4 0 -1.8690897455120488e-06
GD_12_5 b_12 NI_12 NA_5 0 1.0213243116415748e-05
GD_12_6 b_12 NI_12 NA_6 0 -6.7055789012208793e-06
GD_12_7 b_12 NI_12 NA_7 0 2.4542728724291990e-06
GD_12_8 b_12 NI_12 NA_8 0 3.8645531297458971e-06
GD_12_9 b_12 NI_12 NA_9 0 5.9084122161429022e-04
GD_12_10 b_12 NI_12 NA_10 0 1.3006424217651833e-02
GD_12_11 b_12 NI_12 NA_11 0 -4.2260067342107148e-03
GD_12_12 b_12 NI_12 NA_12 0 -8.8592637656548946e-03
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 1.2857601077426406e+01
GS_1_1 0 NS_1 NA_1 0 4.4027142044246531e-01
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 1.7282831464635029e+02
GS_2_1 0 NS_2 NA_1 0 4.4027142044246531e-01
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 5.5743135126264733e+03
GS_3_1 0 NS_3 NA_1 0 4.4027142044246531e-01
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 1.3594126013480764e+03
GS_4_1 0 NS_4 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 1.7904812183888848e+02
RS_6 NS_6 0 1.7904812183888848e+02
GL_5 0 NS_5 NS_6 0 2.6007898045516648e-01
GL_6 0 NS_6 NS_5 0 -2.6007898045516648e-01
GS_5_1 0 NS_5 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 1.2615541320340381e+02
RS_8 NS_8 0 1.2615541320340381e+02
GL_7 0 NS_7 NS_8 0 2.5243684762014923e-01
GL_8 0 NS_8 NS_7 0 -2.5243684762014923e-01
GS_7_1 0 NS_7 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 1.0219948841586964e+02
RS_10 NS_10 0 1.0219948841586965e+02
GL_9 0 NS_9 NS_10 0 2.4690226903121384e-01
GL_10 0 NS_10 NS_9 0 -2.4690226903121384e-01
GS_9_1 0 NS_9 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 1.1002436853144543e+02
RS_12 NS_12 0 1.1002436853144542e+02
GL_11 0 NS_11 NS_12 0 2.4293768067729948e-01
GL_12 0 NS_12 NS_11 0 -2.4293768067729948e-01
GS_11_1 0 NS_11 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 1.0553430908077024e+02
RS_14 NS_14 0 1.0553430908077026e+02
GL_13 0 NS_13 NS_14 0 2.3600513224442521e-01
GL_14 0 NS_14 NS_13 0 -2.3600513224442521e-01
GS_13_1 0 NS_13 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 1.0759915098440327e+02
RS_16 NS_16 0 1.0759915098440327e+02
GL_15 0 NS_15 NS_16 0 2.3090539914362113e-01
GL_16 0 NS_16 NS_15 0 -2.3090539914362113e-01
GS_15_1 0 NS_15 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 1.3295415758774385e+02
RS_18 NS_18 0 1.3295415758774385e+02
GL_17 0 NS_17 NS_18 0 2.3030066292345727e-01
GL_18 0 NS_18 NS_17 0 -2.3030066292345727e-01
GS_17_1 0 NS_17 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 1.1432186998941940e+02
RS_20 NS_20 0 1.1432186998941938e+02
GL_19 0 NS_19 NS_20 0 2.2451058023508991e-01
GL_20 0 NS_20 NS_19 0 -2.2451058023508991e-01
GS_19_1 0 NS_19 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 9.0812703249943667e+01
RS_22 NS_22 0 9.0812703249943652e+01
GL_21 0 NS_21 NS_22 0 2.1702628900531115e-01
GL_22 0 NS_22 NS_21 0 -2.1702628900531115e-01
GS_21_1 0 NS_21 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 9.5643803662064585e+01
RS_24 NS_24 0 9.5643803662064585e+01
GL_23 0 NS_23 NS_24 0 2.1448200383207913e-01
GL_24 0 NS_24 NS_23 0 -2.1448200383207913e-01
GS_23_1 0 NS_23 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 1.0631957479149644e+02
RS_26 NS_26 0 1.0631957479149644e+02
GL_25 0 NS_25 NS_26 0 2.0655001587884311e-01
GL_26 0 NS_26 NS_25 0 -2.0655001587884311e-01
GS_25_1 0 NS_25 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 7.9907264643295406e+01
RS_28 NS_28 0 7.9907264643295420e+01
GL_27 0 NS_27 NS_28 0 2.0133773147328893e-01
GL_28 0 NS_28 NS_27 0 -2.0133773147328893e-01
GS_27_1 0 NS_27 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 1.0625506887893997e+02
RS_30 NS_30 0 1.0625506887893997e+02
GL_29 0 NS_29 NS_30 0 1.9628877333023340e-01
GL_30 0 NS_30 NS_29 0 -1.9628877333023340e-01
GS_29_1 0 NS_29 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 9.6115312638592201e+01
RS_32 NS_32 0 9.6115312638592201e+01
GL_31 0 NS_31 NS_32 0 1.8794816712418483e-01
GL_32 0 NS_32 NS_31 0 -1.8794816712418483e-01
GS_31_1 0 NS_31 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 8.5212696574118169e+01
RS_34 NS_34 0 8.5212696574118169e+01
GL_33 0 NS_33 NS_34 0 1.8572140881490298e-01
GL_34 0 NS_34 NS_33 0 -1.8572140881490298e-01
GS_33_1 0 NS_33 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 1.0905026103375434e+02
RS_36 NS_36 0 1.0905026103375432e+02
GL_35 0 NS_35 NS_36 0 1.7785621200284463e-01
GL_36 0 NS_36 NS_35 0 -1.7785621200284463e-01
GS_35_1 0 NS_35 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 8.3024437910787526e+01
RS_38 NS_38 0 8.3024437910787526e+01
GL_37 0 NS_37 NS_38 0 1.7164509875911016e-01
GL_38 0 NS_38 NS_37 0 -1.7164509875911016e-01
GS_37_1 0 NS_37 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 1.0548793856392000e+02
RS_40 NS_40 0 1.0548793856392000e+02
GL_39 0 NS_39 NS_40 0 1.6750370916002649e-01
GL_40 0 NS_40 NS_39 0 -1.6750370916002649e-01
GS_39_1 0 NS_39 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 1.0753754351502513e+02
RS_42 NS_42 0 1.0753754351502513e+02
GL_41 0 NS_41 NS_42 0 1.5942172238060490e-01
GL_42 0 NS_42 NS_41 0 -1.5942172238060490e-01
GS_41_1 0 NS_41 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 8.6961097797504721e+01
RS_44 NS_44 0 8.6961097797504721e+01
GL_43 0 NS_43 NS_44 0 1.5553892891442009e-01
GL_44 0 NS_44 NS_43 0 -1.5553892891442009e-01
GS_43_1 0 NS_43 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 1.1549771364055694e+02
RS_46 NS_46 0 1.1549771364055692e+02
GL_45 0 NS_45 NS_46 0 1.4899166019107438e-01
GL_46 0 NS_46 NS_45 0 -1.4899166019107438e-01
GS_45_1 0 NS_45 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 9.7194462506038604e+01
RS_48 NS_48 0 9.7194462506038604e+01
GL_47 0 NS_47 NS_48 0 1.4180400817347408e-01
GL_48 0 NS_48 NS_47 0 -1.4180400817347408e-01
GS_47_1 0 NS_47 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 1.0682825030924828e+02
RS_50 NS_50 0 1.0682825030924828e+02
GL_49 0 NS_49 NS_50 0 1.3872377519751058e-01
GL_50 0 NS_50 NS_49 0 -1.3872377519751058e-01
GS_49_1 0 NS_49 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 1.2559585119344567e+02
RS_52 NS_52 0 1.2559585119344568e+02
GL_51 0 NS_51 NS_52 0 1.3097721803321302e-01
GL_52 0 NS_52 NS_51 0 -1.3097721803321302e-01
GS_51_1 0 NS_51 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 1.0417660462554996e+02
RS_54 NS_54 0 1.0417660462554996e+02
GL_53 0 NS_53 NS_54 0 1.2625832867930367e-01
GL_54 0 NS_54 NS_53 0 -1.2625832867930367e-01
GS_53_1 0 NS_53 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 1.3317333532177352e+02
RS_56 NS_56 0 1.3317333532177352e+02
GL_55 0 NS_55 NS_56 0 1.2123672752714061e-01
GL_56 0 NS_56 NS_55 0 -1.2123672752714061e-01
GS_55_1 0 NS_55 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 1.2967831681616519e+02
RS_58 NS_58 0 1.2967831681616519e+02
GL_57 0 NS_57 NS_58 0 1.1651127865768855e-01
GL_58 0 NS_58 NS_57 0 -1.1651127865768855e-01
GS_57_1 0 NS_57 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 1.2999764374401394e+02
RS_60 NS_60 0 1.2999764374401394e+02
GL_59 0 NS_59 NS_60 0 1.1100247696987056e-01
GL_60 0 NS_60 NS_59 0 -1.1100247696987056e-01
GS_59_1 0 NS_59 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 1.2458814074636419e+02
RS_62 NS_62 0 1.2458814074636419e+02
GL_61 0 NS_61 NS_62 0 1.0660000212580591e-01
GL_62 0 NS_62 NS_61 0 -1.0660000212580591e-01
GS_61_1 0 NS_61 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 1.4677191614557748e+02
RS_64 NS_64 0 1.4677191614557748e+02
GL_63 0 NS_63 NS_64 0 1.0224733343325158e-01
GL_64 0 NS_64 NS_63 0 -1.0224733343325158e-01
GS_63_1 0 NS_63 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 1.3445989223131798e+02
RS_66 NS_66 0 1.3445989223131798e+02
GL_65 0 NS_65 NS_66 0 9.8177836948086503e-02
GL_66 0 NS_66 NS_65 0 -9.8177836948086503e-02
GS_65_1 0 NS_65 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 1.3187119040723775e+02
RS_68 NS_68 0 1.3187119040723772e+02
GL_67 0 NS_67 NS_68 0 9.2640196004122682e-02
GL_68 0 NS_68 NS_67 0 -9.2640196004122682e-02
GS_67_1 0 NS_67 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 1.2288401421230557e+02
RS_70 NS_70 0 1.2288401421230557e+02
GL_69 0 NS_69 NS_70 0 8.8704723748248199e-02
GL_70 0 NS_70 NS_69 0 -8.8704723748248199e-02
GS_69_1 0 NS_69 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 1.4123955654153085e+02
RS_72 NS_72 0 1.4123955654153082e+02
GL_71 0 NS_71 NS_72 0 8.4112474498892476e-02
GL_72 0 NS_72 NS_71 0 -8.4112474498892476e-02
GS_71_1 0 NS_71 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 1.2539447312269779e+02
RS_74 NS_74 0 1.2539447312269778e+02
GL_73 0 NS_73 NS_74 0 8.0007658848305588e-02
GL_74 0 NS_74 NS_73 0 -8.0007658848305588e-02
GS_73_1 0 NS_73 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 1.3219601779966965e+02
RS_76 NS_76 0 1.3219601779966968e+02
GL_75 0 NS_75 NS_76 0 7.4373183806052026e-02
GL_76 0 NS_76 NS_75 0 -7.4373183806052026e-02
GS_75_1 0 NS_75 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 1.1951371640958898e+02
RS_78 NS_78 0 1.1951371640958898e+02
GL_77 0 NS_77 NS_78 0 7.1003860961129844e-02
GL_78 0 NS_78 NS_77 0 -7.1003860961129844e-02
GS_77_1 0 NS_77 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 1.3491941875045018e+02
RS_80 NS_80 0 1.3491941875045018e+02
GL_79 0 NS_79 NS_80 0 6.5922080709048564e-02
GL_80 0 NS_80 NS_79 0 -6.5922080709048564e-02
GS_79_1 0 NS_79 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 1.2290405859347165e+02
RS_82 NS_82 0 1.2290405859347166e+02
GL_81 0 NS_81 NS_82 0 6.2340152915784278e-02
GL_82 0 NS_82 NS_81 0 -6.2340152915784278e-02
GS_81_1 0 NS_81 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 1.3258923845358959e+02
RS_84 NS_84 0 1.3258923845358959e+02
GL_83 0 NS_83 NS_84 0 5.6431081088718790e-02
GL_84 0 NS_84 NS_83 0 -5.6431081088718790e-02
GS_83_1 0 NS_83 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 1.0026704639246873e+02
RS_86 NS_86 0 1.0026704639246873e+02
GL_85 0 NS_85 NS_86 0 3.5068885856298401e-02
GL_86 0 NS_86 NS_85 0 -3.5068885856298401e-02
GS_85_1 0 NS_85 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 1.2740726499710033e+02
RS_88 NS_88 0 1.2740726499710034e+02
GL_87 0 NS_87 NS_88 0 5.3740629014256171e-02
GL_88 0 NS_88 NS_87 0 -5.3740629014256171e-02
GS_87_1 0 NS_87 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 2.3804688106534087e+02
RS_90 NS_90 0 2.3804688106534090e+02
GL_89 0 NS_89 NS_90 0 5.1425903265699464e-02
GL_90 0 NS_90 NS_89 0 -5.1425903265699464e-02
GS_89_1 0 NS_89 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 1.3728807739915800e+02
RS_92 NS_92 0 1.3728807739915803e+02
GL_91 0 NS_91 NS_92 0 4.8031392820534764e-02
GL_92 0 NS_92 NS_91 0 -4.8031392820534764e-02
GS_91_1 0 NS_91 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 1.3499477893747948e+02
RS_94 NS_94 0 1.3499477893747945e+02
GL_93 0 NS_93 NS_94 0 4.4453170742682194e-02
GL_94 0 NS_94 NS_93 0 -4.4453170742682194e-02
GS_93_1 0 NS_93 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 1.4121821834962651e+02
RS_96 NS_96 0 1.4121821834962651e+02
GL_95 0 NS_95 NS_96 0 3.8464469217755697e-02
GL_96 0 NS_96 NS_95 0 -3.8464469217755697e-02
GS_95_1 0 NS_95 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 1.3946471282741149e+02
RS_98 NS_98 0 1.3946471282741149e+02
GL_97 0 NS_97 NS_98 0 3.5678935079258622e-02
GL_98 0 NS_98 NS_97 0 -3.5678935079258622e-02
GS_97_1 0 NS_97 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 1.5530211191942624e+02
RS_100 NS_100 0 1.5530211191942627e+02
GL_99 0 NS_99 NS_100 0 2.6209890345437525e-02
GL_100 0 NS_100 NS_99 0 -2.6209890345437525e-02
GS_99_1 0 NS_99 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 1.4887428879582419e+02
RS_102 NS_102 0 1.4887428879582419e+02
GL_101 0 NS_101 NS_102 0 3.0330575323949095e-02
GL_102 0 NS_102 NS_101 0 -3.0330575323949095e-02
GS_101_1 0 NS_101 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 1.5087532095170570e+02
RS_104 NS_104 0 1.5087532095170570e+02
GL_103 0 NS_103 NS_104 0 2.0034138441714564e-02
GL_104 0 NS_104 NS_103 0 -2.0034138441714564e-02
GS_103_1 0 NS_103 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 1.4763793449752018e+02
RS_106 NS_106 0 1.4763793449752018e+02
GL_105 0 NS_105 NS_106 0 1.7017170579416537e-02
GL_106 0 NS_106 NS_105 0 -1.7017170579416537e-02
GS_105_1 0 NS_105 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 1.6285515224442304e+02
RS_108 NS_108 0 1.6285515224442304e+02
GL_107 0 NS_107 NS_108 0 1.0897027002452746e-02
GL_108 0 NS_108 NS_107 0 -1.0897027002452746e-02
GS_107_1 0 NS_107 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 1.7239534388116820e+02
RS_110 NS_110 0 1.7239534388116820e+02
GL_109 0 NS_109 NS_110 0 6.1589693699488982e-03
GL_110 0 NS_110 NS_109 0 -6.1589693699488982e-03
GS_109_1 0 NS_109 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 5.9928710578594173e+03
RS_112 NS_112 0 5.9928710578594173e+03
GL_111 0 NS_111 NS_112 0 1.7541178006601681e-03
GL_112 0 NS_112 NS_111 0 -1.7541178006601681e-03
GS_111_1 0 NS_111 NA_1 0 4.4027142044246531e-01
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 8.0762087901330699e+02
RS_114 NS_114 0 8.0762087901330688e+02
GL_113 0 NS_113 NS_114 0 1.7295489372816217e-03
GL_114 0 NS_114 NS_113 0 -1.7295489372816217e-03
GS_113_1 0 NS_113 NA_1 0 4.4027142044246531e-01
*
* Real pole n. 115
CS_115 NS_115 0 9.9999999999999998e-13
RS_115 NS_115 0 1.2857601077426406e+01
GS_115_2 0 NS_115 NA_2 0 4.4027142044246531e-01
*
* Real pole n. 116
CS_116 NS_116 0 9.9999999999999998e-13
RS_116 NS_116 0 1.7282831464635029e+02
GS_116_2 0 NS_116 NA_2 0 4.4027142044246531e-01
*
* Real pole n. 117
CS_117 NS_117 0 9.9999999999999998e-13
RS_117 NS_117 0 5.5743135126264733e+03
GS_117_2 0 NS_117 NA_2 0 4.4027142044246531e-01
*
* Real pole n. 118
CS_118 NS_118 0 9.9999999999999998e-13
RS_118 NS_118 0 1.3594126013480764e+03
GS_118_2 0 NS_118 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 1.7904812183888848e+02
RS_120 NS_120 0 1.7904812183888848e+02
GL_119 0 NS_119 NS_120 0 2.6007898045516648e-01
GL_120 0 NS_120 NS_119 0 -2.6007898045516648e-01
GS_119_2 0 NS_119 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 1.2615541320340381e+02
RS_122 NS_122 0 1.2615541320340381e+02
GL_121 0 NS_121 NS_122 0 2.5243684762014923e-01
GL_122 0 NS_122 NS_121 0 -2.5243684762014923e-01
GS_121_2 0 NS_121 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 1.0219948841586964e+02
RS_124 NS_124 0 1.0219948841586965e+02
GL_123 0 NS_123 NS_124 0 2.4690226903121384e-01
GL_124 0 NS_124 NS_123 0 -2.4690226903121384e-01
GS_123_2 0 NS_123 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 1.1002436853144543e+02
RS_126 NS_126 0 1.1002436853144542e+02
GL_125 0 NS_125 NS_126 0 2.4293768067729948e-01
GL_126 0 NS_126 NS_125 0 -2.4293768067729948e-01
GS_125_2 0 NS_125 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 1.0553430908077024e+02
RS_128 NS_128 0 1.0553430908077026e+02
GL_127 0 NS_127 NS_128 0 2.3600513224442521e-01
GL_128 0 NS_128 NS_127 0 -2.3600513224442521e-01
GS_127_2 0 NS_127 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 1.0759915098440327e+02
RS_130 NS_130 0 1.0759915098440327e+02
GL_129 0 NS_129 NS_130 0 2.3090539914362113e-01
GL_130 0 NS_130 NS_129 0 -2.3090539914362113e-01
GS_129_2 0 NS_129 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 1.3295415758774385e+02
RS_132 NS_132 0 1.3295415758774385e+02
GL_131 0 NS_131 NS_132 0 2.3030066292345727e-01
GL_132 0 NS_132 NS_131 0 -2.3030066292345727e-01
GS_131_2 0 NS_131 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 133/134
CS_133 NS_133 0 9.9999999999999998e-13
CS_134 NS_134 0 9.9999999999999998e-13
RS_133 NS_133 0 1.1432186998941940e+02
RS_134 NS_134 0 1.1432186998941938e+02
GL_133 0 NS_133 NS_134 0 2.2451058023508991e-01
GL_134 0 NS_134 NS_133 0 -2.2451058023508991e-01
GS_133_2 0 NS_133 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 9.0812703249943667e+01
RS_136 NS_136 0 9.0812703249943652e+01
GL_135 0 NS_135 NS_136 0 2.1702628900531115e-01
GL_136 0 NS_136 NS_135 0 -2.1702628900531115e-01
GS_135_2 0 NS_135 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 9.5643803662064585e+01
RS_138 NS_138 0 9.5643803662064585e+01
GL_137 0 NS_137 NS_138 0 2.1448200383207913e-01
GL_138 0 NS_138 NS_137 0 -2.1448200383207913e-01
GS_137_2 0 NS_137 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 1.0631957479149644e+02
RS_140 NS_140 0 1.0631957479149644e+02
GL_139 0 NS_139 NS_140 0 2.0655001587884311e-01
GL_140 0 NS_140 NS_139 0 -2.0655001587884311e-01
GS_139_2 0 NS_139 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 7.9907264643295406e+01
RS_142 NS_142 0 7.9907264643295420e+01
GL_141 0 NS_141 NS_142 0 2.0133773147328893e-01
GL_142 0 NS_142 NS_141 0 -2.0133773147328893e-01
GS_141_2 0 NS_141 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 1.0625506887893997e+02
RS_144 NS_144 0 1.0625506887893997e+02
GL_143 0 NS_143 NS_144 0 1.9628877333023340e-01
GL_144 0 NS_144 NS_143 0 -1.9628877333023340e-01
GS_143_2 0 NS_143 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 9.6115312638592201e+01
RS_146 NS_146 0 9.6115312638592201e+01
GL_145 0 NS_145 NS_146 0 1.8794816712418483e-01
GL_146 0 NS_146 NS_145 0 -1.8794816712418483e-01
GS_145_2 0 NS_145 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 8.5212696574118169e+01
RS_148 NS_148 0 8.5212696574118169e+01
GL_147 0 NS_147 NS_148 0 1.8572140881490298e-01
GL_148 0 NS_148 NS_147 0 -1.8572140881490298e-01
GS_147_2 0 NS_147 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 1.0905026103375434e+02
RS_150 NS_150 0 1.0905026103375432e+02
GL_149 0 NS_149 NS_150 0 1.7785621200284463e-01
GL_150 0 NS_150 NS_149 0 -1.7785621200284463e-01
GS_149_2 0 NS_149 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 8.3024437910787526e+01
RS_152 NS_152 0 8.3024437910787526e+01
GL_151 0 NS_151 NS_152 0 1.7164509875911016e-01
GL_152 0 NS_152 NS_151 0 -1.7164509875911016e-01
GS_151_2 0 NS_151 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 1.0548793856392000e+02
RS_154 NS_154 0 1.0548793856392000e+02
GL_153 0 NS_153 NS_154 0 1.6750370916002649e-01
GL_154 0 NS_154 NS_153 0 -1.6750370916002649e-01
GS_153_2 0 NS_153 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 1.0753754351502513e+02
RS_156 NS_156 0 1.0753754351502513e+02
GL_155 0 NS_155 NS_156 0 1.5942172238060490e-01
GL_156 0 NS_156 NS_155 0 -1.5942172238060490e-01
GS_155_2 0 NS_155 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 8.6961097797504721e+01
RS_158 NS_158 0 8.6961097797504721e+01
GL_157 0 NS_157 NS_158 0 1.5553892891442009e-01
GL_158 0 NS_158 NS_157 0 -1.5553892891442009e-01
GS_157_2 0 NS_157 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 1.1549771364055694e+02
RS_160 NS_160 0 1.1549771364055692e+02
GL_159 0 NS_159 NS_160 0 1.4899166019107438e-01
GL_160 0 NS_160 NS_159 0 -1.4899166019107438e-01
GS_159_2 0 NS_159 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 9.7194462506038604e+01
RS_162 NS_162 0 9.7194462506038604e+01
GL_161 0 NS_161 NS_162 0 1.4180400817347408e-01
GL_162 0 NS_162 NS_161 0 -1.4180400817347408e-01
GS_161_2 0 NS_161 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 163/164
CS_163 NS_163 0 9.9999999999999998e-13
CS_164 NS_164 0 9.9999999999999998e-13
RS_163 NS_163 0 1.0682825030924828e+02
RS_164 NS_164 0 1.0682825030924828e+02
GL_163 0 NS_163 NS_164 0 1.3872377519751058e-01
GL_164 0 NS_164 NS_163 0 -1.3872377519751058e-01
GS_163_2 0 NS_163 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 1.2559585119344567e+02
RS_166 NS_166 0 1.2559585119344568e+02
GL_165 0 NS_165 NS_166 0 1.3097721803321302e-01
GL_166 0 NS_166 NS_165 0 -1.3097721803321302e-01
GS_165_2 0 NS_165 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 1.0417660462554996e+02
RS_168 NS_168 0 1.0417660462554996e+02
GL_167 0 NS_167 NS_168 0 1.2625832867930367e-01
GL_168 0 NS_168 NS_167 0 -1.2625832867930367e-01
GS_167_2 0 NS_167 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 1.3317333532177352e+02
RS_170 NS_170 0 1.3317333532177352e+02
GL_169 0 NS_169 NS_170 0 1.2123672752714061e-01
GL_170 0 NS_170 NS_169 0 -1.2123672752714061e-01
GS_169_2 0 NS_169 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 1.2967831681616519e+02
RS_172 NS_172 0 1.2967831681616519e+02
GL_171 0 NS_171 NS_172 0 1.1651127865768855e-01
GL_172 0 NS_172 NS_171 0 -1.1651127865768855e-01
GS_171_2 0 NS_171 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 1.2999764374401394e+02
RS_174 NS_174 0 1.2999764374401394e+02
GL_173 0 NS_173 NS_174 0 1.1100247696987056e-01
GL_174 0 NS_174 NS_173 0 -1.1100247696987056e-01
GS_173_2 0 NS_173 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 1.2458814074636419e+02
RS_176 NS_176 0 1.2458814074636419e+02
GL_175 0 NS_175 NS_176 0 1.0660000212580591e-01
GL_176 0 NS_176 NS_175 0 -1.0660000212580591e-01
GS_175_2 0 NS_175 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 1.4677191614557748e+02
RS_178 NS_178 0 1.4677191614557748e+02
GL_177 0 NS_177 NS_178 0 1.0224733343325158e-01
GL_178 0 NS_178 NS_177 0 -1.0224733343325158e-01
GS_177_2 0 NS_177 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 1.3445989223131798e+02
RS_180 NS_180 0 1.3445989223131798e+02
GL_179 0 NS_179 NS_180 0 9.8177836948086503e-02
GL_180 0 NS_180 NS_179 0 -9.8177836948086503e-02
GS_179_2 0 NS_179 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 181/182
CS_181 NS_181 0 9.9999999999999998e-13
CS_182 NS_182 0 9.9999999999999998e-13
RS_181 NS_181 0 1.3187119040723775e+02
RS_182 NS_182 0 1.3187119040723772e+02
GL_181 0 NS_181 NS_182 0 9.2640196004122682e-02
GL_182 0 NS_182 NS_181 0 -9.2640196004122682e-02
GS_181_2 0 NS_181 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 183/184
CS_183 NS_183 0 9.9999999999999998e-13
CS_184 NS_184 0 9.9999999999999998e-13
RS_183 NS_183 0 1.2288401421230557e+02
RS_184 NS_184 0 1.2288401421230557e+02
GL_183 0 NS_183 NS_184 0 8.8704723748248199e-02
GL_184 0 NS_184 NS_183 0 -8.8704723748248199e-02
GS_183_2 0 NS_183 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 1.4123955654153085e+02
RS_186 NS_186 0 1.4123955654153082e+02
GL_185 0 NS_185 NS_186 0 8.4112474498892476e-02
GL_186 0 NS_186 NS_185 0 -8.4112474498892476e-02
GS_185_2 0 NS_185 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 1.2539447312269779e+02
RS_188 NS_188 0 1.2539447312269778e+02
GL_187 0 NS_187 NS_188 0 8.0007658848305588e-02
GL_188 0 NS_188 NS_187 0 -8.0007658848305588e-02
GS_187_2 0 NS_187 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 1.3219601779966965e+02
RS_190 NS_190 0 1.3219601779966968e+02
GL_189 0 NS_189 NS_190 0 7.4373183806052026e-02
GL_190 0 NS_190 NS_189 0 -7.4373183806052026e-02
GS_189_2 0 NS_189 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 1.1951371640958898e+02
RS_192 NS_192 0 1.1951371640958898e+02
GL_191 0 NS_191 NS_192 0 7.1003860961129844e-02
GL_192 0 NS_192 NS_191 0 -7.1003860961129844e-02
GS_191_2 0 NS_191 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 1.3491941875045018e+02
RS_194 NS_194 0 1.3491941875045018e+02
GL_193 0 NS_193 NS_194 0 6.5922080709048564e-02
GL_194 0 NS_194 NS_193 0 -6.5922080709048564e-02
GS_193_2 0 NS_193 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 1.2290405859347165e+02
RS_196 NS_196 0 1.2290405859347166e+02
GL_195 0 NS_195 NS_196 0 6.2340152915784278e-02
GL_196 0 NS_196 NS_195 0 -6.2340152915784278e-02
GS_195_2 0 NS_195 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 1.3258923845358959e+02
RS_198 NS_198 0 1.3258923845358959e+02
GL_197 0 NS_197 NS_198 0 5.6431081088718790e-02
GL_198 0 NS_198 NS_197 0 -5.6431081088718790e-02
GS_197_2 0 NS_197 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 1.0026704639246873e+02
RS_200 NS_200 0 1.0026704639246873e+02
GL_199 0 NS_199 NS_200 0 3.5068885856298401e-02
GL_200 0 NS_200 NS_199 0 -3.5068885856298401e-02
GS_199_2 0 NS_199 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 201/202
CS_201 NS_201 0 9.9999999999999998e-13
CS_202 NS_202 0 9.9999999999999998e-13
RS_201 NS_201 0 1.2740726499710033e+02
RS_202 NS_202 0 1.2740726499710034e+02
GL_201 0 NS_201 NS_202 0 5.3740629014256171e-02
GL_202 0 NS_202 NS_201 0 -5.3740629014256171e-02
GS_201_2 0 NS_201 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 203/204
CS_203 NS_203 0 9.9999999999999998e-13
CS_204 NS_204 0 9.9999999999999998e-13
RS_203 NS_203 0 2.3804688106534087e+02
RS_204 NS_204 0 2.3804688106534090e+02
GL_203 0 NS_203 NS_204 0 5.1425903265699464e-02
GL_204 0 NS_204 NS_203 0 -5.1425903265699464e-02
GS_203_2 0 NS_203 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 1.3728807739915800e+02
RS_206 NS_206 0 1.3728807739915803e+02
GL_205 0 NS_205 NS_206 0 4.8031392820534764e-02
GL_206 0 NS_206 NS_205 0 -4.8031392820534764e-02
GS_205_2 0 NS_205 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 1.3499477893747948e+02
RS_208 NS_208 0 1.3499477893747945e+02
GL_207 0 NS_207 NS_208 0 4.4453170742682194e-02
GL_208 0 NS_208 NS_207 0 -4.4453170742682194e-02
GS_207_2 0 NS_207 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 1.4121821834962651e+02
RS_210 NS_210 0 1.4121821834962651e+02
GL_209 0 NS_209 NS_210 0 3.8464469217755697e-02
GL_210 0 NS_210 NS_209 0 -3.8464469217755697e-02
GS_209_2 0 NS_209 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 1.3946471282741149e+02
RS_212 NS_212 0 1.3946471282741149e+02
GL_211 0 NS_211 NS_212 0 3.5678935079258622e-02
GL_212 0 NS_212 NS_211 0 -3.5678935079258622e-02
GS_211_2 0 NS_211 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 1.5530211191942624e+02
RS_214 NS_214 0 1.5530211191942627e+02
GL_213 0 NS_213 NS_214 0 2.6209890345437525e-02
GL_214 0 NS_214 NS_213 0 -2.6209890345437525e-02
GS_213_2 0 NS_213 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 1.4887428879582419e+02
RS_216 NS_216 0 1.4887428879582419e+02
GL_215 0 NS_215 NS_216 0 3.0330575323949095e-02
GL_216 0 NS_216 NS_215 0 -3.0330575323949095e-02
GS_215_2 0 NS_215 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 1.5087532095170570e+02
RS_218 NS_218 0 1.5087532095170570e+02
GL_217 0 NS_217 NS_218 0 2.0034138441714564e-02
GL_218 0 NS_218 NS_217 0 -2.0034138441714564e-02
GS_217_2 0 NS_217 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 1.4763793449752018e+02
RS_220 NS_220 0 1.4763793449752018e+02
GL_219 0 NS_219 NS_220 0 1.7017170579416537e-02
GL_220 0 NS_220 NS_219 0 -1.7017170579416537e-02
GS_219_2 0 NS_219 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 221/222
CS_221 NS_221 0 9.9999999999999998e-13
CS_222 NS_222 0 9.9999999999999998e-13
RS_221 NS_221 0 1.6285515224442304e+02
RS_222 NS_222 0 1.6285515224442304e+02
GL_221 0 NS_221 NS_222 0 1.0897027002452746e-02
GL_222 0 NS_222 NS_221 0 -1.0897027002452746e-02
GS_221_2 0 NS_221 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 223/224
CS_223 NS_223 0 9.9999999999999998e-13
CS_224 NS_224 0 9.9999999999999998e-13
RS_223 NS_223 0 1.7239534388116820e+02
RS_224 NS_224 0 1.7239534388116820e+02
GL_223 0 NS_223 NS_224 0 6.1589693699488982e-03
GL_224 0 NS_224 NS_223 0 -6.1589693699488982e-03
GS_223_2 0 NS_223 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 225/226
CS_225 NS_225 0 9.9999999999999998e-13
CS_226 NS_226 0 9.9999999999999998e-13
RS_225 NS_225 0 5.9928710578594173e+03
RS_226 NS_226 0 5.9928710578594173e+03
GL_225 0 NS_225 NS_226 0 1.7541178006601681e-03
GL_226 0 NS_226 NS_225 0 -1.7541178006601681e-03
GS_225_2 0 NS_225 NA_2 0 4.4027142044246531e-01
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 8.0762087901330699e+02
RS_228 NS_228 0 8.0762087901330688e+02
GL_227 0 NS_227 NS_228 0 1.7295489372816217e-03
GL_228 0 NS_228 NS_227 0 -1.7295489372816217e-03
GS_227_2 0 NS_227 NA_2 0 4.4027142044246531e-01
*
* Real pole n. 229
CS_229 NS_229 0 9.9999999999999998e-13
RS_229 NS_229 0 1.2857601077426406e+01
GS_229_3 0 NS_229 NA_3 0 4.4027142044246531e-01
*
* Real pole n. 230
CS_230 NS_230 0 9.9999999999999998e-13
RS_230 NS_230 0 1.7282831464635029e+02
GS_230_3 0 NS_230 NA_3 0 4.4027142044246531e-01
*
* Real pole n. 231
CS_231 NS_231 0 9.9999999999999998e-13
RS_231 NS_231 0 5.5743135126264733e+03
GS_231_3 0 NS_231 NA_3 0 4.4027142044246531e-01
*
* Real pole n. 232
CS_232 NS_232 0 9.9999999999999998e-13
RS_232 NS_232 0 1.3594126013480764e+03
GS_232_3 0 NS_232 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 1.7904812183888848e+02
RS_234 NS_234 0 1.7904812183888848e+02
GL_233 0 NS_233 NS_234 0 2.6007898045516648e-01
GL_234 0 NS_234 NS_233 0 -2.6007898045516648e-01
GS_233_3 0 NS_233 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 1.2615541320340381e+02
RS_236 NS_236 0 1.2615541320340381e+02
GL_235 0 NS_235 NS_236 0 2.5243684762014923e-01
GL_236 0 NS_236 NS_235 0 -2.5243684762014923e-01
GS_235_3 0 NS_235 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 1.0219948841586964e+02
RS_238 NS_238 0 1.0219948841586965e+02
GL_237 0 NS_237 NS_238 0 2.4690226903121384e-01
GL_238 0 NS_238 NS_237 0 -2.4690226903121384e-01
GS_237_3 0 NS_237 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 1.1002436853144543e+02
RS_240 NS_240 0 1.1002436853144542e+02
GL_239 0 NS_239 NS_240 0 2.4293768067729948e-01
GL_240 0 NS_240 NS_239 0 -2.4293768067729948e-01
GS_239_3 0 NS_239 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 241/242
CS_241 NS_241 0 9.9999999999999998e-13
CS_242 NS_242 0 9.9999999999999998e-13
RS_241 NS_241 0 1.0553430908077024e+02
RS_242 NS_242 0 1.0553430908077026e+02
GL_241 0 NS_241 NS_242 0 2.3600513224442521e-01
GL_242 0 NS_242 NS_241 0 -2.3600513224442521e-01
GS_241_3 0 NS_241 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 243/244
CS_243 NS_243 0 9.9999999999999998e-13
CS_244 NS_244 0 9.9999999999999998e-13
RS_243 NS_243 0 1.0759915098440327e+02
RS_244 NS_244 0 1.0759915098440327e+02
GL_243 0 NS_243 NS_244 0 2.3090539914362113e-01
GL_244 0 NS_244 NS_243 0 -2.3090539914362113e-01
GS_243_3 0 NS_243 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 245/246
CS_245 NS_245 0 9.9999999999999998e-13
CS_246 NS_246 0 9.9999999999999998e-13
RS_245 NS_245 0 1.3295415758774385e+02
RS_246 NS_246 0 1.3295415758774385e+02
GL_245 0 NS_245 NS_246 0 2.3030066292345727e-01
GL_246 0 NS_246 NS_245 0 -2.3030066292345727e-01
GS_245_3 0 NS_245 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 247/248
CS_247 NS_247 0 9.9999999999999998e-13
CS_248 NS_248 0 9.9999999999999998e-13
RS_247 NS_247 0 1.1432186998941940e+02
RS_248 NS_248 0 1.1432186998941938e+02
GL_247 0 NS_247 NS_248 0 2.2451058023508991e-01
GL_248 0 NS_248 NS_247 0 -2.2451058023508991e-01
GS_247_3 0 NS_247 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 249/250
CS_249 NS_249 0 9.9999999999999998e-13
CS_250 NS_250 0 9.9999999999999998e-13
RS_249 NS_249 0 9.0812703249943667e+01
RS_250 NS_250 0 9.0812703249943652e+01
GL_249 0 NS_249 NS_250 0 2.1702628900531115e-01
GL_250 0 NS_250 NS_249 0 -2.1702628900531115e-01
GS_249_3 0 NS_249 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 251/252
CS_251 NS_251 0 9.9999999999999998e-13
CS_252 NS_252 0 9.9999999999999998e-13
RS_251 NS_251 0 9.5643803662064585e+01
RS_252 NS_252 0 9.5643803662064585e+01
GL_251 0 NS_251 NS_252 0 2.1448200383207913e-01
GL_252 0 NS_252 NS_251 0 -2.1448200383207913e-01
GS_251_3 0 NS_251 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 253/254
CS_253 NS_253 0 9.9999999999999998e-13
CS_254 NS_254 0 9.9999999999999998e-13
RS_253 NS_253 0 1.0631957479149644e+02
RS_254 NS_254 0 1.0631957479149644e+02
GL_253 0 NS_253 NS_254 0 2.0655001587884311e-01
GL_254 0 NS_254 NS_253 0 -2.0655001587884311e-01
GS_253_3 0 NS_253 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 255/256
CS_255 NS_255 0 9.9999999999999998e-13
CS_256 NS_256 0 9.9999999999999998e-13
RS_255 NS_255 0 7.9907264643295406e+01
RS_256 NS_256 0 7.9907264643295420e+01
GL_255 0 NS_255 NS_256 0 2.0133773147328893e-01
GL_256 0 NS_256 NS_255 0 -2.0133773147328893e-01
GS_255_3 0 NS_255 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 257/258
CS_257 NS_257 0 9.9999999999999998e-13
CS_258 NS_258 0 9.9999999999999998e-13
RS_257 NS_257 0 1.0625506887893997e+02
RS_258 NS_258 0 1.0625506887893997e+02
GL_257 0 NS_257 NS_258 0 1.9628877333023340e-01
GL_258 0 NS_258 NS_257 0 -1.9628877333023340e-01
GS_257_3 0 NS_257 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 259/260
CS_259 NS_259 0 9.9999999999999998e-13
CS_260 NS_260 0 9.9999999999999998e-13
RS_259 NS_259 0 9.6115312638592201e+01
RS_260 NS_260 0 9.6115312638592201e+01
GL_259 0 NS_259 NS_260 0 1.8794816712418483e-01
GL_260 0 NS_260 NS_259 0 -1.8794816712418483e-01
GS_259_3 0 NS_259 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 261/262
CS_261 NS_261 0 9.9999999999999998e-13
CS_262 NS_262 0 9.9999999999999998e-13
RS_261 NS_261 0 8.5212696574118169e+01
RS_262 NS_262 0 8.5212696574118169e+01
GL_261 0 NS_261 NS_262 0 1.8572140881490298e-01
GL_262 0 NS_262 NS_261 0 -1.8572140881490298e-01
GS_261_3 0 NS_261 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 263/264
CS_263 NS_263 0 9.9999999999999998e-13
CS_264 NS_264 0 9.9999999999999998e-13
RS_263 NS_263 0 1.0905026103375434e+02
RS_264 NS_264 0 1.0905026103375432e+02
GL_263 0 NS_263 NS_264 0 1.7785621200284463e-01
GL_264 0 NS_264 NS_263 0 -1.7785621200284463e-01
GS_263_3 0 NS_263 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 265/266
CS_265 NS_265 0 9.9999999999999998e-13
CS_266 NS_266 0 9.9999999999999998e-13
RS_265 NS_265 0 8.3024437910787526e+01
RS_266 NS_266 0 8.3024437910787526e+01
GL_265 0 NS_265 NS_266 0 1.7164509875911016e-01
GL_266 0 NS_266 NS_265 0 -1.7164509875911016e-01
GS_265_3 0 NS_265 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 267/268
CS_267 NS_267 0 9.9999999999999998e-13
CS_268 NS_268 0 9.9999999999999998e-13
RS_267 NS_267 0 1.0548793856392000e+02
RS_268 NS_268 0 1.0548793856392000e+02
GL_267 0 NS_267 NS_268 0 1.6750370916002649e-01
GL_268 0 NS_268 NS_267 0 -1.6750370916002649e-01
GS_267_3 0 NS_267 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 269/270
CS_269 NS_269 0 9.9999999999999998e-13
CS_270 NS_270 0 9.9999999999999998e-13
RS_269 NS_269 0 1.0753754351502513e+02
RS_270 NS_270 0 1.0753754351502513e+02
GL_269 0 NS_269 NS_270 0 1.5942172238060490e-01
GL_270 0 NS_270 NS_269 0 -1.5942172238060490e-01
GS_269_3 0 NS_269 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 271/272
CS_271 NS_271 0 9.9999999999999998e-13
CS_272 NS_272 0 9.9999999999999998e-13
RS_271 NS_271 0 8.6961097797504721e+01
RS_272 NS_272 0 8.6961097797504721e+01
GL_271 0 NS_271 NS_272 0 1.5553892891442009e-01
GL_272 0 NS_272 NS_271 0 -1.5553892891442009e-01
GS_271_3 0 NS_271 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 273/274
CS_273 NS_273 0 9.9999999999999998e-13
CS_274 NS_274 0 9.9999999999999998e-13
RS_273 NS_273 0 1.1549771364055694e+02
RS_274 NS_274 0 1.1549771364055692e+02
GL_273 0 NS_273 NS_274 0 1.4899166019107438e-01
GL_274 0 NS_274 NS_273 0 -1.4899166019107438e-01
GS_273_3 0 NS_273 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 275/276
CS_275 NS_275 0 9.9999999999999998e-13
CS_276 NS_276 0 9.9999999999999998e-13
RS_275 NS_275 0 9.7194462506038604e+01
RS_276 NS_276 0 9.7194462506038604e+01
GL_275 0 NS_275 NS_276 0 1.4180400817347408e-01
GL_276 0 NS_276 NS_275 0 -1.4180400817347408e-01
GS_275_3 0 NS_275 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 277/278
CS_277 NS_277 0 9.9999999999999998e-13
CS_278 NS_278 0 9.9999999999999998e-13
RS_277 NS_277 0 1.0682825030924828e+02
RS_278 NS_278 0 1.0682825030924828e+02
GL_277 0 NS_277 NS_278 0 1.3872377519751058e-01
GL_278 0 NS_278 NS_277 0 -1.3872377519751058e-01
GS_277_3 0 NS_277 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 279/280
CS_279 NS_279 0 9.9999999999999998e-13
CS_280 NS_280 0 9.9999999999999998e-13
RS_279 NS_279 0 1.2559585119344567e+02
RS_280 NS_280 0 1.2559585119344568e+02
GL_279 0 NS_279 NS_280 0 1.3097721803321302e-01
GL_280 0 NS_280 NS_279 0 -1.3097721803321302e-01
GS_279_3 0 NS_279 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 281/282
CS_281 NS_281 0 9.9999999999999998e-13
CS_282 NS_282 0 9.9999999999999998e-13
RS_281 NS_281 0 1.0417660462554996e+02
RS_282 NS_282 0 1.0417660462554996e+02
GL_281 0 NS_281 NS_282 0 1.2625832867930367e-01
GL_282 0 NS_282 NS_281 0 -1.2625832867930367e-01
GS_281_3 0 NS_281 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 283/284
CS_283 NS_283 0 9.9999999999999998e-13
CS_284 NS_284 0 9.9999999999999998e-13
RS_283 NS_283 0 1.3317333532177352e+02
RS_284 NS_284 0 1.3317333532177352e+02
GL_283 0 NS_283 NS_284 0 1.2123672752714061e-01
GL_284 0 NS_284 NS_283 0 -1.2123672752714061e-01
GS_283_3 0 NS_283 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 285/286
CS_285 NS_285 0 9.9999999999999998e-13
CS_286 NS_286 0 9.9999999999999998e-13
RS_285 NS_285 0 1.2967831681616519e+02
RS_286 NS_286 0 1.2967831681616519e+02
GL_285 0 NS_285 NS_286 0 1.1651127865768855e-01
GL_286 0 NS_286 NS_285 0 -1.1651127865768855e-01
GS_285_3 0 NS_285 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 287/288
CS_287 NS_287 0 9.9999999999999998e-13
CS_288 NS_288 0 9.9999999999999998e-13
RS_287 NS_287 0 1.2999764374401394e+02
RS_288 NS_288 0 1.2999764374401394e+02
GL_287 0 NS_287 NS_288 0 1.1100247696987056e-01
GL_288 0 NS_288 NS_287 0 -1.1100247696987056e-01
GS_287_3 0 NS_287 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 289/290
CS_289 NS_289 0 9.9999999999999998e-13
CS_290 NS_290 0 9.9999999999999998e-13
RS_289 NS_289 0 1.2458814074636419e+02
RS_290 NS_290 0 1.2458814074636419e+02
GL_289 0 NS_289 NS_290 0 1.0660000212580591e-01
GL_290 0 NS_290 NS_289 0 -1.0660000212580591e-01
GS_289_3 0 NS_289 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 291/292
CS_291 NS_291 0 9.9999999999999998e-13
CS_292 NS_292 0 9.9999999999999998e-13
RS_291 NS_291 0 1.4677191614557748e+02
RS_292 NS_292 0 1.4677191614557748e+02
GL_291 0 NS_291 NS_292 0 1.0224733343325158e-01
GL_292 0 NS_292 NS_291 0 -1.0224733343325158e-01
GS_291_3 0 NS_291 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 293/294
CS_293 NS_293 0 9.9999999999999998e-13
CS_294 NS_294 0 9.9999999999999998e-13
RS_293 NS_293 0 1.3445989223131798e+02
RS_294 NS_294 0 1.3445989223131798e+02
GL_293 0 NS_293 NS_294 0 9.8177836948086503e-02
GL_294 0 NS_294 NS_293 0 -9.8177836948086503e-02
GS_293_3 0 NS_293 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 295/296
CS_295 NS_295 0 9.9999999999999998e-13
CS_296 NS_296 0 9.9999999999999998e-13
RS_295 NS_295 0 1.3187119040723775e+02
RS_296 NS_296 0 1.3187119040723772e+02
GL_295 0 NS_295 NS_296 0 9.2640196004122682e-02
GL_296 0 NS_296 NS_295 0 -9.2640196004122682e-02
GS_295_3 0 NS_295 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 297/298
CS_297 NS_297 0 9.9999999999999998e-13
CS_298 NS_298 0 9.9999999999999998e-13
RS_297 NS_297 0 1.2288401421230557e+02
RS_298 NS_298 0 1.2288401421230557e+02
GL_297 0 NS_297 NS_298 0 8.8704723748248199e-02
GL_298 0 NS_298 NS_297 0 -8.8704723748248199e-02
GS_297_3 0 NS_297 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 299/300
CS_299 NS_299 0 9.9999999999999998e-13
CS_300 NS_300 0 9.9999999999999998e-13
RS_299 NS_299 0 1.4123955654153085e+02
RS_300 NS_300 0 1.4123955654153082e+02
GL_299 0 NS_299 NS_300 0 8.4112474498892476e-02
GL_300 0 NS_300 NS_299 0 -8.4112474498892476e-02
GS_299_3 0 NS_299 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 301/302
CS_301 NS_301 0 9.9999999999999998e-13
CS_302 NS_302 0 9.9999999999999998e-13
RS_301 NS_301 0 1.2539447312269779e+02
RS_302 NS_302 0 1.2539447312269778e+02
GL_301 0 NS_301 NS_302 0 8.0007658848305588e-02
GL_302 0 NS_302 NS_301 0 -8.0007658848305588e-02
GS_301_3 0 NS_301 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 303/304
CS_303 NS_303 0 9.9999999999999998e-13
CS_304 NS_304 0 9.9999999999999998e-13
RS_303 NS_303 0 1.3219601779966965e+02
RS_304 NS_304 0 1.3219601779966968e+02
GL_303 0 NS_303 NS_304 0 7.4373183806052026e-02
GL_304 0 NS_304 NS_303 0 -7.4373183806052026e-02
GS_303_3 0 NS_303 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 305/306
CS_305 NS_305 0 9.9999999999999998e-13
CS_306 NS_306 0 9.9999999999999998e-13
RS_305 NS_305 0 1.1951371640958898e+02
RS_306 NS_306 0 1.1951371640958898e+02
GL_305 0 NS_305 NS_306 0 7.1003860961129844e-02
GL_306 0 NS_306 NS_305 0 -7.1003860961129844e-02
GS_305_3 0 NS_305 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 307/308
CS_307 NS_307 0 9.9999999999999998e-13
CS_308 NS_308 0 9.9999999999999998e-13
RS_307 NS_307 0 1.3491941875045018e+02
RS_308 NS_308 0 1.3491941875045018e+02
GL_307 0 NS_307 NS_308 0 6.5922080709048564e-02
GL_308 0 NS_308 NS_307 0 -6.5922080709048564e-02
GS_307_3 0 NS_307 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 309/310
CS_309 NS_309 0 9.9999999999999998e-13
CS_310 NS_310 0 9.9999999999999998e-13
RS_309 NS_309 0 1.2290405859347165e+02
RS_310 NS_310 0 1.2290405859347166e+02
GL_309 0 NS_309 NS_310 0 6.2340152915784278e-02
GL_310 0 NS_310 NS_309 0 -6.2340152915784278e-02
GS_309_3 0 NS_309 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 311/312
CS_311 NS_311 0 9.9999999999999998e-13
CS_312 NS_312 0 9.9999999999999998e-13
RS_311 NS_311 0 1.3258923845358959e+02
RS_312 NS_312 0 1.3258923845358959e+02
GL_311 0 NS_311 NS_312 0 5.6431081088718790e-02
GL_312 0 NS_312 NS_311 0 -5.6431081088718790e-02
GS_311_3 0 NS_311 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 313/314
CS_313 NS_313 0 9.9999999999999998e-13
CS_314 NS_314 0 9.9999999999999998e-13
RS_313 NS_313 0 1.0026704639246873e+02
RS_314 NS_314 0 1.0026704639246873e+02
GL_313 0 NS_313 NS_314 0 3.5068885856298401e-02
GL_314 0 NS_314 NS_313 0 -3.5068885856298401e-02
GS_313_3 0 NS_313 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 315/316
CS_315 NS_315 0 9.9999999999999998e-13
CS_316 NS_316 0 9.9999999999999998e-13
RS_315 NS_315 0 1.2740726499710033e+02
RS_316 NS_316 0 1.2740726499710034e+02
GL_315 0 NS_315 NS_316 0 5.3740629014256171e-02
GL_316 0 NS_316 NS_315 0 -5.3740629014256171e-02
GS_315_3 0 NS_315 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 317/318
CS_317 NS_317 0 9.9999999999999998e-13
CS_318 NS_318 0 9.9999999999999998e-13
RS_317 NS_317 0 2.3804688106534087e+02
RS_318 NS_318 0 2.3804688106534090e+02
GL_317 0 NS_317 NS_318 0 5.1425903265699464e-02
GL_318 0 NS_318 NS_317 0 -5.1425903265699464e-02
GS_317_3 0 NS_317 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 319/320
CS_319 NS_319 0 9.9999999999999998e-13
CS_320 NS_320 0 9.9999999999999998e-13
RS_319 NS_319 0 1.3728807739915800e+02
RS_320 NS_320 0 1.3728807739915803e+02
GL_319 0 NS_319 NS_320 0 4.8031392820534764e-02
GL_320 0 NS_320 NS_319 0 -4.8031392820534764e-02
GS_319_3 0 NS_319 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 321/322
CS_321 NS_321 0 9.9999999999999998e-13
CS_322 NS_322 0 9.9999999999999998e-13
RS_321 NS_321 0 1.3499477893747948e+02
RS_322 NS_322 0 1.3499477893747945e+02
GL_321 0 NS_321 NS_322 0 4.4453170742682194e-02
GL_322 0 NS_322 NS_321 0 -4.4453170742682194e-02
GS_321_3 0 NS_321 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 323/324
CS_323 NS_323 0 9.9999999999999998e-13
CS_324 NS_324 0 9.9999999999999998e-13
RS_323 NS_323 0 1.4121821834962651e+02
RS_324 NS_324 0 1.4121821834962651e+02
GL_323 0 NS_323 NS_324 0 3.8464469217755697e-02
GL_324 0 NS_324 NS_323 0 -3.8464469217755697e-02
GS_323_3 0 NS_323 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 325/326
CS_325 NS_325 0 9.9999999999999998e-13
CS_326 NS_326 0 9.9999999999999998e-13
RS_325 NS_325 0 1.3946471282741149e+02
RS_326 NS_326 0 1.3946471282741149e+02
GL_325 0 NS_325 NS_326 0 3.5678935079258622e-02
GL_326 0 NS_326 NS_325 0 -3.5678935079258622e-02
GS_325_3 0 NS_325 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 327/328
CS_327 NS_327 0 9.9999999999999998e-13
CS_328 NS_328 0 9.9999999999999998e-13
RS_327 NS_327 0 1.5530211191942624e+02
RS_328 NS_328 0 1.5530211191942627e+02
GL_327 0 NS_327 NS_328 0 2.6209890345437525e-02
GL_328 0 NS_328 NS_327 0 -2.6209890345437525e-02
GS_327_3 0 NS_327 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 329/330
CS_329 NS_329 0 9.9999999999999998e-13
CS_330 NS_330 0 9.9999999999999998e-13
RS_329 NS_329 0 1.4887428879582419e+02
RS_330 NS_330 0 1.4887428879582419e+02
GL_329 0 NS_329 NS_330 0 3.0330575323949095e-02
GL_330 0 NS_330 NS_329 0 -3.0330575323949095e-02
GS_329_3 0 NS_329 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 331/332
CS_331 NS_331 0 9.9999999999999998e-13
CS_332 NS_332 0 9.9999999999999998e-13
RS_331 NS_331 0 1.5087532095170570e+02
RS_332 NS_332 0 1.5087532095170570e+02
GL_331 0 NS_331 NS_332 0 2.0034138441714564e-02
GL_332 0 NS_332 NS_331 0 -2.0034138441714564e-02
GS_331_3 0 NS_331 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 333/334
CS_333 NS_333 0 9.9999999999999998e-13
CS_334 NS_334 0 9.9999999999999998e-13
RS_333 NS_333 0 1.4763793449752018e+02
RS_334 NS_334 0 1.4763793449752018e+02
GL_333 0 NS_333 NS_334 0 1.7017170579416537e-02
GL_334 0 NS_334 NS_333 0 -1.7017170579416537e-02
GS_333_3 0 NS_333 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 335/336
CS_335 NS_335 0 9.9999999999999998e-13
CS_336 NS_336 0 9.9999999999999998e-13
RS_335 NS_335 0 1.6285515224442304e+02
RS_336 NS_336 0 1.6285515224442304e+02
GL_335 0 NS_335 NS_336 0 1.0897027002452746e-02
GL_336 0 NS_336 NS_335 0 -1.0897027002452746e-02
GS_335_3 0 NS_335 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 337/338
CS_337 NS_337 0 9.9999999999999998e-13
CS_338 NS_338 0 9.9999999999999998e-13
RS_337 NS_337 0 1.7239534388116820e+02
RS_338 NS_338 0 1.7239534388116820e+02
GL_337 0 NS_337 NS_338 0 6.1589693699488982e-03
GL_338 0 NS_338 NS_337 0 -6.1589693699488982e-03
GS_337_3 0 NS_337 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 339/340
CS_339 NS_339 0 9.9999999999999998e-13
CS_340 NS_340 0 9.9999999999999998e-13
RS_339 NS_339 0 5.9928710578594173e+03
RS_340 NS_340 0 5.9928710578594173e+03
GL_339 0 NS_339 NS_340 0 1.7541178006601681e-03
GL_340 0 NS_340 NS_339 0 -1.7541178006601681e-03
GS_339_3 0 NS_339 NA_3 0 4.4027142044246531e-01
*
* Complex pair n. 341/342
CS_341 NS_341 0 9.9999999999999998e-13
CS_342 NS_342 0 9.9999999999999998e-13
RS_341 NS_341 0 8.0762087901330699e+02
RS_342 NS_342 0 8.0762087901330688e+02
GL_341 0 NS_341 NS_342 0 1.7295489372816217e-03
GL_342 0 NS_342 NS_341 0 -1.7295489372816217e-03
GS_341_3 0 NS_341 NA_3 0 4.4027142044246531e-01
*
* Real pole n. 343
CS_343 NS_343 0 9.9999999999999998e-13
RS_343 NS_343 0 1.2857601077426406e+01
GS_343_4 0 NS_343 NA_4 0 4.4027142044246531e-01
*
* Real pole n. 344
CS_344 NS_344 0 9.9999999999999998e-13
RS_344 NS_344 0 1.7282831464635029e+02
GS_344_4 0 NS_344 NA_4 0 4.4027142044246531e-01
*
* Real pole n. 345
CS_345 NS_345 0 9.9999999999999998e-13
RS_345 NS_345 0 5.5743135126264733e+03
GS_345_4 0 NS_345 NA_4 0 4.4027142044246531e-01
*
* Real pole n. 346
CS_346 NS_346 0 9.9999999999999998e-13
RS_346 NS_346 0 1.3594126013480764e+03
GS_346_4 0 NS_346 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 347/348
CS_347 NS_347 0 9.9999999999999998e-13
CS_348 NS_348 0 9.9999999999999998e-13
RS_347 NS_347 0 1.7904812183888848e+02
RS_348 NS_348 0 1.7904812183888848e+02
GL_347 0 NS_347 NS_348 0 2.6007898045516648e-01
GL_348 0 NS_348 NS_347 0 -2.6007898045516648e-01
GS_347_4 0 NS_347 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 349/350
CS_349 NS_349 0 9.9999999999999998e-13
CS_350 NS_350 0 9.9999999999999998e-13
RS_349 NS_349 0 1.2615541320340381e+02
RS_350 NS_350 0 1.2615541320340381e+02
GL_349 0 NS_349 NS_350 0 2.5243684762014923e-01
GL_350 0 NS_350 NS_349 0 -2.5243684762014923e-01
GS_349_4 0 NS_349 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 351/352
CS_351 NS_351 0 9.9999999999999998e-13
CS_352 NS_352 0 9.9999999999999998e-13
RS_351 NS_351 0 1.0219948841586964e+02
RS_352 NS_352 0 1.0219948841586965e+02
GL_351 0 NS_351 NS_352 0 2.4690226903121384e-01
GL_352 0 NS_352 NS_351 0 -2.4690226903121384e-01
GS_351_4 0 NS_351 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 353/354
CS_353 NS_353 0 9.9999999999999998e-13
CS_354 NS_354 0 9.9999999999999998e-13
RS_353 NS_353 0 1.1002436853144543e+02
RS_354 NS_354 0 1.1002436853144542e+02
GL_353 0 NS_353 NS_354 0 2.4293768067729948e-01
GL_354 0 NS_354 NS_353 0 -2.4293768067729948e-01
GS_353_4 0 NS_353 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 355/356
CS_355 NS_355 0 9.9999999999999998e-13
CS_356 NS_356 0 9.9999999999999998e-13
RS_355 NS_355 0 1.0553430908077024e+02
RS_356 NS_356 0 1.0553430908077026e+02
GL_355 0 NS_355 NS_356 0 2.3600513224442521e-01
GL_356 0 NS_356 NS_355 0 -2.3600513224442521e-01
GS_355_4 0 NS_355 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 357/358
CS_357 NS_357 0 9.9999999999999998e-13
CS_358 NS_358 0 9.9999999999999998e-13
RS_357 NS_357 0 1.0759915098440327e+02
RS_358 NS_358 0 1.0759915098440327e+02
GL_357 0 NS_357 NS_358 0 2.3090539914362113e-01
GL_358 0 NS_358 NS_357 0 -2.3090539914362113e-01
GS_357_4 0 NS_357 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 359/360
CS_359 NS_359 0 9.9999999999999998e-13
CS_360 NS_360 0 9.9999999999999998e-13
RS_359 NS_359 0 1.3295415758774385e+02
RS_360 NS_360 0 1.3295415758774385e+02
GL_359 0 NS_359 NS_360 0 2.3030066292345727e-01
GL_360 0 NS_360 NS_359 0 -2.3030066292345727e-01
GS_359_4 0 NS_359 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 361/362
CS_361 NS_361 0 9.9999999999999998e-13
CS_362 NS_362 0 9.9999999999999998e-13
RS_361 NS_361 0 1.1432186998941940e+02
RS_362 NS_362 0 1.1432186998941938e+02
GL_361 0 NS_361 NS_362 0 2.2451058023508991e-01
GL_362 0 NS_362 NS_361 0 -2.2451058023508991e-01
GS_361_4 0 NS_361 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 363/364
CS_363 NS_363 0 9.9999999999999998e-13
CS_364 NS_364 0 9.9999999999999998e-13
RS_363 NS_363 0 9.0812703249943667e+01
RS_364 NS_364 0 9.0812703249943652e+01
GL_363 0 NS_363 NS_364 0 2.1702628900531115e-01
GL_364 0 NS_364 NS_363 0 -2.1702628900531115e-01
GS_363_4 0 NS_363 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 365/366
CS_365 NS_365 0 9.9999999999999998e-13
CS_366 NS_366 0 9.9999999999999998e-13
RS_365 NS_365 0 9.5643803662064585e+01
RS_366 NS_366 0 9.5643803662064585e+01
GL_365 0 NS_365 NS_366 0 2.1448200383207913e-01
GL_366 0 NS_366 NS_365 0 -2.1448200383207913e-01
GS_365_4 0 NS_365 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 367/368
CS_367 NS_367 0 9.9999999999999998e-13
CS_368 NS_368 0 9.9999999999999998e-13
RS_367 NS_367 0 1.0631957479149644e+02
RS_368 NS_368 0 1.0631957479149644e+02
GL_367 0 NS_367 NS_368 0 2.0655001587884311e-01
GL_368 0 NS_368 NS_367 0 -2.0655001587884311e-01
GS_367_4 0 NS_367 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 369/370
CS_369 NS_369 0 9.9999999999999998e-13
CS_370 NS_370 0 9.9999999999999998e-13
RS_369 NS_369 0 7.9907264643295406e+01
RS_370 NS_370 0 7.9907264643295420e+01
GL_369 0 NS_369 NS_370 0 2.0133773147328893e-01
GL_370 0 NS_370 NS_369 0 -2.0133773147328893e-01
GS_369_4 0 NS_369 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 371/372
CS_371 NS_371 0 9.9999999999999998e-13
CS_372 NS_372 0 9.9999999999999998e-13
RS_371 NS_371 0 1.0625506887893997e+02
RS_372 NS_372 0 1.0625506887893997e+02
GL_371 0 NS_371 NS_372 0 1.9628877333023340e-01
GL_372 0 NS_372 NS_371 0 -1.9628877333023340e-01
GS_371_4 0 NS_371 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 373/374
CS_373 NS_373 0 9.9999999999999998e-13
CS_374 NS_374 0 9.9999999999999998e-13
RS_373 NS_373 0 9.6115312638592201e+01
RS_374 NS_374 0 9.6115312638592201e+01
GL_373 0 NS_373 NS_374 0 1.8794816712418483e-01
GL_374 0 NS_374 NS_373 0 -1.8794816712418483e-01
GS_373_4 0 NS_373 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 375/376
CS_375 NS_375 0 9.9999999999999998e-13
CS_376 NS_376 0 9.9999999999999998e-13
RS_375 NS_375 0 8.5212696574118169e+01
RS_376 NS_376 0 8.5212696574118169e+01
GL_375 0 NS_375 NS_376 0 1.8572140881490298e-01
GL_376 0 NS_376 NS_375 0 -1.8572140881490298e-01
GS_375_4 0 NS_375 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 377/378
CS_377 NS_377 0 9.9999999999999998e-13
CS_378 NS_378 0 9.9999999999999998e-13
RS_377 NS_377 0 1.0905026103375434e+02
RS_378 NS_378 0 1.0905026103375432e+02
GL_377 0 NS_377 NS_378 0 1.7785621200284463e-01
GL_378 0 NS_378 NS_377 0 -1.7785621200284463e-01
GS_377_4 0 NS_377 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 379/380
CS_379 NS_379 0 9.9999999999999998e-13
CS_380 NS_380 0 9.9999999999999998e-13
RS_379 NS_379 0 8.3024437910787526e+01
RS_380 NS_380 0 8.3024437910787526e+01
GL_379 0 NS_379 NS_380 0 1.7164509875911016e-01
GL_380 0 NS_380 NS_379 0 -1.7164509875911016e-01
GS_379_4 0 NS_379 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 381/382
CS_381 NS_381 0 9.9999999999999998e-13
CS_382 NS_382 0 9.9999999999999998e-13
RS_381 NS_381 0 1.0548793856392000e+02
RS_382 NS_382 0 1.0548793856392000e+02
GL_381 0 NS_381 NS_382 0 1.6750370916002649e-01
GL_382 0 NS_382 NS_381 0 -1.6750370916002649e-01
GS_381_4 0 NS_381 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 383/384
CS_383 NS_383 0 9.9999999999999998e-13
CS_384 NS_384 0 9.9999999999999998e-13
RS_383 NS_383 0 1.0753754351502513e+02
RS_384 NS_384 0 1.0753754351502513e+02
GL_383 0 NS_383 NS_384 0 1.5942172238060490e-01
GL_384 0 NS_384 NS_383 0 -1.5942172238060490e-01
GS_383_4 0 NS_383 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 385/386
CS_385 NS_385 0 9.9999999999999998e-13
CS_386 NS_386 0 9.9999999999999998e-13
RS_385 NS_385 0 8.6961097797504721e+01
RS_386 NS_386 0 8.6961097797504721e+01
GL_385 0 NS_385 NS_386 0 1.5553892891442009e-01
GL_386 0 NS_386 NS_385 0 -1.5553892891442009e-01
GS_385_4 0 NS_385 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 387/388
CS_387 NS_387 0 9.9999999999999998e-13
CS_388 NS_388 0 9.9999999999999998e-13
RS_387 NS_387 0 1.1549771364055694e+02
RS_388 NS_388 0 1.1549771364055692e+02
GL_387 0 NS_387 NS_388 0 1.4899166019107438e-01
GL_388 0 NS_388 NS_387 0 -1.4899166019107438e-01
GS_387_4 0 NS_387 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 389/390
CS_389 NS_389 0 9.9999999999999998e-13
CS_390 NS_390 0 9.9999999999999998e-13
RS_389 NS_389 0 9.7194462506038604e+01
RS_390 NS_390 0 9.7194462506038604e+01
GL_389 0 NS_389 NS_390 0 1.4180400817347408e-01
GL_390 0 NS_390 NS_389 0 -1.4180400817347408e-01
GS_389_4 0 NS_389 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 391/392
CS_391 NS_391 0 9.9999999999999998e-13
CS_392 NS_392 0 9.9999999999999998e-13
RS_391 NS_391 0 1.0682825030924828e+02
RS_392 NS_392 0 1.0682825030924828e+02
GL_391 0 NS_391 NS_392 0 1.3872377519751058e-01
GL_392 0 NS_392 NS_391 0 -1.3872377519751058e-01
GS_391_4 0 NS_391 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 393/394
CS_393 NS_393 0 9.9999999999999998e-13
CS_394 NS_394 0 9.9999999999999998e-13
RS_393 NS_393 0 1.2559585119344567e+02
RS_394 NS_394 0 1.2559585119344568e+02
GL_393 0 NS_393 NS_394 0 1.3097721803321302e-01
GL_394 0 NS_394 NS_393 0 -1.3097721803321302e-01
GS_393_4 0 NS_393 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 395/396
CS_395 NS_395 0 9.9999999999999998e-13
CS_396 NS_396 0 9.9999999999999998e-13
RS_395 NS_395 0 1.0417660462554996e+02
RS_396 NS_396 0 1.0417660462554996e+02
GL_395 0 NS_395 NS_396 0 1.2625832867930367e-01
GL_396 0 NS_396 NS_395 0 -1.2625832867930367e-01
GS_395_4 0 NS_395 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 397/398
CS_397 NS_397 0 9.9999999999999998e-13
CS_398 NS_398 0 9.9999999999999998e-13
RS_397 NS_397 0 1.3317333532177352e+02
RS_398 NS_398 0 1.3317333532177352e+02
GL_397 0 NS_397 NS_398 0 1.2123672752714061e-01
GL_398 0 NS_398 NS_397 0 -1.2123672752714061e-01
GS_397_4 0 NS_397 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 399/400
CS_399 NS_399 0 9.9999999999999998e-13
CS_400 NS_400 0 9.9999999999999998e-13
RS_399 NS_399 0 1.2967831681616519e+02
RS_400 NS_400 0 1.2967831681616519e+02
GL_399 0 NS_399 NS_400 0 1.1651127865768855e-01
GL_400 0 NS_400 NS_399 0 -1.1651127865768855e-01
GS_399_4 0 NS_399 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 401/402
CS_401 NS_401 0 9.9999999999999998e-13
CS_402 NS_402 0 9.9999999999999998e-13
RS_401 NS_401 0 1.2999764374401394e+02
RS_402 NS_402 0 1.2999764374401394e+02
GL_401 0 NS_401 NS_402 0 1.1100247696987056e-01
GL_402 0 NS_402 NS_401 0 -1.1100247696987056e-01
GS_401_4 0 NS_401 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 403/404
CS_403 NS_403 0 9.9999999999999998e-13
CS_404 NS_404 0 9.9999999999999998e-13
RS_403 NS_403 0 1.2458814074636419e+02
RS_404 NS_404 0 1.2458814074636419e+02
GL_403 0 NS_403 NS_404 0 1.0660000212580591e-01
GL_404 0 NS_404 NS_403 0 -1.0660000212580591e-01
GS_403_4 0 NS_403 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 405/406
CS_405 NS_405 0 9.9999999999999998e-13
CS_406 NS_406 0 9.9999999999999998e-13
RS_405 NS_405 0 1.4677191614557748e+02
RS_406 NS_406 0 1.4677191614557748e+02
GL_405 0 NS_405 NS_406 0 1.0224733343325158e-01
GL_406 0 NS_406 NS_405 0 -1.0224733343325158e-01
GS_405_4 0 NS_405 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 407/408
CS_407 NS_407 0 9.9999999999999998e-13
CS_408 NS_408 0 9.9999999999999998e-13
RS_407 NS_407 0 1.3445989223131798e+02
RS_408 NS_408 0 1.3445989223131798e+02
GL_407 0 NS_407 NS_408 0 9.8177836948086503e-02
GL_408 0 NS_408 NS_407 0 -9.8177836948086503e-02
GS_407_4 0 NS_407 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 409/410
CS_409 NS_409 0 9.9999999999999998e-13
CS_410 NS_410 0 9.9999999999999998e-13
RS_409 NS_409 0 1.3187119040723775e+02
RS_410 NS_410 0 1.3187119040723772e+02
GL_409 0 NS_409 NS_410 0 9.2640196004122682e-02
GL_410 0 NS_410 NS_409 0 -9.2640196004122682e-02
GS_409_4 0 NS_409 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 411/412
CS_411 NS_411 0 9.9999999999999998e-13
CS_412 NS_412 0 9.9999999999999998e-13
RS_411 NS_411 0 1.2288401421230557e+02
RS_412 NS_412 0 1.2288401421230557e+02
GL_411 0 NS_411 NS_412 0 8.8704723748248199e-02
GL_412 0 NS_412 NS_411 0 -8.8704723748248199e-02
GS_411_4 0 NS_411 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 413/414
CS_413 NS_413 0 9.9999999999999998e-13
CS_414 NS_414 0 9.9999999999999998e-13
RS_413 NS_413 0 1.4123955654153085e+02
RS_414 NS_414 0 1.4123955654153082e+02
GL_413 0 NS_413 NS_414 0 8.4112474498892476e-02
GL_414 0 NS_414 NS_413 0 -8.4112474498892476e-02
GS_413_4 0 NS_413 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 415/416
CS_415 NS_415 0 9.9999999999999998e-13
CS_416 NS_416 0 9.9999999999999998e-13
RS_415 NS_415 0 1.2539447312269779e+02
RS_416 NS_416 0 1.2539447312269778e+02
GL_415 0 NS_415 NS_416 0 8.0007658848305588e-02
GL_416 0 NS_416 NS_415 0 -8.0007658848305588e-02
GS_415_4 0 NS_415 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 417/418
CS_417 NS_417 0 9.9999999999999998e-13
CS_418 NS_418 0 9.9999999999999998e-13
RS_417 NS_417 0 1.3219601779966965e+02
RS_418 NS_418 0 1.3219601779966968e+02
GL_417 0 NS_417 NS_418 0 7.4373183806052026e-02
GL_418 0 NS_418 NS_417 0 -7.4373183806052026e-02
GS_417_4 0 NS_417 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 419/420
CS_419 NS_419 0 9.9999999999999998e-13
CS_420 NS_420 0 9.9999999999999998e-13
RS_419 NS_419 0 1.1951371640958898e+02
RS_420 NS_420 0 1.1951371640958898e+02
GL_419 0 NS_419 NS_420 0 7.1003860961129844e-02
GL_420 0 NS_420 NS_419 0 -7.1003860961129844e-02
GS_419_4 0 NS_419 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 421/422
CS_421 NS_421 0 9.9999999999999998e-13
CS_422 NS_422 0 9.9999999999999998e-13
RS_421 NS_421 0 1.3491941875045018e+02
RS_422 NS_422 0 1.3491941875045018e+02
GL_421 0 NS_421 NS_422 0 6.5922080709048564e-02
GL_422 0 NS_422 NS_421 0 -6.5922080709048564e-02
GS_421_4 0 NS_421 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 423/424
CS_423 NS_423 0 9.9999999999999998e-13
CS_424 NS_424 0 9.9999999999999998e-13
RS_423 NS_423 0 1.2290405859347165e+02
RS_424 NS_424 0 1.2290405859347166e+02
GL_423 0 NS_423 NS_424 0 6.2340152915784278e-02
GL_424 0 NS_424 NS_423 0 -6.2340152915784278e-02
GS_423_4 0 NS_423 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 425/426
CS_425 NS_425 0 9.9999999999999998e-13
CS_426 NS_426 0 9.9999999999999998e-13
RS_425 NS_425 0 1.3258923845358959e+02
RS_426 NS_426 0 1.3258923845358959e+02
GL_425 0 NS_425 NS_426 0 5.6431081088718790e-02
GL_426 0 NS_426 NS_425 0 -5.6431081088718790e-02
GS_425_4 0 NS_425 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 427/428
CS_427 NS_427 0 9.9999999999999998e-13
CS_428 NS_428 0 9.9999999999999998e-13
RS_427 NS_427 0 1.0026704639246873e+02
RS_428 NS_428 0 1.0026704639246873e+02
GL_427 0 NS_427 NS_428 0 3.5068885856298401e-02
GL_428 0 NS_428 NS_427 0 -3.5068885856298401e-02
GS_427_4 0 NS_427 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 429/430
CS_429 NS_429 0 9.9999999999999998e-13
CS_430 NS_430 0 9.9999999999999998e-13
RS_429 NS_429 0 1.2740726499710033e+02
RS_430 NS_430 0 1.2740726499710034e+02
GL_429 0 NS_429 NS_430 0 5.3740629014256171e-02
GL_430 0 NS_430 NS_429 0 -5.3740629014256171e-02
GS_429_4 0 NS_429 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 431/432
CS_431 NS_431 0 9.9999999999999998e-13
CS_432 NS_432 0 9.9999999999999998e-13
RS_431 NS_431 0 2.3804688106534087e+02
RS_432 NS_432 0 2.3804688106534090e+02
GL_431 0 NS_431 NS_432 0 5.1425903265699464e-02
GL_432 0 NS_432 NS_431 0 -5.1425903265699464e-02
GS_431_4 0 NS_431 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 433/434
CS_433 NS_433 0 9.9999999999999998e-13
CS_434 NS_434 0 9.9999999999999998e-13
RS_433 NS_433 0 1.3728807739915800e+02
RS_434 NS_434 0 1.3728807739915803e+02
GL_433 0 NS_433 NS_434 0 4.8031392820534764e-02
GL_434 0 NS_434 NS_433 0 -4.8031392820534764e-02
GS_433_4 0 NS_433 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 435/436
CS_435 NS_435 0 9.9999999999999998e-13
CS_436 NS_436 0 9.9999999999999998e-13
RS_435 NS_435 0 1.3499477893747948e+02
RS_436 NS_436 0 1.3499477893747945e+02
GL_435 0 NS_435 NS_436 0 4.4453170742682194e-02
GL_436 0 NS_436 NS_435 0 -4.4453170742682194e-02
GS_435_4 0 NS_435 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 437/438
CS_437 NS_437 0 9.9999999999999998e-13
CS_438 NS_438 0 9.9999999999999998e-13
RS_437 NS_437 0 1.4121821834962651e+02
RS_438 NS_438 0 1.4121821834962651e+02
GL_437 0 NS_437 NS_438 0 3.8464469217755697e-02
GL_438 0 NS_438 NS_437 0 -3.8464469217755697e-02
GS_437_4 0 NS_437 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 439/440
CS_439 NS_439 0 9.9999999999999998e-13
CS_440 NS_440 0 9.9999999999999998e-13
RS_439 NS_439 0 1.3946471282741149e+02
RS_440 NS_440 0 1.3946471282741149e+02
GL_439 0 NS_439 NS_440 0 3.5678935079258622e-02
GL_440 0 NS_440 NS_439 0 -3.5678935079258622e-02
GS_439_4 0 NS_439 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 441/442
CS_441 NS_441 0 9.9999999999999998e-13
CS_442 NS_442 0 9.9999999999999998e-13
RS_441 NS_441 0 1.5530211191942624e+02
RS_442 NS_442 0 1.5530211191942627e+02
GL_441 0 NS_441 NS_442 0 2.6209890345437525e-02
GL_442 0 NS_442 NS_441 0 -2.6209890345437525e-02
GS_441_4 0 NS_441 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 443/444
CS_443 NS_443 0 9.9999999999999998e-13
CS_444 NS_444 0 9.9999999999999998e-13
RS_443 NS_443 0 1.4887428879582419e+02
RS_444 NS_444 0 1.4887428879582419e+02
GL_443 0 NS_443 NS_444 0 3.0330575323949095e-02
GL_444 0 NS_444 NS_443 0 -3.0330575323949095e-02
GS_443_4 0 NS_443 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 445/446
CS_445 NS_445 0 9.9999999999999998e-13
CS_446 NS_446 0 9.9999999999999998e-13
RS_445 NS_445 0 1.5087532095170570e+02
RS_446 NS_446 0 1.5087532095170570e+02
GL_445 0 NS_445 NS_446 0 2.0034138441714564e-02
GL_446 0 NS_446 NS_445 0 -2.0034138441714564e-02
GS_445_4 0 NS_445 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 447/448
CS_447 NS_447 0 9.9999999999999998e-13
CS_448 NS_448 0 9.9999999999999998e-13
RS_447 NS_447 0 1.4763793449752018e+02
RS_448 NS_448 0 1.4763793449752018e+02
GL_447 0 NS_447 NS_448 0 1.7017170579416537e-02
GL_448 0 NS_448 NS_447 0 -1.7017170579416537e-02
GS_447_4 0 NS_447 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 449/450
CS_449 NS_449 0 9.9999999999999998e-13
CS_450 NS_450 0 9.9999999999999998e-13
RS_449 NS_449 0 1.6285515224442304e+02
RS_450 NS_450 0 1.6285515224442304e+02
GL_449 0 NS_449 NS_450 0 1.0897027002452746e-02
GL_450 0 NS_450 NS_449 0 -1.0897027002452746e-02
GS_449_4 0 NS_449 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 451/452
CS_451 NS_451 0 9.9999999999999998e-13
CS_452 NS_452 0 9.9999999999999998e-13
RS_451 NS_451 0 1.7239534388116820e+02
RS_452 NS_452 0 1.7239534388116820e+02
GL_451 0 NS_451 NS_452 0 6.1589693699488982e-03
GL_452 0 NS_452 NS_451 0 -6.1589693699488982e-03
GS_451_4 0 NS_451 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 453/454
CS_453 NS_453 0 9.9999999999999998e-13
CS_454 NS_454 0 9.9999999999999998e-13
RS_453 NS_453 0 5.9928710578594173e+03
RS_454 NS_454 0 5.9928710578594173e+03
GL_453 0 NS_453 NS_454 0 1.7541178006601681e-03
GL_454 0 NS_454 NS_453 0 -1.7541178006601681e-03
GS_453_4 0 NS_453 NA_4 0 4.4027142044246531e-01
*
* Complex pair n. 455/456
CS_455 NS_455 0 9.9999999999999998e-13
CS_456 NS_456 0 9.9999999999999998e-13
RS_455 NS_455 0 8.0762087901330699e+02
RS_456 NS_456 0 8.0762087901330688e+02
GL_455 0 NS_455 NS_456 0 1.7295489372816217e-03
GL_456 0 NS_456 NS_455 0 -1.7295489372816217e-03
GS_455_4 0 NS_455 NA_4 0 4.4027142044246531e-01
*
* Real pole n. 457
CS_457 NS_457 0 9.9999999999999998e-13
RS_457 NS_457 0 1.2857601077426406e+01
GS_457_5 0 NS_457 NA_5 0 4.4027142044246531e-01
*
* Real pole n. 458
CS_458 NS_458 0 9.9999999999999998e-13
RS_458 NS_458 0 1.7282831464635029e+02
GS_458_5 0 NS_458 NA_5 0 4.4027142044246531e-01
*
* Real pole n. 459
CS_459 NS_459 0 9.9999999999999998e-13
RS_459 NS_459 0 5.5743135126264733e+03
GS_459_5 0 NS_459 NA_5 0 4.4027142044246531e-01
*
* Real pole n. 460
CS_460 NS_460 0 9.9999999999999998e-13
RS_460 NS_460 0 1.3594126013480764e+03
GS_460_5 0 NS_460 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 461/462
CS_461 NS_461 0 9.9999999999999998e-13
CS_462 NS_462 0 9.9999999999999998e-13
RS_461 NS_461 0 1.7904812183888848e+02
RS_462 NS_462 0 1.7904812183888848e+02
GL_461 0 NS_461 NS_462 0 2.6007898045516648e-01
GL_462 0 NS_462 NS_461 0 -2.6007898045516648e-01
GS_461_5 0 NS_461 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 463/464
CS_463 NS_463 0 9.9999999999999998e-13
CS_464 NS_464 0 9.9999999999999998e-13
RS_463 NS_463 0 1.2615541320340381e+02
RS_464 NS_464 0 1.2615541320340381e+02
GL_463 0 NS_463 NS_464 0 2.5243684762014923e-01
GL_464 0 NS_464 NS_463 0 -2.5243684762014923e-01
GS_463_5 0 NS_463 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 465/466
CS_465 NS_465 0 9.9999999999999998e-13
CS_466 NS_466 0 9.9999999999999998e-13
RS_465 NS_465 0 1.0219948841586964e+02
RS_466 NS_466 0 1.0219948841586965e+02
GL_465 0 NS_465 NS_466 0 2.4690226903121384e-01
GL_466 0 NS_466 NS_465 0 -2.4690226903121384e-01
GS_465_5 0 NS_465 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 467/468
CS_467 NS_467 0 9.9999999999999998e-13
CS_468 NS_468 0 9.9999999999999998e-13
RS_467 NS_467 0 1.1002436853144543e+02
RS_468 NS_468 0 1.1002436853144542e+02
GL_467 0 NS_467 NS_468 0 2.4293768067729948e-01
GL_468 0 NS_468 NS_467 0 -2.4293768067729948e-01
GS_467_5 0 NS_467 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 469/470
CS_469 NS_469 0 9.9999999999999998e-13
CS_470 NS_470 0 9.9999999999999998e-13
RS_469 NS_469 0 1.0553430908077024e+02
RS_470 NS_470 0 1.0553430908077026e+02
GL_469 0 NS_469 NS_470 0 2.3600513224442521e-01
GL_470 0 NS_470 NS_469 0 -2.3600513224442521e-01
GS_469_5 0 NS_469 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 471/472
CS_471 NS_471 0 9.9999999999999998e-13
CS_472 NS_472 0 9.9999999999999998e-13
RS_471 NS_471 0 1.0759915098440327e+02
RS_472 NS_472 0 1.0759915098440327e+02
GL_471 0 NS_471 NS_472 0 2.3090539914362113e-01
GL_472 0 NS_472 NS_471 0 -2.3090539914362113e-01
GS_471_5 0 NS_471 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 473/474
CS_473 NS_473 0 9.9999999999999998e-13
CS_474 NS_474 0 9.9999999999999998e-13
RS_473 NS_473 0 1.3295415758774385e+02
RS_474 NS_474 0 1.3295415758774385e+02
GL_473 0 NS_473 NS_474 0 2.3030066292345727e-01
GL_474 0 NS_474 NS_473 0 -2.3030066292345727e-01
GS_473_5 0 NS_473 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 475/476
CS_475 NS_475 0 9.9999999999999998e-13
CS_476 NS_476 0 9.9999999999999998e-13
RS_475 NS_475 0 1.1432186998941940e+02
RS_476 NS_476 0 1.1432186998941938e+02
GL_475 0 NS_475 NS_476 0 2.2451058023508991e-01
GL_476 0 NS_476 NS_475 0 -2.2451058023508991e-01
GS_475_5 0 NS_475 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 477/478
CS_477 NS_477 0 9.9999999999999998e-13
CS_478 NS_478 0 9.9999999999999998e-13
RS_477 NS_477 0 9.0812703249943667e+01
RS_478 NS_478 0 9.0812703249943652e+01
GL_477 0 NS_477 NS_478 0 2.1702628900531115e-01
GL_478 0 NS_478 NS_477 0 -2.1702628900531115e-01
GS_477_5 0 NS_477 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 479/480
CS_479 NS_479 0 9.9999999999999998e-13
CS_480 NS_480 0 9.9999999999999998e-13
RS_479 NS_479 0 9.5643803662064585e+01
RS_480 NS_480 0 9.5643803662064585e+01
GL_479 0 NS_479 NS_480 0 2.1448200383207913e-01
GL_480 0 NS_480 NS_479 0 -2.1448200383207913e-01
GS_479_5 0 NS_479 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 481/482
CS_481 NS_481 0 9.9999999999999998e-13
CS_482 NS_482 0 9.9999999999999998e-13
RS_481 NS_481 0 1.0631957479149644e+02
RS_482 NS_482 0 1.0631957479149644e+02
GL_481 0 NS_481 NS_482 0 2.0655001587884311e-01
GL_482 0 NS_482 NS_481 0 -2.0655001587884311e-01
GS_481_5 0 NS_481 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 483/484
CS_483 NS_483 0 9.9999999999999998e-13
CS_484 NS_484 0 9.9999999999999998e-13
RS_483 NS_483 0 7.9907264643295406e+01
RS_484 NS_484 0 7.9907264643295420e+01
GL_483 0 NS_483 NS_484 0 2.0133773147328893e-01
GL_484 0 NS_484 NS_483 0 -2.0133773147328893e-01
GS_483_5 0 NS_483 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 485/486
CS_485 NS_485 0 9.9999999999999998e-13
CS_486 NS_486 0 9.9999999999999998e-13
RS_485 NS_485 0 1.0625506887893997e+02
RS_486 NS_486 0 1.0625506887893997e+02
GL_485 0 NS_485 NS_486 0 1.9628877333023340e-01
GL_486 0 NS_486 NS_485 0 -1.9628877333023340e-01
GS_485_5 0 NS_485 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 487/488
CS_487 NS_487 0 9.9999999999999998e-13
CS_488 NS_488 0 9.9999999999999998e-13
RS_487 NS_487 0 9.6115312638592201e+01
RS_488 NS_488 0 9.6115312638592201e+01
GL_487 0 NS_487 NS_488 0 1.8794816712418483e-01
GL_488 0 NS_488 NS_487 0 -1.8794816712418483e-01
GS_487_5 0 NS_487 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 489/490
CS_489 NS_489 0 9.9999999999999998e-13
CS_490 NS_490 0 9.9999999999999998e-13
RS_489 NS_489 0 8.5212696574118169e+01
RS_490 NS_490 0 8.5212696574118169e+01
GL_489 0 NS_489 NS_490 0 1.8572140881490298e-01
GL_490 0 NS_490 NS_489 0 -1.8572140881490298e-01
GS_489_5 0 NS_489 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 491/492
CS_491 NS_491 0 9.9999999999999998e-13
CS_492 NS_492 0 9.9999999999999998e-13
RS_491 NS_491 0 1.0905026103375434e+02
RS_492 NS_492 0 1.0905026103375432e+02
GL_491 0 NS_491 NS_492 0 1.7785621200284463e-01
GL_492 0 NS_492 NS_491 0 -1.7785621200284463e-01
GS_491_5 0 NS_491 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 493/494
CS_493 NS_493 0 9.9999999999999998e-13
CS_494 NS_494 0 9.9999999999999998e-13
RS_493 NS_493 0 8.3024437910787526e+01
RS_494 NS_494 0 8.3024437910787526e+01
GL_493 0 NS_493 NS_494 0 1.7164509875911016e-01
GL_494 0 NS_494 NS_493 0 -1.7164509875911016e-01
GS_493_5 0 NS_493 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 495/496
CS_495 NS_495 0 9.9999999999999998e-13
CS_496 NS_496 0 9.9999999999999998e-13
RS_495 NS_495 0 1.0548793856392000e+02
RS_496 NS_496 0 1.0548793856392000e+02
GL_495 0 NS_495 NS_496 0 1.6750370916002649e-01
GL_496 0 NS_496 NS_495 0 -1.6750370916002649e-01
GS_495_5 0 NS_495 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 497/498
CS_497 NS_497 0 9.9999999999999998e-13
CS_498 NS_498 0 9.9999999999999998e-13
RS_497 NS_497 0 1.0753754351502513e+02
RS_498 NS_498 0 1.0753754351502513e+02
GL_497 0 NS_497 NS_498 0 1.5942172238060490e-01
GL_498 0 NS_498 NS_497 0 -1.5942172238060490e-01
GS_497_5 0 NS_497 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 499/500
CS_499 NS_499 0 9.9999999999999998e-13
CS_500 NS_500 0 9.9999999999999998e-13
RS_499 NS_499 0 8.6961097797504721e+01
RS_500 NS_500 0 8.6961097797504721e+01
GL_499 0 NS_499 NS_500 0 1.5553892891442009e-01
GL_500 0 NS_500 NS_499 0 -1.5553892891442009e-01
GS_499_5 0 NS_499 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 501/502
CS_501 NS_501 0 9.9999999999999998e-13
CS_502 NS_502 0 9.9999999999999998e-13
RS_501 NS_501 0 1.1549771364055694e+02
RS_502 NS_502 0 1.1549771364055692e+02
GL_501 0 NS_501 NS_502 0 1.4899166019107438e-01
GL_502 0 NS_502 NS_501 0 -1.4899166019107438e-01
GS_501_5 0 NS_501 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 503/504
CS_503 NS_503 0 9.9999999999999998e-13
CS_504 NS_504 0 9.9999999999999998e-13
RS_503 NS_503 0 9.7194462506038604e+01
RS_504 NS_504 0 9.7194462506038604e+01
GL_503 0 NS_503 NS_504 0 1.4180400817347408e-01
GL_504 0 NS_504 NS_503 0 -1.4180400817347408e-01
GS_503_5 0 NS_503 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 505/506
CS_505 NS_505 0 9.9999999999999998e-13
CS_506 NS_506 0 9.9999999999999998e-13
RS_505 NS_505 0 1.0682825030924828e+02
RS_506 NS_506 0 1.0682825030924828e+02
GL_505 0 NS_505 NS_506 0 1.3872377519751058e-01
GL_506 0 NS_506 NS_505 0 -1.3872377519751058e-01
GS_505_5 0 NS_505 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 507/508
CS_507 NS_507 0 9.9999999999999998e-13
CS_508 NS_508 0 9.9999999999999998e-13
RS_507 NS_507 0 1.2559585119344567e+02
RS_508 NS_508 0 1.2559585119344568e+02
GL_507 0 NS_507 NS_508 0 1.3097721803321302e-01
GL_508 0 NS_508 NS_507 0 -1.3097721803321302e-01
GS_507_5 0 NS_507 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 509/510
CS_509 NS_509 0 9.9999999999999998e-13
CS_510 NS_510 0 9.9999999999999998e-13
RS_509 NS_509 0 1.0417660462554996e+02
RS_510 NS_510 0 1.0417660462554996e+02
GL_509 0 NS_509 NS_510 0 1.2625832867930367e-01
GL_510 0 NS_510 NS_509 0 -1.2625832867930367e-01
GS_509_5 0 NS_509 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 511/512
CS_511 NS_511 0 9.9999999999999998e-13
CS_512 NS_512 0 9.9999999999999998e-13
RS_511 NS_511 0 1.3317333532177352e+02
RS_512 NS_512 0 1.3317333532177352e+02
GL_511 0 NS_511 NS_512 0 1.2123672752714061e-01
GL_512 0 NS_512 NS_511 0 -1.2123672752714061e-01
GS_511_5 0 NS_511 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 513/514
CS_513 NS_513 0 9.9999999999999998e-13
CS_514 NS_514 0 9.9999999999999998e-13
RS_513 NS_513 0 1.2967831681616519e+02
RS_514 NS_514 0 1.2967831681616519e+02
GL_513 0 NS_513 NS_514 0 1.1651127865768855e-01
GL_514 0 NS_514 NS_513 0 -1.1651127865768855e-01
GS_513_5 0 NS_513 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 515/516
CS_515 NS_515 0 9.9999999999999998e-13
CS_516 NS_516 0 9.9999999999999998e-13
RS_515 NS_515 0 1.2999764374401394e+02
RS_516 NS_516 0 1.2999764374401394e+02
GL_515 0 NS_515 NS_516 0 1.1100247696987056e-01
GL_516 0 NS_516 NS_515 0 -1.1100247696987056e-01
GS_515_5 0 NS_515 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 517/518
CS_517 NS_517 0 9.9999999999999998e-13
CS_518 NS_518 0 9.9999999999999998e-13
RS_517 NS_517 0 1.2458814074636419e+02
RS_518 NS_518 0 1.2458814074636419e+02
GL_517 0 NS_517 NS_518 0 1.0660000212580591e-01
GL_518 0 NS_518 NS_517 0 -1.0660000212580591e-01
GS_517_5 0 NS_517 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 519/520
CS_519 NS_519 0 9.9999999999999998e-13
CS_520 NS_520 0 9.9999999999999998e-13
RS_519 NS_519 0 1.4677191614557748e+02
RS_520 NS_520 0 1.4677191614557748e+02
GL_519 0 NS_519 NS_520 0 1.0224733343325158e-01
GL_520 0 NS_520 NS_519 0 -1.0224733343325158e-01
GS_519_5 0 NS_519 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 521/522
CS_521 NS_521 0 9.9999999999999998e-13
CS_522 NS_522 0 9.9999999999999998e-13
RS_521 NS_521 0 1.3445989223131798e+02
RS_522 NS_522 0 1.3445989223131798e+02
GL_521 0 NS_521 NS_522 0 9.8177836948086503e-02
GL_522 0 NS_522 NS_521 0 -9.8177836948086503e-02
GS_521_5 0 NS_521 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 523/524
CS_523 NS_523 0 9.9999999999999998e-13
CS_524 NS_524 0 9.9999999999999998e-13
RS_523 NS_523 0 1.3187119040723775e+02
RS_524 NS_524 0 1.3187119040723772e+02
GL_523 0 NS_523 NS_524 0 9.2640196004122682e-02
GL_524 0 NS_524 NS_523 0 -9.2640196004122682e-02
GS_523_5 0 NS_523 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 525/526
CS_525 NS_525 0 9.9999999999999998e-13
CS_526 NS_526 0 9.9999999999999998e-13
RS_525 NS_525 0 1.2288401421230557e+02
RS_526 NS_526 0 1.2288401421230557e+02
GL_525 0 NS_525 NS_526 0 8.8704723748248199e-02
GL_526 0 NS_526 NS_525 0 -8.8704723748248199e-02
GS_525_5 0 NS_525 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 527/528
CS_527 NS_527 0 9.9999999999999998e-13
CS_528 NS_528 0 9.9999999999999998e-13
RS_527 NS_527 0 1.4123955654153085e+02
RS_528 NS_528 0 1.4123955654153082e+02
GL_527 0 NS_527 NS_528 0 8.4112474498892476e-02
GL_528 0 NS_528 NS_527 0 -8.4112474498892476e-02
GS_527_5 0 NS_527 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 529/530
CS_529 NS_529 0 9.9999999999999998e-13
CS_530 NS_530 0 9.9999999999999998e-13
RS_529 NS_529 0 1.2539447312269779e+02
RS_530 NS_530 0 1.2539447312269778e+02
GL_529 0 NS_529 NS_530 0 8.0007658848305588e-02
GL_530 0 NS_530 NS_529 0 -8.0007658848305588e-02
GS_529_5 0 NS_529 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 531/532
CS_531 NS_531 0 9.9999999999999998e-13
CS_532 NS_532 0 9.9999999999999998e-13
RS_531 NS_531 0 1.3219601779966965e+02
RS_532 NS_532 0 1.3219601779966968e+02
GL_531 0 NS_531 NS_532 0 7.4373183806052026e-02
GL_532 0 NS_532 NS_531 0 -7.4373183806052026e-02
GS_531_5 0 NS_531 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 533/534
CS_533 NS_533 0 9.9999999999999998e-13
CS_534 NS_534 0 9.9999999999999998e-13
RS_533 NS_533 0 1.1951371640958898e+02
RS_534 NS_534 0 1.1951371640958898e+02
GL_533 0 NS_533 NS_534 0 7.1003860961129844e-02
GL_534 0 NS_534 NS_533 0 -7.1003860961129844e-02
GS_533_5 0 NS_533 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 535/536
CS_535 NS_535 0 9.9999999999999998e-13
CS_536 NS_536 0 9.9999999999999998e-13
RS_535 NS_535 0 1.3491941875045018e+02
RS_536 NS_536 0 1.3491941875045018e+02
GL_535 0 NS_535 NS_536 0 6.5922080709048564e-02
GL_536 0 NS_536 NS_535 0 -6.5922080709048564e-02
GS_535_5 0 NS_535 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 537/538
CS_537 NS_537 0 9.9999999999999998e-13
CS_538 NS_538 0 9.9999999999999998e-13
RS_537 NS_537 0 1.2290405859347165e+02
RS_538 NS_538 0 1.2290405859347166e+02
GL_537 0 NS_537 NS_538 0 6.2340152915784278e-02
GL_538 0 NS_538 NS_537 0 -6.2340152915784278e-02
GS_537_5 0 NS_537 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 539/540
CS_539 NS_539 0 9.9999999999999998e-13
CS_540 NS_540 0 9.9999999999999998e-13
RS_539 NS_539 0 1.3258923845358959e+02
RS_540 NS_540 0 1.3258923845358959e+02
GL_539 0 NS_539 NS_540 0 5.6431081088718790e-02
GL_540 0 NS_540 NS_539 0 -5.6431081088718790e-02
GS_539_5 0 NS_539 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 541/542
CS_541 NS_541 0 9.9999999999999998e-13
CS_542 NS_542 0 9.9999999999999998e-13
RS_541 NS_541 0 1.0026704639246873e+02
RS_542 NS_542 0 1.0026704639246873e+02
GL_541 0 NS_541 NS_542 0 3.5068885856298401e-02
GL_542 0 NS_542 NS_541 0 -3.5068885856298401e-02
GS_541_5 0 NS_541 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 543/544
CS_543 NS_543 0 9.9999999999999998e-13
CS_544 NS_544 0 9.9999999999999998e-13
RS_543 NS_543 0 1.2740726499710033e+02
RS_544 NS_544 0 1.2740726499710034e+02
GL_543 0 NS_543 NS_544 0 5.3740629014256171e-02
GL_544 0 NS_544 NS_543 0 -5.3740629014256171e-02
GS_543_5 0 NS_543 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 545/546
CS_545 NS_545 0 9.9999999999999998e-13
CS_546 NS_546 0 9.9999999999999998e-13
RS_545 NS_545 0 2.3804688106534087e+02
RS_546 NS_546 0 2.3804688106534090e+02
GL_545 0 NS_545 NS_546 0 5.1425903265699464e-02
GL_546 0 NS_546 NS_545 0 -5.1425903265699464e-02
GS_545_5 0 NS_545 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 547/548
CS_547 NS_547 0 9.9999999999999998e-13
CS_548 NS_548 0 9.9999999999999998e-13
RS_547 NS_547 0 1.3728807739915800e+02
RS_548 NS_548 0 1.3728807739915803e+02
GL_547 0 NS_547 NS_548 0 4.8031392820534764e-02
GL_548 0 NS_548 NS_547 0 -4.8031392820534764e-02
GS_547_5 0 NS_547 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 549/550
CS_549 NS_549 0 9.9999999999999998e-13
CS_550 NS_550 0 9.9999999999999998e-13
RS_549 NS_549 0 1.3499477893747948e+02
RS_550 NS_550 0 1.3499477893747945e+02
GL_549 0 NS_549 NS_550 0 4.4453170742682194e-02
GL_550 0 NS_550 NS_549 0 -4.4453170742682194e-02
GS_549_5 0 NS_549 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 551/552
CS_551 NS_551 0 9.9999999999999998e-13
CS_552 NS_552 0 9.9999999999999998e-13
RS_551 NS_551 0 1.4121821834962651e+02
RS_552 NS_552 0 1.4121821834962651e+02
GL_551 0 NS_551 NS_552 0 3.8464469217755697e-02
GL_552 0 NS_552 NS_551 0 -3.8464469217755697e-02
GS_551_5 0 NS_551 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 553/554
CS_553 NS_553 0 9.9999999999999998e-13
CS_554 NS_554 0 9.9999999999999998e-13
RS_553 NS_553 0 1.3946471282741149e+02
RS_554 NS_554 0 1.3946471282741149e+02
GL_553 0 NS_553 NS_554 0 3.5678935079258622e-02
GL_554 0 NS_554 NS_553 0 -3.5678935079258622e-02
GS_553_5 0 NS_553 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 555/556
CS_555 NS_555 0 9.9999999999999998e-13
CS_556 NS_556 0 9.9999999999999998e-13
RS_555 NS_555 0 1.5530211191942624e+02
RS_556 NS_556 0 1.5530211191942627e+02
GL_555 0 NS_555 NS_556 0 2.6209890345437525e-02
GL_556 0 NS_556 NS_555 0 -2.6209890345437525e-02
GS_555_5 0 NS_555 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 557/558
CS_557 NS_557 0 9.9999999999999998e-13
CS_558 NS_558 0 9.9999999999999998e-13
RS_557 NS_557 0 1.4887428879582419e+02
RS_558 NS_558 0 1.4887428879582419e+02
GL_557 0 NS_557 NS_558 0 3.0330575323949095e-02
GL_558 0 NS_558 NS_557 0 -3.0330575323949095e-02
GS_557_5 0 NS_557 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 559/560
CS_559 NS_559 0 9.9999999999999998e-13
CS_560 NS_560 0 9.9999999999999998e-13
RS_559 NS_559 0 1.5087532095170570e+02
RS_560 NS_560 0 1.5087532095170570e+02
GL_559 0 NS_559 NS_560 0 2.0034138441714564e-02
GL_560 0 NS_560 NS_559 0 -2.0034138441714564e-02
GS_559_5 0 NS_559 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 561/562
CS_561 NS_561 0 9.9999999999999998e-13
CS_562 NS_562 0 9.9999999999999998e-13
RS_561 NS_561 0 1.4763793449752018e+02
RS_562 NS_562 0 1.4763793449752018e+02
GL_561 0 NS_561 NS_562 0 1.7017170579416537e-02
GL_562 0 NS_562 NS_561 0 -1.7017170579416537e-02
GS_561_5 0 NS_561 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 563/564
CS_563 NS_563 0 9.9999999999999998e-13
CS_564 NS_564 0 9.9999999999999998e-13
RS_563 NS_563 0 1.6285515224442304e+02
RS_564 NS_564 0 1.6285515224442304e+02
GL_563 0 NS_563 NS_564 0 1.0897027002452746e-02
GL_564 0 NS_564 NS_563 0 -1.0897027002452746e-02
GS_563_5 0 NS_563 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 565/566
CS_565 NS_565 0 9.9999999999999998e-13
CS_566 NS_566 0 9.9999999999999998e-13
RS_565 NS_565 0 1.7239534388116820e+02
RS_566 NS_566 0 1.7239534388116820e+02
GL_565 0 NS_565 NS_566 0 6.1589693699488982e-03
GL_566 0 NS_566 NS_565 0 -6.1589693699488982e-03
GS_565_5 0 NS_565 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 567/568
CS_567 NS_567 0 9.9999999999999998e-13
CS_568 NS_568 0 9.9999999999999998e-13
RS_567 NS_567 0 5.9928710578594173e+03
RS_568 NS_568 0 5.9928710578594173e+03
GL_567 0 NS_567 NS_568 0 1.7541178006601681e-03
GL_568 0 NS_568 NS_567 0 -1.7541178006601681e-03
GS_567_5 0 NS_567 NA_5 0 4.4027142044246531e-01
*
* Complex pair n. 569/570
CS_569 NS_569 0 9.9999999999999998e-13
CS_570 NS_570 0 9.9999999999999998e-13
RS_569 NS_569 0 8.0762087901330699e+02
RS_570 NS_570 0 8.0762087901330688e+02
GL_569 0 NS_569 NS_570 0 1.7295489372816217e-03
GL_570 0 NS_570 NS_569 0 -1.7295489372816217e-03
GS_569_5 0 NS_569 NA_5 0 4.4027142044246531e-01
*
* Real pole n. 571
CS_571 NS_571 0 9.9999999999999998e-13
RS_571 NS_571 0 1.2857601077426406e+01
GS_571_6 0 NS_571 NA_6 0 4.4027142044246531e-01
*
* Real pole n. 572
CS_572 NS_572 0 9.9999999999999998e-13
RS_572 NS_572 0 1.7282831464635029e+02
GS_572_6 0 NS_572 NA_6 0 4.4027142044246531e-01
*
* Real pole n. 573
CS_573 NS_573 0 9.9999999999999998e-13
RS_573 NS_573 0 5.5743135126264733e+03
GS_573_6 0 NS_573 NA_6 0 4.4027142044246531e-01
*
* Real pole n. 574
CS_574 NS_574 0 9.9999999999999998e-13
RS_574 NS_574 0 1.3594126013480764e+03
GS_574_6 0 NS_574 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 575/576
CS_575 NS_575 0 9.9999999999999998e-13
CS_576 NS_576 0 9.9999999999999998e-13
RS_575 NS_575 0 1.7904812183888848e+02
RS_576 NS_576 0 1.7904812183888848e+02
GL_575 0 NS_575 NS_576 0 2.6007898045516648e-01
GL_576 0 NS_576 NS_575 0 -2.6007898045516648e-01
GS_575_6 0 NS_575 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 577/578
CS_577 NS_577 0 9.9999999999999998e-13
CS_578 NS_578 0 9.9999999999999998e-13
RS_577 NS_577 0 1.2615541320340381e+02
RS_578 NS_578 0 1.2615541320340381e+02
GL_577 0 NS_577 NS_578 0 2.5243684762014923e-01
GL_578 0 NS_578 NS_577 0 -2.5243684762014923e-01
GS_577_6 0 NS_577 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 579/580
CS_579 NS_579 0 9.9999999999999998e-13
CS_580 NS_580 0 9.9999999999999998e-13
RS_579 NS_579 0 1.0219948841586964e+02
RS_580 NS_580 0 1.0219948841586965e+02
GL_579 0 NS_579 NS_580 0 2.4690226903121384e-01
GL_580 0 NS_580 NS_579 0 -2.4690226903121384e-01
GS_579_6 0 NS_579 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 581/582
CS_581 NS_581 0 9.9999999999999998e-13
CS_582 NS_582 0 9.9999999999999998e-13
RS_581 NS_581 0 1.1002436853144543e+02
RS_582 NS_582 0 1.1002436853144542e+02
GL_581 0 NS_581 NS_582 0 2.4293768067729948e-01
GL_582 0 NS_582 NS_581 0 -2.4293768067729948e-01
GS_581_6 0 NS_581 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 583/584
CS_583 NS_583 0 9.9999999999999998e-13
CS_584 NS_584 0 9.9999999999999998e-13
RS_583 NS_583 0 1.0553430908077024e+02
RS_584 NS_584 0 1.0553430908077026e+02
GL_583 0 NS_583 NS_584 0 2.3600513224442521e-01
GL_584 0 NS_584 NS_583 0 -2.3600513224442521e-01
GS_583_6 0 NS_583 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 585/586
CS_585 NS_585 0 9.9999999999999998e-13
CS_586 NS_586 0 9.9999999999999998e-13
RS_585 NS_585 0 1.0759915098440327e+02
RS_586 NS_586 0 1.0759915098440327e+02
GL_585 0 NS_585 NS_586 0 2.3090539914362113e-01
GL_586 0 NS_586 NS_585 0 -2.3090539914362113e-01
GS_585_6 0 NS_585 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 587/588
CS_587 NS_587 0 9.9999999999999998e-13
CS_588 NS_588 0 9.9999999999999998e-13
RS_587 NS_587 0 1.3295415758774385e+02
RS_588 NS_588 0 1.3295415758774385e+02
GL_587 0 NS_587 NS_588 0 2.3030066292345727e-01
GL_588 0 NS_588 NS_587 0 -2.3030066292345727e-01
GS_587_6 0 NS_587 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 589/590
CS_589 NS_589 0 9.9999999999999998e-13
CS_590 NS_590 0 9.9999999999999998e-13
RS_589 NS_589 0 1.1432186998941940e+02
RS_590 NS_590 0 1.1432186998941938e+02
GL_589 0 NS_589 NS_590 0 2.2451058023508991e-01
GL_590 0 NS_590 NS_589 0 -2.2451058023508991e-01
GS_589_6 0 NS_589 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 591/592
CS_591 NS_591 0 9.9999999999999998e-13
CS_592 NS_592 0 9.9999999999999998e-13
RS_591 NS_591 0 9.0812703249943667e+01
RS_592 NS_592 0 9.0812703249943652e+01
GL_591 0 NS_591 NS_592 0 2.1702628900531115e-01
GL_592 0 NS_592 NS_591 0 -2.1702628900531115e-01
GS_591_6 0 NS_591 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 593/594
CS_593 NS_593 0 9.9999999999999998e-13
CS_594 NS_594 0 9.9999999999999998e-13
RS_593 NS_593 0 9.5643803662064585e+01
RS_594 NS_594 0 9.5643803662064585e+01
GL_593 0 NS_593 NS_594 0 2.1448200383207913e-01
GL_594 0 NS_594 NS_593 0 -2.1448200383207913e-01
GS_593_6 0 NS_593 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 595/596
CS_595 NS_595 0 9.9999999999999998e-13
CS_596 NS_596 0 9.9999999999999998e-13
RS_595 NS_595 0 1.0631957479149644e+02
RS_596 NS_596 0 1.0631957479149644e+02
GL_595 0 NS_595 NS_596 0 2.0655001587884311e-01
GL_596 0 NS_596 NS_595 0 -2.0655001587884311e-01
GS_595_6 0 NS_595 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 597/598
CS_597 NS_597 0 9.9999999999999998e-13
CS_598 NS_598 0 9.9999999999999998e-13
RS_597 NS_597 0 7.9907264643295406e+01
RS_598 NS_598 0 7.9907264643295420e+01
GL_597 0 NS_597 NS_598 0 2.0133773147328893e-01
GL_598 0 NS_598 NS_597 0 -2.0133773147328893e-01
GS_597_6 0 NS_597 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 599/600
CS_599 NS_599 0 9.9999999999999998e-13
CS_600 NS_600 0 9.9999999999999998e-13
RS_599 NS_599 0 1.0625506887893997e+02
RS_600 NS_600 0 1.0625506887893997e+02
GL_599 0 NS_599 NS_600 0 1.9628877333023340e-01
GL_600 0 NS_600 NS_599 0 -1.9628877333023340e-01
GS_599_6 0 NS_599 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 601/602
CS_601 NS_601 0 9.9999999999999998e-13
CS_602 NS_602 0 9.9999999999999998e-13
RS_601 NS_601 0 9.6115312638592201e+01
RS_602 NS_602 0 9.6115312638592201e+01
GL_601 0 NS_601 NS_602 0 1.8794816712418483e-01
GL_602 0 NS_602 NS_601 0 -1.8794816712418483e-01
GS_601_6 0 NS_601 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 603/604
CS_603 NS_603 0 9.9999999999999998e-13
CS_604 NS_604 0 9.9999999999999998e-13
RS_603 NS_603 0 8.5212696574118169e+01
RS_604 NS_604 0 8.5212696574118169e+01
GL_603 0 NS_603 NS_604 0 1.8572140881490298e-01
GL_604 0 NS_604 NS_603 0 -1.8572140881490298e-01
GS_603_6 0 NS_603 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 605/606
CS_605 NS_605 0 9.9999999999999998e-13
CS_606 NS_606 0 9.9999999999999998e-13
RS_605 NS_605 0 1.0905026103375434e+02
RS_606 NS_606 0 1.0905026103375432e+02
GL_605 0 NS_605 NS_606 0 1.7785621200284463e-01
GL_606 0 NS_606 NS_605 0 -1.7785621200284463e-01
GS_605_6 0 NS_605 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 607/608
CS_607 NS_607 0 9.9999999999999998e-13
CS_608 NS_608 0 9.9999999999999998e-13
RS_607 NS_607 0 8.3024437910787526e+01
RS_608 NS_608 0 8.3024437910787526e+01
GL_607 0 NS_607 NS_608 0 1.7164509875911016e-01
GL_608 0 NS_608 NS_607 0 -1.7164509875911016e-01
GS_607_6 0 NS_607 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 609/610
CS_609 NS_609 0 9.9999999999999998e-13
CS_610 NS_610 0 9.9999999999999998e-13
RS_609 NS_609 0 1.0548793856392000e+02
RS_610 NS_610 0 1.0548793856392000e+02
GL_609 0 NS_609 NS_610 0 1.6750370916002649e-01
GL_610 0 NS_610 NS_609 0 -1.6750370916002649e-01
GS_609_6 0 NS_609 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 611/612
CS_611 NS_611 0 9.9999999999999998e-13
CS_612 NS_612 0 9.9999999999999998e-13
RS_611 NS_611 0 1.0753754351502513e+02
RS_612 NS_612 0 1.0753754351502513e+02
GL_611 0 NS_611 NS_612 0 1.5942172238060490e-01
GL_612 0 NS_612 NS_611 0 -1.5942172238060490e-01
GS_611_6 0 NS_611 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 613/614
CS_613 NS_613 0 9.9999999999999998e-13
CS_614 NS_614 0 9.9999999999999998e-13
RS_613 NS_613 0 8.6961097797504721e+01
RS_614 NS_614 0 8.6961097797504721e+01
GL_613 0 NS_613 NS_614 0 1.5553892891442009e-01
GL_614 0 NS_614 NS_613 0 -1.5553892891442009e-01
GS_613_6 0 NS_613 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 615/616
CS_615 NS_615 0 9.9999999999999998e-13
CS_616 NS_616 0 9.9999999999999998e-13
RS_615 NS_615 0 1.1549771364055694e+02
RS_616 NS_616 0 1.1549771364055692e+02
GL_615 0 NS_615 NS_616 0 1.4899166019107438e-01
GL_616 0 NS_616 NS_615 0 -1.4899166019107438e-01
GS_615_6 0 NS_615 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 617/618
CS_617 NS_617 0 9.9999999999999998e-13
CS_618 NS_618 0 9.9999999999999998e-13
RS_617 NS_617 0 9.7194462506038604e+01
RS_618 NS_618 0 9.7194462506038604e+01
GL_617 0 NS_617 NS_618 0 1.4180400817347408e-01
GL_618 0 NS_618 NS_617 0 -1.4180400817347408e-01
GS_617_6 0 NS_617 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 619/620
CS_619 NS_619 0 9.9999999999999998e-13
CS_620 NS_620 0 9.9999999999999998e-13
RS_619 NS_619 0 1.0682825030924828e+02
RS_620 NS_620 0 1.0682825030924828e+02
GL_619 0 NS_619 NS_620 0 1.3872377519751058e-01
GL_620 0 NS_620 NS_619 0 -1.3872377519751058e-01
GS_619_6 0 NS_619 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 621/622
CS_621 NS_621 0 9.9999999999999998e-13
CS_622 NS_622 0 9.9999999999999998e-13
RS_621 NS_621 0 1.2559585119344567e+02
RS_622 NS_622 0 1.2559585119344568e+02
GL_621 0 NS_621 NS_622 0 1.3097721803321302e-01
GL_622 0 NS_622 NS_621 0 -1.3097721803321302e-01
GS_621_6 0 NS_621 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 623/624
CS_623 NS_623 0 9.9999999999999998e-13
CS_624 NS_624 0 9.9999999999999998e-13
RS_623 NS_623 0 1.0417660462554996e+02
RS_624 NS_624 0 1.0417660462554996e+02
GL_623 0 NS_623 NS_624 0 1.2625832867930367e-01
GL_624 0 NS_624 NS_623 0 -1.2625832867930367e-01
GS_623_6 0 NS_623 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 625/626
CS_625 NS_625 0 9.9999999999999998e-13
CS_626 NS_626 0 9.9999999999999998e-13
RS_625 NS_625 0 1.3317333532177352e+02
RS_626 NS_626 0 1.3317333532177352e+02
GL_625 0 NS_625 NS_626 0 1.2123672752714061e-01
GL_626 0 NS_626 NS_625 0 -1.2123672752714061e-01
GS_625_6 0 NS_625 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 627/628
CS_627 NS_627 0 9.9999999999999998e-13
CS_628 NS_628 0 9.9999999999999998e-13
RS_627 NS_627 0 1.2967831681616519e+02
RS_628 NS_628 0 1.2967831681616519e+02
GL_627 0 NS_627 NS_628 0 1.1651127865768855e-01
GL_628 0 NS_628 NS_627 0 -1.1651127865768855e-01
GS_627_6 0 NS_627 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 629/630
CS_629 NS_629 0 9.9999999999999998e-13
CS_630 NS_630 0 9.9999999999999998e-13
RS_629 NS_629 0 1.2999764374401394e+02
RS_630 NS_630 0 1.2999764374401394e+02
GL_629 0 NS_629 NS_630 0 1.1100247696987056e-01
GL_630 0 NS_630 NS_629 0 -1.1100247696987056e-01
GS_629_6 0 NS_629 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 631/632
CS_631 NS_631 0 9.9999999999999998e-13
CS_632 NS_632 0 9.9999999999999998e-13
RS_631 NS_631 0 1.2458814074636419e+02
RS_632 NS_632 0 1.2458814074636419e+02
GL_631 0 NS_631 NS_632 0 1.0660000212580591e-01
GL_632 0 NS_632 NS_631 0 -1.0660000212580591e-01
GS_631_6 0 NS_631 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 633/634
CS_633 NS_633 0 9.9999999999999998e-13
CS_634 NS_634 0 9.9999999999999998e-13
RS_633 NS_633 0 1.4677191614557748e+02
RS_634 NS_634 0 1.4677191614557748e+02
GL_633 0 NS_633 NS_634 0 1.0224733343325158e-01
GL_634 0 NS_634 NS_633 0 -1.0224733343325158e-01
GS_633_6 0 NS_633 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 635/636
CS_635 NS_635 0 9.9999999999999998e-13
CS_636 NS_636 0 9.9999999999999998e-13
RS_635 NS_635 0 1.3445989223131798e+02
RS_636 NS_636 0 1.3445989223131798e+02
GL_635 0 NS_635 NS_636 0 9.8177836948086503e-02
GL_636 0 NS_636 NS_635 0 -9.8177836948086503e-02
GS_635_6 0 NS_635 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 637/638
CS_637 NS_637 0 9.9999999999999998e-13
CS_638 NS_638 0 9.9999999999999998e-13
RS_637 NS_637 0 1.3187119040723775e+02
RS_638 NS_638 0 1.3187119040723772e+02
GL_637 0 NS_637 NS_638 0 9.2640196004122682e-02
GL_638 0 NS_638 NS_637 0 -9.2640196004122682e-02
GS_637_6 0 NS_637 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 639/640
CS_639 NS_639 0 9.9999999999999998e-13
CS_640 NS_640 0 9.9999999999999998e-13
RS_639 NS_639 0 1.2288401421230557e+02
RS_640 NS_640 0 1.2288401421230557e+02
GL_639 0 NS_639 NS_640 0 8.8704723748248199e-02
GL_640 0 NS_640 NS_639 0 -8.8704723748248199e-02
GS_639_6 0 NS_639 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 641/642
CS_641 NS_641 0 9.9999999999999998e-13
CS_642 NS_642 0 9.9999999999999998e-13
RS_641 NS_641 0 1.4123955654153085e+02
RS_642 NS_642 0 1.4123955654153082e+02
GL_641 0 NS_641 NS_642 0 8.4112474498892476e-02
GL_642 0 NS_642 NS_641 0 -8.4112474498892476e-02
GS_641_6 0 NS_641 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 643/644
CS_643 NS_643 0 9.9999999999999998e-13
CS_644 NS_644 0 9.9999999999999998e-13
RS_643 NS_643 0 1.2539447312269779e+02
RS_644 NS_644 0 1.2539447312269778e+02
GL_643 0 NS_643 NS_644 0 8.0007658848305588e-02
GL_644 0 NS_644 NS_643 0 -8.0007658848305588e-02
GS_643_6 0 NS_643 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 645/646
CS_645 NS_645 0 9.9999999999999998e-13
CS_646 NS_646 0 9.9999999999999998e-13
RS_645 NS_645 0 1.3219601779966965e+02
RS_646 NS_646 0 1.3219601779966968e+02
GL_645 0 NS_645 NS_646 0 7.4373183806052026e-02
GL_646 0 NS_646 NS_645 0 -7.4373183806052026e-02
GS_645_6 0 NS_645 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 647/648
CS_647 NS_647 0 9.9999999999999998e-13
CS_648 NS_648 0 9.9999999999999998e-13
RS_647 NS_647 0 1.1951371640958898e+02
RS_648 NS_648 0 1.1951371640958898e+02
GL_647 0 NS_647 NS_648 0 7.1003860961129844e-02
GL_648 0 NS_648 NS_647 0 -7.1003860961129844e-02
GS_647_6 0 NS_647 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 649/650
CS_649 NS_649 0 9.9999999999999998e-13
CS_650 NS_650 0 9.9999999999999998e-13
RS_649 NS_649 0 1.3491941875045018e+02
RS_650 NS_650 0 1.3491941875045018e+02
GL_649 0 NS_649 NS_650 0 6.5922080709048564e-02
GL_650 0 NS_650 NS_649 0 -6.5922080709048564e-02
GS_649_6 0 NS_649 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 651/652
CS_651 NS_651 0 9.9999999999999998e-13
CS_652 NS_652 0 9.9999999999999998e-13
RS_651 NS_651 0 1.2290405859347165e+02
RS_652 NS_652 0 1.2290405859347166e+02
GL_651 0 NS_651 NS_652 0 6.2340152915784278e-02
GL_652 0 NS_652 NS_651 0 -6.2340152915784278e-02
GS_651_6 0 NS_651 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 653/654
CS_653 NS_653 0 9.9999999999999998e-13
CS_654 NS_654 0 9.9999999999999998e-13
RS_653 NS_653 0 1.3258923845358959e+02
RS_654 NS_654 0 1.3258923845358959e+02
GL_653 0 NS_653 NS_654 0 5.6431081088718790e-02
GL_654 0 NS_654 NS_653 0 -5.6431081088718790e-02
GS_653_6 0 NS_653 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 655/656
CS_655 NS_655 0 9.9999999999999998e-13
CS_656 NS_656 0 9.9999999999999998e-13
RS_655 NS_655 0 1.0026704639246873e+02
RS_656 NS_656 0 1.0026704639246873e+02
GL_655 0 NS_655 NS_656 0 3.5068885856298401e-02
GL_656 0 NS_656 NS_655 0 -3.5068885856298401e-02
GS_655_6 0 NS_655 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 657/658
CS_657 NS_657 0 9.9999999999999998e-13
CS_658 NS_658 0 9.9999999999999998e-13
RS_657 NS_657 0 1.2740726499710033e+02
RS_658 NS_658 0 1.2740726499710034e+02
GL_657 0 NS_657 NS_658 0 5.3740629014256171e-02
GL_658 0 NS_658 NS_657 0 -5.3740629014256171e-02
GS_657_6 0 NS_657 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 659/660
CS_659 NS_659 0 9.9999999999999998e-13
CS_660 NS_660 0 9.9999999999999998e-13
RS_659 NS_659 0 2.3804688106534087e+02
RS_660 NS_660 0 2.3804688106534090e+02
GL_659 0 NS_659 NS_660 0 5.1425903265699464e-02
GL_660 0 NS_660 NS_659 0 -5.1425903265699464e-02
GS_659_6 0 NS_659 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 661/662
CS_661 NS_661 0 9.9999999999999998e-13
CS_662 NS_662 0 9.9999999999999998e-13
RS_661 NS_661 0 1.3728807739915800e+02
RS_662 NS_662 0 1.3728807739915803e+02
GL_661 0 NS_661 NS_662 0 4.8031392820534764e-02
GL_662 0 NS_662 NS_661 0 -4.8031392820534764e-02
GS_661_6 0 NS_661 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 663/664
CS_663 NS_663 0 9.9999999999999998e-13
CS_664 NS_664 0 9.9999999999999998e-13
RS_663 NS_663 0 1.3499477893747948e+02
RS_664 NS_664 0 1.3499477893747945e+02
GL_663 0 NS_663 NS_664 0 4.4453170742682194e-02
GL_664 0 NS_664 NS_663 0 -4.4453170742682194e-02
GS_663_6 0 NS_663 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 665/666
CS_665 NS_665 0 9.9999999999999998e-13
CS_666 NS_666 0 9.9999999999999998e-13
RS_665 NS_665 0 1.4121821834962651e+02
RS_666 NS_666 0 1.4121821834962651e+02
GL_665 0 NS_665 NS_666 0 3.8464469217755697e-02
GL_666 0 NS_666 NS_665 0 -3.8464469217755697e-02
GS_665_6 0 NS_665 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 667/668
CS_667 NS_667 0 9.9999999999999998e-13
CS_668 NS_668 0 9.9999999999999998e-13
RS_667 NS_667 0 1.3946471282741149e+02
RS_668 NS_668 0 1.3946471282741149e+02
GL_667 0 NS_667 NS_668 0 3.5678935079258622e-02
GL_668 0 NS_668 NS_667 0 -3.5678935079258622e-02
GS_667_6 0 NS_667 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 669/670
CS_669 NS_669 0 9.9999999999999998e-13
CS_670 NS_670 0 9.9999999999999998e-13
RS_669 NS_669 0 1.5530211191942624e+02
RS_670 NS_670 0 1.5530211191942627e+02
GL_669 0 NS_669 NS_670 0 2.6209890345437525e-02
GL_670 0 NS_670 NS_669 0 -2.6209890345437525e-02
GS_669_6 0 NS_669 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 671/672
CS_671 NS_671 0 9.9999999999999998e-13
CS_672 NS_672 0 9.9999999999999998e-13
RS_671 NS_671 0 1.4887428879582419e+02
RS_672 NS_672 0 1.4887428879582419e+02
GL_671 0 NS_671 NS_672 0 3.0330575323949095e-02
GL_672 0 NS_672 NS_671 0 -3.0330575323949095e-02
GS_671_6 0 NS_671 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 673/674
CS_673 NS_673 0 9.9999999999999998e-13
CS_674 NS_674 0 9.9999999999999998e-13
RS_673 NS_673 0 1.5087532095170570e+02
RS_674 NS_674 0 1.5087532095170570e+02
GL_673 0 NS_673 NS_674 0 2.0034138441714564e-02
GL_674 0 NS_674 NS_673 0 -2.0034138441714564e-02
GS_673_6 0 NS_673 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 675/676
CS_675 NS_675 0 9.9999999999999998e-13
CS_676 NS_676 0 9.9999999999999998e-13
RS_675 NS_675 0 1.4763793449752018e+02
RS_676 NS_676 0 1.4763793449752018e+02
GL_675 0 NS_675 NS_676 0 1.7017170579416537e-02
GL_676 0 NS_676 NS_675 0 -1.7017170579416537e-02
GS_675_6 0 NS_675 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 677/678
CS_677 NS_677 0 9.9999999999999998e-13
CS_678 NS_678 0 9.9999999999999998e-13
RS_677 NS_677 0 1.6285515224442304e+02
RS_678 NS_678 0 1.6285515224442304e+02
GL_677 0 NS_677 NS_678 0 1.0897027002452746e-02
GL_678 0 NS_678 NS_677 0 -1.0897027002452746e-02
GS_677_6 0 NS_677 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 679/680
CS_679 NS_679 0 9.9999999999999998e-13
CS_680 NS_680 0 9.9999999999999998e-13
RS_679 NS_679 0 1.7239534388116820e+02
RS_680 NS_680 0 1.7239534388116820e+02
GL_679 0 NS_679 NS_680 0 6.1589693699488982e-03
GL_680 0 NS_680 NS_679 0 -6.1589693699488982e-03
GS_679_6 0 NS_679 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 681/682
CS_681 NS_681 0 9.9999999999999998e-13
CS_682 NS_682 0 9.9999999999999998e-13
RS_681 NS_681 0 5.9928710578594173e+03
RS_682 NS_682 0 5.9928710578594173e+03
GL_681 0 NS_681 NS_682 0 1.7541178006601681e-03
GL_682 0 NS_682 NS_681 0 -1.7541178006601681e-03
GS_681_6 0 NS_681 NA_6 0 4.4027142044246531e-01
*
* Complex pair n. 683/684
CS_683 NS_683 0 9.9999999999999998e-13
CS_684 NS_684 0 9.9999999999999998e-13
RS_683 NS_683 0 8.0762087901330699e+02
RS_684 NS_684 0 8.0762087901330688e+02
GL_683 0 NS_683 NS_684 0 1.7295489372816217e-03
GL_684 0 NS_684 NS_683 0 -1.7295489372816217e-03
GS_683_6 0 NS_683 NA_6 0 4.4027142044246531e-01
*
* Real pole n. 685
CS_685 NS_685 0 9.9999999999999998e-13
RS_685 NS_685 0 1.2857601077426406e+01
GS_685_7 0 NS_685 NA_7 0 4.4027142044246531e-01
*
* Real pole n. 686
CS_686 NS_686 0 9.9999999999999998e-13
RS_686 NS_686 0 1.7282831464635029e+02
GS_686_7 0 NS_686 NA_7 0 4.4027142044246531e-01
*
* Real pole n. 687
CS_687 NS_687 0 9.9999999999999998e-13
RS_687 NS_687 0 5.5743135126264733e+03
GS_687_7 0 NS_687 NA_7 0 4.4027142044246531e-01
*
* Real pole n. 688
CS_688 NS_688 0 9.9999999999999998e-13
RS_688 NS_688 0 1.3594126013480764e+03
GS_688_7 0 NS_688 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 689/690
CS_689 NS_689 0 9.9999999999999998e-13
CS_690 NS_690 0 9.9999999999999998e-13
RS_689 NS_689 0 1.7904812183888848e+02
RS_690 NS_690 0 1.7904812183888848e+02
GL_689 0 NS_689 NS_690 0 2.6007898045516648e-01
GL_690 0 NS_690 NS_689 0 -2.6007898045516648e-01
GS_689_7 0 NS_689 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 691/692
CS_691 NS_691 0 9.9999999999999998e-13
CS_692 NS_692 0 9.9999999999999998e-13
RS_691 NS_691 0 1.2615541320340381e+02
RS_692 NS_692 0 1.2615541320340381e+02
GL_691 0 NS_691 NS_692 0 2.5243684762014923e-01
GL_692 0 NS_692 NS_691 0 -2.5243684762014923e-01
GS_691_7 0 NS_691 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 693/694
CS_693 NS_693 0 9.9999999999999998e-13
CS_694 NS_694 0 9.9999999999999998e-13
RS_693 NS_693 0 1.0219948841586964e+02
RS_694 NS_694 0 1.0219948841586965e+02
GL_693 0 NS_693 NS_694 0 2.4690226903121384e-01
GL_694 0 NS_694 NS_693 0 -2.4690226903121384e-01
GS_693_7 0 NS_693 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 695/696
CS_695 NS_695 0 9.9999999999999998e-13
CS_696 NS_696 0 9.9999999999999998e-13
RS_695 NS_695 0 1.1002436853144543e+02
RS_696 NS_696 0 1.1002436853144542e+02
GL_695 0 NS_695 NS_696 0 2.4293768067729948e-01
GL_696 0 NS_696 NS_695 0 -2.4293768067729948e-01
GS_695_7 0 NS_695 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 697/698
CS_697 NS_697 0 9.9999999999999998e-13
CS_698 NS_698 0 9.9999999999999998e-13
RS_697 NS_697 0 1.0553430908077024e+02
RS_698 NS_698 0 1.0553430908077026e+02
GL_697 0 NS_697 NS_698 0 2.3600513224442521e-01
GL_698 0 NS_698 NS_697 0 -2.3600513224442521e-01
GS_697_7 0 NS_697 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 699/700
CS_699 NS_699 0 9.9999999999999998e-13
CS_700 NS_700 0 9.9999999999999998e-13
RS_699 NS_699 0 1.0759915098440327e+02
RS_700 NS_700 0 1.0759915098440327e+02
GL_699 0 NS_699 NS_700 0 2.3090539914362113e-01
GL_700 0 NS_700 NS_699 0 -2.3090539914362113e-01
GS_699_7 0 NS_699 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 701/702
CS_701 NS_701 0 9.9999999999999998e-13
CS_702 NS_702 0 9.9999999999999998e-13
RS_701 NS_701 0 1.3295415758774385e+02
RS_702 NS_702 0 1.3295415758774385e+02
GL_701 0 NS_701 NS_702 0 2.3030066292345727e-01
GL_702 0 NS_702 NS_701 0 -2.3030066292345727e-01
GS_701_7 0 NS_701 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 703/704
CS_703 NS_703 0 9.9999999999999998e-13
CS_704 NS_704 0 9.9999999999999998e-13
RS_703 NS_703 0 1.1432186998941940e+02
RS_704 NS_704 0 1.1432186998941938e+02
GL_703 0 NS_703 NS_704 0 2.2451058023508991e-01
GL_704 0 NS_704 NS_703 0 -2.2451058023508991e-01
GS_703_7 0 NS_703 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 705/706
CS_705 NS_705 0 9.9999999999999998e-13
CS_706 NS_706 0 9.9999999999999998e-13
RS_705 NS_705 0 9.0812703249943667e+01
RS_706 NS_706 0 9.0812703249943652e+01
GL_705 0 NS_705 NS_706 0 2.1702628900531115e-01
GL_706 0 NS_706 NS_705 0 -2.1702628900531115e-01
GS_705_7 0 NS_705 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 707/708
CS_707 NS_707 0 9.9999999999999998e-13
CS_708 NS_708 0 9.9999999999999998e-13
RS_707 NS_707 0 9.5643803662064585e+01
RS_708 NS_708 0 9.5643803662064585e+01
GL_707 0 NS_707 NS_708 0 2.1448200383207913e-01
GL_708 0 NS_708 NS_707 0 -2.1448200383207913e-01
GS_707_7 0 NS_707 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 709/710
CS_709 NS_709 0 9.9999999999999998e-13
CS_710 NS_710 0 9.9999999999999998e-13
RS_709 NS_709 0 1.0631957479149644e+02
RS_710 NS_710 0 1.0631957479149644e+02
GL_709 0 NS_709 NS_710 0 2.0655001587884311e-01
GL_710 0 NS_710 NS_709 0 -2.0655001587884311e-01
GS_709_7 0 NS_709 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 711/712
CS_711 NS_711 0 9.9999999999999998e-13
CS_712 NS_712 0 9.9999999999999998e-13
RS_711 NS_711 0 7.9907264643295406e+01
RS_712 NS_712 0 7.9907264643295420e+01
GL_711 0 NS_711 NS_712 0 2.0133773147328893e-01
GL_712 0 NS_712 NS_711 0 -2.0133773147328893e-01
GS_711_7 0 NS_711 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 713/714
CS_713 NS_713 0 9.9999999999999998e-13
CS_714 NS_714 0 9.9999999999999998e-13
RS_713 NS_713 0 1.0625506887893997e+02
RS_714 NS_714 0 1.0625506887893997e+02
GL_713 0 NS_713 NS_714 0 1.9628877333023340e-01
GL_714 0 NS_714 NS_713 0 -1.9628877333023340e-01
GS_713_7 0 NS_713 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 715/716
CS_715 NS_715 0 9.9999999999999998e-13
CS_716 NS_716 0 9.9999999999999998e-13
RS_715 NS_715 0 9.6115312638592201e+01
RS_716 NS_716 0 9.6115312638592201e+01
GL_715 0 NS_715 NS_716 0 1.8794816712418483e-01
GL_716 0 NS_716 NS_715 0 -1.8794816712418483e-01
GS_715_7 0 NS_715 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 717/718
CS_717 NS_717 0 9.9999999999999998e-13
CS_718 NS_718 0 9.9999999999999998e-13
RS_717 NS_717 0 8.5212696574118169e+01
RS_718 NS_718 0 8.5212696574118169e+01
GL_717 0 NS_717 NS_718 0 1.8572140881490298e-01
GL_718 0 NS_718 NS_717 0 -1.8572140881490298e-01
GS_717_7 0 NS_717 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 719/720
CS_719 NS_719 0 9.9999999999999998e-13
CS_720 NS_720 0 9.9999999999999998e-13
RS_719 NS_719 0 1.0905026103375434e+02
RS_720 NS_720 0 1.0905026103375432e+02
GL_719 0 NS_719 NS_720 0 1.7785621200284463e-01
GL_720 0 NS_720 NS_719 0 -1.7785621200284463e-01
GS_719_7 0 NS_719 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 721/722
CS_721 NS_721 0 9.9999999999999998e-13
CS_722 NS_722 0 9.9999999999999998e-13
RS_721 NS_721 0 8.3024437910787526e+01
RS_722 NS_722 0 8.3024437910787526e+01
GL_721 0 NS_721 NS_722 0 1.7164509875911016e-01
GL_722 0 NS_722 NS_721 0 -1.7164509875911016e-01
GS_721_7 0 NS_721 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 723/724
CS_723 NS_723 0 9.9999999999999998e-13
CS_724 NS_724 0 9.9999999999999998e-13
RS_723 NS_723 0 1.0548793856392000e+02
RS_724 NS_724 0 1.0548793856392000e+02
GL_723 0 NS_723 NS_724 0 1.6750370916002649e-01
GL_724 0 NS_724 NS_723 0 -1.6750370916002649e-01
GS_723_7 0 NS_723 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 725/726
CS_725 NS_725 0 9.9999999999999998e-13
CS_726 NS_726 0 9.9999999999999998e-13
RS_725 NS_725 0 1.0753754351502513e+02
RS_726 NS_726 0 1.0753754351502513e+02
GL_725 0 NS_725 NS_726 0 1.5942172238060490e-01
GL_726 0 NS_726 NS_725 0 -1.5942172238060490e-01
GS_725_7 0 NS_725 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 727/728
CS_727 NS_727 0 9.9999999999999998e-13
CS_728 NS_728 0 9.9999999999999998e-13
RS_727 NS_727 0 8.6961097797504721e+01
RS_728 NS_728 0 8.6961097797504721e+01
GL_727 0 NS_727 NS_728 0 1.5553892891442009e-01
GL_728 0 NS_728 NS_727 0 -1.5553892891442009e-01
GS_727_7 0 NS_727 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 729/730
CS_729 NS_729 0 9.9999999999999998e-13
CS_730 NS_730 0 9.9999999999999998e-13
RS_729 NS_729 0 1.1549771364055694e+02
RS_730 NS_730 0 1.1549771364055692e+02
GL_729 0 NS_729 NS_730 0 1.4899166019107438e-01
GL_730 0 NS_730 NS_729 0 -1.4899166019107438e-01
GS_729_7 0 NS_729 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 731/732
CS_731 NS_731 0 9.9999999999999998e-13
CS_732 NS_732 0 9.9999999999999998e-13
RS_731 NS_731 0 9.7194462506038604e+01
RS_732 NS_732 0 9.7194462506038604e+01
GL_731 0 NS_731 NS_732 0 1.4180400817347408e-01
GL_732 0 NS_732 NS_731 0 -1.4180400817347408e-01
GS_731_7 0 NS_731 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 733/734
CS_733 NS_733 0 9.9999999999999998e-13
CS_734 NS_734 0 9.9999999999999998e-13
RS_733 NS_733 0 1.0682825030924828e+02
RS_734 NS_734 0 1.0682825030924828e+02
GL_733 0 NS_733 NS_734 0 1.3872377519751058e-01
GL_734 0 NS_734 NS_733 0 -1.3872377519751058e-01
GS_733_7 0 NS_733 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 735/736
CS_735 NS_735 0 9.9999999999999998e-13
CS_736 NS_736 0 9.9999999999999998e-13
RS_735 NS_735 0 1.2559585119344567e+02
RS_736 NS_736 0 1.2559585119344568e+02
GL_735 0 NS_735 NS_736 0 1.3097721803321302e-01
GL_736 0 NS_736 NS_735 0 -1.3097721803321302e-01
GS_735_7 0 NS_735 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 737/738
CS_737 NS_737 0 9.9999999999999998e-13
CS_738 NS_738 0 9.9999999999999998e-13
RS_737 NS_737 0 1.0417660462554996e+02
RS_738 NS_738 0 1.0417660462554996e+02
GL_737 0 NS_737 NS_738 0 1.2625832867930367e-01
GL_738 0 NS_738 NS_737 0 -1.2625832867930367e-01
GS_737_7 0 NS_737 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 739/740
CS_739 NS_739 0 9.9999999999999998e-13
CS_740 NS_740 0 9.9999999999999998e-13
RS_739 NS_739 0 1.3317333532177352e+02
RS_740 NS_740 0 1.3317333532177352e+02
GL_739 0 NS_739 NS_740 0 1.2123672752714061e-01
GL_740 0 NS_740 NS_739 0 -1.2123672752714061e-01
GS_739_7 0 NS_739 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 741/742
CS_741 NS_741 0 9.9999999999999998e-13
CS_742 NS_742 0 9.9999999999999998e-13
RS_741 NS_741 0 1.2967831681616519e+02
RS_742 NS_742 0 1.2967831681616519e+02
GL_741 0 NS_741 NS_742 0 1.1651127865768855e-01
GL_742 0 NS_742 NS_741 0 -1.1651127865768855e-01
GS_741_7 0 NS_741 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 743/744
CS_743 NS_743 0 9.9999999999999998e-13
CS_744 NS_744 0 9.9999999999999998e-13
RS_743 NS_743 0 1.2999764374401394e+02
RS_744 NS_744 0 1.2999764374401394e+02
GL_743 0 NS_743 NS_744 0 1.1100247696987056e-01
GL_744 0 NS_744 NS_743 0 -1.1100247696987056e-01
GS_743_7 0 NS_743 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 745/746
CS_745 NS_745 0 9.9999999999999998e-13
CS_746 NS_746 0 9.9999999999999998e-13
RS_745 NS_745 0 1.2458814074636419e+02
RS_746 NS_746 0 1.2458814074636419e+02
GL_745 0 NS_745 NS_746 0 1.0660000212580591e-01
GL_746 0 NS_746 NS_745 0 -1.0660000212580591e-01
GS_745_7 0 NS_745 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 747/748
CS_747 NS_747 0 9.9999999999999998e-13
CS_748 NS_748 0 9.9999999999999998e-13
RS_747 NS_747 0 1.4677191614557748e+02
RS_748 NS_748 0 1.4677191614557748e+02
GL_747 0 NS_747 NS_748 0 1.0224733343325158e-01
GL_748 0 NS_748 NS_747 0 -1.0224733343325158e-01
GS_747_7 0 NS_747 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 749/750
CS_749 NS_749 0 9.9999999999999998e-13
CS_750 NS_750 0 9.9999999999999998e-13
RS_749 NS_749 0 1.3445989223131798e+02
RS_750 NS_750 0 1.3445989223131798e+02
GL_749 0 NS_749 NS_750 0 9.8177836948086503e-02
GL_750 0 NS_750 NS_749 0 -9.8177836948086503e-02
GS_749_7 0 NS_749 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 751/752
CS_751 NS_751 0 9.9999999999999998e-13
CS_752 NS_752 0 9.9999999999999998e-13
RS_751 NS_751 0 1.3187119040723775e+02
RS_752 NS_752 0 1.3187119040723772e+02
GL_751 0 NS_751 NS_752 0 9.2640196004122682e-02
GL_752 0 NS_752 NS_751 0 -9.2640196004122682e-02
GS_751_7 0 NS_751 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 753/754
CS_753 NS_753 0 9.9999999999999998e-13
CS_754 NS_754 0 9.9999999999999998e-13
RS_753 NS_753 0 1.2288401421230557e+02
RS_754 NS_754 0 1.2288401421230557e+02
GL_753 0 NS_753 NS_754 0 8.8704723748248199e-02
GL_754 0 NS_754 NS_753 0 -8.8704723748248199e-02
GS_753_7 0 NS_753 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 755/756
CS_755 NS_755 0 9.9999999999999998e-13
CS_756 NS_756 0 9.9999999999999998e-13
RS_755 NS_755 0 1.4123955654153085e+02
RS_756 NS_756 0 1.4123955654153082e+02
GL_755 0 NS_755 NS_756 0 8.4112474498892476e-02
GL_756 0 NS_756 NS_755 0 -8.4112474498892476e-02
GS_755_7 0 NS_755 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 757/758
CS_757 NS_757 0 9.9999999999999998e-13
CS_758 NS_758 0 9.9999999999999998e-13
RS_757 NS_757 0 1.2539447312269779e+02
RS_758 NS_758 0 1.2539447312269778e+02
GL_757 0 NS_757 NS_758 0 8.0007658848305588e-02
GL_758 0 NS_758 NS_757 0 -8.0007658848305588e-02
GS_757_7 0 NS_757 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 759/760
CS_759 NS_759 0 9.9999999999999998e-13
CS_760 NS_760 0 9.9999999999999998e-13
RS_759 NS_759 0 1.3219601779966965e+02
RS_760 NS_760 0 1.3219601779966968e+02
GL_759 0 NS_759 NS_760 0 7.4373183806052026e-02
GL_760 0 NS_760 NS_759 0 -7.4373183806052026e-02
GS_759_7 0 NS_759 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 761/762
CS_761 NS_761 0 9.9999999999999998e-13
CS_762 NS_762 0 9.9999999999999998e-13
RS_761 NS_761 0 1.1951371640958898e+02
RS_762 NS_762 0 1.1951371640958898e+02
GL_761 0 NS_761 NS_762 0 7.1003860961129844e-02
GL_762 0 NS_762 NS_761 0 -7.1003860961129844e-02
GS_761_7 0 NS_761 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 763/764
CS_763 NS_763 0 9.9999999999999998e-13
CS_764 NS_764 0 9.9999999999999998e-13
RS_763 NS_763 0 1.3491941875045018e+02
RS_764 NS_764 0 1.3491941875045018e+02
GL_763 0 NS_763 NS_764 0 6.5922080709048564e-02
GL_764 0 NS_764 NS_763 0 -6.5922080709048564e-02
GS_763_7 0 NS_763 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 765/766
CS_765 NS_765 0 9.9999999999999998e-13
CS_766 NS_766 0 9.9999999999999998e-13
RS_765 NS_765 0 1.2290405859347165e+02
RS_766 NS_766 0 1.2290405859347166e+02
GL_765 0 NS_765 NS_766 0 6.2340152915784278e-02
GL_766 0 NS_766 NS_765 0 -6.2340152915784278e-02
GS_765_7 0 NS_765 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 767/768
CS_767 NS_767 0 9.9999999999999998e-13
CS_768 NS_768 0 9.9999999999999998e-13
RS_767 NS_767 0 1.3258923845358959e+02
RS_768 NS_768 0 1.3258923845358959e+02
GL_767 0 NS_767 NS_768 0 5.6431081088718790e-02
GL_768 0 NS_768 NS_767 0 -5.6431081088718790e-02
GS_767_7 0 NS_767 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 769/770
CS_769 NS_769 0 9.9999999999999998e-13
CS_770 NS_770 0 9.9999999999999998e-13
RS_769 NS_769 0 1.0026704639246873e+02
RS_770 NS_770 0 1.0026704639246873e+02
GL_769 0 NS_769 NS_770 0 3.5068885856298401e-02
GL_770 0 NS_770 NS_769 0 -3.5068885856298401e-02
GS_769_7 0 NS_769 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 771/772
CS_771 NS_771 0 9.9999999999999998e-13
CS_772 NS_772 0 9.9999999999999998e-13
RS_771 NS_771 0 1.2740726499710033e+02
RS_772 NS_772 0 1.2740726499710034e+02
GL_771 0 NS_771 NS_772 0 5.3740629014256171e-02
GL_772 0 NS_772 NS_771 0 -5.3740629014256171e-02
GS_771_7 0 NS_771 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 773/774
CS_773 NS_773 0 9.9999999999999998e-13
CS_774 NS_774 0 9.9999999999999998e-13
RS_773 NS_773 0 2.3804688106534087e+02
RS_774 NS_774 0 2.3804688106534090e+02
GL_773 0 NS_773 NS_774 0 5.1425903265699464e-02
GL_774 0 NS_774 NS_773 0 -5.1425903265699464e-02
GS_773_7 0 NS_773 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 775/776
CS_775 NS_775 0 9.9999999999999998e-13
CS_776 NS_776 0 9.9999999999999998e-13
RS_775 NS_775 0 1.3728807739915800e+02
RS_776 NS_776 0 1.3728807739915803e+02
GL_775 0 NS_775 NS_776 0 4.8031392820534764e-02
GL_776 0 NS_776 NS_775 0 -4.8031392820534764e-02
GS_775_7 0 NS_775 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 777/778
CS_777 NS_777 0 9.9999999999999998e-13
CS_778 NS_778 0 9.9999999999999998e-13
RS_777 NS_777 0 1.3499477893747948e+02
RS_778 NS_778 0 1.3499477893747945e+02
GL_777 0 NS_777 NS_778 0 4.4453170742682194e-02
GL_778 0 NS_778 NS_777 0 -4.4453170742682194e-02
GS_777_7 0 NS_777 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 779/780
CS_779 NS_779 0 9.9999999999999998e-13
CS_780 NS_780 0 9.9999999999999998e-13
RS_779 NS_779 0 1.4121821834962651e+02
RS_780 NS_780 0 1.4121821834962651e+02
GL_779 0 NS_779 NS_780 0 3.8464469217755697e-02
GL_780 0 NS_780 NS_779 0 -3.8464469217755697e-02
GS_779_7 0 NS_779 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 781/782
CS_781 NS_781 0 9.9999999999999998e-13
CS_782 NS_782 0 9.9999999999999998e-13
RS_781 NS_781 0 1.3946471282741149e+02
RS_782 NS_782 0 1.3946471282741149e+02
GL_781 0 NS_781 NS_782 0 3.5678935079258622e-02
GL_782 0 NS_782 NS_781 0 -3.5678935079258622e-02
GS_781_7 0 NS_781 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 783/784
CS_783 NS_783 0 9.9999999999999998e-13
CS_784 NS_784 0 9.9999999999999998e-13
RS_783 NS_783 0 1.5530211191942624e+02
RS_784 NS_784 0 1.5530211191942627e+02
GL_783 0 NS_783 NS_784 0 2.6209890345437525e-02
GL_784 0 NS_784 NS_783 0 -2.6209890345437525e-02
GS_783_7 0 NS_783 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 785/786
CS_785 NS_785 0 9.9999999999999998e-13
CS_786 NS_786 0 9.9999999999999998e-13
RS_785 NS_785 0 1.4887428879582419e+02
RS_786 NS_786 0 1.4887428879582419e+02
GL_785 0 NS_785 NS_786 0 3.0330575323949095e-02
GL_786 0 NS_786 NS_785 0 -3.0330575323949095e-02
GS_785_7 0 NS_785 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 787/788
CS_787 NS_787 0 9.9999999999999998e-13
CS_788 NS_788 0 9.9999999999999998e-13
RS_787 NS_787 0 1.5087532095170570e+02
RS_788 NS_788 0 1.5087532095170570e+02
GL_787 0 NS_787 NS_788 0 2.0034138441714564e-02
GL_788 0 NS_788 NS_787 0 -2.0034138441714564e-02
GS_787_7 0 NS_787 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 789/790
CS_789 NS_789 0 9.9999999999999998e-13
CS_790 NS_790 0 9.9999999999999998e-13
RS_789 NS_789 0 1.4763793449752018e+02
RS_790 NS_790 0 1.4763793449752018e+02
GL_789 0 NS_789 NS_790 0 1.7017170579416537e-02
GL_790 0 NS_790 NS_789 0 -1.7017170579416537e-02
GS_789_7 0 NS_789 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 791/792
CS_791 NS_791 0 9.9999999999999998e-13
CS_792 NS_792 0 9.9999999999999998e-13
RS_791 NS_791 0 1.6285515224442304e+02
RS_792 NS_792 0 1.6285515224442304e+02
GL_791 0 NS_791 NS_792 0 1.0897027002452746e-02
GL_792 0 NS_792 NS_791 0 -1.0897027002452746e-02
GS_791_7 0 NS_791 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 793/794
CS_793 NS_793 0 9.9999999999999998e-13
CS_794 NS_794 0 9.9999999999999998e-13
RS_793 NS_793 0 1.7239534388116820e+02
RS_794 NS_794 0 1.7239534388116820e+02
GL_793 0 NS_793 NS_794 0 6.1589693699488982e-03
GL_794 0 NS_794 NS_793 0 -6.1589693699488982e-03
GS_793_7 0 NS_793 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 795/796
CS_795 NS_795 0 9.9999999999999998e-13
CS_796 NS_796 0 9.9999999999999998e-13
RS_795 NS_795 0 5.9928710578594173e+03
RS_796 NS_796 0 5.9928710578594173e+03
GL_795 0 NS_795 NS_796 0 1.7541178006601681e-03
GL_796 0 NS_796 NS_795 0 -1.7541178006601681e-03
GS_795_7 0 NS_795 NA_7 0 4.4027142044246531e-01
*
* Complex pair n. 797/798
CS_797 NS_797 0 9.9999999999999998e-13
CS_798 NS_798 0 9.9999999999999998e-13
RS_797 NS_797 0 8.0762087901330699e+02
RS_798 NS_798 0 8.0762087901330688e+02
GL_797 0 NS_797 NS_798 0 1.7295489372816217e-03
GL_798 0 NS_798 NS_797 0 -1.7295489372816217e-03
GS_797_7 0 NS_797 NA_7 0 4.4027142044246531e-01
*
* Real pole n. 799
CS_799 NS_799 0 9.9999999999999998e-13
RS_799 NS_799 0 1.2857601077426406e+01
GS_799_8 0 NS_799 NA_8 0 4.4027142044246531e-01
*
* Real pole n. 800
CS_800 NS_800 0 9.9999999999999998e-13
RS_800 NS_800 0 1.7282831464635029e+02
GS_800_8 0 NS_800 NA_8 0 4.4027142044246531e-01
*
* Real pole n. 801
CS_801 NS_801 0 9.9999999999999998e-13
RS_801 NS_801 0 5.5743135126264733e+03
GS_801_8 0 NS_801 NA_8 0 4.4027142044246531e-01
*
* Real pole n. 802
CS_802 NS_802 0 9.9999999999999998e-13
RS_802 NS_802 0 1.3594126013480764e+03
GS_802_8 0 NS_802 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 803/804
CS_803 NS_803 0 9.9999999999999998e-13
CS_804 NS_804 0 9.9999999999999998e-13
RS_803 NS_803 0 1.7904812183888848e+02
RS_804 NS_804 0 1.7904812183888848e+02
GL_803 0 NS_803 NS_804 0 2.6007898045516648e-01
GL_804 0 NS_804 NS_803 0 -2.6007898045516648e-01
GS_803_8 0 NS_803 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 805/806
CS_805 NS_805 0 9.9999999999999998e-13
CS_806 NS_806 0 9.9999999999999998e-13
RS_805 NS_805 0 1.2615541320340381e+02
RS_806 NS_806 0 1.2615541320340381e+02
GL_805 0 NS_805 NS_806 0 2.5243684762014923e-01
GL_806 0 NS_806 NS_805 0 -2.5243684762014923e-01
GS_805_8 0 NS_805 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 807/808
CS_807 NS_807 0 9.9999999999999998e-13
CS_808 NS_808 0 9.9999999999999998e-13
RS_807 NS_807 0 1.0219948841586964e+02
RS_808 NS_808 0 1.0219948841586965e+02
GL_807 0 NS_807 NS_808 0 2.4690226903121384e-01
GL_808 0 NS_808 NS_807 0 -2.4690226903121384e-01
GS_807_8 0 NS_807 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 809/810
CS_809 NS_809 0 9.9999999999999998e-13
CS_810 NS_810 0 9.9999999999999998e-13
RS_809 NS_809 0 1.1002436853144543e+02
RS_810 NS_810 0 1.1002436853144542e+02
GL_809 0 NS_809 NS_810 0 2.4293768067729948e-01
GL_810 0 NS_810 NS_809 0 -2.4293768067729948e-01
GS_809_8 0 NS_809 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 811/812
CS_811 NS_811 0 9.9999999999999998e-13
CS_812 NS_812 0 9.9999999999999998e-13
RS_811 NS_811 0 1.0553430908077024e+02
RS_812 NS_812 0 1.0553430908077026e+02
GL_811 0 NS_811 NS_812 0 2.3600513224442521e-01
GL_812 0 NS_812 NS_811 0 -2.3600513224442521e-01
GS_811_8 0 NS_811 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 813/814
CS_813 NS_813 0 9.9999999999999998e-13
CS_814 NS_814 0 9.9999999999999998e-13
RS_813 NS_813 0 1.0759915098440327e+02
RS_814 NS_814 0 1.0759915098440327e+02
GL_813 0 NS_813 NS_814 0 2.3090539914362113e-01
GL_814 0 NS_814 NS_813 0 -2.3090539914362113e-01
GS_813_8 0 NS_813 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 815/816
CS_815 NS_815 0 9.9999999999999998e-13
CS_816 NS_816 0 9.9999999999999998e-13
RS_815 NS_815 0 1.3295415758774385e+02
RS_816 NS_816 0 1.3295415758774385e+02
GL_815 0 NS_815 NS_816 0 2.3030066292345727e-01
GL_816 0 NS_816 NS_815 0 -2.3030066292345727e-01
GS_815_8 0 NS_815 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 817/818
CS_817 NS_817 0 9.9999999999999998e-13
CS_818 NS_818 0 9.9999999999999998e-13
RS_817 NS_817 0 1.1432186998941940e+02
RS_818 NS_818 0 1.1432186998941938e+02
GL_817 0 NS_817 NS_818 0 2.2451058023508991e-01
GL_818 0 NS_818 NS_817 0 -2.2451058023508991e-01
GS_817_8 0 NS_817 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 819/820
CS_819 NS_819 0 9.9999999999999998e-13
CS_820 NS_820 0 9.9999999999999998e-13
RS_819 NS_819 0 9.0812703249943667e+01
RS_820 NS_820 0 9.0812703249943652e+01
GL_819 0 NS_819 NS_820 0 2.1702628900531115e-01
GL_820 0 NS_820 NS_819 0 -2.1702628900531115e-01
GS_819_8 0 NS_819 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 821/822
CS_821 NS_821 0 9.9999999999999998e-13
CS_822 NS_822 0 9.9999999999999998e-13
RS_821 NS_821 0 9.5643803662064585e+01
RS_822 NS_822 0 9.5643803662064585e+01
GL_821 0 NS_821 NS_822 0 2.1448200383207913e-01
GL_822 0 NS_822 NS_821 0 -2.1448200383207913e-01
GS_821_8 0 NS_821 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 823/824
CS_823 NS_823 0 9.9999999999999998e-13
CS_824 NS_824 0 9.9999999999999998e-13
RS_823 NS_823 0 1.0631957479149644e+02
RS_824 NS_824 0 1.0631957479149644e+02
GL_823 0 NS_823 NS_824 0 2.0655001587884311e-01
GL_824 0 NS_824 NS_823 0 -2.0655001587884311e-01
GS_823_8 0 NS_823 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 825/826
CS_825 NS_825 0 9.9999999999999998e-13
CS_826 NS_826 0 9.9999999999999998e-13
RS_825 NS_825 0 7.9907264643295406e+01
RS_826 NS_826 0 7.9907264643295420e+01
GL_825 0 NS_825 NS_826 0 2.0133773147328893e-01
GL_826 0 NS_826 NS_825 0 -2.0133773147328893e-01
GS_825_8 0 NS_825 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 827/828
CS_827 NS_827 0 9.9999999999999998e-13
CS_828 NS_828 0 9.9999999999999998e-13
RS_827 NS_827 0 1.0625506887893997e+02
RS_828 NS_828 0 1.0625506887893997e+02
GL_827 0 NS_827 NS_828 0 1.9628877333023340e-01
GL_828 0 NS_828 NS_827 0 -1.9628877333023340e-01
GS_827_8 0 NS_827 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 829/830
CS_829 NS_829 0 9.9999999999999998e-13
CS_830 NS_830 0 9.9999999999999998e-13
RS_829 NS_829 0 9.6115312638592201e+01
RS_830 NS_830 0 9.6115312638592201e+01
GL_829 0 NS_829 NS_830 0 1.8794816712418483e-01
GL_830 0 NS_830 NS_829 0 -1.8794816712418483e-01
GS_829_8 0 NS_829 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 831/832
CS_831 NS_831 0 9.9999999999999998e-13
CS_832 NS_832 0 9.9999999999999998e-13
RS_831 NS_831 0 8.5212696574118169e+01
RS_832 NS_832 0 8.5212696574118169e+01
GL_831 0 NS_831 NS_832 0 1.8572140881490298e-01
GL_832 0 NS_832 NS_831 0 -1.8572140881490298e-01
GS_831_8 0 NS_831 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 833/834
CS_833 NS_833 0 9.9999999999999998e-13
CS_834 NS_834 0 9.9999999999999998e-13
RS_833 NS_833 0 1.0905026103375434e+02
RS_834 NS_834 0 1.0905026103375432e+02
GL_833 0 NS_833 NS_834 0 1.7785621200284463e-01
GL_834 0 NS_834 NS_833 0 -1.7785621200284463e-01
GS_833_8 0 NS_833 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 835/836
CS_835 NS_835 0 9.9999999999999998e-13
CS_836 NS_836 0 9.9999999999999998e-13
RS_835 NS_835 0 8.3024437910787526e+01
RS_836 NS_836 0 8.3024437910787526e+01
GL_835 0 NS_835 NS_836 0 1.7164509875911016e-01
GL_836 0 NS_836 NS_835 0 -1.7164509875911016e-01
GS_835_8 0 NS_835 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 837/838
CS_837 NS_837 0 9.9999999999999998e-13
CS_838 NS_838 0 9.9999999999999998e-13
RS_837 NS_837 0 1.0548793856392000e+02
RS_838 NS_838 0 1.0548793856392000e+02
GL_837 0 NS_837 NS_838 0 1.6750370916002649e-01
GL_838 0 NS_838 NS_837 0 -1.6750370916002649e-01
GS_837_8 0 NS_837 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 839/840
CS_839 NS_839 0 9.9999999999999998e-13
CS_840 NS_840 0 9.9999999999999998e-13
RS_839 NS_839 0 1.0753754351502513e+02
RS_840 NS_840 0 1.0753754351502513e+02
GL_839 0 NS_839 NS_840 0 1.5942172238060490e-01
GL_840 0 NS_840 NS_839 0 -1.5942172238060490e-01
GS_839_8 0 NS_839 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 841/842
CS_841 NS_841 0 9.9999999999999998e-13
CS_842 NS_842 0 9.9999999999999998e-13
RS_841 NS_841 0 8.6961097797504721e+01
RS_842 NS_842 0 8.6961097797504721e+01
GL_841 0 NS_841 NS_842 0 1.5553892891442009e-01
GL_842 0 NS_842 NS_841 0 -1.5553892891442009e-01
GS_841_8 0 NS_841 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 843/844
CS_843 NS_843 0 9.9999999999999998e-13
CS_844 NS_844 0 9.9999999999999998e-13
RS_843 NS_843 0 1.1549771364055694e+02
RS_844 NS_844 0 1.1549771364055692e+02
GL_843 0 NS_843 NS_844 0 1.4899166019107438e-01
GL_844 0 NS_844 NS_843 0 -1.4899166019107438e-01
GS_843_8 0 NS_843 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 845/846
CS_845 NS_845 0 9.9999999999999998e-13
CS_846 NS_846 0 9.9999999999999998e-13
RS_845 NS_845 0 9.7194462506038604e+01
RS_846 NS_846 0 9.7194462506038604e+01
GL_845 0 NS_845 NS_846 0 1.4180400817347408e-01
GL_846 0 NS_846 NS_845 0 -1.4180400817347408e-01
GS_845_8 0 NS_845 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 847/848
CS_847 NS_847 0 9.9999999999999998e-13
CS_848 NS_848 0 9.9999999999999998e-13
RS_847 NS_847 0 1.0682825030924828e+02
RS_848 NS_848 0 1.0682825030924828e+02
GL_847 0 NS_847 NS_848 0 1.3872377519751058e-01
GL_848 0 NS_848 NS_847 0 -1.3872377519751058e-01
GS_847_8 0 NS_847 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 849/850
CS_849 NS_849 0 9.9999999999999998e-13
CS_850 NS_850 0 9.9999999999999998e-13
RS_849 NS_849 0 1.2559585119344567e+02
RS_850 NS_850 0 1.2559585119344568e+02
GL_849 0 NS_849 NS_850 0 1.3097721803321302e-01
GL_850 0 NS_850 NS_849 0 -1.3097721803321302e-01
GS_849_8 0 NS_849 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 851/852
CS_851 NS_851 0 9.9999999999999998e-13
CS_852 NS_852 0 9.9999999999999998e-13
RS_851 NS_851 0 1.0417660462554996e+02
RS_852 NS_852 0 1.0417660462554996e+02
GL_851 0 NS_851 NS_852 0 1.2625832867930367e-01
GL_852 0 NS_852 NS_851 0 -1.2625832867930367e-01
GS_851_8 0 NS_851 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 853/854
CS_853 NS_853 0 9.9999999999999998e-13
CS_854 NS_854 0 9.9999999999999998e-13
RS_853 NS_853 0 1.3317333532177352e+02
RS_854 NS_854 0 1.3317333532177352e+02
GL_853 0 NS_853 NS_854 0 1.2123672752714061e-01
GL_854 0 NS_854 NS_853 0 -1.2123672752714061e-01
GS_853_8 0 NS_853 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 855/856
CS_855 NS_855 0 9.9999999999999998e-13
CS_856 NS_856 0 9.9999999999999998e-13
RS_855 NS_855 0 1.2967831681616519e+02
RS_856 NS_856 0 1.2967831681616519e+02
GL_855 0 NS_855 NS_856 0 1.1651127865768855e-01
GL_856 0 NS_856 NS_855 0 -1.1651127865768855e-01
GS_855_8 0 NS_855 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 857/858
CS_857 NS_857 0 9.9999999999999998e-13
CS_858 NS_858 0 9.9999999999999998e-13
RS_857 NS_857 0 1.2999764374401394e+02
RS_858 NS_858 0 1.2999764374401394e+02
GL_857 0 NS_857 NS_858 0 1.1100247696987056e-01
GL_858 0 NS_858 NS_857 0 -1.1100247696987056e-01
GS_857_8 0 NS_857 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 859/860
CS_859 NS_859 0 9.9999999999999998e-13
CS_860 NS_860 0 9.9999999999999998e-13
RS_859 NS_859 0 1.2458814074636419e+02
RS_860 NS_860 0 1.2458814074636419e+02
GL_859 0 NS_859 NS_860 0 1.0660000212580591e-01
GL_860 0 NS_860 NS_859 0 -1.0660000212580591e-01
GS_859_8 0 NS_859 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 861/862
CS_861 NS_861 0 9.9999999999999998e-13
CS_862 NS_862 0 9.9999999999999998e-13
RS_861 NS_861 0 1.4677191614557748e+02
RS_862 NS_862 0 1.4677191614557748e+02
GL_861 0 NS_861 NS_862 0 1.0224733343325158e-01
GL_862 0 NS_862 NS_861 0 -1.0224733343325158e-01
GS_861_8 0 NS_861 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 863/864
CS_863 NS_863 0 9.9999999999999998e-13
CS_864 NS_864 0 9.9999999999999998e-13
RS_863 NS_863 0 1.3445989223131798e+02
RS_864 NS_864 0 1.3445989223131798e+02
GL_863 0 NS_863 NS_864 0 9.8177836948086503e-02
GL_864 0 NS_864 NS_863 0 -9.8177836948086503e-02
GS_863_8 0 NS_863 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 865/866
CS_865 NS_865 0 9.9999999999999998e-13
CS_866 NS_866 0 9.9999999999999998e-13
RS_865 NS_865 0 1.3187119040723775e+02
RS_866 NS_866 0 1.3187119040723772e+02
GL_865 0 NS_865 NS_866 0 9.2640196004122682e-02
GL_866 0 NS_866 NS_865 0 -9.2640196004122682e-02
GS_865_8 0 NS_865 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 867/868
CS_867 NS_867 0 9.9999999999999998e-13
CS_868 NS_868 0 9.9999999999999998e-13
RS_867 NS_867 0 1.2288401421230557e+02
RS_868 NS_868 0 1.2288401421230557e+02
GL_867 0 NS_867 NS_868 0 8.8704723748248199e-02
GL_868 0 NS_868 NS_867 0 -8.8704723748248199e-02
GS_867_8 0 NS_867 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 869/870
CS_869 NS_869 0 9.9999999999999998e-13
CS_870 NS_870 0 9.9999999999999998e-13
RS_869 NS_869 0 1.4123955654153085e+02
RS_870 NS_870 0 1.4123955654153082e+02
GL_869 0 NS_869 NS_870 0 8.4112474498892476e-02
GL_870 0 NS_870 NS_869 0 -8.4112474498892476e-02
GS_869_8 0 NS_869 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 871/872
CS_871 NS_871 0 9.9999999999999998e-13
CS_872 NS_872 0 9.9999999999999998e-13
RS_871 NS_871 0 1.2539447312269779e+02
RS_872 NS_872 0 1.2539447312269778e+02
GL_871 0 NS_871 NS_872 0 8.0007658848305588e-02
GL_872 0 NS_872 NS_871 0 -8.0007658848305588e-02
GS_871_8 0 NS_871 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 873/874
CS_873 NS_873 0 9.9999999999999998e-13
CS_874 NS_874 0 9.9999999999999998e-13
RS_873 NS_873 0 1.3219601779966965e+02
RS_874 NS_874 0 1.3219601779966968e+02
GL_873 0 NS_873 NS_874 0 7.4373183806052026e-02
GL_874 0 NS_874 NS_873 0 -7.4373183806052026e-02
GS_873_8 0 NS_873 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 875/876
CS_875 NS_875 0 9.9999999999999998e-13
CS_876 NS_876 0 9.9999999999999998e-13
RS_875 NS_875 0 1.1951371640958898e+02
RS_876 NS_876 0 1.1951371640958898e+02
GL_875 0 NS_875 NS_876 0 7.1003860961129844e-02
GL_876 0 NS_876 NS_875 0 -7.1003860961129844e-02
GS_875_8 0 NS_875 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 877/878
CS_877 NS_877 0 9.9999999999999998e-13
CS_878 NS_878 0 9.9999999999999998e-13
RS_877 NS_877 0 1.3491941875045018e+02
RS_878 NS_878 0 1.3491941875045018e+02
GL_877 0 NS_877 NS_878 0 6.5922080709048564e-02
GL_878 0 NS_878 NS_877 0 -6.5922080709048564e-02
GS_877_8 0 NS_877 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 879/880
CS_879 NS_879 0 9.9999999999999998e-13
CS_880 NS_880 0 9.9999999999999998e-13
RS_879 NS_879 0 1.2290405859347165e+02
RS_880 NS_880 0 1.2290405859347166e+02
GL_879 0 NS_879 NS_880 0 6.2340152915784278e-02
GL_880 0 NS_880 NS_879 0 -6.2340152915784278e-02
GS_879_8 0 NS_879 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 881/882
CS_881 NS_881 0 9.9999999999999998e-13
CS_882 NS_882 0 9.9999999999999998e-13
RS_881 NS_881 0 1.3258923845358959e+02
RS_882 NS_882 0 1.3258923845358959e+02
GL_881 0 NS_881 NS_882 0 5.6431081088718790e-02
GL_882 0 NS_882 NS_881 0 -5.6431081088718790e-02
GS_881_8 0 NS_881 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 883/884
CS_883 NS_883 0 9.9999999999999998e-13
CS_884 NS_884 0 9.9999999999999998e-13
RS_883 NS_883 0 1.0026704639246873e+02
RS_884 NS_884 0 1.0026704639246873e+02
GL_883 0 NS_883 NS_884 0 3.5068885856298401e-02
GL_884 0 NS_884 NS_883 0 -3.5068885856298401e-02
GS_883_8 0 NS_883 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 885/886
CS_885 NS_885 0 9.9999999999999998e-13
CS_886 NS_886 0 9.9999999999999998e-13
RS_885 NS_885 0 1.2740726499710033e+02
RS_886 NS_886 0 1.2740726499710034e+02
GL_885 0 NS_885 NS_886 0 5.3740629014256171e-02
GL_886 0 NS_886 NS_885 0 -5.3740629014256171e-02
GS_885_8 0 NS_885 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 887/888
CS_887 NS_887 0 9.9999999999999998e-13
CS_888 NS_888 0 9.9999999999999998e-13
RS_887 NS_887 0 2.3804688106534087e+02
RS_888 NS_888 0 2.3804688106534090e+02
GL_887 0 NS_887 NS_888 0 5.1425903265699464e-02
GL_888 0 NS_888 NS_887 0 -5.1425903265699464e-02
GS_887_8 0 NS_887 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 889/890
CS_889 NS_889 0 9.9999999999999998e-13
CS_890 NS_890 0 9.9999999999999998e-13
RS_889 NS_889 0 1.3728807739915800e+02
RS_890 NS_890 0 1.3728807739915803e+02
GL_889 0 NS_889 NS_890 0 4.8031392820534764e-02
GL_890 0 NS_890 NS_889 0 -4.8031392820534764e-02
GS_889_8 0 NS_889 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 891/892
CS_891 NS_891 0 9.9999999999999998e-13
CS_892 NS_892 0 9.9999999999999998e-13
RS_891 NS_891 0 1.3499477893747948e+02
RS_892 NS_892 0 1.3499477893747945e+02
GL_891 0 NS_891 NS_892 0 4.4453170742682194e-02
GL_892 0 NS_892 NS_891 0 -4.4453170742682194e-02
GS_891_8 0 NS_891 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 893/894
CS_893 NS_893 0 9.9999999999999998e-13
CS_894 NS_894 0 9.9999999999999998e-13
RS_893 NS_893 0 1.4121821834962651e+02
RS_894 NS_894 0 1.4121821834962651e+02
GL_893 0 NS_893 NS_894 0 3.8464469217755697e-02
GL_894 0 NS_894 NS_893 0 -3.8464469217755697e-02
GS_893_8 0 NS_893 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 895/896
CS_895 NS_895 0 9.9999999999999998e-13
CS_896 NS_896 0 9.9999999999999998e-13
RS_895 NS_895 0 1.3946471282741149e+02
RS_896 NS_896 0 1.3946471282741149e+02
GL_895 0 NS_895 NS_896 0 3.5678935079258622e-02
GL_896 0 NS_896 NS_895 0 -3.5678935079258622e-02
GS_895_8 0 NS_895 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 897/898
CS_897 NS_897 0 9.9999999999999998e-13
CS_898 NS_898 0 9.9999999999999998e-13
RS_897 NS_897 0 1.5530211191942624e+02
RS_898 NS_898 0 1.5530211191942627e+02
GL_897 0 NS_897 NS_898 0 2.6209890345437525e-02
GL_898 0 NS_898 NS_897 0 -2.6209890345437525e-02
GS_897_8 0 NS_897 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 899/900
CS_899 NS_899 0 9.9999999999999998e-13
CS_900 NS_900 0 9.9999999999999998e-13
RS_899 NS_899 0 1.4887428879582419e+02
RS_900 NS_900 0 1.4887428879582419e+02
GL_899 0 NS_899 NS_900 0 3.0330575323949095e-02
GL_900 0 NS_900 NS_899 0 -3.0330575323949095e-02
GS_899_8 0 NS_899 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 901/902
CS_901 NS_901 0 9.9999999999999998e-13
CS_902 NS_902 0 9.9999999999999998e-13
RS_901 NS_901 0 1.5087532095170570e+02
RS_902 NS_902 0 1.5087532095170570e+02
GL_901 0 NS_901 NS_902 0 2.0034138441714564e-02
GL_902 0 NS_902 NS_901 0 -2.0034138441714564e-02
GS_901_8 0 NS_901 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 903/904
CS_903 NS_903 0 9.9999999999999998e-13
CS_904 NS_904 0 9.9999999999999998e-13
RS_903 NS_903 0 1.4763793449752018e+02
RS_904 NS_904 0 1.4763793449752018e+02
GL_903 0 NS_903 NS_904 0 1.7017170579416537e-02
GL_904 0 NS_904 NS_903 0 -1.7017170579416537e-02
GS_903_8 0 NS_903 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 905/906
CS_905 NS_905 0 9.9999999999999998e-13
CS_906 NS_906 0 9.9999999999999998e-13
RS_905 NS_905 0 1.6285515224442304e+02
RS_906 NS_906 0 1.6285515224442304e+02
GL_905 0 NS_905 NS_906 0 1.0897027002452746e-02
GL_906 0 NS_906 NS_905 0 -1.0897027002452746e-02
GS_905_8 0 NS_905 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 907/908
CS_907 NS_907 0 9.9999999999999998e-13
CS_908 NS_908 0 9.9999999999999998e-13
RS_907 NS_907 0 1.7239534388116820e+02
RS_908 NS_908 0 1.7239534388116820e+02
GL_907 0 NS_907 NS_908 0 6.1589693699488982e-03
GL_908 0 NS_908 NS_907 0 -6.1589693699488982e-03
GS_907_8 0 NS_907 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 909/910
CS_909 NS_909 0 9.9999999999999998e-13
CS_910 NS_910 0 9.9999999999999998e-13
RS_909 NS_909 0 5.9928710578594173e+03
RS_910 NS_910 0 5.9928710578594173e+03
GL_909 0 NS_909 NS_910 0 1.7541178006601681e-03
GL_910 0 NS_910 NS_909 0 -1.7541178006601681e-03
GS_909_8 0 NS_909 NA_8 0 4.4027142044246531e-01
*
* Complex pair n. 911/912
CS_911 NS_911 0 9.9999999999999998e-13
CS_912 NS_912 0 9.9999999999999998e-13
RS_911 NS_911 0 8.0762087901330699e+02
RS_912 NS_912 0 8.0762087901330688e+02
GL_911 0 NS_911 NS_912 0 1.7295489372816217e-03
GL_912 0 NS_912 NS_911 0 -1.7295489372816217e-03
GS_911_8 0 NS_911 NA_8 0 4.4027142044246531e-01
*
* Real pole n. 913
CS_913 NS_913 0 9.9999999999999998e-13
RS_913 NS_913 0 1.2857601077426406e+01
GS_913_9 0 NS_913 NA_9 0 4.4027142044246531e-01
*
* Real pole n. 914
CS_914 NS_914 0 9.9999999999999998e-13
RS_914 NS_914 0 1.7282831464635029e+02
GS_914_9 0 NS_914 NA_9 0 4.4027142044246531e-01
*
* Real pole n. 915
CS_915 NS_915 0 9.9999999999999998e-13
RS_915 NS_915 0 5.5743135126264733e+03
GS_915_9 0 NS_915 NA_9 0 4.4027142044246531e-01
*
* Real pole n. 916
CS_916 NS_916 0 9.9999999999999998e-13
RS_916 NS_916 0 1.3594126013480764e+03
GS_916_9 0 NS_916 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 917/918
CS_917 NS_917 0 9.9999999999999998e-13
CS_918 NS_918 0 9.9999999999999998e-13
RS_917 NS_917 0 1.7904812183888848e+02
RS_918 NS_918 0 1.7904812183888848e+02
GL_917 0 NS_917 NS_918 0 2.6007898045516648e-01
GL_918 0 NS_918 NS_917 0 -2.6007898045516648e-01
GS_917_9 0 NS_917 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 919/920
CS_919 NS_919 0 9.9999999999999998e-13
CS_920 NS_920 0 9.9999999999999998e-13
RS_919 NS_919 0 1.2615541320340381e+02
RS_920 NS_920 0 1.2615541320340381e+02
GL_919 0 NS_919 NS_920 0 2.5243684762014923e-01
GL_920 0 NS_920 NS_919 0 -2.5243684762014923e-01
GS_919_9 0 NS_919 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 921/922
CS_921 NS_921 0 9.9999999999999998e-13
CS_922 NS_922 0 9.9999999999999998e-13
RS_921 NS_921 0 1.0219948841586964e+02
RS_922 NS_922 0 1.0219948841586965e+02
GL_921 0 NS_921 NS_922 0 2.4690226903121384e-01
GL_922 0 NS_922 NS_921 0 -2.4690226903121384e-01
GS_921_9 0 NS_921 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 923/924
CS_923 NS_923 0 9.9999999999999998e-13
CS_924 NS_924 0 9.9999999999999998e-13
RS_923 NS_923 0 1.1002436853144543e+02
RS_924 NS_924 0 1.1002436853144542e+02
GL_923 0 NS_923 NS_924 0 2.4293768067729948e-01
GL_924 0 NS_924 NS_923 0 -2.4293768067729948e-01
GS_923_9 0 NS_923 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 925/926
CS_925 NS_925 0 9.9999999999999998e-13
CS_926 NS_926 0 9.9999999999999998e-13
RS_925 NS_925 0 1.0553430908077024e+02
RS_926 NS_926 0 1.0553430908077026e+02
GL_925 0 NS_925 NS_926 0 2.3600513224442521e-01
GL_926 0 NS_926 NS_925 0 -2.3600513224442521e-01
GS_925_9 0 NS_925 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 927/928
CS_927 NS_927 0 9.9999999999999998e-13
CS_928 NS_928 0 9.9999999999999998e-13
RS_927 NS_927 0 1.0759915098440327e+02
RS_928 NS_928 0 1.0759915098440327e+02
GL_927 0 NS_927 NS_928 0 2.3090539914362113e-01
GL_928 0 NS_928 NS_927 0 -2.3090539914362113e-01
GS_927_9 0 NS_927 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 929/930
CS_929 NS_929 0 9.9999999999999998e-13
CS_930 NS_930 0 9.9999999999999998e-13
RS_929 NS_929 0 1.3295415758774385e+02
RS_930 NS_930 0 1.3295415758774385e+02
GL_929 0 NS_929 NS_930 0 2.3030066292345727e-01
GL_930 0 NS_930 NS_929 0 -2.3030066292345727e-01
GS_929_9 0 NS_929 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 931/932
CS_931 NS_931 0 9.9999999999999998e-13
CS_932 NS_932 0 9.9999999999999998e-13
RS_931 NS_931 0 1.1432186998941940e+02
RS_932 NS_932 0 1.1432186998941938e+02
GL_931 0 NS_931 NS_932 0 2.2451058023508991e-01
GL_932 0 NS_932 NS_931 0 -2.2451058023508991e-01
GS_931_9 0 NS_931 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 933/934
CS_933 NS_933 0 9.9999999999999998e-13
CS_934 NS_934 0 9.9999999999999998e-13
RS_933 NS_933 0 9.0812703249943667e+01
RS_934 NS_934 0 9.0812703249943652e+01
GL_933 0 NS_933 NS_934 0 2.1702628900531115e-01
GL_934 0 NS_934 NS_933 0 -2.1702628900531115e-01
GS_933_9 0 NS_933 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 935/936
CS_935 NS_935 0 9.9999999999999998e-13
CS_936 NS_936 0 9.9999999999999998e-13
RS_935 NS_935 0 9.5643803662064585e+01
RS_936 NS_936 0 9.5643803662064585e+01
GL_935 0 NS_935 NS_936 0 2.1448200383207913e-01
GL_936 0 NS_936 NS_935 0 -2.1448200383207913e-01
GS_935_9 0 NS_935 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 937/938
CS_937 NS_937 0 9.9999999999999998e-13
CS_938 NS_938 0 9.9999999999999998e-13
RS_937 NS_937 0 1.0631957479149644e+02
RS_938 NS_938 0 1.0631957479149644e+02
GL_937 0 NS_937 NS_938 0 2.0655001587884311e-01
GL_938 0 NS_938 NS_937 0 -2.0655001587884311e-01
GS_937_9 0 NS_937 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 939/940
CS_939 NS_939 0 9.9999999999999998e-13
CS_940 NS_940 0 9.9999999999999998e-13
RS_939 NS_939 0 7.9907264643295406e+01
RS_940 NS_940 0 7.9907264643295420e+01
GL_939 0 NS_939 NS_940 0 2.0133773147328893e-01
GL_940 0 NS_940 NS_939 0 -2.0133773147328893e-01
GS_939_9 0 NS_939 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 941/942
CS_941 NS_941 0 9.9999999999999998e-13
CS_942 NS_942 0 9.9999999999999998e-13
RS_941 NS_941 0 1.0625506887893997e+02
RS_942 NS_942 0 1.0625506887893997e+02
GL_941 0 NS_941 NS_942 0 1.9628877333023340e-01
GL_942 0 NS_942 NS_941 0 -1.9628877333023340e-01
GS_941_9 0 NS_941 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 943/944
CS_943 NS_943 0 9.9999999999999998e-13
CS_944 NS_944 0 9.9999999999999998e-13
RS_943 NS_943 0 9.6115312638592201e+01
RS_944 NS_944 0 9.6115312638592201e+01
GL_943 0 NS_943 NS_944 0 1.8794816712418483e-01
GL_944 0 NS_944 NS_943 0 -1.8794816712418483e-01
GS_943_9 0 NS_943 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 945/946
CS_945 NS_945 0 9.9999999999999998e-13
CS_946 NS_946 0 9.9999999999999998e-13
RS_945 NS_945 0 8.5212696574118169e+01
RS_946 NS_946 0 8.5212696574118169e+01
GL_945 0 NS_945 NS_946 0 1.8572140881490298e-01
GL_946 0 NS_946 NS_945 0 -1.8572140881490298e-01
GS_945_9 0 NS_945 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 947/948
CS_947 NS_947 0 9.9999999999999998e-13
CS_948 NS_948 0 9.9999999999999998e-13
RS_947 NS_947 0 1.0905026103375434e+02
RS_948 NS_948 0 1.0905026103375432e+02
GL_947 0 NS_947 NS_948 0 1.7785621200284463e-01
GL_948 0 NS_948 NS_947 0 -1.7785621200284463e-01
GS_947_9 0 NS_947 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 949/950
CS_949 NS_949 0 9.9999999999999998e-13
CS_950 NS_950 0 9.9999999999999998e-13
RS_949 NS_949 0 8.3024437910787526e+01
RS_950 NS_950 0 8.3024437910787526e+01
GL_949 0 NS_949 NS_950 0 1.7164509875911016e-01
GL_950 0 NS_950 NS_949 0 -1.7164509875911016e-01
GS_949_9 0 NS_949 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 951/952
CS_951 NS_951 0 9.9999999999999998e-13
CS_952 NS_952 0 9.9999999999999998e-13
RS_951 NS_951 0 1.0548793856392000e+02
RS_952 NS_952 0 1.0548793856392000e+02
GL_951 0 NS_951 NS_952 0 1.6750370916002649e-01
GL_952 0 NS_952 NS_951 0 -1.6750370916002649e-01
GS_951_9 0 NS_951 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 953/954
CS_953 NS_953 0 9.9999999999999998e-13
CS_954 NS_954 0 9.9999999999999998e-13
RS_953 NS_953 0 1.0753754351502513e+02
RS_954 NS_954 0 1.0753754351502513e+02
GL_953 0 NS_953 NS_954 0 1.5942172238060490e-01
GL_954 0 NS_954 NS_953 0 -1.5942172238060490e-01
GS_953_9 0 NS_953 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 955/956
CS_955 NS_955 0 9.9999999999999998e-13
CS_956 NS_956 0 9.9999999999999998e-13
RS_955 NS_955 0 8.6961097797504721e+01
RS_956 NS_956 0 8.6961097797504721e+01
GL_955 0 NS_955 NS_956 0 1.5553892891442009e-01
GL_956 0 NS_956 NS_955 0 -1.5553892891442009e-01
GS_955_9 0 NS_955 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 957/958
CS_957 NS_957 0 9.9999999999999998e-13
CS_958 NS_958 0 9.9999999999999998e-13
RS_957 NS_957 0 1.1549771364055694e+02
RS_958 NS_958 0 1.1549771364055692e+02
GL_957 0 NS_957 NS_958 0 1.4899166019107438e-01
GL_958 0 NS_958 NS_957 0 -1.4899166019107438e-01
GS_957_9 0 NS_957 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 959/960
CS_959 NS_959 0 9.9999999999999998e-13
CS_960 NS_960 0 9.9999999999999998e-13
RS_959 NS_959 0 9.7194462506038604e+01
RS_960 NS_960 0 9.7194462506038604e+01
GL_959 0 NS_959 NS_960 0 1.4180400817347408e-01
GL_960 0 NS_960 NS_959 0 -1.4180400817347408e-01
GS_959_9 0 NS_959 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 961/962
CS_961 NS_961 0 9.9999999999999998e-13
CS_962 NS_962 0 9.9999999999999998e-13
RS_961 NS_961 0 1.0682825030924828e+02
RS_962 NS_962 0 1.0682825030924828e+02
GL_961 0 NS_961 NS_962 0 1.3872377519751058e-01
GL_962 0 NS_962 NS_961 0 -1.3872377519751058e-01
GS_961_9 0 NS_961 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 963/964
CS_963 NS_963 0 9.9999999999999998e-13
CS_964 NS_964 0 9.9999999999999998e-13
RS_963 NS_963 0 1.2559585119344567e+02
RS_964 NS_964 0 1.2559585119344568e+02
GL_963 0 NS_963 NS_964 0 1.3097721803321302e-01
GL_964 0 NS_964 NS_963 0 -1.3097721803321302e-01
GS_963_9 0 NS_963 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 965/966
CS_965 NS_965 0 9.9999999999999998e-13
CS_966 NS_966 0 9.9999999999999998e-13
RS_965 NS_965 0 1.0417660462554996e+02
RS_966 NS_966 0 1.0417660462554996e+02
GL_965 0 NS_965 NS_966 0 1.2625832867930367e-01
GL_966 0 NS_966 NS_965 0 -1.2625832867930367e-01
GS_965_9 0 NS_965 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 967/968
CS_967 NS_967 0 9.9999999999999998e-13
CS_968 NS_968 0 9.9999999999999998e-13
RS_967 NS_967 0 1.3317333532177352e+02
RS_968 NS_968 0 1.3317333532177352e+02
GL_967 0 NS_967 NS_968 0 1.2123672752714061e-01
GL_968 0 NS_968 NS_967 0 -1.2123672752714061e-01
GS_967_9 0 NS_967 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 969/970
CS_969 NS_969 0 9.9999999999999998e-13
CS_970 NS_970 0 9.9999999999999998e-13
RS_969 NS_969 0 1.2967831681616519e+02
RS_970 NS_970 0 1.2967831681616519e+02
GL_969 0 NS_969 NS_970 0 1.1651127865768855e-01
GL_970 0 NS_970 NS_969 0 -1.1651127865768855e-01
GS_969_9 0 NS_969 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 971/972
CS_971 NS_971 0 9.9999999999999998e-13
CS_972 NS_972 0 9.9999999999999998e-13
RS_971 NS_971 0 1.2999764374401394e+02
RS_972 NS_972 0 1.2999764374401394e+02
GL_971 0 NS_971 NS_972 0 1.1100247696987056e-01
GL_972 0 NS_972 NS_971 0 -1.1100247696987056e-01
GS_971_9 0 NS_971 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 973/974
CS_973 NS_973 0 9.9999999999999998e-13
CS_974 NS_974 0 9.9999999999999998e-13
RS_973 NS_973 0 1.2458814074636419e+02
RS_974 NS_974 0 1.2458814074636419e+02
GL_973 0 NS_973 NS_974 0 1.0660000212580591e-01
GL_974 0 NS_974 NS_973 0 -1.0660000212580591e-01
GS_973_9 0 NS_973 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 975/976
CS_975 NS_975 0 9.9999999999999998e-13
CS_976 NS_976 0 9.9999999999999998e-13
RS_975 NS_975 0 1.4677191614557748e+02
RS_976 NS_976 0 1.4677191614557748e+02
GL_975 0 NS_975 NS_976 0 1.0224733343325158e-01
GL_976 0 NS_976 NS_975 0 -1.0224733343325158e-01
GS_975_9 0 NS_975 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 977/978
CS_977 NS_977 0 9.9999999999999998e-13
CS_978 NS_978 0 9.9999999999999998e-13
RS_977 NS_977 0 1.3445989223131798e+02
RS_978 NS_978 0 1.3445989223131798e+02
GL_977 0 NS_977 NS_978 0 9.8177836948086503e-02
GL_978 0 NS_978 NS_977 0 -9.8177836948086503e-02
GS_977_9 0 NS_977 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 979/980
CS_979 NS_979 0 9.9999999999999998e-13
CS_980 NS_980 0 9.9999999999999998e-13
RS_979 NS_979 0 1.3187119040723775e+02
RS_980 NS_980 0 1.3187119040723772e+02
GL_979 0 NS_979 NS_980 0 9.2640196004122682e-02
GL_980 0 NS_980 NS_979 0 -9.2640196004122682e-02
GS_979_9 0 NS_979 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 981/982
CS_981 NS_981 0 9.9999999999999998e-13
CS_982 NS_982 0 9.9999999999999998e-13
RS_981 NS_981 0 1.2288401421230557e+02
RS_982 NS_982 0 1.2288401421230557e+02
GL_981 0 NS_981 NS_982 0 8.8704723748248199e-02
GL_982 0 NS_982 NS_981 0 -8.8704723748248199e-02
GS_981_9 0 NS_981 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 983/984
CS_983 NS_983 0 9.9999999999999998e-13
CS_984 NS_984 0 9.9999999999999998e-13
RS_983 NS_983 0 1.4123955654153085e+02
RS_984 NS_984 0 1.4123955654153082e+02
GL_983 0 NS_983 NS_984 0 8.4112474498892476e-02
GL_984 0 NS_984 NS_983 0 -8.4112474498892476e-02
GS_983_9 0 NS_983 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 985/986
CS_985 NS_985 0 9.9999999999999998e-13
CS_986 NS_986 0 9.9999999999999998e-13
RS_985 NS_985 0 1.2539447312269779e+02
RS_986 NS_986 0 1.2539447312269778e+02
GL_985 0 NS_985 NS_986 0 8.0007658848305588e-02
GL_986 0 NS_986 NS_985 0 -8.0007658848305588e-02
GS_985_9 0 NS_985 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 987/988
CS_987 NS_987 0 9.9999999999999998e-13
CS_988 NS_988 0 9.9999999999999998e-13
RS_987 NS_987 0 1.3219601779966965e+02
RS_988 NS_988 0 1.3219601779966968e+02
GL_987 0 NS_987 NS_988 0 7.4373183806052026e-02
GL_988 0 NS_988 NS_987 0 -7.4373183806052026e-02
GS_987_9 0 NS_987 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 989/990
CS_989 NS_989 0 9.9999999999999998e-13
CS_990 NS_990 0 9.9999999999999998e-13
RS_989 NS_989 0 1.1951371640958898e+02
RS_990 NS_990 0 1.1951371640958898e+02
GL_989 0 NS_989 NS_990 0 7.1003860961129844e-02
GL_990 0 NS_990 NS_989 0 -7.1003860961129844e-02
GS_989_9 0 NS_989 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 991/992
CS_991 NS_991 0 9.9999999999999998e-13
CS_992 NS_992 0 9.9999999999999998e-13
RS_991 NS_991 0 1.3491941875045018e+02
RS_992 NS_992 0 1.3491941875045018e+02
GL_991 0 NS_991 NS_992 0 6.5922080709048564e-02
GL_992 0 NS_992 NS_991 0 -6.5922080709048564e-02
GS_991_9 0 NS_991 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 993/994
CS_993 NS_993 0 9.9999999999999998e-13
CS_994 NS_994 0 9.9999999999999998e-13
RS_993 NS_993 0 1.2290405859347165e+02
RS_994 NS_994 0 1.2290405859347166e+02
GL_993 0 NS_993 NS_994 0 6.2340152915784278e-02
GL_994 0 NS_994 NS_993 0 -6.2340152915784278e-02
GS_993_9 0 NS_993 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 995/996
CS_995 NS_995 0 9.9999999999999998e-13
CS_996 NS_996 0 9.9999999999999998e-13
RS_995 NS_995 0 1.3258923845358959e+02
RS_996 NS_996 0 1.3258923845358959e+02
GL_995 0 NS_995 NS_996 0 5.6431081088718790e-02
GL_996 0 NS_996 NS_995 0 -5.6431081088718790e-02
GS_995_9 0 NS_995 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 997/998
CS_997 NS_997 0 9.9999999999999998e-13
CS_998 NS_998 0 9.9999999999999998e-13
RS_997 NS_997 0 1.0026704639246873e+02
RS_998 NS_998 0 1.0026704639246873e+02
GL_997 0 NS_997 NS_998 0 3.5068885856298401e-02
GL_998 0 NS_998 NS_997 0 -3.5068885856298401e-02
GS_997_9 0 NS_997 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 999/1000
CS_999 NS_999 0 9.9999999999999998e-13
CS_1000 NS_1000 0 9.9999999999999998e-13
RS_999 NS_999 0 1.2740726499710033e+02
RS_1000 NS_1000 0 1.2740726499710034e+02
GL_999 0 NS_999 NS_1000 0 5.3740629014256171e-02
GL_1000 0 NS_1000 NS_999 0 -5.3740629014256171e-02
GS_999_9 0 NS_999 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1001/1002
CS_1001 NS_1001 0 9.9999999999999998e-13
CS_1002 NS_1002 0 9.9999999999999998e-13
RS_1001 NS_1001 0 2.3804688106534087e+02
RS_1002 NS_1002 0 2.3804688106534090e+02
GL_1001 0 NS_1001 NS_1002 0 5.1425903265699464e-02
GL_1002 0 NS_1002 NS_1001 0 -5.1425903265699464e-02
GS_1001_9 0 NS_1001 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1003/1004
CS_1003 NS_1003 0 9.9999999999999998e-13
CS_1004 NS_1004 0 9.9999999999999998e-13
RS_1003 NS_1003 0 1.3728807739915800e+02
RS_1004 NS_1004 0 1.3728807739915803e+02
GL_1003 0 NS_1003 NS_1004 0 4.8031392820534764e-02
GL_1004 0 NS_1004 NS_1003 0 -4.8031392820534764e-02
GS_1003_9 0 NS_1003 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1005/1006
CS_1005 NS_1005 0 9.9999999999999998e-13
CS_1006 NS_1006 0 9.9999999999999998e-13
RS_1005 NS_1005 0 1.3499477893747948e+02
RS_1006 NS_1006 0 1.3499477893747945e+02
GL_1005 0 NS_1005 NS_1006 0 4.4453170742682194e-02
GL_1006 0 NS_1006 NS_1005 0 -4.4453170742682194e-02
GS_1005_9 0 NS_1005 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1007/1008
CS_1007 NS_1007 0 9.9999999999999998e-13
CS_1008 NS_1008 0 9.9999999999999998e-13
RS_1007 NS_1007 0 1.4121821834962651e+02
RS_1008 NS_1008 0 1.4121821834962651e+02
GL_1007 0 NS_1007 NS_1008 0 3.8464469217755697e-02
GL_1008 0 NS_1008 NS_1007 0 -3.8464469217755697e-02
GS_1007_9 0 NS_1007 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1009/1010
CS_1009 NS_1009 0 9.9999999999999998e-13
CS_1010 NS_1010 0 9.9999999999999998e-13
RS_1009 NS_1009 0 1.3946471282741149e+02
RS_1010 NS_1010 0 1.3946471282741149e+02
GL_1009 0 NS_1009 NS_1010 0 3.5678935079258622e-02
GL_1010 0 NS_1010 NS_1009 0 -3.5678935079258622e-02
GS_1009_9 0 NS_1009 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1011/1012
CS_1011 NS_1011 0 9.9999999999999998e-13
CS_1012 NS_1012 0 9.9999999999999998e-13
RS_1011 NS_1011 0 1.5530211191942624e+02
RS_1012 NS_1012 0 1.5530211191942627e+02
GL_1011 0 NS_1011 NS_1012 0 2.6209890345437525e-02
GL_1012 0 NS_1012 NS_1011 0 -2.6209890345437525e-02
GS_1011_9 0 NS_1011 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1013/1014
CS_1013 NS_1013 0 9.9999999999999998e-13
CS_1014 NS_1014 0 9.9999999999999998e-13
RS_1013 NS_1013 0 1.4887428879582419e+02
RS_1014 NS_1014 0 1.4887428879582419e+02
GL_1013 0 NS_1013 NS_1014 0 3.0330575323949095e-02
GL_1014 0 NS_1014 NS_1013 0 -3.0330575323949095e-02
GS_1013_9 0 NS_1013 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1015/1016
CS_1015 NS_1015 0 9.9999999999999998e-13
CS_1016 NS_1016 0 9.9999999999999998e-13
RS_1015 NS_1015 0 1.5087532095170570e+02
RS_1016 NS_1016 0 1.5087532095170570e+02
GL_1015 0 NS_1015 NS_1016 0 2.0034138441714564e-02
GL_1016 0 NS_1016 NS_1015 0 -2.0034138441714564e-02
GS_1015_9 0 NS_1015 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1017/1018
CS_1017 NS_1017 0 9.9999999999999998e-13
CS_1018 NS_1018 0 9.9999999999999998e-13
RS_1017 NS_1017 0 1.4763793449752018e+02
RS_1018 NS_1018 0 1.4763793449752018e+02
GL_1017 0 NS_1017 NS_1018 0 1.7017170579416537e-02
GL_1018 0 NS_1018 NS_1017 0 -1.7017170579416537e-02
GS_1017_9 0 NS_1017 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1019/1020
CS_1019 NS_1019 0 9.9999999999999998e-13
CS_1020 NS_1020 0 9.9999999999999998e-13
RS_1019 NS_1019 0 1.6285515224442304e+02
RS_1020 NS_1020 0 1.6285515224442304e+02
GL_1019 0 NS_1019 NS_1020 0 1.0897027002452746e-02
GL_1020 0 NS_1020 NS_1019 0 -1.0897027002452746e-02
GS_1019_9 0 NS_1019 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1021/1022
CS_1021 NS_1021 0 9.9999999999999998e-13
CS_1022 NS_1022 0 9.9999999999999998e-13
RS_1021 NS_1021 0 1.7239534388116820e+02
RS_1022 NS_1022 0 1.7239534388116820e+02
GL_1021 0 NS_1021 NS_1022 0 6.1589693699488982e-03
GL_1022 0 NS_1022 NS_1021 0 -6.1589693699488982e-03
GS_1021_9 0 NS_1021 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1023/1024
CS_1023 NS_1023 0 9.9999999999999998e-13
CS_1024 NS_1024 0 9.9999999999999998e-13
RS_1023 NS_1023 0 5.9928710578594173e+03
RS_1024 NS_1024 0 5.9928710578594173e+03
GL_1023 0 NS_1023 NS_1024 0 1.7541178006601681e-03
GL_1024 0 NS_1024 NS_1023 0 -1.7541178006601681e-03
GS_1023_9 0 NS_1023 NA_9 0 4.4027142044246531e-01
*
* Complex pair n. 1025/1026
CS_1025 NS_1025 0 9.9999999999999998e-13
CS_1026 NS_1026 0 9.9999999999999998e-13
RS_1025 NS_1025 0 8.0762087901330699e+02
RS_1026 NS_1026 0 8.0762087901330688e+02
GL_1025 0 NS_1025 NS_1026 0 1.7295489372816217e-03
GL_1026 0 NS_1026 NS_1025 0 -1.7295489372816217e-03
GS_1025_9 0 NS_1025 NA_9 0 4.4027142044246531e-01
*
* Real pole n. 1027
CS_1027 NS_1027 0 9.9999999999999998e-13
RS_1027 NS_1027 0 1.2857601077426406e+01
GS_1027_10 0 NS_1027 NA_10 0 4.4027142044246531e-01
*
* Real pole n. 1028
CS_1028 NS_1028 0 9.9999999999999998e-13
RS_1028 NS_1028 0 1.7282831464635029e+02
GS_1028_10 0 NS_1028 NA_10 0 4.4027142044246531e-01
*
* Real pole n. 1029
CS_1029 NS_1029 0 9.9999999999999998e-13
RS_1029 NS_1029 0 5.5743135126264733e+03
GS_1029_10 0 NS_1029 NA_10 0 4.4027142044246531e-01
*
* Real pole n. 1030
CS_1030 NS_1030 0 9.9999999999999998e-13
RS_1030 NS_1030 0 1.3594126013480764e+03
GS_1030_10 0 NS_1030 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1031/1032
CS_1031 NS_1031 0 9.9999999999999998e-13
CS_1032 NS_1032 0 9.9999999999999998e-13
RS_1031 NS_1031 0 1.7904812183888848e+02
RS_1032 NS_1032 0 1.7904812183888848e+02
GL_1031 0 NS_1031 NS_1032 0 2.6007898045516648e-01
GL_1032 0 NS_1032 NS_1031 0 -2.6007898045516648e-01
GS_1031_10 0 NS_1031 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1033/1034
CS_1033 NS_1033 0 9.9999999999999998e-13
CS_1034 NS_1034 0 9.9999999999999998e-13
RS_1033 NS_1033 0 1.2615541320340381e+02
RS_1034 NS_1034 0 1.2615541320340381e+02
GL_1033 0 NS_1033 NS_1034 0 2.5243684762014923e-01
GL_1034 0 NS_1034 NS_1033 0 -2.5243684762014923e-01
GS_1033_10 0 NS_1033 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1035/1036
CS_1035 NS_1035 0 9.9999999999999998e-13
CS_1036 NS_1036 0 9.9999999999999998e-13
RS_1035 NS_1035 0 1.0219948841586964e+02
RS_1036 NS_1036 0 1.0219948841586965e+02
GL_1035 0 NS_1035 NS_1036 0 2.4690226903121384e-01
GL_1036 0 NS_1036 NS_1035 0 -2.4690226903121384e-01
GS_1035_10 0 NS_1035 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1037/1038
CS_1037 NS_1037 0 9.9999999999999998e-13
CS_1038 NS_1038 0 9.9999999999999998e-13
RS_1037 NS_1037 0 1.1002436853144543e+02
RS_1038 NS_1038 0 1.1002436853144542e+02
GL_1037 0 NS_1037 NS_1038 0 2.4293768067729948e-01
GL_1038 0 NS_1038 NS_1037 0 -2.4293768067729948e-01
GS_1037_10 0 NS_1037 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1039/1040
CS_1039 NS_1039 0 9.9999999999999998e-13
CS_1040 NS_1040 0 9.9999999999999998e-13
RS_1039 NS_1039 0 1.0553430908077024e+02
RS_1040 NS_1040 0 1.0553430908077026e+02
GL_1039 0 NS_1039 NS_1040 0 2.3600513224442521e-01
GL_1040 0 NS_1040 NS_1039 0 -2.3600513224442521e-01
GS_1039_10 0 NS_1039 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1041/1042
CS_1041 NS_1041 0 9.9999999999999998e-13
CS_1042 NS_1042 0 9.9999999999999998e-13
RS_1041 NS_1041 0 1.0759915098440327e+02
RS_1042 NS_1042 0 1.0759915098440327e+02
GL_1041 0 NS_1041 NS_1042 0 2.3090539914362113e-01
GL_1042 0 NS_1042 NS_1041 0 -2.3090539914362113e-01
GS_1041_10 0 NS_1041 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1043/1044
CS_1043 NS_1043 0 9.9999999999999998e-13
CS_1044 NS_1044 0 9.9999999999999998e-13
RS_1043 NS_1043 0 1.3295415758774385e+02
RS_1044 NS_1044 0 1.3295415758774385e+02
GL_1043 0 NS_1043 NS_1044 0 2.3030066292345727e-01
GL_1044 0 NS_1044 NS_1043 0 -2.3030066292345727e-01
GS_1043_10 0 NS_1043 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1045/1046
CS_1045 NS_1045 0 9.9999999999999998e-13
CS_1046 NS_1046 0 9.9999999999999998e-13
RS_1045 NS_1045 0 1.1432186998941940e+02
RS_1046 NS_1046 0 1.1432186998941938e+02
GL_1045 0 NS_1045 NS_1046 0 2.2451058023508991e-01
GL_1046 0 NS_1046 NS_1045 0 -2.2451058023508991e-01
GS_1045_10 0 NS_1045 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1047/1048
CS_1047 NS_1047 0 9.9999999999999998e-13
CS_1048 NS_1048 0 9.9999999999999998e-13
RS_1047 NS_1047 0 9.0812703249943667e+01
RS_1048 NS_1048 0 9.0812703249943652e+01
GL_1047 0 NS_1047 NS_1048 0 2.1702628900531115e-01
GL_1048 0 NS_1048 NS_1047 0 -2.1702628900531115e-01
GS_1047_10 0 NS_1047 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1049/1050
CS_1049 NS_1049 0 9.9999999999999998e-13
CS_1050 NS_1050 0 9.9999999999999998e-13
RS_1049 NS_1049 0 9.5643803662064585e+01
RS_1050 NS_1050 0 9.5643803662064585e+01
GL_1049 0 NS_1049 NS_1050 0 2.1448200383207913e-01
GL_1050 0 NS_1050 NS_1049 0 -2.1448200383207913e-01
GS_1049_10 0 NS_1049 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1051/1052
CS_1051 NS_1051 0 9.9999999999999998e-13
CS_1052 NS_1052 0 9.9999999999999998e-13
RS_1051 NS_1051 0 1.0631957479149644e+02
RS_1052 NS_1052 0 1.0631957479149644e+02
GL_1051 0 NS_1051 NS_1052 0 2.0655001587884311e-01
GL_1052 0 NS_1052 NS_1051 0 -2.0655001587884311e-01
GS_1051_10 0 NS_1051 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1053/1054
CS_1053 NS_1053 0 9.9999999999999998e-13
CS_1054 NS_1054 0 9.9999999999999998e-13
RS_1053 NS_1053 0 7.9907264643295406e+01
RS_1054 NS_1054 0 7.9907264643295420e+01
GL_1053 0 NS_1053 NS_1054 0 2.0133773147328893e-01
GL_1054 0 NS_1054 NS_1053 0 -2.0133773147328893e-01
GS_1053_10 0 NS_1053 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1055/1056
CS_1055 NS_1055 0 9.9999999999999998e-13
CS_1056 NS_1056 0 9.9999999999999998e-13
RS_1055 NS_1055 0 1.0625506887893997e+02
RS_1056 NS_1056 0 1.0625506887893997e+02
GL_1055 0 NS_1055 NS_1056 0 1.9628877333023340e-01
GL_1056 0 NS_1056 NS_1055 0 -1.9628877333023340e-01
GS_1055_10 0 NS_1055 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1057/1058
CS_1057 NS_1057 0 9.9999999999999998e-13
CS_1058 NS_1058 0 9.9999999999999998e-13
RS_1057 NS_1057 0 9.6115312638592201e+01
RS_1058 NS_1058 0 9.6115312638592201e+01
GL_1057 0 NS_1057 NS_1058 0 1.8794816712418483e-01
GL_1058 0 NS_1058 NS_1057 0 -1.8794816712418483e-01
GS_1057_10 0 NS_1057 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1059/1060
CS_1059 NS_1059 0 9.9999999999999998e-13
CS_1060 NS_1060 0 9.9999999999999998e-13
RS_1059 NS_1059 0 8.5212696574118169e+01
RS_1060 NS_1060 0 8.5212696574118169e+01
GL_1059 0 NS_1059 NS_1060 0 1.8572140881490298e-01
GL_1060 0 NS_1060 NS_1059 0 -1.8572140881490298e-01
GS_1059_10 0 NS_1059 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1061/1062
CS_1061 NS_1061 0 9.9999999999999998e-13
CS_1062 NS_1062 0 9.9999999999999998e-13
RS_1061 NS_1061 0 1.0905026103375434e+02
RS_1062 NS_1062 0 1.0905026103375432e+02
GL_1061 0 NS_1061 NS_1062 0 1.7785621200284463e-01
GL_1062 0 NS_1062 NS_1061 0 -1.7785621200284463e-01
GS_1061_10 0 NS_1061 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1063/1064
CS_1063 NS_1063 0 9.9999999999999998e-13
CS_1064 NS_1064 0 9.9999999999999998e-13
RS_1063 NS_1063 0 8.3024437910787526e+01
RS_1064 NS_1064 0 8.3024437910787526e+01
GL_1063 0 NS_1063 NS_1064 0 1.7164509875911016e-01
GL_1064 0 NS_1064 NS_1063 0 -1.7164509875911016e-01
GS_1063_10 0 NS_1063 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1065/1066
CS_1065 NS_1065 0 9.9999999999999998e-13
CS_1066 NS_1066 0 9.9999999999999998e-13
RS_1065 NS_1065 0 1.0548793856392000e+02
RS_1066 NS_1066 0 1.0548793856392000e+02
GL_1065 0 NS_1065 NS_1066 0 1.6750370916002649e-01
GL_1066 0 NS_1066 NS_1065 0 -1.6750370916002649e-01
GS_1065_10 0 NS_1065 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1067/1068
CS_1067 NS_1067 0 9.9999999999999998e-13
CS_1068 NS_1068 0 9.9999999999999998e-13
RS_1067 NS_1067 0 1.0753754351502513e+02
RS_1068 NS_1068 0 1.0753754351502513e+02
GL_1067 0 NS_1067 NS_1068 0 1.5942172238060490e-01
GL_1068 0 NS_1068 NS_1067 0 -1.5942172238060490e-01
GS_1067_10 0 NS_1067 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1069/1070
CS_1069 NS_1069 0 9.9999999999999998e-13
CS_1070 NS_1070 0 9.9999999999999998e-13
RS_1069 NS_1069 0 8.6961097797504721e+01
RS_1070 NS_1070 0 8.6961097797504721e+01
GL_1069 0 NS_1069 NS_1070 0 1.5553892891442009e-01
GL_1070 0 NS_1070 NS_1069 0 -1.5553892891442009e-01
GS_1069_10 0 NS_1069 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1071/1072
CS_1071 NS_1071 0 9.9999999999999998e-13
CS_1072 NS_1072 0 9.9999999999999998e-13
RS_1071 NS_1071 0 1.1549771364055694e+02
RS_1072 NS_1072 0 1.1549771364055692e+02
GL_1071 0 NS_1071 NS_1072 0 1.4899166019107438e-01
GL_1072 0 NS_1072 NS_1071 0 -1.4899166019107438e-01
GS_1071_10 0 NS_1071 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1073/1074
CS_1073 NS_1073 0 9.9999999999999998e-13
CS_1074 NS_1074 0 9.9999999999999998e-13
RS_1073 NS_1073 0 9.7194462506038604e+01
RS_1074 NS_1074 0 9.7194462506038604e+01
GL_1073 0 NS_1073 NS_1074 0 1.4180400817347408e-01
GL_1074 0 NS_1074 NS_1073 0 -1.4180400817347408e-01
GS_1073_10 0 NS_1073 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1075/1076
CS_1075 NS_1075 0 9.9999999999999998e-13
CS_1076 NS_1076 0 9.9999999999999998e-13
RS_1075 NS_1075 0 1.0682825030924828e+02
RS_1076 NS_1076 0 1.0682825030924828e+02
GL_1075 0 NS_1075 NS_1076 0 1.3872377519751058e-01
GL_1076 0 NS_1076 NS_1075 0 -1.3872377519751058e-01
GS_1075_10 0 NS_1075 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1077/1078
CS_1077 NS_1077 0 9.9999999999999998e-13
CS_1078 NS_1078 0 9.9999999999999998e-13
RS_1077 NS_1077 0 1.2559585119344567e+02
RS_1078 NS_1078 0 1.2559585119344568e+02
GL_1077 0 NS_1077 NS_1078 0 1.3097721803321302e-01
GL_1078 0 NS_1078 NS_1077 0 -1.3097721803321302e-01
GS_1077_10 0 NS_1077 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1079/1080
CS_1079 NS_1079 0 9.9999999999999998e-13
CS_1080 NS_1080 0 9.9999999999999998e-13
RS_1079 NS_1079 0 1.0417660462554996e+02
RS_1080 NS_1080 0 1.0417660462554996e+02
GL_1079 0 NS_1079 NS_1080 0 1.2625832867930367e-01
GL_1080 0 NS_1080 NS_1079 0 -1.2625832867930367e-01
GS_1079_10 0 NS_1079 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1081/1082
CS_1081 NS_1081 0 9.9999999999999998e-13
CS_1082 NS_1082 0 9.9999999999999998e-13
RS_1081 NS_1081 0 1.3317333532177352e+02
RS_1082 NS_1082 0 1.3317333532177352e+02
GL_1081 0 NS_1081 NS_1082 0 1.2123672752714061e-01
GL_1082 0 NS_1082 NS_1081 0 -1.2123672752714061e-01
GS_1081_10 0 NS_1081 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1083/1084
CS_1083 NS_1083 0 9.9999999999999998e-13
CS_1084 NS_1084 0 9.9999999999999998e-13
RS_1083 NS_1083 0 1.2967831681616519e+02
RS_1084 NS_1084 0 1.2967831681616519e+02
GL_1083 0 NS_1083 NS_1084 0 1.1651127865768855e-01
GL_1084 0 NS_1084 NS_1083 0 -1.1651127865768855e-01
GS_1083_10 0 NS_1083 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1085/1086
CS_1085 NS_1085 0 9.9999999999999998e-13
CS_1086 NS_1086 0 9.9999999999999998e-13
RS_1085 NS_1085 0 1.2999764374401394e+02
RS_1086 NS_1086 0 1.2999764374401394e+02
GL_1085 0 NS_1085 NS_1086 0 1.1100247696987056e-01
GL_1086 0 NS_1086 NS_1085 0 -1.1100247696987056e-01
GS_1085_10 0 NS_1085 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1087/1088
CS_1087 NS_1087 0 9.9999999999999998e-13
CS_1088 NS_1088 0 9.9999999999999998e-13
RS_1087 NS_1087 0 1.2458814074636419e+02
RS_1088 NS_1088 0 1.2458814074636419e+02
GL_1087 0 NS_1087 NS_1088 0 1.0660000212580591e-01
GL_1088 0 NS_1088 NS_1087 0 -1.0660000212580591e-01
GS_1087_10 0 NS_1087 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1089/1090
CS_1089 NS_1089 0 9.9999999999999998e-13
CS_1090 NS_1090 0 9.9999999999999998e-13
RS_1089 NS_1089 0 1.4677191614557748e+02
RS_1090 NS_1090 0 1.4677191614557748e+02
GL_1089 0 NS_1089 NS_1090 0 1.0224733343325158e-01
GL_1090 0 NS_1090 NS_1089 0 -1.0224733343325158e-01
GS_1089_10 0 NS_1089 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1091/1092
CS_1091 NS_1091 0 9.9999999999999998e-13
CS_1092 NS_1092 0 9.9999999999999998e-13
RS_1091 NS_1091 0 1.3445989223131798e+02
RS_1092 NS_1092 0 1.3445989223131798e+02
GL_1091 0 NS_1091 NS_1092 0 9.8177836948086503e-02
GL_1092 0 NS_1092 NS_1091 0 -9.8177836948086503e-02
GS_1091_10 0 NS_1091 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1093/1094
CS_1093 NS_1093 0 9.9999999999999998e-13
CS_1094 NS_1094 0 9.9999999999999998e-13
RS_1093 NS_1093 0 1.3187119040723775e+02
RS_1094 NS_1094 0 1.3187119040723772e+02
GL_1093 0 NS_1093 NS_1094 0 9.2640196004122682e-02
GL_1094 0 NS_1094 NS_1093 0 -9.2640196004122682e-02
GS_1093_10 0 NS_1093 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1095/1096
CS_1095 NS_1095 0 9.9999999999999998e-13
CS_1096 NS_1096 0 9.9999999999999998e-13
RS_1095 NS_1095 0 1.2288401421230557e+02
RS_1096 NS_1096 0 1.2288401421230557e+02
GL_1095 0 NS_1095 NS_1096 0 8.8704723748248199e-02
GL_1096 0 NS_1096 NS_1095 0 -8.8704723748248199e-02
GS_1095_10 0 NS_1095 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1097/1098
CS_1097 NS_1097 0 9.9999999999999998e-13
CS_1098 NS_1098 0 9.9999999999999998e-13
RS_1097 NS_1097 0 1.4123955654153085e+02
RS_1098 NS_1098 0 1.4123955654153082e+02
GL_1097 0 NS_1097 NS_1098 0 8.4112474498892476e-02
GL_1098 0 NS_1098 NS_1097 0 -8.4112474498892476e-02
GS_1097_10 0 NS_1097 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1099/1100
CS_1099 NS_1099 0 9.9999999999999998e-13
CS_1100 NS_1100 0 9.9999999999999998e-13
RS_1099 NS_1099 0 1.2539447312269779e+02
RS_1100 NS_1100 0 1.2539447312269778e+02
GL_1099 0 NS_1099 NS_1100 0 8.0007658848305588e-02
GL_1100 0 NS_1100 NS_1099 0 -8.0007658848305588e-02
GS_1099_10 0 NS_1099 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1101/1102
CS_1101 NS_1101 0 9.9999999999999998e-13
CS_1102 NS_1102 0 9.9999999999999998e-13
RS_1101 NS_1101 0 1.3219601779966965e+02
RS_1102 NS_1102 0 1.3219601779966968e+02
GL_1101 0 NS_1101 NS_1102 0 7.4373183806052026e-02
GL_1102 0 NS_1102 NS_1101 0 -7.4373183806052026e-02
GS_1101_10 0 NS_1101 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1103/1104
CS_1103 NS_1103 0 9.9999999999999998e-13
CS_1104 NS_1104 0 9.9999999999999998e-13
RS_1103 NS_1103 0 1.1951371640958898e+02
RS_1104 NS_1104 0 1.1951371640958898e+02
GL_1103 0 NS_1103 NS_1104 0 7.1003860961129844e-02
GL_1104 0 NS_1104 NS_1103 0 -7.1003860961129844e-02
GS_1103_10 0 NS_1103 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1105/1106
CS_1105 NS_1105 0 9.9999999999999998e-13
CS_1106 NS_1106 0 9.9999999999999998e-13
RS_1105 NS_1105 0 1.3491941875045018e+02
RS_1106 NS_1106 0 1.3491941875045018e+02
GL_1105 0 NS_1105 NS_1106 0 6.5922080709048564e-02
GL_1106 0 NS_1106 NS_1105 0 -6.5922080709048564e-02
GS_1105_10 0 NS_1105 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1107/1108
CS_1107 NS_1107 0 9.9999999999999998e-13
CS_1108 NS_1108 0 9.9999999999999998e-13
RS_1107 NS_1107 0 1.2290405859347165e+02
RS_1108 NS_1108 0 1.2290405859347166e+02
GL_1107 0 NS_1107 NS_1108 0 6.2340152915784278e-02
GL_1108 0 NS_1108 NS_1107 0 -6.2340152915784278e-02
GS_1107_10 0 NS_1107 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1109/1110
CS_1109 NS_1109 0 9.9999999999999998e-13
CS_1110 NS_1110 0 9.9999999999999998e-13
RS_1109 NS_1109 0 1.3258923845358959e+02
RS_1110 NS_1110 0 1.3258923845358959e+02
GL_1109 0 NS_1109 NS_1110 0 5.6431081088718790e-02
GL_1110 0 NS_1110 NS_1109 0 -5.6431081088718790e-02
GS_1109_10 0 NS_1109 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1111/1112
CS_1111 NS_1111 0 9.9999999999999998e-13
CS_1112 NS_1112 0 9.9999999999999998e-13
RS_1111 NS_1111 0 1.0026704639246873e+02
RS_1112 NS_1112 0 1.0026704639246873e+02
GL_1111 0 NS_1111 NS_1112 0 3.5068885856298401e-02
GL_1112 0 NS_1112 NS_1111 0 -3.5068885856298401e-02
GS_1111_10 0 NS_1111 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1113/1114
CS_1113 NS_1113 0 9.9999999999999998e-13
CS_1114 NS_1114 0 9.9999999999999998e-13
RS_1113 NS_1113 0 1.2740726499710033e+02
RS_1114 NS_1114 0 1.2740726499710034e+02
GL_1113 0 NS_1113 NS_1114 0 5.3740629014256171e-02
GL_1114 0 NS_1114 NS_1113 0 -5.3740629014256171e-02
GS_1113_10 0 NS_1113 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1115/1116
CS_1115 NS_1115 0 9.9999999999999998e-13
CS_1116 NS_1116 0 9.9999999999999998e-13
RS_1115 NS_1115 0 2.3804688106534087e+02
RS_1116 NS_1116 0 2.3804688106534090e+02
GL_1115 0 NS_1115 NS_1116 0 5.1425903265699464e-02
GL_1116 0 NS_1116 NS_1115 0 -5.1425903265699464e-02
GS_1115_10 0 NS_1115 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1117/1118
CS_1117 NS_1117 0 9.9999999999999998e-13
CS_1118 NS_1118 0 9.9999999999999998e-13
RS_1117 NS_1117 0 1.3728807739915800e+02
RS_1118 NS_1118 0 1.3728807739915803e+02
GL_1117 0 NS_1117 NS_1118 0 4.8031392820534764e-02
GL_1118 0 NS_1118 NS_1117 0 -4.8031392820534764e-02
GS_1117_10 0 NS_1117 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1119/1120
CS_1119 NS_1119 0 9.9999999999999998e-13
CS_1120 NS_1120 0 9.9999999999999998e-13
RS_1119 NS_1119 0 1.3499477893747948e+02
RS_1120 NS_1120 0 1.3499477893747945e+02
GL_1119 0 NS_1119 NS_1120 0 4.4453170742682194e-02
GL_1120 0 NS_1120 NS_1119 0 -4.4453170742682194e-02
GS_1119_10 0 NS_1119 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1121/1122
CS_1121 NS_1121 0 9.9999999999999998e-13
CS_1122 NS_1122 0 9.9999999999999998e-13
RS_1121 NS_1121 0 1.4121821834962651e+02
RS_1122 NS_1122 0 1.4121821834962651e+02
GL_1121 0 NS_1121 NS_1122 0 3.8464469217755697e-02
GL_1122 0 NS_1122 NS_1121 0 -3.8464469217755697e-02
GS_1121_10 0 NS_1121 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1123/1124
CS_1123 NS_1123 0 9.9999999999999998e-13
CS_1124 NS_1124 0 9.9999999999999998e-13
RS_1123 NS_1123 0 1.3946471282741149e+02
RS_1124 NS_1124 0 1.3946471282741149e+02
GL_1123 0 NS_1123 NS_1124 0 3.5678935079258622e-02
GL_1124 0 NS_1124 NS_1123 0 -3.5678935079258622e-02
GS_1123_10 0 NS_1123 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1125/1126
CS_1125 NS_1125 0 9.9999999999999998e-13
CS_1126 NS_1126 0 9.9999999999999998e-13
RS_1125 NS_1125 0 1.5530211191942624e+02
RS_1126 NS_1126 0 1.5530211191942627e+02
GL_1125 0 NS_1125 NS_1126 0 2.6209890345437525e-02
GL_1126 0 NS_1126 NS_1125 0 -2.6209890345437525e-02
GS_1125_10 0 NS_1125 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1127/1128
CS_1127 NS_1127 0 9.9999999999999998e-13
CS_1128 NS_1128 0 9.9999999999999998e-13
RS_1127 NS_1127 0 1.4887428879582419e+02
RS_1128 NS_1128 0 1.4887428879582419e+02
GL_1127 0 NS_1127 NS_1128 0 3.0330575323949095e-02
GL_1128 0 NS_1128 NS_1127 0 -3.0330575323949095e-02
GS_1127_10 0 NS_1127 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1129/1130
CS_1129 NS_1129 0 9.9999999999999998e-13
CS_1130 NS_1130 0 9.9999999999999998e-13
RS_1129 NS_1129 0 1.5087532095170570e+02
RS_1130 NS_1130 0 1.5087532095170570e+02
GL_1129 0 NS_1129 NS_1130 0 2.0034138441714564e-02
GL_1130 0 NS_1130 NS_1129 0 -2.0034138441714564e-02
GS_1129_10 0 NS_1129 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1131/1132
CS_1131 NS_1131 0 9.9999999999999998e-13
CS_1132 NS_1132 0 9.9999999999999998e-13
RS_1131 NS_1131 0 1.4763793449752018e+02
RS_1132 NS_1132 0 1.4763793449752018e+02
GL_1131 0 NS_1131 NS_1132 0 1.7017170579416537e-02
GL_1132 0 NS_1132 NS_1131 0 -1.7017170579416537e-02
GS_1131_10 0 NS_1131 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1133/1134
CS_1133 NS_1133 0 9.9999999999999998e-13
CS_1134 NS_1134 0 9.9999999999999998e-13
RS_1133 NS_1133 0 1.6285515224442304e+02
RS_1134 NS_1134 0 1.6285515224442304e+02
GL_1133 0 NS_1133 NS_1134 0 1.0897027002452746e-02
GL_1134 0 NS_1134 NS_1133 0 -1.0897027002452746e-02
GS_1133_10 0 NS_1133 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1135/1136
CS_1135 NS_1135 0 9.9999999999999998e-13
CS_1136 NS_1136 0 9.9999999999999998e-13
RS_1135 NS_1135 0 1.7239534388116820e+02
RS_1136 NS_1136 0 1.7239534388116820e+02
GL_1135 0 NS_1135 NS_1136 0 6.1589693699488982e-03
GL_1136 0 NS_1136 NS_1135 0 -6.1589693699488982e-03
GS_1135_10 0 NS_1135 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1137/1138
CS_1137 NS_1137 0 9.9999999999999998e-13
CS_1138 NS_1138 0 9.9999999999999998e-13
RS_1137 NS_1137 0 5.9928710578594173e+03
RS_1138 NS_1138 0 5.9928710578594173e+03
GL_1137 0 NS_1137 NS_1138 0 1.7541178006601681e-03
GL_1138 0 NS_1138 NS_1137 0 -1.7541178006601681e-03
GS_1137_10 0 NS_1137 NA_10 0 4.4027142044246531e-01
*
* Complex pair n. 1139/1140
CS_1139 NS_1139 0 9.9999999999999998e-13
CS_1140 NS_1140 0 9.9999999999999998e-13
RS_1139 NS_1139 0 8.0762087901330699e+02
RS_1140 NS_1140 0 8.0762087901330688e+02
GL_1139 0 NS_1139 NS_1140 0 1.7295489372816217e-03
GL_1140 0 NS_1140 NS_1139 0 -1.7295489372816217e-03
GS_1139_10 0 NS_1139 NA_10 0 4.4027142044246531e-01
*
* Real pole n. 1141
CS_1141 NS_1141 0 9.9999999999999998e-13
RS_1141 NS_1141 0 1.2857601077426406e+01
GS_1141_11 0 NS_1141 NA_11 0 4.4027142044246531e-01
*
* Real pole n. 1142
CS_1142 NS_1142 0 9.9999999999999998e-13
RS_1142 NS_1142 0 1.7282831464635029e+02
GS_1142_11 0 NS_1142 NA_11 0 4.4027142044246531e-01
*
* Real pole n. 1143
CS_1143 NS_1143 0 9.9999999999999998e-13
RS_1143 NS_1143 0 5.5743135126264733e+03
GS_1143_11 0 NS_1143 NA_11 0 4.4027142044246531e-01
*
* Real pole n. 1144
CS_1144 NS_1144 0 9.9999999999999998e-13
RS_1144 NS_1144 0 1.3594126013480764e+03
GS_1144_11 0 NS_1144 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1145/1146
CS_1145 NS_1145 0 9.9999999999999998e-13
CS_1146 NS_1146 0 9.9999999999999998e-13
RS_1145 NS_1145 0 1.7904812183888848e+02
RS_1146 NS_1146 0 1.7904812183888848e+02
GL_1145 0 NS_1145 NS_1146 0 2.6007898045516648e-01
GL_1146 0 NS_1146 NS_1145 0 -2.6007898045516648e-01
GS_1145_11 0 NS_1145 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1147/1148
CS_1147 NS_1147 0 9.9999999999999998e-13
CS_1148 NS_1148 0 9.9999999999999998e-13
RS_1147 NS_1147 0 1.2615541320340381e+02
RS_1148 NS_1148 0 1.2615541320340381e+02
GL_1147 0 NS_1147 NS_1148 0 2.5243684762014923e-01
GL_1148 0 NS_1148 NS_1147 0 -2.5243684762014923e-01
GS_1147_11 0 NS_1147 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1149/1150
CS_1149 NS_1149 0 9.9999999999999998e-13
CS_1150 NS_1150 0 9.9999999999999998e-13
RS_1149 NS_1149 0 1.0219948841586964e+02
RS_1150 NS_1150 0 1.0219948841586965e+02
GL_1149 0 NS_1149 NS_1150 0 2.4690226903121384e-01
GL_1150 0 NS_1150 NS_1149 0 -2.4690226903121384e-01
GS_1149_11 0 NS_1149 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1151/1152
CS_1151 NS_1151 0 9.9999999999999998e-13
CS_1152 NS_1152 0 9.9999999999999998e-13
RS_1151 NS_1151 0 1.1002436853144543e+02
RS_1152 NS_1152 0 1.1002436853144542e+02
GL_1151 0 NS_1151 NS_1152 0 2.4293768067729948e-01
GL_1152 0 NS_1152 NS_1151 0 -2.4293768067729948e-01
GS_1151_11 0 NS_1151 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1153/1154
CS_1153 NS_1153 0 9.9999999999999998e-13
CS_1154 NS_1154 0 9.9999999999999998e-13
RS_1153 NS_1153 0 1.0553430908077024e+02
RS_1154 NS_1154 0 1.0553430908077026e+02
GL_1153 0 NS_1153 NS_1154 0 2.3600513224442521e-01
GL_1154 0 NS_1154 NS_1153 0 -2.3600513224442521e-01
GS_1153_11 0 NS_1153 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1155/1156
CS_1155 NS_1155 0 9.9999999999999998e-13
CS_1156 NS_1156 0 9.9999999999999998e-13
RS_1155 NS_1155 0 1.0759915098440327e+02
RS_1156 NS_1156 0 1.0759915098440327e+02
GL_1155 0 NS_1155 NS_1156 0 2.3090539914362113e-01
GL_1156 0 NS_1156 NS_1155 0 -2.3090539914362113e-01
GS_1155_11 0 NS_1155 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1157/1158
CS_1157 NS_1157 0 9.9999999999999998e-13
CS_1158 NS_1158 0 9.9999999999999998e-13
RS_1157 NS_1157 0 1.3295415758774385e+02
RS_1158 NS_1158 0 1.3295415758774385e+02
GL_1157 0 NS_1157 NS_1158 0 2.3030066292345727e-01
GL_1158 0 NS_1158 NS_1157 0 -2.3030066292345727e-01
GS_1157_11 0 NS_1157 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1159/1160
CS_1159 NS_1159 0 9.9999999999999998e-13
CS_1160 NS_1160 0 9.9999999999999998e-13
RS_1159 NS_1159 0 1.1432186998941940e+02
RS_1160 NS_1160 0 1.1432186998941938e+02
GL_1159 0 NS_1159 NS_1160 0 2.2451058023508991e-01
GL_1160 0 NS_1160 NS_1159 0 -2.2451058023508991e-01
GS_1159_11 0 NS_1159 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1161/1162
CS_1161 NS_1161 0 9.9999999999999998e-13
CS_1162 NS_1162 0 9.9999999999999998e-13
RS_1161 NS_1161 0 9.0812703249943667e+01
RS_1162 NS_1162 0 9.0812703249943652e+01
GL_1161 0 NS_1161 NS_1162 0 2.1702628900531115e-01
GL_1162 0 NS_1162 NS_1161 0 -2.1702628900531115e-01
GS_1161_11 0 NS_1161 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1163/1164
CS_1163 NS_1163 0 9.9999999999999998e-13
CS_1164 NS_1164 0 9.9999999999999998e-13
RS_1163 NS_1163 0 9.5643803662064585e+01
RS_1164 NS_1164 0 9.5643803662064585e+01
GL_1163 0 NS_1163 NS_1164 0 2.1448200383207913e-01
GL_1164 0 NS_1164 NS_1163 0 -2.1448200383207913e-01
GS_1163_11 0 NS_1163 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1165/1166
CS_1165 NS_1165 0 9.9999999999999998e-13
CS_1166 NS_1166 0 9.9999999999999998e-13
RS_1165 NS_1165 0 1.0631957479149644e+02
RS_1166 NS_1166 0 1.0631957479149644e+02
GL_1165 0 NS_1165 NS_1166 0 2.0655001587884311e-01
GL_1166 0 NS_1166 NS_1165 0 -2.0655001587884311e-01
GS_1165_11 0 NS_1165 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1167/1168
CS_1167 NS_1167 0 9.9999999999999998e-13
CS_1168 NS_1168 0 9.9999999999999998e-13
RS_1167 NS_1167 0 7.9907264643295406e+01
RS_1168 NS_1168 0 7.9907264643295420e+01
GL_1167 0 NS_1167 NS_1168 0 2.0133773147328893e-01
GL_1168 0 NS_1168 NS_1167 0 -2.0133773147328893e-01
GS_1167_11 0 NS_1167 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1169/1170
CS_1169 NS_1169 0 9.9999999999999998e-13
CS_1170 NS_1170 0 9.9999999999999998e-13
RS_1169 NS_1169 0 1.0625506887893997e+02
RS_1170 NS_1170 0 1.0625506887893997e+02
GL_1169 0 NS_1169 NS_1170 0 1.9628877333023340e-01
GL_1170 0 NS_1170 NS_1169 0 -1.9628877333023340e-01
GS_1169_11 0 NS_1169 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1171/1172
CS_1171 NS_1171 0 9.9999999999999998e-13
CS_1172 NS_1172 0 9.9999999999999998e-13
RS_1171 NS_1171 0 9.6115312638592201e+01
RS_1172 NS_1172 0 9.6115312638592201e+01
GL_1171 0 NS_1171 NS_1172 0 1.8794816712418483e-01
GL_1172 0 NS_1172 NS_1171 0 -1.8794816712418483e-01
GS_1171_11 0 NS_1171 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1173/1174
CS_1173 NS_1173 0 9.9999999999999998e-13
CS_1174 NS_1174 0 9.9999999999999998e-13
RS_1173 NS_1173 0 8.5212696574118169e+01
RS_1174 NS_1174 0 8.5212696574118169e+01
GL_1173 0 NS_1173 NS_1174 0 1.8572140881490298e-01
GL_1174 0 NS_1174 NS_1173 0 -1.8572140881490298e-01
GS_1173_11 0 NS_1173 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1175/1176
CS_1175 NS_1175 0 9.9999999999999998e-13
CS_1176 NS_1176 0 9.9999999999999998e-13
RS_1175 NS_1175 0 1.0905026103375434e+02
RS_1176 NS_1176 0 1.0905026103375432e+02
GL_1175 0 NS_1175 NS_1176 0 1.7785621200284463e-01
GL_1176 0 NS_1176 NS_1175 0 -1.7785621200284463e-01
GS_1175_11 0 NS_1175 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1177/1178
CS_1177 NS_1177 0 9.9999999999999998e-13
CS_1178 NS_1178 0 9.9999999999999998e-13
RS_1177 NS_1177 0 8.3024437910787526e+01
RS_1178 NS_1178 0 8.3024437910787526e+01
GL_1177 0 NS_1177 NS_1178 0 1.7164509875911016e-01
GL_1178 0 NS_1178 NS_1177 0 -1.7164509875911016e-01
GS_1177_11 0 NS_1177 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1179/1180
CS_1179 NS_1179 0 9.9999999999999998e-13
CS_1180 NS_1180 0 9.9999999999999998e-13
RS_1179 NS_1179 0 1.0548793856392000e+02
RS_1180 NS_1180 0 1.0548793856392000e+02
GL_1179 0 NS_1179 NS_1180 0 1.6750370916002649e-01
GL_1180 0 NS_1180 NS_1179 0 -1.6750370916002649e-01
GS_1179_11 0 NS_1179 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1181/1182
CS_1181 NS_1181 0 9.9999999999999998e-13
CS_1182 NS_1182 0 9.9999999999999998e-13
RS_1181 NS_1181 0 1.0753754351502513e+02
RS_1182 NS_1182 0 1.0753754351502513e+02
GL_1181 0 NS_1181 NS_1182 0 1.5942172238060490e-01
GL_1182 0 NS_1182 NS_1181 0 -1.5942172238060490e-01
GS_1181_11 0 NS_1181 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1183/1184
CS_1183 NS_1183 0 9.9999999999999998e-13
CS_1184 NS_1184 0 9.9999999999999998e-13
RS_1183 NS_1183 0 8.6961097797504721e+01
RS_1184 NS_1184 0 8.6961097797504721e+01
GL_1183 0 NS_1183 NS_1184 0 1.5553892891442009e-01
GL_1184 0 NS_1184 NS_1183 0 -1.5553892891442009e-01
GS_1183_11 0 NS_1183 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1185/1186
CS_1185 NS_1185 0 9.9999999999999998e-13
CS_1186 NS_1186 0 9.9999999999999998e-13
RS_1185 NS_1185 0 1.1549771364055694e+02
RS_1186 NS_1186 0 1.1549771364055692e+02
GL_1185 0 NS_1185 NS_1186 0 1.4899166019107438e-01
GL_1186 0 NS_1186 NS_1185 0 -1.4899166019107438e-01
GS_1185_11 0 NS_1185 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1187/1188
CS_1187 NS_1187 0 9.9999999999999998e-13
CS_1188 NS_1188 0 9.9999999999999998e-13
RS_1187 NS_1187 0 9.7194462506038604e+01
RS_1188 NS_1188 0 9.7194462506038604e+01
GL_1187 0 NS_1187 NS_1188 0 1.4180400817347408e-01
GL_1188 0 NS_1188 NS_1187 0 -1.4180400817347408e-01
GS_1187_11 0 NS_1187 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1189/1190
CS_1189 NS_1189 0 9.9999999999999998e-13
CS_1190 NS_1190 0 9.9999999999999998e-13
RS_1189 NS_1189 0 1.0682825030924828e+02
RS_1190 NS_1190 0 1.0682825030924828e+02
GL_1189 0 NS_1189 NS_1190 0 1.3872377519751058e-01
GL_1190 0 NS_1190 NS_1189 0 -1.3872377519751058e-01
GS_1189_11 0 NS_1189 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1191/1192
CS_1191 NS_1191 0 9.9999999999999998e-13
CS_1192 NS_1192 0 9.9999999999999998e-13
RS_1191 NS_1191 0 1.2559585119344567e+02
RS_1192 NS_1192 0 1.2559585119344568e+02
GL_1191 0 NS_1191 NS_1192 0 1.3097721803321302e-01
GL_1192 0 NS_1192 NS_1191 0 -1.3097721803321302e-01
GS_1191_11 0 NS_1191 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1193/1194
CS_1193 NS_1193 0 9.9999999999999998e-13
CS_1194 NS_1194 0 9.9999999999999998e-13
RS_1193 NS_1193 0 1.0417660462554996e+02
RS_1194 NS_1194 0 1.0417660462554996e+02
GL_1193 0 NS_1193 NS_1194 0 1.2625832867930367e-01
GL_1194 0 NS_1194 NS_1193 0 -1.2625832867930367e-01
GS_1193_11 0 NS_1193 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1195/1196
CS_1195 NS_1195 0 9.9999999999999998e-13
CS_1196 NS_1196 0 9.9999999999999998e-13
RS_1195 NS_1195 0 1.3317333532177352e+02
RS_1196 NS_1196 0 1.3317333532177352e+02
GL_1195 0 NS_1195 NS_1196 0 1.2123672752714061e-01
GL_1196 0 NS_1196 NS_1195 0 -1.2123672752714061e-01
GS_1195_11 0 NS_1195 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1197/1198
CS_1197 NS_1197 0 9.9999999999999998e-13
CS_1198 NS_1198 0 9.9999999999999998e-13
RS_1197 NS_1197 0 1.2967831681616519e+02
RS_1198 NS_1198 0 1.2967831681616519e+02
GL_1197 0 NS_1197 NS_1198 0 1.1651127865768855e-01
GL_1198 0 NS_1198 NS_1197 0 -1.1651127865768855e-01
GS_1197_11 0 NS_1197 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1199/1200
CS_1199 NS_1199 0 9.9999999999999998e-13
CS_1200 NS_1200 0 9.9999999999999998e-13
RS_1199 NS_1199 0 1.2999764374401394e+02
RS_1200 NS_1200 0 1.2999764374401394e+02
GL_1199 0 NS_1199 NS_1200 0 1.1100247696987056e-01
GL_1200 0 NS_1200 NS_1199 0 -1.1100247696987056e-01
GS_1199_11 0 NS_1199 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1201/1202
CS_1201 NS_1201 0 9.9999999999999998e-13
CS_1202 NS_1202 0 9.9999999999999998e-13
RS_1201 NS_1201 0 1.2458814074636419e+02
RS_1202 NS_1202 0 1.2458814074636419e+02
GL_1201 0 NS_1201 NS_1202 0 1.0660000212580591e-01
GL_1202 0 NS_1202 NS_1201 0 -1.0660000212580591e-01
GS_1201_11 0 NS_1201 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1203/1204
CS_1203 NS_1203 0 9.9999999999999998e-13
CS_1204 NS_1204 0 9.9999999999999998e-13
RS_1203 NS_1203 0 1.4677191614557748e+02
RS_1204 NS_1204 0 1.4677191614557748e+02
GL_1203 0 NS_1203 NS_1204 0 1.0224733343325158e-01
GL_1204 0 NS_1204 NS_1203 0 -1.0224733343325158e-01
GS_1203_11 0 NS_1203 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1205/1206
CS_1205 NS_1205 0 9.9999999999999998e-13
CS_1206 NS_1206 0 9.9999999999999998e-13
RS_1205 NS_1205 0 1.3445989223131798e+02
RS_1206 NS_1206 0 1.3445989223131798e+02
GL_1205 0 NS_1205 NS_1206 0 9.8177836948086503e-02
GL_1206 0 NS_1206 NS_1205 0 -9.8177836948086503e-02
GS_1205_11 0 NS_1205 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1207/1208
CS_1207 NS_1207 0 9.9999999999999998e-13
CS_1208 NS_1208 0 9.9999999999999998e-13
RS_1207 NS_1207 0 1.3187119040723775e+02
RS_1208 NS_1208 0 1.3187119040723772e+02
GL_1207 0 NS_1207 NS_1208 0 9.2640196004122682e-02
GL_1208 0 NS_1208 NS_1207 0 -9.2640196004122682e-02
GS_1207_11 0 NS_1207 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1209/1210
CS_1209 NS_1209 0 9.9999999999999998e-13
CS_1210 NS_1210 0 9.9999999999999998e-13
RS_1209 NS_1209 0 1.2288401421230557e+02
RS_1210 NS_1210 0 1.2288401421230557e+02
GL_1209 0 NS_1209 NS_1210 0 8.8704723748248199e-02
GL_1210 0 NS_1210 NS_1209 0 -8.8704723748248199e-02
GS_1209_11 0 NS_1209 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1211/1212
CS_1211 NS_1211 0 9.9999999999999998e-13
CS_1212 NS_1212 0 9.9999999999999998e-13
RS_1211 NS_1211 0 1.4123955654153085e+02
RS_1212 NS_1212 0 1.4123955654153082e+02
GL_1211 0 NS_1211 NS_1212 0 8.4112474498892476e-02
GL_1212 0 NS_1212 NS_1211 0 -8.4112474498892476e-02
GS_1211_11 0 NS_1211 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1213/1214
CS_1213 NS_1213 0 9.9999999999999998e-13
CS_1214 NS_1214 0 9.9999999999999998e-13
RS_1213 NS_1213 0 1.2539447312269779e+02
RS_1214 NS_1214 0 1.2539447312269778e+02
GL_1213 0 NS_1213 NS_1214 0 8.0007658848305588e-02
GL_1214 0 NS_1214 NS_1213 0 -8.0007658848305588e-02
GS_1213_11 0 NS_1213 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1215/1216
CS_1215 NS_1215 0 9.9999999999999998e-13
CS_1216 NS_1216 0 9.9999999999999998e-13
RS_1215 NS_1215 0 1.3219601779966965e+02
RS_1216 NS_1216 0 1.3219601779966968e+02
GL_1215 0 NS_1215 NS_1216 0 7.4373183806052026e-02
GL_1216 0 NS_1216 NS_1215 0 -7.4373183806052026e-02
GS_1215_11 0 NS_1215 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1217/1218
CS_1217 NS_1217 0 9.9999999999999998e-13
CS_1218 NS_1218 0 9.9999999999999998e-13
RS_1217 NS_1217 0 1.1951371640958898e+02
RS_1218 NS_1218 0 1.1951371640958898e+02
GL_1217 0 NS_1217 NS_1218 0 7.1003860961129844e-02
GL_1218 0 NS_1218 NS_1217 0 -7.1003860961129844e-02
GS_1217_11 0 NS_1217 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1219/1220
CS_1219 NS_1219 0 9.9999999999999998e-13
CS_1220 NS_1220 0 9.9999999999999998e-13
RS_1219 NS_1219 0 1.3491941875045018e+02
RS_1220 NS_1220 0 1.3491941875045018e+02
GL_1219 0 NS_1219 NS_1220 0 6.5922080709048564e-02
GL_1220 0 NS_1220 NS_1219 0 -6.5922080709048564e-02
GS_1219_11 0 NS_1219 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1221/1222
CS_1221 NS_1221 0 9.9999999999999998e-13
CS_1222 NS_1222 0 9.9999999999999998e-13
RS_1221 NS_1221 0 1.2290405859347165e+02
RS_1222 NS_1222 0 1.2290405859347166e+02
GL_1221 0 NS_1221 NS_1222 0 6.2340152915784278e-02
GL_1222 0 NS_1222 NS_1221 0 -6.2340152915784278e-02
GS_1221_11 0 NS_1221 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1223/1224
CS_1223 NS_1223 0 9.9999999999999998e-13
CS_1224 NS_1224 0 9.9999999999999998e-13
RS_1223 NS_1223 0 1.3258923845358959e+02
RS_1224 NS_1224 0 1.3258923845358959e+02
GL_1223 0 NS_1223 NS_1224 0 5.6431081088718790e-02
GL_1224 0 NS_1224 NS_1223 0 -5.6431081088718790e-02
GS_1223_11 0 NS_1223 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1225/1226
CS_1225 NS_1225 0 9.9999999999999998e-13
CS_1226 NS_1226 0 9.9999999999999998e-13
RS_1225 NS_1225 0 1.0026704639246873e+02
RS_1226 NS_1226 0 1.0026704639246873e+02
GL_1225 0 NS_1225 NS_1226 0 3.5068885856298401e-02
GL_1226 0 NS_1226 NS_1225 0 -3.5068885856298401e-02
GS_1225_11 0 NS_1225 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1227/1228
CS_1227 NS_1227 0 9.9999999999999998e-13
CS_1228 NS_1228 0 9.9999999999999998e-13
RS_1227 NS_1227 0 1.2740726499710033e+02
RS_1228 NS_1228 0 1.2740726499710034e+02
GL_1227 0 NS_1227 NS_1228 0 5.3740629014256171e-02
GL_1228 0 NS_1228 NS_1227 0 -5.3740629014256171e-02
GS_1227_11 0 NS_1227 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1229/1230
CS_1229 NS_1229 0 9.9999999999999998e-13
CS_1230 NS_1230 0 9.9999999999999998e-13
RS_1229 NS_1229 0 2.3804688106534087e+02
RS_1230 NS_1230 0 2.3804688106534090e+02
GL_1229 0 NS_1229 NS_1230 0 5.1425903265699464e-02
GL_1230 0 NS_1230 NS_1229 0 -5.1425903265699464e-02
GS_1229_11 0 NS_1229 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1231/1232
CS_1231 NS_1231 0 9.9999999999999998e-13
CS_1232 NS_1232 0 9.9999999999999998e-13
RS_1231 NS_1231 0 1.3728807739915800e+02
RS_1232 NS_1232 0 1.3728807739915803e+02
GL_1231 0 NS_1231 NS_1232 0 4.8031392820534764e-02
GL_1232 0 NS_1232 NS_1231 0 -4.8031392820534764e-02
GS_1231_11 0 NS_1231 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1233/1234
CS_1233 NS_1233 0 9.9999999999999998e-13
CS_1234 NS_1234 0 9.9999999999999998e-13
RS_1233 NS_1233 0 1.3499477893747948e+02
RS_1234 NS_1234 0 1.3499477893747945e+02
GL_1233 0 NS_1233 NS_1234 0 4.4453170742682194e-02
GL_1234 0 NS_1234 NS_1233 0 -4.4453170742682194e-02
GS_1233_11 0 NS_1233 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1235/1236
CS_1235 NS_1235 0 9.9999999999999998e-13
CS_1236 NS_1236 0 9.9999999999999998e-13
RS_1235 NS_1235 0 1.4121821834962651e+02
RS_1236 NS_1236 0 1.4121821834962651e+02
GL_1235 0 NS_1235 NS_1236 0 3.8464469217755697e-02
GL_1236 0 NS_1236 NS_1235 0 -3.8464469217755697e-02
GS_1235_11 0 NS_1235 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1237/1238
CS_1237 NS_1237 0 9.9999999999999998e-13
CS_1238 NS_1238 0 9.9999999999999998e-13
RS_1237 NS_1237 0 1.3946471282741149e+02
RS_1238 NS_1238 0 1.3946471282741149e+02
GL_1237 0 NS_1237 NS_1238 0 3.5678935079258622e-02
GL_1238 0 NS_1238 NS_1237 0 -3.5678935079258622e-02
GS_1237_11 0 NS_1237 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1239/1240
CS_1239 NS_1239 0 9.9999999999999998e-13
CS_1240 NS_1240 0 9.9999999999999998e-13
RS_1239 NS_1239 0 1.5530211191942624e+02
RS_1240 NS_1240 0 1.5530211191942627e+02
GL_1239 0 NS_1239 NS_1240 0 2.6209890345437525e-02
GL_1240 0 NS_1240 NS_1239 0 -2.6209890345437525e-02
GS_1239_11 0 NS_1239 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1241/1242
CS_1241 NS_1241 0 9.9999999999999998e-13
CS_1242 NS_1242 0 9.9999999999999998e-13
RS_1241 NS_1241 0 1.4887428879582419e+02
RS_1242 NS_1242 0 1.4887428879582419e+02
GL_1241 0 NS_1241 NS_1242 0 3.0330575323949095e-02
GL_1242 0 NS_1242 NS_1241 0 -3.0330575323949095e-02
GS_1241_11 0 NS_1241 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1243/1244
CS_1243 NS_1243 0 9.9999999999999998e-13
CS_1244 NS_1244 0 9.9999999999999998e-13
RS_1243 NS_1243 0 1.5087532095170570e+02
RS_1244 NS_1244 0 1.5087532095170570e+02
GL_1243 0 NS_1243 NS_1244 0 2.0034138441714564e-02
GL_1244 0 NS_1244 NS_1243 0 -2.0034138441714564e-02
GS_1243_11 0 NS_1243 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1245/1246
CS_1245 NS_1245 0 9.9999999999999998e-13
CS_1246 NS_1246 0 9.9999999999999998e-13
RS_1245 NS_1245 0 1.4763793449752018e+02
RS_1246 NS_1246 0 1.4763793449752018e+02
GL_1245 0 NS_1245 NS_1246 0 1.7017170579416537e-02
GL_1246 0 NS_1246 NS_1245 0 -1.7017170579416537e-02
GS_1245_11 0 NS_1245 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1247/1248
CS_1247 NS_1247 0 9.9999999999999998e-13
CS_1248 NS_1248 0 9.9999999999999998e-13
RS_1247 NS_1247 0 1.6285515224442304e+02
RS_1248 NS_1248 0 1.6285515224442304e+02
GL_1247 0 NS_1247 NS_1248 0 1.0897027002452746e-02
GL_1248 0 NS_1248 NS_1247 0 -1.0897027002452746e-02
GS_1247_11 0 NS_1247 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1249/1250
CS_1249 NS_1249 0 9.9999999999999998e-13
CS_1250 NS_1250 0 9.9999999999999998e-13
RS_1249 NS_1249 0 1.7239534388116820e+02
RS_1250 NS_1250 0 1.7239534388116820e+02
GL_1249 0 NS_1249 NS_1250 0 6.1589693699488982e-03
GL_1250 0 NS_1250 NS_1249 0 -6.1589693699488982e-03
GS_1249_11 0 NS_1249 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1251/1252
CS_1251 NS_1251 0 9.9999999999999998e-13
CS_1252 NS_1252 0 9.9999999999999998e-13
RS_1251 NS_1251 0 5.9928710578594173e+03
RS_1252 NS_1252 0 5.9928710578594173e+03
GL_1251 0 NS_1251 NS_1252 0 1.7541178006601681e-03
GL_1252 0 NS_1252 NS_1251 0 -1.7541178006601681e-03
GS_1251_11 0 NS_1251 NA_11 0 4.4027142044246531e-01
*
* Complex pair n. 1253/1254
CS_1253 NS_1253 0 9.9999999999999998e-13
CS_1254 NS_1254 0 9.9999999999999998e-13
RS_1253 NS_1253 0 8.0762087901330699e+02
RS_1254 NS_1254 0 8.0762087901330688e+02
GL_1253 0 NS_1253 NS_1254 0 1.7295489372816217e-03
GL_1254 0 NS_1254 NS_1253 0 -1.7295489372816217e-03
GS_1253_11 0 NS_1253 NA_11 0 4.4027142044246531e-01
*
* Real pole n. 1255
CS_1255 NS_1255 0 9.9999999999999998e-13
RS_1255 NS_1255 0 1.2857601077426406e+01
GS_1255_12 0 NS_1255 NA_12 0 4.4027142044246531e-01
*
* Real pole n. 1256
CS_1256 NS_1256 0 9.9999999999999998e-13
RS_1256 NS_1256 0 1.7282831464635029e+02
GS_1256_12 0 NS_1256 NA_12 0 4.4027142044246531e-01
*
* Real pole n. 1257
CS_1257 NS_1257 0 9.9999999999999998e-13
RS_1257 NS_1257 0 5.5743135126264733e+03
GS_1257_12 0 NS_1257 NA_12 0 4.4027142044246531e-01
*
* Real pole n. 1258
CS_1258 NS_1258 0 9.9999999999999998e-13
RS_1258 NS_1258 0 1.3594126013480764e+03
GS_1258_12 0 NS_1258 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1259/1260
CS_1259 NS_1259 0 9.9999999999999998e-13
CS_1260 NS_1260 0 9.9999999999999998e-13
RS_1259 NS_1259 0 1.7904812183888848e+02
RS_1260 NS_1260 0 1.7904812183888848e+02
GL_1259 0 NS_1259 NS_1260 0 2.6007898045516648e-01
GL_1260 0 NS_1260 NS_1259 0 -2.6007898045516648e-01
GS_1259_12 0 NS_1259 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1261/1262
CS_1261 NS_1261 0 9.9999999999999998e-13
CS_1262 NS_1262 0 9.9999999999999998e-13
RS_1261 NS_1261 0 1.2615541320340381e+02
RS_1262 NS_1262 0 1.2615541320340381e+02
GL_1261 0 NS_1261 NS_1262 0 2.5243684762014923e-01
GL_1262 0 NS_1262 NS_1261 0 -2.5243684762014923e-01
GS_1261_12 0 NS_1261 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1263/1264
CS_1263 NS_1263 0 9.9999999999999998e-13
CS_1264 NS_1264 0 9.9999999999999998e-13
RS_1263 NS_1263 0 1.0219948841586964e+02
RS_1264 NS_1264 0 1.0219948841586965e+02
GL_1263 0 NS_1263 NS_1264 0 2.4690226903121384e-01
GL_1264 0 NS_1264 NS_1263 0 -2.4690226903121384e-01
GS_1263_12 0 NS_1263 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1265/1266
CS_1265 NS_1265 0 9.9999999999999998e-13
CS_1266 NS_1266 0 9.9999999999999998e-13
RS_1265 NS_1265 0 1.1002436853144543e+02
RS_1266 NS_1266 0 1.1002436853144542e+02
GL_1265 0 NS_1265 NS_1266 0 2.4293768067729948e-01
GL_1266 0 NS_1266 NS_1265 0 -2.4293768067729948e-01
GS_1265_12 0 NS_1265 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1267/1268
CS_1267 NS_1267 0 9.9999999999999998e-13
CS_1268 NS_1268 0 9.9999999999999998e-13
RS_1267 NS_1267 0 1.0553430908077024e+02
RS_1268 NS_1268 0 1.0553430908077026e+02
GL_1267 0 NS_1267 NS_1268 0 2.3600513224442521e-01
GL_1268 0 NS_1268 NS_1267 0 -2.3600513224442521e-01
GS_1267_12 0 NS_1267 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1269/1270
CS_1269 NS_1269 0 9.9999999999999998e-13
CS_1270 NS_1270 0 9.9999999999999998e-13
RS_1269 NS_1269 0 1.0759915098440327e+02
RS_1270 NS_1270 0 1.0759915098440327e+02
GL_1269 0 NS_1269 NS_1270 0 2.3090539914362113e-01
GL_1270 0 NS_1270 NS_1269 0 -2.3090539914362113e-01
GS_1269_12 0 NS_1269 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1271/1272
CS_1271 NS_1271 0 9.9999999999999998e-13
CS_1272 NS_1272 0 9.9999999999999998e-13
RS_1271 NS_1271 0 1.3295415758774385e+02
RS_1272 NS_1272 0 1.3295415758774385e+02
GL_1271 0 NS_1271 NS_1272 0 2.3030066292345727e-01
GL_1272 0 NS_1272 NS_1271 0 -2.3030066292345727e-01
GS_1271_12 0 NS_1271 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1273/1274
CS_1273 NS_1273 0 9.9999999999999998e-13
CS_1274 NS_1274 0 9.9999999999999998e-13
RS_1273 NS_1273 0 1.1432186998941940e+02
RS_1274 NS_1274 0 1.1432186998941938e+02
GL_1273 0 NS_1273 NS_1274 0 2.2451058023508991e-01
GL_1274 0 NS_1274 NS_1273 0 -2.2451058023508991e-01
GS_1273_12 0 NS_1273 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1275/1276
CS_1275 NS_1275 0 9.9999999999999998e-13
CS_1276 NS_1276 0 9.9999999999999998e-13
RS_1275 NS_1275 0 9.0812703249943667e+01
RS_1276 NS_1276 0 9.0812703249943652e+01
GL_1275 0 NS_1275 NS_1276 0 2.1702628900531115e-01
GL_1276 0 NS_1276 NS_1275 0 -2.1702628900531115e-01
GS_1275_12 0 NS_1275 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1277/1278
CS_1277 NS_1277 0 9.9999999999999998e-13
CS_1278 NS_1278 0 9.9999999999999998e-13
RS_1277 NS_1277 0 9.5643803662064585e+01
RS_1278 NS_1278 0 9.5643803662064585e+01
GL_1277 0 NS_1277 NS_1278 0 2.1448200383207913e-01
GL_1278 0 NS_1278 NS_1277 0 -2.1448200383207913e-01
GS_1277_12 0 NS_1277 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1279/1280
CS_1279 NS_1279 0 9.9999999999999998e-13
CS_1280 NS_1280 0 9.9999999999999998e-13
RS_1279 NS_1279 0 1.0631957479149644e+02
RS_1280 NS_1280 0 1.0631957479149644e+02
GL_1279 0 NS_1279 NS_1280 0 2.0655001587884311e-01
GL_1280 0 NS_1280 NS_1279 0 -2.0655001587884311e-01
GS_1279_12 0 NS_1279 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1281/1282
CS_1281 NS_1281 0 9.9999999999999998e-13
CS_1282 NS_1282 0 9.9999999999999998e-13
RS_1281 NS_1281 0 7.9907264643295406e+01
RS_1282 NS_1282 0 7.9907264643295420e+01
GL_1281 0 NS_1281 NS_1282 0 2.0133773147328893e-01
GL_1282 0 NS_1282 NS_1281 0 -2.0133773147328893e-01
GS_1281_12 0 NS_1281 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1283/1284
CS_1283 NS_1283 0 9.9999999999999998e-13
CS_1284 NS_1284 0 9.9999999999999998e-13
RS_1283 NS_1283 0 1.0625506887893997e+02
RS_1284 NS_1284 0 1.0625506887893997e+02
GL_1283 0 NS_1283 NS_1284 0 1.9628877333023340e-01
GL_1284 0 NS_1284 NS_1283 0 -1.9628877333023340e-01
GS_1283_12 0 NS_1283 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1285/1286
CS_1285 NS_1285 0 9.9999999999999998e-13
CS_1286 NS_1286 0 9.9999999999999998e-13
RS_1285 NS_1285 0 9.6115312638592201e+01
RS_1286 NS_1286 0 9.6115312638592201e+01
GL_1285 0 NS_1285 NS_1286 0 1.8794816712418483e-01
GL_1286 0 NS_1286 NS_1285 0 -1.8794816712418483e-01
GS_1285_12 0 NS_1285 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1287/1288
CS_1287 NS_1287 0 9.9999999999999998e-13
CS_1288 NS_1288 0 9.9999999999999998e-13
RS_1287 NS_1287 0 8.5212696574118169e+01
RS_1288 NS_1288 0 8.5212696574118169e+01
GL_1287 0 NS_1287 NS_1288 0 1.8572140881490298e-01
GL_1288 0 NS_1288 NS_1287 0 -1.8572140881490298e-01
GS_1287_12 0 NS_1287 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1289/1290
CS_1289 NS_1289 0 9.9999999999999998e-13
CS_1290 NS_1290 0 9.9999999999999998e-13
RS_1289 NS_1289 0 1.0905026103375434e+02
RS_1290 NS_1290 0 1.0905026103375432e+02
GL_1289 0 NS_1289 NS_1290 0 1.7785621200284463e-01
GL_1290 0 NS_1290 NS_1289 0 -1.7785621200284463e-01
GS_1289_12 0 NS_1289 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1291/1292
CS_1291 NS_1291 0 9.9999999999999998e-13
CS_1292 NS_1292 0 9.9999999999999998e-13
RS_1291 NS_1291 0 8.3024437910787526e+01
RS_1292 NS_1292 0 8.3024437910787526e+01
GL_1291 0 NS_1291 NS_1292 0 1.7164509875911016e-01
GL_1292 0 NS_1292 NS_1291 0 -1.7164509875911016e-01
GS_1291_12 0 NS_1291 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1293/1294
CS_1293 NS_1293 0 9.9999999999999998e-13
CS_1294 NS_1294 0 9.9999999999999998e-13
RS_1293 NS_1293 0 1.0548793856392000e+02
RS_1294 NS_1294 0 1.0548793856392000e+02
GL_1293 0 NS_1293 NS_1294 0 1.6750370916002649e-01
GL_1294 0 NS_1294 NS_1293 0 -1.6750370916002649e-01
GS_1293_12 0 NS_1293 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1295/1296
CS_1295 NS_1295 0 9.9999999999999998e-13
CS_1296 NS_1296 0 9.9999999999999998e-13
RS_1295 NS_1295 0 1.0753754351502513e+02
RS_1296 NS_1296 0 1.0753754351502513e+02
GL_1295 0 NS_1295 NS_1296 0 1.5942172238060490e-01
GL_1296 0 NS_1296 NS_1295 0 -1.5942172238060490e-01
GS_1295_12 0 NS_1295 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1297/1298
CS_1297 NS_1297 0 9.9999999999999998e-13
CS_1298 NS_1298 0 9.9999999999999998e-13
RS_1297 NS_1297 0 8.6961097797504721e+01
RS_1298 NS_1298 0 8.6961097797504721e+01
GL_1297 0 NS_1297 NS_1298 0 1.5553892891442009e-01
GL_1298 0 NS_1298 NS_1297 0 -1.5553892891442009e-01
GS_1297_12 0 NS_1297 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1299/1300
CS_1299 NS_1299 0 9.9999999999999998e-13
CS_1300 NS_1300 0 9.9999999999999998e-13
RS_1299 NS_1299 0 1.1549771364055694e+02
RS_1300 NS_1300 0 1.1549771364055692e+02
GL_1299 0 NS_1299 NS_1300 0 1.4899166019107438e-01
GL_1300 0 NS_1300 NS_1299 0 -1.4899166019107438e-01
GS_1299_12 0 NS_1299 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1301/1302
CS_1301 NS_1301 0 9.9999999999999998e-13
CS_1302 NS_1302 0 9.9999999999999998e-13
RS_1301 NS_1301 0 9.7194462506038604e+01
RS_1302 NS_1302 0 9.7194462506038604e+01
GL_1301 0 NS_1301 NS_1302 0 1.4180400817347408e-01
GL_1302 0 NS_1302 NS_1301 0 -1.4180400817347408e-01
GS_1301_12 0 NS_1301 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1303/1304
CS_1303 NS_1303 0 9.9999999999999998e-13
CS_1304 NS_1304 0 9.9999999999999998e-13
RS_1303 NS_1303 0 1.0682825030924828e+02
RS_1304 NS_1304 0 1.0682825030924828e+02
GL_1303 0 NS_1303 NS_1304 0 1.3872377519751058e-01
GL_1304 0 NS_1304 NS_1303 0 -1.3872377519751058e-01
GS_1303_12 0 NS_1303 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1305/1306
CS_1305 NS_1305 0 9.9999999999999998e-13
CS_1306 NS_1306 0 9.9999999999999998e-13
RS_1305 NS_1305 0 1.2559585119344567e+02
RS_1306 NS_1306 0 1.2559585119344568e+02
GL_1305 0 NS_1305 NS_1306 0 1.3097721803321302e-01
GL_1306 0 NS_1306 NS_1305 0 -1.3097721803321302e-01
GS_1305_12 0 NS_1305 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1307/1308
CS_1307 NS_1307 0 9.9999999999999998e-13
CS_1308 NS_1308 0 9.9999999999999998e-13
RS_1307 NS_1307 0 1.0417660462554996e+02
RS_1308 NS_1308 0 1.0417660462554996e+02
GL_1307 0 NS_1307 NS_1308 0 1.2625832867930367e-01
GL_1308 0 NS_1308 NS_1307 0 -1.2625832867930367e-01
GS_1307_12 0 NS_1307 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1309/1310
CS_1309 NS_1309 0 9.9999999999999998e-13
CS_1310 NS_1310 0 9.9999999999999998e-13
RS_1309 NS_1309 0 1.3317333532177352e+02
RS_1310 NS_1310 0 1.3317333532177352e+02
GL_1309 0 NS_1309 NS_1310 0 1.2123672752714061e-01
GL_1310 0 NS_1310 NS_1309 0 -1.2123672752714061e-01
GS_1309_12 0 NS_1309 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1311/1312
CS_1311 NS_1311 0 9.9999999999999998e-13
CS_1312 NS_1312 0 9.9999999999999998e-13
RS_1311 NS_1311 0 1.2967831681616519e+02
RS_1312 NS_1312 0 1.2967831681616519e+02
GL_1311 0 NS_1311 NS_1312 0 1.1651127865768855e-01
GL_1312 0 NS_1312 NS_1311 0 -1.1651127865768855e-01
GS_1311_12 0 NS_1311 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1313/1314
CS_1313 NS_1313 0 9.9999999999999998e-13
CS_1314 NS_1314 0 9.9999999999999998e-13
RS_1313 NS_1313 0 1.2999764374401394e+02
RS_1314 NS_1314 0 1.2999764374401394e+02
GL_1313 0 NS_1313 NS_1314 0 1.1100247696987056e-01
GL_1314 0 NS_1314 NS_1313 0 -1.1100247696987056e-01
GS_1313_12 0 NS_1313 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1315/1316
CS_1315 NS_1315 0 9.9999999999999998e-13
CS_1316 NS_1316 0 9.9999999999999998e-13
RS_1315 NS_1315 0 1.2458814074636419e+02
RS_1316 NS_1316 0 1.2458814074636419e+02
GL_1315 0 NS_1315 NS_1316 0 1.0660000212580591e-01
GL_1316 0 NS_1316 NS_1315 0 -1.0660000212580591e-01
GS_1315_12 0 NS_1315 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1317/1318
CS_1317 NS_1317 0 9.9999999999999998e-13
CS_1318 NS_1318 0 9.9999999999999998e-13
RS_1317 NS_1317 0 1.4677191614557748e+02
RS_1318 NS_1318 0 1.4677191614557748e+02
GL_1317 0 NS_1317 NS_1318 0 1.0224733343325158e-01
GL_1318 0 NS_1318 NS_1317 0 -1.0224733343325158e-01
GS_1317_12 0 NS_1317 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1319/1320
CS_1319 NS_1319 0 9.9999999999999998e-13
CS_1320 NS_1320 0 9.9999999999999998e-13
RS_1319 NS_1319 0 1.3445989223131798e+02
RS_1320 NS_1320 0 1.3445989223131798e+02
GL_1319 0 NS_1319 NS_1320 0 9.8177836948086503e-02
GL_1320 0 NS_1320 NS_1319 0 -9.8177836948086503e-02
GS_1319_12 0 NS_1319 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1321/1322
CS_1321 NS_1321 0 9.9999999999999998e-13
CS_1322 NS_1322 0 9.9999999999999998e-13
RS_1321 NS_1321 0 1.3187119040723775e+02
RS_1322 NS_1322 0 1.3187119040723772e+02
GL_1321 0 NS_1321 NS_1322 0 9.2640196004122682e-02
GL_1322 0 NS_1322 NS_1321 0 -9.2640196004122682e-02
GS_1321_12 0 NS_1321 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1323/1324
CS_1323 NS_1323 0 9.9999999999999998e-13
CS_1324 NS_1324 0 9.9999999999999998e-13
RS_1323 NS_1323 0 1.2288401421230557e+02
RS_1324 NS_1324 0 1.2288401421230557e+02
GL_1323 0 NS_1323 NS_1324 0 8.8704723748248199e-02
GL_1324 0 NS_1324 NS_1323 0 -8.8704723748248199e-02
GS_1323_12 0 NS_1323 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1325/1326
CS_1325 NS_1325 0 9.9999999999999998e-13
CS_1326 NS_1326 0 9.9999999999999998e-13
RS_1325 NS_1325 0 1.4123955654153085e+02
RS_1326 NS_1326 0 1.4123955654153082e+02
GL_1325 0 NS_1325 NS_1326 0 8.4112474498892476e-02
GL_1326 0 NS_1326 NS_1325 0 -8.4112474498892476e-02
GS_1325_12 0 NS_1325 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1327/1328
CS_1327 NS_1327 0 9.9999999999999998e-13
CS_1328 NS_1328 0 9.9999999999999998e-13
RS_1327 NS_1327 0 1.2539447312269779e+02
RS_1328 NS_1328 0 1.2539447312269778e+02
GL_1327 0 NS_1327 NS_1328 0 8.0007658848305588e-02
GL_1328 0 NS_1328 NS_1327 0 -8.0007658848305588e-02
GS_1327_12 0 NS_1327 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1329/1330
CS_1329 NS_1329 0 9.9999999999999998e-13
CS_1330 NS_1330 0 9.9999999999999998e-13
RS_1329 NS_1329 0 1.3219601779966965e+02
RS_1330 NS_1330 0 1.3219601779966968e+02
GL_1329 0 NS_1329 NS_1330 0 7.4373183806052026e-02
GL_1330 0 NS_1330 NS_1329 0 -7.4373183806052026e-02
GS_1329_12 0 NS_1329 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1331/1332
CS_1331 NS_1331 0 9.9999999999999998e-13
CS_1332 NS_1332 0 9.9999999999999998e-13
RS_1331 NS_1331 0 1.1951371640958898e+02
RS_1332 NS_1332 0 1.1951371640958898e+02
GL_1331 0 NS_1331 NS_1332 0 7.1003860961129844e-02
GL_1332 0 NS_1332 NS_1331 0 -7.1003860961129844e-02
GS_1331_12 0 NS_1331 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1333/1334
CS_1333 NS_1333 0 9.9999999999999998e-13
CS_1334 NS_1334 0 9.9999999999999998e-13
RS_1333 NS_1333 0 1.3491941875045018e+02
RS_1334 NS_1334 0 1.3491941875045018e+02
GL_1333 0 NS_1333 NS_1334 0 6.5922080709048564e-02
GL_1334 0 NS_1334 NS_1333 0 -6.5922080709048564e-02
GS_1333_12 0 NS_1333 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1335/1336
CS_1335 NS_1335 0 9.9999999999999998e-13
CS_1336 NS_1336 0 9.9999999999999998e-13
RS_1335 NS_1335 0 1.2290405859347165e+02
RS_1336 NS_1336 0 1.2290405859347166e+02
GL_1335 0 NS_1335 NS_1336 0 6.2340152915784278e-02
GL_1336 0 NS_1336 NS_1335 0 -6.2340152915784278e-02
GS_1335_12 0 NS_1335 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1337/1338
CS_1337 NS_1337 0 9.9999999999999998e-13
CS_1338 NS_1338 0 9.9999999999999998e-13
RS_1337 NS_1337 0 1.3258923845358959e+02
RS_1338 NS_1338 0 1.3258923845358959e+02
GL_1337 0 NS_1337 NS_1338 0 5.6431081088718790e-02
GL_1338 0 NS_1338 NS_1337 0 -5.6431081088718790e-02
GS_1337_12 0 NS_1337 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1339/1340
CS_1339 NS_1339 0 9.9999999999999998e-13
CS_1340 NS_1340 0 9.9999999999999998e-13
RS_1339 NS_1339 0 1.0026704639246873e+02
RS_1340 NS_1340 0 1.0026704639246873e+02
GL_1339 0 NS_1339 NS_1340 0 3.5068885856298401e-02
GL_1340 0 NS_1340 NS_1339 0 -3.5068885856298401e-02
GS_1339_12 0 NS_1339 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1341/1342
CS_1341 NS_1341 0 9.9999999999999998e-13
CS_1342 NS_1342 0 9.9999999999999998e-13
RS_1341 NS_1341 0 1.2740726499710033e+02
RS_1342 NS_1342 0 1.2740726499710034e+02
GL_1341 0 NS_1341 NS_1342 0 5.3740629014256171e-02
GL_1342 0 NS_1342 NS_1341 0 -5.3740629014256171e-02
GS_1341_12 0 NS_1341 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1343/1344
CS_1343 NS_1343 0 9.9999999999999998e-13
CS_1344 NS_1344 0 9.9999999999999998e-13
RS_1343 NS_1343 0 2.3804688106534087e+02
RS_1344 NS_1344 0 2.3804688106534090e+02
GL_1343 0 NS_1343 NS_1344 0 5.1425903265699464e-02
GL_1344 0 NS_1344 NS_1343 0 -5.1425903265699464e-02
GS_1343_12 0 NS_1343 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1345/1346
CS_1345 NS_1345 0 9.9999999999999998e-13
CS_1346 NS_1346 0 9.9999999999999998e-13
RS_1345 NS_1345 0 1.3728807739915800e+02
RS_1346 NS_1346 0 1.3728807739915803e+02
GL_1345 0 NS_1345 NS_1346 0 4.8031392820534764e-02
GL_1346 0 NS_1346 NS_1345 0 -4.8031392820534764e-02
GS_1345_12 0 NS_1345 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1347/1348
CS_1347 NS_1347 0 9.9999999999999998e-13
CS_1348 NS_1348 0 9.9999999999999998e-13
RS_1347 NS_1347 0 1.3499477893747948e+02
RS_1348 NS_1348 0 1.3499477893747945e+02
GL_1347 0 NS_1347 NS_1348 0 4.4453170742682194e-02
GL_1348 0 NS_1348 NS_1347 0 -4.4453170742682194e-02
GS_1347_12 0 NS_1347 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1349/1350
CS_1349 NS_1349 0 9.9999999999999998e-13
CS_1350 NS_1350 0 9.9999999999999998e-13
RS_1349 NS_1349 0 1.4121821834962651e+02
RS_1350 NS_1350 0 1.4121821834962651e+02
GL_1349 0 NS_1349 NS_1350 0 3.8464469217755697e-02
GL_1350 0 NS_1350 NS_1349 0 -3.8464469217755697e-02
GS_1349_12 0 NS_1349 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1351/1352
CS_1351 NS_1351 0 9.9999999999999998e-13
CS_1352 NS_1352 0 9.9999999999999998e-13
RS_1351 NS_1351 0 1.3946471282741149e+02
RS_1352 NS_1352 0 1.3946471282741149e+02
GL_1351 0 NS_1351 NS_1352 0 3.5678935079258622e-02
GL_1352 0 NS_1352 NS_1351 0 -3.5678935079258622e-02
GS_1351_12 0 NS_1351 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1353/1354
CS_1353 NS_1353 0 9.9999999999999998e-13
CS_1354 NS_1354 0 9.9999999999999998e-13
RS_1353 NS_1353 0 1.5530211191942624e+02
RS_1354 NS_1354 0 1.5530211191942627e+02
GL_1353 0 NS_1353 NS_1354 0 2.6209890345437525e-02
GL_1354 0 NS_1354 NS_1353 0 -2.6209890345437525e-02
GS_1353_12 0 NS_1353 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1355/1356
CS_1355 NS_1355 0 9.9999999999999998e-13
CS_1356 NS_1356 0 9.9999999999999998e-13
RS_1355 NS_1355 0 1.4887428879582419e+02
RS_1356 NS_1356 0 1.4887428879582419e+02
GL_1355 0 NS_1355 NS_1356 0 3.0330575323949095e-02
GL_1356 0 NS_1356 NS_1355 0 -3.0330575323949095e-02
GS_1355_12 0 NS_1355 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1357/1358
CS_1357 NS_1357 0 9.9999999999999998e-13
CS_1358 NS_1358 0 9.9999999999999998e-13
RS_1357 NS_1357 0 1.5087532095170570e+02
RS_1358 NS_1358 0 1.5087532095170570e+02
GL_1357 0 NS_1357 NS_1358 0 2.0034138441714564e-02
GL_1358 0 NS_1358 NS_1357 0 -2.0034138441714564e-02
GS_1357_12 0 NS_1357 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1359/1360
CS_1359 NS_1359 0 9.9999999999999998e-13
CS_1360 NS_1360 0 9.9999999999999998e-13
RS_1359 NS_1359 0 1.4763793449752018e+02
RS_1360 NS_1360 0 1.4763793449752018e+02
GL_1359 0 NS_1359 NS_1360 0 1.7017170579416537e-02
GL_1360 0 NS_1360 NS_1359 0 -1.7017170579416537e-02
GS_1359_12 0 NS_1359 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1361/1362
CS_1361 NS_1361 0 9.9999999999999998e-13
CS_1362 NS_1362 0 9.9999999999999998e-13
RS_1361 NS_1361 0 1.6285515224442304e+02
RS_1362 NS_1362 0 1.6285515224442304e+02
GL_1361 0 NS_1361 NS_1362 0 1.0897027002452746e-02
GL_1362 0 NS_1362 NS_1361 0 -1.0897027002452746e-02
GS_1361_12 0 NS_1361 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1363/1364
CS_1363 NS_1363 0 9.9999999999999998e-13
CS_1364 NS_1364 0 9.9999999999999998e-13
RS_1363 NS_1363 0 1.7239534388116820e+02
RS_1364 NS_1364 0 1.7239534388116820e+02
GL_1363 0 NS_1363 NS_1364 0 6.1589693699488982e-03
GL_1364 0 NS_1364 NS_1363 0 -6.1589693699488982e-03
GS_1363_12 0 NS_1363 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1365/1366
CS_1365 NS_1365 0 9.9999999999999998e-13
CS_1366 NS_1366 0 9.9999999999999998e-13
RS_1365 NS_1365 0 5.9928710578594173e+03
RS_1366 NS_1366 0 5.9928710578594173e+03
GL_1365 0 NS_1365 NS_1366 0 1.7541178006601681e-03
GL_1366 0 NS_1366 NS_1365 0 -1.7541178006601681e-03
GS_1365_12 0 NS_1365 NA_12 0 4.4027142044246531e-01
*
* Complex pair n. 1367/1368
CS_1367 NS_1367 0 9.9999999999999998e-13
CS_1368 NS_1368 0 9.9999999999999998e-13
RS_1367 NS_1367 0 8.0762087901330699e+02
RS_1368 NS_1368 0 8.0762087901330688e+02
GL_1367 0 NS_1367 NS_1368 0 1.7295489372816217e-03
GL_1368 0 NS_1368 NS_1367 0 -1.7295489372816217e-03
GS_1367_12 0 NS_1367 NA_12 0 4.4027142044246531e-01
*
******************************


.ends
*******************
* End of subcircuit
*******************
