**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 5.0000e+10 Hz
** Order: [6 4 32] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** n/a - passivity was not enforced
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_11_Module_wire_5mm_lowloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 1.2526108569063432e-01
GC_1_2 b_1 NI_1 NS_2 0 -9.7551738268519157e-03
GC_1_3 b_1 NI_1 NS_3 0 -2.1879140150518010e-05
GC_1_4 b_1 NI_1 NS_4 0 -3.7984593841402384e-06
GC_1_5 b_1 NI_1 NS_5 0 -8.0420603776076398e-03
GC_1_6 b_1 NI_1 NS_6 0 6.5371474564688615e-04
GC_1_7 b_1 NI_1 NS_7 0 -1.9771749923377080e-03
GC_1_8 b_1 NI_1 NS_8 0 1.0156944859433434e-04
GC_1_9 b_1 NI_1 NS_9 0 -1.2487317258108406e-02
GC_1_10 b_1 NI_1 NS_10 0 8.2382539291840137e-03
GC_1_11 b_1 NI_1 NS_11 0 -1.0111830234426761e-02
GC_1_12 b_1 NI_1 NS_12 0 -5.9611418424683211e-04
GC_1_13 b_1 NI_1 NS_13 0 -3.4891091292881932e-03
GC_1_14 b_1 NI_1 NS_14 0 1.6807110978405138e-02
GC_1_15 b_1 NI_1 NS_15 0 -7.7156973516644602e-03
GC_1_16 b_1 NI_1 NS_16 0 1.3269796070236673e-02
GC_1_17 b_1 NI_1 NS_17 0 -3.8876518720963598e-03
GC_1_18 b_1 NI_1 NS_18 0 6.8943385148697483e-03
GC_1_19 b_1 NI_1 NS_19 0 -2.7117302567003297e-03
GC_1_20 b_1 NI_1 NS_20 0 1.2199575250037460e-02
GC_1_21 b_1 NI_1 NS_21 0 -2.2742233491917594e-02
GC_1_22 b_1 NI_1 NS_22 0 5.9617102582374785e-03
GC_1_23 b_1 NI_1 NS_23 0 -8.4148567214239979e-04
GC_1_24 b_1 NI_1 NS_24 0 8.1300274134813182e-04
GC_1_25 b_1 NI_1 NS_25 0 -5.1564584094578177e-04
GC_1_26 b_1 NI_1 NS_26 0 -4.3051992490342449e-04
GC_1_27 b_1 NI_1 NS_27 0 -5.9275332955223228e-08
GC_1_28 b_1 NI_1 NS_28 0 -1.8756500527532273e-07
GC_1_29 b_1 NI_1 NS_29 0 -3.3579646716802352e-09
GC_1_30 b_1 NI_1 NS_30 0 5.3365681839066293e-09
GC_1_31 b_1 NI_1 NS_31 0 -7.0424920157876200e-02
GC_1_32 b_1 NI_1 NS_32 0 2.4192877757459548e-02
GC_1_33 b_1 NI_1 NS_33 0 2.2092711031652662e-05
GC_1_34 b_1 NI_1 NS_34 0 5.3186652035091707e-06
GC_1_35 b_1 NI_1 NS_35 0 1.8108338331854382e-02
GC_1_36 b_1 NI_1 NS_36 0 2.7946288947457463e-02
GC_1_37 b_1 NI_1 NS_37 0 -1.9395012070035831e-02
GC_1_38 b_1 NI_1 NS_38 0 8.3724642966768736e-03
GC_1_39 b_1 NI_1 NS_39 0 -5.8925695965379504e-03
GC_1_40 b_1 NI_1 NS_40 0 -2.2930859702124197e-02
GC_1_41 b_1 NI_1 NS_41 0 2.6387231825091097e-02
GC_1_42 b_1 NI_1 NS_42 0 -1.4337550170623494e-02
GC_1_43 b_1 NI_1 NS_43 0 3.4164772289171058e-02
GC_1_44 b_1 NI_1 NS_44 0 5.2157221280880245e-03
GC_1_45 b_1 NI_1 NS_45 0 9.5147596731506509e-03
GC_1_46 b_1 NI_1 NS_46 0 1.4168166331716017e-02
GC_1_47 b_1 NI_1 NS_47 0 -1.2626473784182198e-02
GC_1_48 b_1 NI_1 NS_48 0 1.1356489442714170e-02
GC_1_49 b_1 NI_1 NS_49 0 -1.1978297075822058e-02
GC_1_50 b_1 NI_1 NS_50 0 -1.1686204389078069e-02
GC_1_51 b_1 NI_1 NS_51 0 1.9051214451824543e-02
GC_1_52 b_1 NI_1 NS_52 0 -2.5965268339774330e-02
GC_1_53 b_1 NI_1 NS_53 0 9.0695177020609207e-04
GC_1_54 b_1 NI_1 NS_54 0 -1.0849123686524557e-03
GC_1_55 b_1 NI_1 NS_55 0 6.2679895242324316e-04
GC_1_56 b_1 NI_1 NS_56 0 3.2176426318909692e-04
GC_1_57 b_1 NI_1 NS_57 0 9.0179869225616734e-08
GC_1_58 b_1 NI_1 NS_58 0 4.0615057593027028e-07
GC_1_59 b_1 NI_1 NS_59 0 -9.1806595449948917e-09
GC_1_60 b_1 NI_1 NS_60 0 -1.8630956836277454e-08
GC_1_61 b_1 NI_1 NS_61 0 -5.5801074585759038e-04
GC_1_62 b_1 NI_1 NS_62 0 -2.9007616243774429e-03
GC_1_63 b_1 NI_1 NS_63 0 -6.1510250245751212e-06
GC_1_64 b_1 NI_1 NS_64 0 -3.8641528467974879e-07
GC_1_65 b_1 NI_1 NS_65 0 2.6869528711996630e-03
GC_1_66 b_1 NI_1 NS_66 0 -1.9871035345262055e-03
GC_1_67 b_1 NI_1 NS_67 0 -6.1985251461648553e-03
GC_1_68 b_1 NI_1 NS_68 0 1.7528631976777577e-03
GC_1_69 b_1 NI_1 NS_69 0 4.7654008991355893e-03
GC_1_70 b_1 NI_1 NS_70 0 -5.5287242487481996e-03
GC_1_71 b_1 NI_1 NS_71 0 -2.4763103518418749e-04
GC_1_72 b_1 NI_1 NS_72 0 7.2490216894756324e-03
GC_1_73 b_1 NI_1 NS_73 0 -6.3151021330544272e-03
GC_1_74 b_1 NI_1 NS_74 0 -5.0558253063660010e-03
GC_1_75 b_1 NI_1 NS_75 0 4.5028162175350956e-03
GC_1_76 b_1 NI_1 NS_76 0 -1.7122915625087667e-03
GC_1_77 b_1 NI_1 NS_77 0 -5.9096753128089067e-04
GC_1_78 b_1 NI_1 NS_78 0 6.9470776365120812e-03
GC_1_79 b_1 NI_1 NS_79 0 -3.4358105681738574e-03
GC_1_80 b_1 NI_1 NS_80 0 -3.6826697954909131e-03
GC_1_81 b_1 NI_1 NS_81 0 5.9256580380199313e-03
GC_1_82 b_1 NI_1 NS_82 0 3.9686148946459308e-04
GC_1_83 b_1 NI_1 NS_83 0 6.3856041305008845e-05
GC_1_84 b_1 NI_1 NS_84 0 8.4381967270728538e-06
GC_1_85 b_1 NI_1 NS_85 0 1.5113680855539863e-05
GC_1_86 b_1 NI_1 NS_86 0 3.9976674192848513e-05
GC_1_87 b_1 NI_1 NS_87 0 7.1156028022053443e-09
GC_1_88 b_1 NI_1 NS_88 0 -2.9351516618552961e-08
GC_1_89 b_1 NI_1 NS_89 0 -1.8855648137921119e-09
GC_1_90 b_1 NI_1 NS_90 0 -5.6002683984234213e-10
GC_1_91 b_1 NI_1 NS_91 0 1.3560957424002648e-03
GC_1_92 b_1 NI_1 NS_92 0 -1.2038969319481860e-03
GC_1_93 b_1 NI_1 NS_93 0 3.7358059729846304e-06
GC_1_94 b_1 NI_1 NS_94 0 2.8902002006203510e-07
GC_1_95 b_1 NI_1 NS_95 0 1.2295927453638333e-04
GC_1_96 b_1 NI_1 NS_96 0 8.9417218272067978e-04
GC_1_97 b_1 NI_1 NS_97 0 1.8425109579822123e-03
GC_1_98 b_1 NI_1 NS_98 0 -8.6745731587439150e-04
GC_1_99 b_1 NI_1 NS_99 0 -2.9666009049716812e-03
GC_1_100 b_1 NI_1 NS_100 0 -1.6486043793047156e-03
GC_1_101 b_1 NI_1 NS_101 0 2.2194918517918802e-03
GC_1_102 b_1 NI_1 NS_102 0 2.6689302751265239e-03
GC_1_103 b_1 NI_1 NS_103 0 -1.4401400996335413e-03
GC_1_104 b_1 NI_1 NS_104 0 -2.9129078615486347e-03
GC_1_105 b_1 NI_1 NS_105 0 1.0698829994959188e-03
GC_1_106 b_1 NI_1 NS_106 0 2.2566979184930878e-03
GC_1_107 b_1 NI_1 NS_107 0 -1.6275462029623866e-03
GC_1_108 b_1 NI_1 NS_108 0 -2.1363605820791894e-03
GC_1_109 b_1 NI_1 NS_109 0 4.2046424181054322e-04
GC_1_110 b_1 NI_1 NS_110 0 2.0118561347711372e-03
GC_1_111 b_1 NI_1 NS_111 0 2.1506913134739471e-04
GC_1_112 b_1 NI_1 NS_112 0 -2.1102665149562109e-03
GC_1_113 b_1 NI_1 NS_113 0 -4.3297326345120761e-06
GC_1_114 b_1 NI_1 NS_114 0 4.3533494645864053e-06
GC_1_115 b_1 NI_1 NS_115 0 -7.8987647927371315e-07
GC_1_116 b_1 NI_1 NS_116 0 -3.5253666127663393e-06
GC_1_117 b_1 NI_1 NS_117 0 -7.5480260267779697e-09
GC_1_118 b_1 NI_1 NS_118 0 2.2567511316039984e-08
GC_1_119 b_1 NI_1 NS_119 0 2.3359255862190867e-09
GC_1_120 b_1 NI_1 NS_120 0 1.5101864268763741e-09
GC_1_121 b_1 NI_1 NS_121 0 1.4263880551265674e-04
GC_1_122 b_1 NI_1 NS_122 0 1.2397282119280829e-06
GC_1_123 b_1 NI_1 NS_123 0 -2.0479871692038686e-07
GC_1_124 b_1 NI_1 NS_124 0 -9.2517561068432064e-09
GC_1_125 b_1 NI_1 NS_125 0 4.9822047746826239e-05
GC_1_126 b_1 NI_1 NS_126 0 -2.0166476261031301e-06
GC_1_127 b_1 NI_1 NS_127 0 2.5357888591234080e-05
GC_1_128 b_1 NI_1 NS_128 0 -7.6229365003372955e-06
GC_1_129 b_1 NI_1 NS_129 0 2.2183853306492134e-05
GC_1_130 b_1 NI_1 NS_130 0 -2.6867991396468764e-04
GC_1_131 b_1 NI_1 NS_131 0 -2.9255258094330113e-04
GC_1_132 b_1 NI_1 NS_132 0 4.0714051694092986e-05
GC_1_133 b_1 NI_1 NS_133 0 -5.5577241280132159e-05
GC_1_134 b_1 NI_1 NS_134 0 2.2174315922405632e-04
GC_1_135 b_1 NI_1 NS_135 0 1.6780985312118407e-04
GC_1_136 b_1 NI_1 NS_136 0 -1.0454530625694145e-04
GC_1_137 b_1 NI_1 NS_137 0 -1.8111484364178790e-04
GC_1_138 b_1 NI_1 NS_138 0 6.2085961448376438e-05
GC_1_139 b_1 NI_1 NS_139 0 -5.0743164978243793e-05
GC_1_140 b_1 NI_1 NS_140 0 1.2107951032006854e-04
GC_1_141 b_1 NI_1 NS_141 0 1.3633682349464837e-04
GC_1_142 b_1 NI_1 NS_142 0 7.1243819608447431e-05
GC_1_143 b_1 NI_1 NS_143 0 -9.2884414606083208e-08
GC_1_144 b_1 NI_1 NS_144 0 4.4336493969468755e-06
GC_1_145 b_1 NI_1 NS_145 0 -2.0707155077367479e-06
GC_1_146 b_1 NI_1 NS_146 0 1.1473724863465880e-08
GC_1_147 b_1 NI_1 NS_147 0 6.2405873647293122e-10
GC_1_148 b_1 NI_1 NS_148 0 -6.3535516627720578e-10
GC_1_149 b_1 NI_1 NS_149 0 -1.5179185687246724e-10
GC_1_150 b_1 NI_1 NS_150 0 -1.2381860134912864e-09
GC_1_151 b_1 NI_1 NS_151 0 4.7532302495608042e-05
GC_1_152 b_1 NI_1 NS_152 0 9.2489060326326726e-05
GC_1_153 b_1 NI_1 NS_153 0 2.8963098674808707e-07
GC_1_154 b_1 NI_1 NS_154 0 8.4382804081398386e-09
GC_1_155 b_1 NI_1 NS_155 0 -3.9637600902170396e-05
GC_1_156 b_1 NI_1 NS_156 0 -8.5805859938133149e-05
GC_1_157 b_1 NI_1 NS_157 0 -2.2607906933834939e-04
GC_1_158 b_1 NI_1 NS_158 0 9.6527610894751769e-05
GC_1_159 b_1 NI_1 NS_159 0 2.8256934487319021e-04
GC_1_160 b_1 NI_1 NS_160 0 1.5421120011208897e-04
GC_1_161 b_1 NI_1 NS_161 0 -3.0587235898538303e-04
GC_1_162 b_1 NI_1 NS_162 0 -2.0977069118951854e-04
GC_1_163 b_1 NI_1 NS_163 0 1.8405493224260970e-04
GC_1_164 b_1 NI_1 NS_164 0 3.8935394711262601e-04
GC_1_165 b_1 NI_1 NS_165 0 -9.5573096313403963e-05
GC_1_166 b_1 NI_1 NS_166 0 -1.5669757790313975e-04
GC_1_167 b_1 NI_1 NS_167 0 2.3688406284309840e-04
GC_1_168 b_1 NI_1 NS_168 0 2.1604672907658801e-04
GC_1_169 b_1 NI_1 NS_169 0 -5.9367851293225056e-05
GC_1_170 b_1 NI_1 NS_170 0 -2.0749584370072797e-04
GC_1_171 b_1 NI_1 NS_171 0 -1.3067238855365497e-06
GC_1_172 b_1 NI_1 NS_172 0 2.1379961213818804e-04
GC_1_173 b_1 NI_1 NS_173 0 -2.2338732722259515e-06
GC_1_174 b_1 NI_1 NS_174 0 -4.4288826154165652e-08
GC_1_175 b_1 NI_1 NS_175 0 -4.0520404906195207e-07
GC_1_176 b_1 NI_1 NS_176 0 -4.3742218187353717e-07
GC_1_177 b_1 NI_1 NS_177 0 -7.4128427003811198e-10
GC_1_178 b_1 NI_1 NS_178 0 5.0839393853508331e-10
GC_1_179 b_1 NI_1 NS_179 0 1.5218539449255427e-10
GC_1_180 b_1 NI_1 NS_180 0 1.2347106299852556e-09
GC_1_181 b_1 NI_1 NS_181 0 -4.8030165494245016e-05
GC_1_182 b_1 NI_1 NS_182 0 -6.2106765977532692e-06
GC_1_183 b_1 NI_1 NS_183 0 -5.0822324214157624e-08
GC_1_184 b_1 NI_1 NS_184 0 -6.2461229807028533e-10
GC_1_185 b_1 NI_1 NS_185 0 -7.2122566014816763e-06
GC_1_186 b_1 NI_1 NS_186 0 -5.3858960035276435e-06
GC_1_187 b_1 NI_1 NS_187 0 -3.2447467578923798e-05
GC_1_188 b_1 NI_1 NS_188 0 1.3398731150196164e-05
GC_1_189 b_1 NI_1 NS_189 0 1.9868488015255909e-05
GC_1_190 b_1 NI_1 NS_190 0 6.7344523783714072e-05
GC_1_191 b_1 NI_1 NS_191 0 9.5695706376606416e-05
GC_1_192 b_1 NI_1 NS_192 0 5.2354545406303797e-06
GC_1_193 b_1 NI_1 NS_193 0 -1.6522317451739621e-05
GC_1_194 b_1 NI_1 NS_194 0 -8.9248189255793420e-05
GC_1_195 b_1 NI_1 NS_195 0 -2.8891588383810032e-05
GC_1_196 b_1 NI_1 NS_196 0 3.4604100334440696e-05
GC_1_197 b_1 NI_1 NS_197 0 5.9453625508822583e-05
GC_1_198 b_1 NI_1 NS_198 0 -3.6932691003253775e-06
GC_1_199 b_1 NI_1 NS_199 0 -5.0298066873603150e-06
GC_1_200 b_1 NI_1 NS_200 0 -5.5556149487564649e-05
GC_1_201 b_1 NI_1 NS_201 0 -2.4338392976761649e-05
GC_1_202 b_1 NI_1 NS_202 0 -1.2670122059159569e-05
GC_1_203 b_1 NI_1 NS_203 0 5.7847744909666445e-07
GC_1_204 b_1 NI_1 NS_204 0 -6.2045995145258772e-07
GC_1_205 b_1 NI_1 NS_205 0 3.4415518204085189e-07
GC_1_206 b_1 NI_1 NS_206 0 1.0348433095811233e-07
GC_1_207 b_1 NI_1 NS_207 0 1.6603308182730933e-10
GC_1_208 b_1 NI_1 NS_208 0 -8.2919294637014571e-11
GC_1_209 b_1 NI_1 NS_209 0 -7.1939834810748987e-11
GC_1_210 b_1 NI_1 NS_210 0 -4.3735873399216048e-10
GC_1_211 b_1 NI_1 NS_211 0 9.9930229858361322e-05
GC_1_212 b_1 NI_1 NS_212 0 -2.5739247203627146e-07
GC_1_213 b_1 NI_1 NS_213 0 3.9431183166667662e-08
GC_1_214 b_1 NI_1 NS_214 0 6.8131648852553780e-10
GC_1_215 b_1 NI_1 NS_215 0 2.6782821366412917e-07
GC_1_216 b_1 NI_1 NS_216 0 -1.4818922345471805e-06
GC_1_217 b_1 NI_1 NS_217 0 -9.2953824929448453e-06
GC_1_218 b_1 NI_1 NS_218 0 2.4293152255426223e-05
GC_1_219 b_1 NI_1 NS_219 0 7.9303136001844738e-05
GC_1_220 b_1 NI_1 NS_220 0 8.7579688584126695e-06
GC_1_221 b_1 NI_1 NS_221 0 1.1180701426662704e-05
GC_1_222 b_1 NI_1 NS_222 0 -7.9803303614140863e-05
GC_1_223 b_1 NI_1 NS_223 0 -7.1787625874350799e-06
GC_1_224 b_1 NI_1 NS_224 0 -4.3358678496788322e-05
GC_1_225 b_1 NI_1 NS_225 0 -9.5157367135186005e-05
GC_1_226 b_1 NI_1 NS_226 0 -5.4098637776844110e-05
GC_1_227 b_1 NI_1 NS_227 0 -4.5957061041972963e-05
GC_1_228 b_1 NI_1 NS_228 0 5.3040645741054880e-05
GC_1_229 b_1 NI_1 NS_229 0 -3.1272897361819280e-05
GC_1_230 b_1 NI_1 NS_230 0 1.2847064624797766e-05
GC_1_231 b_1 NI_1 NS_231 0 -1.6072317526480767e-05
GC_1_232 b_1 NI_1 NS_232 0 4.9857337097149633e-05
GC_1_233 b_1 NI_1 NS_233 0 -7.4582987532229643e-07
GC_1_234 b_1 NI_1 NS_234 0 -4.3446859565703741e-07
GC_1_235 b_1 NI_1 NS_235 0 1.2918952731890074e-07
GC_1_236 b_1 NI_1 NS_236 0 -3.6965427990487062e-07
GC_1_237 b_1 NI_1 NS_237 0 -1.5102428144675171e-10
GC_1_238 b_1 NI_1 NS_238 0 9.1264401285216907e-11
GC_1_239 b_1 NI_1 NS_239 0 7.1484117947439684e-11
GC_1_240 b_1 NI_1 NS_240 0 4.3623181910386343e-10
GC_1_241 b_1 NI_1 NS_241 0 1.8182625212720791e-05
GC_1_242 b_1 NI_1 NS_242 0 -2.5901336057782799e-06
GC_1_243 b_1 NI_1 NS_243 0 1.0334193042149505e-08
GC_1_244 b_1 NI_1 NS_244 0 -2.6700209463035799e-10
GC_1_245 b_1 NI_1 NS_245 0 -1.2561972122238310e-06
GC_1_246 b_1 NI_1 NS_246 0 -1.1110382636917718e-06
GC_1_247 b_1 NI_1 NS_247 0 -2.4938859599919018e-06
GC_1_248 b_1 NI_1 NS_248 0 5.3481704497596538e-07
GC_1_249 b_1 NI_1 NS_249 0 -1.2776559247790226e-06
GC_1_250 b_1 NI_1 NS_250 0 2.6875757557267938e-06
GC_1_251 b_1 NI_1 NS_251 0 1.8066986621114676e-06
GC_1_252 b_1 NI_1 NS_252 0 7.9089583455092584e-07
GC_1_253 b_1 NI_1 NS_253 0 -2.7692143574901110e-06
GC_1_254 b_1 NI_1 NS_254 0 -1.3482200148191698e-06
GC_1_255 b_1 NI_1 NS_255 0 -2.1726548319226219e-06
GC_1_256 b_1 NI_1 NS_256 0 3.4750576977494943e-06
GC_1_257 b_1 NI_1 NS_257 0 1.2557147979045646e-06
GC_1_258 b_1 NI_1 NS_258 0 2.3797765001328960e-06
GC_1_259 b_1 NI_1 NS_259 0 -9.2223765867157320e-07
GC_1_260 b_1 NI_1 NS_260 0 -3.7752720202538635e-07
GC_1_261 b_1 NI_1 NS_261 0 -3.3379670611664461e-06
GC_1_262 b_1 NI_1 NS_262 0 6.3278240379373288e-07
GC_1_263 b_1 NI_1 NS_263 0 -1.4338068586508528e-07
GC_1_264 b_1 NI_1 NS_264 0 -7.6374260657740297e-08
GC_1_265 b_1 NI_1 NS_265 0 2.3067702960128693e-08
GC_1_266 b_1 NI_1 NS_266 0 -5.2057472065136429e-08
GC_1_267 b_1 NI_1 NS_267 0 -1.8003829267488215e-11
GC_1_268 b_1 NI_1 NS_268 0 -1.0118382283199071e-10
GC_1_269 b_1 NI_1 NS_269 0 -3.8104000299223816e-11
GC_1_270 b_1 NI_1 NS_270 0 -1.6272437085525247e-10
GC_1_271 b_1 NI_1 NS_271 0 -3.1794850001861703e-05
GC_1_272 b_1 NI_1 NS_272 0 3.5425559380123644e-06
GC_1_273 b_1 NI_1 NS_273 0 -1.3247268645226713e-08
GC_1_274 b_1 NI_1 NS_274 0 3.4619745659529338e-10
GC_1_275 b_1 NI_1 NS_275 0 2.0232773863559903e-06
GC_1_276 b_1 NI_1 NS_276 0 2.9214615071111607e-07
GC_1_277 b_1 NI_1 NS_277 0 1.7680035523468812e-06
GC_1_278 b_1 NI_1 NS_278 0 -1.7931868606344991e-06
GC_1_279 b_1 NI_1 NS_279 0 2.2222057082724778e-06
GC_1_280 b_1 NI_1 NS_280 0 -1.9596522354926773e-06
GC_1_281 b_1 NI_1 NS_281 0 1.2037875421192283e-06
GC_1_282 b_1 NI_1 NS_282 0 -1.4895734197171997e-06
GC_1_283 b_1 NI_1 NS_283 0 1.6529677244294450e-06
GC_1_284 b_1 NI_1 NS_284 0 -1.3654354542635612e-06
GC_1_285 b_1 NI_1 NS_285 0 1.7718816347546757e-06
GC_1_286 b_1 NI_1 NS_286 0 -3.2631842367615317e-06
GC_1_287 b_1 NI_1 NS_287 0 1.9918739984064681e-06
GC_1_288 b_1 NI_1 NS_288 0 -3.6176766849437601e-06
GC_1_289 b_1 NI_1 NS_289 0 7.3166891044326505e-07
GC_1_290 b_1 NI_1 NS_290 0 -3.2936828329093863e-06
GC_1_291 b_1 NI_1 NS_291 0 3.3991695936595275e-06
GC_1_292 b_1 NI_1 NS_292 0 -1.4916170300591602e-06
GC_1_293 b_1 NI_1 NS_293 0 2.6898773438681725e-07
GC_1_294 b_1 NI_1 NS_294 0 3.2027539901819584e-08
GC_1_295 b_1 NI_1 NS_295 0 1.3104225981326649e-08
GC_1_296 b_1 NI_1 NS_296 0 1.2281583388441014e-07
GC_1_297 b_1 NI_1 NS_297 0 2.5320408897344669e-11
GC_1_298 b_1 NI_1 NS_298 0 1.2029654794175411e-10
GC_1_299 b_1 NI_1 NS_299 0 3.7619725736881019e-11
GC_1_300 b_1 NI_1 NS_300 0 1.6471728009536804e-10
GC_1_301 b_1 NI_1 NS_301 0 -3.0823041159463641e-05
GC_1_302 b_1 NI_1 NS_302 0 4.3669469206544884e-06
GC_1_303 b_1 NI_1 NS_303 0 -1.9330742639840092e-08
GC_1_304 b_1 NI_1 NS_304 0 3.1701659074088982e-10
GC_1_305 b_1 NI_1 NS_305 0 1.4873081353908588e-06
GC_1_306 b_1 NI_1 NS_306 0 4.2936621737491370e-07
GC_1_307 b_1 NI_1 NS_307 0 1.3518705165209421e-06
GC_1_308 b_1 NI_1 NS_308 0 -4.6259406423695931e-07
GC_1_309 b_1 NI_1 NS_309 0 2.0702782626877476e-06
GC_1_310 b_1 NI_1 NS_310 0 -5.7993616505246919e-07
GC_1_311 b_1 NI_1 NS_311 0 2.2939801237439134e-06
GC_1_312 b_1 NI_1 NS_312 0 -9.4232589017833131e-07
GC_1_313 b_1 NI_1 NS_313 0 1.8336067200804371e-06
GC_1_314 b_1 NI_1 NS_314 0 -2.7426509942743725e-06
GC_1_315 b_1 NI_1 NS_315 0 9.1063621933386100e-07
GC_1_316 b_1 NI_1 NS_316 0 -2.2463638816117886e-06
GC_1_317 b_1 NI_1 NS_317 0 1.6377156658388929e-06
GC_1_318 b_1 NI_1 NS_318 0 -2.1620951539659531e-06
GC_1_319 b_1 NI_1 NS_319 0 1.5040100244500240e-06
GC_1_320 b_1 NI_1 NS_320 0 -1.7688846752749136e-06
GC_1_321 b_1 NI_1 NS_321 0 5.2307160855944447e-06
GC_1_322 b_1 NI_1 NS_322 0 -4.1141527227809607e-07
GC_1_323 b_1 NI_1 NS_323 0 3.8001754836372970e-07
GC_1_324 b_1 NI_1 NS_324 0 -1.9134699893845350e-08
GC_1_325 b_1 NI_1 NS_325 0 3.5322962729343012e-08
GC_1_326 b_1 NI_1 NS_326 0 1.6834348811765540e-07
GC_1_327 b_1 NI_1 NS_327 0 8.1397044866661010e-11
GC_1_328 b_1 NI_1 NS_328 0 -1.5436046543742493e-12
GC_1_329 b_1 NI_1 NS_329 0 -4.0249851792097435e-11
GC_1_330 b_1 NI_1 NS_330 0 -1.3801730243923780e-10
GC_1_331 b_1 NI_1 NS_331 0 -1.5473891009724389e-05
GC_1_332 b_1 NI_1 NS_332 0 5.0273919491687584e-07
GC_1_333 b_1 NI_1 NS_333 0 9.6893760062598422e-09
GC_1_334 b_1 NI_1 NS_334 0 -7.3056667979487944e-11
GC_1_335 b_1 NI_1 NS_335 0 1.1231109018942431e-06
GC_1_336 b_1 NI_1 NS_336 0 2.1488802263240310e-07
GC_1_337 b_1 NI_1 NS_337 0 1.1947568618812426e-06
GC_1_338 b_1 NI_1 NS_338 0 -1.3852148686748370e-07
GC_1_339 b_1 NI_1 NS_339 0 9.0379842315313543e-07
GC_1_340 b_1 NI_1 NS_340 0 -1.0516121061574309e-06
GC_1_341 b_1 NI_1 NS_341 0 8.4623776183425452e-07
GC_1_342 b_1 NI_1 NS_342 0 -4.8065438920568379e-07
GC_1_343 b_1 NI_1 NS_343 0 1.5417938274263870e-06
GC_1_344 b_1 NI_1 NS_344 0 -9.6405338861935125e-07
GC_1_345 b_1 NI_1 NS_345 0 1.0933707110777042e-06
GC_1_346 b_1 NI_1 NS_346 0 -1.7255575062250296e-06
GC_1_347 b_1 NI_1 NS_347 0 1.0576547076433122e-06
GC_1_348 b_1 NI_1 NS_348 0 -2.2497661051703504e-06
GC_1_349 b_1 NI_1 NS_349 0 6.5021034836509512e-07
GC_1_350 b_1 NI_1 NS_350 0 -1.7357122085014962e-06
GC_1_351 b_1 NI_1 NS_351 0 1.7290801823499282e-06
GC_1_352 b_1 NI_1 NS_352 0 -2.0366571167603228e-06
GC_1_353 b_1 NI_1 NS_353 0 1.1291332138200713e-09
GC_1_354 b_1 NI_1 NS_354 0 -2.3439243502814946e-07
GC_1_355 b_1 NI_1 NS_355 0 1.1724055544102185e-07
GC_1_356 b_1 NI_1 NS_356 0 2.0287778198687974e-08
GC_1_357 b_1 NI_1 NS_357 0 -7.0700042972473101e-11
GC_1_358 b_1 NI_1 NS_358 0 5.3485835597488332e-11
GC_1_359 b_1 NI_1 NS_359 0 3.3464773786076912e-11
GC_1_360 b_1 NI_1 NS_360 0 1.2644123521570174e-10
GD_1_1 b_1 NI_1 NA_1 0 -4.0049975508414160e-02
GD_1_2 b_1 NI_1 NA_2 0 -1.0827014056013235e-02
GD_1_3 b_1 NI_1 NA_3 0 1.6056004849533949e-02
GD_1_4 b_1 NI_1 NA_4 0 -9.1340175096391680e-05
GD_1_5 b_1 NI_1 NA_5 0 1.6881266759458048e-04
GD_1_6 b_1 NI_1 NA_6 0 -6.0788962078540493e-05
GD_1_7 b_1 NI_1 NA_7 0 2.0534845509270064e-06
GD_1_8 b_1 NI_1 NA_8 0 8.3717107010715086e-06
GD_1_9 b_1 NI_1 NA_9 0 -1.7399465073016224e-06
GD_1_10 b_1 NI_1 NA_10 0 7.7104331759435749e-06
GD_1_11 b_1 NI_1 NA_11 0 5.1394395385474123e-06
GD_1_12 b_1 NI_1 NA_12 0 2.7202904986132240e-06
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 -7.0424727392403116e-02
GC_2_2 b_2 NI_2 NS_2 0 2.4192834837785771e-02
GC_2_3 b_2 NI_2 NS_3 0 2.2092933769820189e-05
GC_2_4 b_2 NI_2 NS_4 0 5.3186599157114162e-06
GC_2_5 b_2 NI_2 NS_5 0 1.8108338849417645e-02
GC_2_6 b_2 NI_2 NS_6 0 2.7946335353168480e-02
GC_2_7 b_2 NI_2 NS_7 0 -1.9395058756833134e-02
GC_2_8 b_2 NI_2 NS_8 0 8.3724949376921438e-03
GC_2_9 b_2 NI_2 NS_9 0 -5.8925728120722181e-03
GC_2_10 b_2 NI_2 NS_10 0 -2.2930897953348291e-02
GC_2_11 b_2 NI_2 NS_11 0 2.6387189303234193e-02
GC_2_12 b_2 NI_2 NS_12 0 -1.4337489845710682e-02
GC_2_13 b_2 NI_2 NS_13 0 3.4164839587030066e-02
GC_2_14 b_2 NI_2 NS_14 0 5.2157736701611236e-03
GC_2_15 b_2 NI_2 NS_15 0 9.5147632681178082e-03
GC_2_16 b_2 NI_2 NS_16 0 1.4168224215240445e-02
GC_2_17 b_2 NI_2 NS_17 0 -1.2626416207372298e-02
GC_2_18 b_2 NI_2 NS_18 0 1.1356483334400721e-02
GC_2_19 b_2 NI_2 NS_19 0 -1.1978307960545557e-02
GC_2_20 b_2 NI_2 NS_20 0 -1.1686227616094910e-02
GC_2_21 b_2 NI_2 NS_21 0 1.9051198532209733e-02
GC_2_22 b_2 NI_2 NS_22 0 -2.5965294083176136e-02
GC_2_23 b_2 NI_2 NS_23 0 9.0694545815386829e-04
GC_2_24 b_2 NI_2 NS_24 0 -1.0849119409543234e-03
GC_2_25 b_2 NI_2 NS_25 0 6.2679747823162673e-04
GC_2_26 b_2 NI_2 NS_26 0 3.2175984387846517e-04
GC_2_27 b_2 NI_2 NS_27 0 9.0179349467595180e-08
GC_2_28 b_2 NI_2 NS_28 0 4.0614943939421670e-07
GC_2_29 b_2 NI_2 NS_29 0 -9.1805817910990836e-09
GC_2_30 b_2 NI_2 NS_30 0 -1.8631085292257708e-08
GC_2_31 b_2 NI_2 NS_31 0 1.2526108569063468e-01
GC_2_32 b_2 NI_2 NS_32 0 -9.7551738268520007e-03
GC_2_33 b_2 NI_2 NS_33 0 -2.1879140150518190e-05
GC_2_34 b_2 NI_2 NS_34 0 -3.7984593841401867e-06
GC_2_35 b_2 NI_2 NS_35 0 -8.0420603776076450e-03
GC_2_36 b_2 NI_2 NS_36 0 6.5371474564688496e-04
GC_2_37 b_2 NI_2 NS_37 0 -1.9771749923377119e-03
GC_2_38 b_2 NI_2 NS_38 0 1.0156944859432946e-04
GC_2_39 b_2 NI_2 NS_39 0 -1.2487317258108407e-02
GC_2_40 b_2 NI_2 NS_40 0 8.2382539291840032e-03
GC_2_41 b_2 NI_2 NS_41 0 -1.0111830234426761e-02
GC_2_42 b_2 NI_2 NS_42 0 -5.9611418424684534e-04
GC_2_43 b_2 NI_2 NS_43 0 -3.4891091292882166e-03
GC_2_44 b_2 NI_2 NS_44 0 1.6807110978405121e-02
GC_2_45 b_2 NI_2 NS_45 0 -7.7156973516644958e-03
GC_2_46 b_2 NI_2 NS_46 0 1.3269796070236668e-02
GC_2_47 b_2 NI_2 NS_47 0 -3.8876518720964018e-03
GC_2_48 b_2 NI_2 NS_48 0 6.8943385148697483e-03
GC_2_49 b_2 NI_2 NS_49 0 -2.7117302567003744e-03
GC_2_50 b_2 NI_2 NS_50 0 1.2199575250037462e-02
GC_2_51 b_2 NI_2 NS_51 0 -2.2742233491917691e-02
GC_2_52 b_2 NI_2 NS_52 0 5.9617102582374543e-03
GC_2_53 b_2 NI_2 NS_53 0 -8.4148567214240868e-04
GC_2_54 b_2 NI_2 NS_54 0 8.1300274134813279e-04
GC_2_55 b_2 NI_2 NS_55 0 -5.1564584094578253e-04
GC_2_56 b_2 NI_2 NS_56 0 -4.3051992490342899e-04
GC_2_57 b_2 NI_2 NS_57 0 -5.9275332955220085e-08
GC_2_58 b_2 NI_2 NS_58 0 -1.8756500527532776e-07
GC_2_59 b_2 NI_2 NS_59 0 -3.3579646716791644e-09
GC_2_60 b_2 NI_2 NS_60 0 5.3365681839077154e-09
GC_2_61 b_2 NI_2 NS_61 0 1.3559977266744913e-03
GC_2_62 b_2 NI_2 NS_62 0 -1.2038876436075252e-03
GC_2_63 b_2 NI_2 NS_63 0 3.7357899062376710e-06
GC_2_64 b_2 NI_2 NS_64 0 2.8902025643849504e-07
GC_2_65 b_2 NI_2 NS_65 0 1.2297103897554874e-04
GC_2_66 b_2 NI_2 NS_66 0 8.9417681564479302e-04
GC_2_67 b_2 NI_2 NS_67 0 1.8425181613901315e-03
GC_2_68 b_2 NI_2 NS_68 0 -8.6745204795828318e-04
GC_2_69 b_2 NI_2 NS_69 0 -2.9665984448699568e-03
GC_2_70 b_2 NI_2 NS_70 0 -1.6486215866938043e-03
GC_2_71 b_2 NI_2 NS_71 0 2.2194995090932318e-03
GC_2_72 b_2 NI_2 NS_72 0 2.6689300497476057e-03
GC_2_73 b_2 NI_2 NS_73 0 -1.4401272077413688e-03
GC_2_74 b_2 NI_2 NS_74 0 -2.9129239481826830e-03
GC_2_75 b_2 NI_2 NS_75 0 1.0698835745838750e-03
GC_2_76 b_2 NI_2 NS_76 0 2.2566924764752961e-03
GC_2_77 b_2 NI_2 NS_77 0 -1.6275425023276815e-03
GC_2_78 b_2 NI_2 NS_78 0 -2.1363730378469023e-03
GC_2_79 b_2 NI_2 NS_79 0 4.2046566768591022e-04
GC_2_80 b_2 NI_2 NS_80 0 2.0118498158383678e-03
GC_2_81 b_2 NI_2 NS_81 0 2.1508326771149073e-04
GC_2_82 b_2 NI_2 NS_82 0 -2.1102726803263836e-03
GC_2_83 b_2 NI_2 NS_83 0 -4.3290758021215855e-06
GC_2_84 b_2 NI_2 NS_84 0 4.3528691030183871e-06
GC_2_85 b_2 NI_2 NS_85 0 -7.8953772068273550e-07
GC_2_86 b_2 NI_2 NS_86 0 -3.5250190153439896e-06
GC_2_87 b_2 NI_2 NS_87 0 -7.5479910794323688e-09
GC_2_88 b_2 NI_2 NS_88 0 2.2567545206182170e-08
GC_2_89 b_2 NI_2 NS_89 0 2.3359230281103038e-09
GC_2_90 b_2 NI_2 NS_90 0 1.5101849077683507e-09
GC_2_91 b_2 NI_2 NS_91 0 -5.4930026805724032e-04
GC_2_92 b_2 NI_2 NS_92 0 -2.9018693022416259e-03
GC_2_93 b_2 NI_2 NS_93 0 -6.1489190989427876e-06
GC_2_94 b_2 NI_2 NS_94 0 -3.8642013610523104e-07
GC_2_95 b_2 NI_2 NS_95 0 2.6865571608067529e-03
GC_2_96 b_2 NI_2 NS_96 0 -1.9871345790794521e-03
GC_2_97 b_2 NI_2 NS_97 0 -6.1989446682094110e-03
GC_2_98 b_2 NI_2 NS_98 0 1.7530826878390327e-03
GC_2_99 b_2 NI_2 NS_99 0 4.7648950909667783e-03
GC_2_100 b_2 NI_2 NS_100 0 -5.5284542855493076e-03
GC_2_101 b_2 NI_2 NS_101 0 -2.4813945917554571e-04
GC_2_102 b_2 NI_2 NS_102 0 7.2493802967724440e-03
GC_2_103 b_2 NI_2 NS_103 0 -6.3155980978114139e-03
GC_2_104 b_2 NI_2 NS_104 0 -5.0550518692204045e-03
GC_2_105 b_2 NI_2 NS_105 0 4.5025743711784817e-03
GC_2_106 b_2 NI_2 NS_106 0 -1.7116291151872489e-03
GC_2_107 b_2 NI_2 NS_107 0 -5.9124273565084099e-04
GC_2_108 b_2 NI_2 NS_108 0 6.9477768462132428e-03
GC_2_109 b_2 NI_2 NS_109 0 -3.4362381852351101e-03
GC_2_110 b_2 NI_2 NS_110 0 -3.6821939951053985e-03
GC_2_111 b_2 NI_2 NS_111 0 5.9242818960603310e-03
GC_2_112 b_2 NI_2 NS_112 0 3.9701299788723587e-04
GC_2_113 b_2 NI_2 NS_113 0 6.3747582452007386e-05
GC_2_114 b_2 NI_2 NS_114 0 8.4790923774572153e-06
GC_2_115 b_2 NI_2 NS_115 0 1.5085785272717732e-05
GC_2_116 b_2 NI_2 NS_116 0 3.9927089988350551e-05
GC_2_117 b_2 NI_2 NS_117 0 7.1121045721118138e-09
GC_2_118 b_2 NI_2 NS_118 0 -2.9352073930738686e-08
GC_2_119 b_2 NI_2 NS_119 0 -1.8854152519877874e-09
GC_2_120 b_2 NI_2 NS_120 0 -5.6020820707838304e-10
GC_2_121 b_2 NI_2 NS_121 0 4.7529413165484524e-05
GC_2_122 b_2 NI_2 NS_122 0 9.2489244857228448e-05
GC_2_123 b_2 NI_2 NS_123 0 2.8963834630997502e-07
GC_2_124 b_2 NI_2 NS_124 0 8.4383170805671048e-09
GC_2_125 b_2 NI_2 NS_125 0 -3.9637640075695551e-05
GC_2_126 b_2 NI_2 NS_126 0 -8.5800994876814569e-05
GC_2_127 b_2 NI_2 NS_127 0 -2.2608169023087221e-04
GC_2_128 b_2 NI_2 NS_128 0 9.6531803376803655e-05
GC_2_129 b_2 NI_2 NS_129 0 2.8257314186657214e-04
GC_2_130 b_2 NI_2 NS_130 0 1.5420735095425704e-04
GC_2_131 b_2 NI_2 NS_131 0 -3.0587341643104467e-04
GC_2_132 b_2 NI_2 NS_132 0 -2.0976792741888266e-04
GC_2_133 b_2 NI_2 NS_133 0 1.8406147562467147e-04
GC_2_134 b_2 NI_2 NS_134 0 3.8935567160207693e-04
GC_2_135 b_2 NI_2 NS_135 0 -9.5573712235923154e-05
GC_2_136 b_2 NI_2 NS_136 0 -1.5669664060308678e-04
GC_2_137 b_2 NI_2 NS_137 0 2.3688714571948406e-04
GC_2_138 b_2 NI_2 NS_138 0 2.1604584921773519e-04
GC_2_139 b_2 NI_2 NS_139 0 -5.9368011903499912e-05
GC_2_140 b_2 NI_2 NS_140 0 -2.0749699594071669e-04
GC_2_141 b_2 NI_2 NS_141 0 -1.3040378654955030e-06
GC_2_142 b_2 NI_2 NS_142 0 2.1379953079372620e-04
GC_2_143 b_2 NI_2 NS_143 0 -2.2339329408223775e-06
GC_2_144 b_2 NI_2 NS_144 0 -4.4443803625378544e-08
GC_2_145 b_2 NI_2 NS_145 0 -4.0519947981923578e-07
GC_2_146 b_2 NI_2 NS_146 0 -4.3752055683372772e-07
GC_2_147 b_2 NI_2 NS_147 0 -7.4130864852889069e-10
GC_2_148 b_2 NI_2 NS_148 0 5.0839010624250623e-10
GC_2_149 b_2 NI_2 NS_149 0 1.5218849424757864e-10
GC_2_150 b_2 NI_2 NS_150 0 1.2347152275016276e-09
GC_2_151 b_2 NI_2 NS_151 0 1.2794855192473160e-04
GC_2_152 b_2 NI_2 NS_152 0 2.8895182655522254e-06
GC_2_153 b_2 NI_2 NS_153 0 -2.0789759231299858e-07
GC_2_154 b_2 NI_2 NS_154 0 -9.2148621634976437e-09
GC_2_155 b_2 NI_2 NS_155 0 5.0391238638772716e-05
GC_2_156 b_2 NI_2 NS_156 0 -1.8561640247832048e-06
GC_2_157 b_2 NI_2 NS_157 0 2.6276469853080685e-05
GC_2_158 b_2 NI_2 NS_158 0 -7.5099482206127105e-06
GC_2_159 b_2 NI_2 NS_159 0 2.3050776493658090e-05
GC_2_160 b_2 NI_2 NS_160 0 -2.6914133535686124e-04
GC_2_161 b_2 NI_2 NS_161 0 -2.9117457361226880e-04
GC_2_162 b_2 NI_2 NS_162 0 4.0238017781552404e-05
GC_2_163 b_2 NI_2 NS_163 0 -5.4545161838428489e-05
GC_2_164 b_2 NI_2 NS_164 0 2.2062130375134488e-04
GC_2_165 b_2 NI_2 NS_165 0 1.6841453183222339e-04
GC_2_166 b_2 NI_2 NS_166 0 -1.0598925854589854e-04
GC_2_167 b_2 NI_2 NS_167 0 -1.8032968810932095e-04
GC_2_168 b_2 NI_2 NS_168 0 6.0705395711715805e-05
GC_2_169 b_2 NI_2 NS_169 0 -5.0071063353889852e-05
GC_2_170 b_2 NI_2 NS_170 0 1.2013387923837640e-04
GC_2_171 b_2 NI_2 NS_171 0 1.3866115967268544e-04
GC_2_172 b_2 NI_2 NS_172 0 7.0602025123805637e-05
GC_2_173 b_2 NI_2 NS_173 0 4.2957807930818278e-08
GC_2_174 b_2 NI_2 NS_174 0 4.3451731169801397e-06
GC_2_175 b_2 NI_2 NS_175 0 -2.0150898600880364e-06
GC_2_176 b_2 NI_2 NS_176 0 7.7203156428997177e-08
GC_2_177 b_2 NI_2 NS_177 0 6.2847951574025054e-10
GC_2_178 b_2 NI_2 NS_178 0 -6.3035852452798058e-10
GC_2_179 b_2 NI_2 NS_179 0 -1.5189613838040431e-10
GC_2_180 b_2 NI_2 NS_180 0 -1.2381203643571034e-09
GC_2_181 b_2 NI_2 NS_181 0 9.8877785070643459e-05
GC_2_182 b_2 NI_2 NS_182 0 -1.7560093488485004e-07
GC_2_183 b_2 NI_2 NS_183 0 3.9323538744480882e-08
GC_2_184 b_2 NI_2 NS_184 0 6.8242717487886893e-10
GC_2_185 b_2 NI_2 NS_185 0 4.2701071249617115e-07
GC_2_186 b_2 NI_2 NS_186 0 -1.4257167325828964e-06
GC_2_187 b_2 NI_2 NS_187 0 -9.1784462901672188e-06
GC_2_188 b_2 NI_2 NS_188 0 2.4322921242336077e-05
GC_2_189 b_2 NI_2 NS_189 0 7.9325301335251921e-05
GC_2_190 b_2 NI_2 NS_190 0 8.5014431698911742e-06
GC_2_191 b_2 NI_2 NS_191 0 1.1235555374812648e-05
GC_2_192 b_2 NI_2 NS_192 0 -7.9840732395680488e-05
GC_2_193 b_2 NI_2 NS_193 0 -7.0607541942039519e-06
GC_2_194 b_2 NI_2 NS_194 0 -4.3550072088876475e-05
GC_2_195 b_2 NI_2 NS_195 0 -9.5183559073734342e-05
GC_2_196 b_2 NI_2 NS_196 0 -5.4168023905006704e-05
GC_2_197 b_2 NI_2 NS_197 0 -4.5943856432065576e-05
GC_2_198 b_2 NI_2 NS_198 0 5.2906450068040912e-05
GC_2_199 b_2 NI_2 NS_199 0 -3.1270743479699501e-05
GC_2_200 b_2 NI_2 NS_200 0 1.2779481423219312e-05
GC_2_201 b_2 NI_2 NS_201 0 -1.5940311237708078e-05
GC_2_202 b_2 NI_2 NS_202 0 4.9776955278230399e-05
GC_2_203 b_2 NI_2 NS_203 0 -7.4154433515940611e-07
GC_2_204 b_2 NI_2 NS_204 0 -4.3929230201024221e-07
GC_2_205 b_2 NI_2 NS_205 0 1.3271427074365062e-07
GC_2_206 b_2 NI_2 NS_206 0 -3.6747240861395457e-07
GC_2_207 b_2 NI_2 NS_207 0 -1.5075739537554006e-10
GC_2_208 b_2 NI_2 NS_208 0 9.1441434255970572e-11
GC_2_209 b_2 NI_2 NS_209 0 7.1476092619088932e-11
GC_2_210 b_2 NI_2 NS_210 0 4.3621313986425694e-10
GC_2_211 b_2 NI_2 NS_211 0 -4.8135714769825500e-05
GC_2_212 b_2 NI_2 NS_212 0 -6.1994511271867682e-06
GC_2_213 b_2 NI_2 NS_213 0 -5.0843099261702141e-08
GC_2_214 b_2 NI_2 NS_214 0 -6.2431981832288768e-10
GC_2_215 b_2 NI_2 NS_215 0 -7.2065667795029314e-06
GC_2_216 b_2 NI_2 NS_216 0 -5.3857708434163281e-06
GC_2_217 b_2 NI_2 NS_217 0 -3.2442024648178950e-05
GC_2_218 b_2 NI_2 NS_218 0 1.3398299595943438e-05
GC_2_219 b_2 NI_2 NS_219 0 1.9876528156601649e-05
GC_2_220 b_2 NI_2 NS_220 0 6.7339623922866361e-05
GC_2_221 b_2 NI_2 NS_221 0 9.5704756287069608e-05
GC_2_222 b_2 NI_2 NS_222 0 5.2308314636381354e-06
GC_2_223 b_2 NI_2 NS_223 0 -1.6517241259511441e-05
GC_2_224 b_2 NI_2 NS_224 0 -8.9259113655620255e-05
GC_2_225 b_2 NI_2 NS_225 0 -2.8888132894773618e-05
GC_2_226 b_2 NI_2 NS_226 0 3.4594520379346589e-05
GC_2_227 b_2 NI_2 NS_227 0 5.9457511346590108e-05
GC_2_228 b_2 NI_2 NS_228 0 -3.7031010423944560e-06
GC_2_229 b_2 NI_2 NS_229 0 -5.0255516147133633e-06
GC_2_230 b_2 NI_2 NS_230 0 -5.5563156298473177e-05
GC_2_231 b_2 NI_2 NS_231 0 -2.4322595421449320e-05
GC_2_232 b_2 NI_2 NS_232 0 -1.2674779114447670e-05
GC_2_233 b_2 NI_2 NS_233 0 5.7935587685385404e-07
GC_2_234 b_2 NI_2 NS_234 0 -6.2107067174505409e-07
GC_2_235 b_2 NI_2 NS_235 0 3.4453230455533446e-07
GC_2_236 b_2 NI_2 NS_236 0 1.0390765899563617e-07
GC_2_237 b_2 NI_2 NS_237 0 1.6608214093380748e-10
GC_2_238 b_2 NI_2 NS_238 0 -8.2866585860421686e-11
GC_2_239 b_2 NI_2 NS_239 0 -7.1942980316782607e-11
GC_2_240 b_2 NI_2 NS_240 0 -4.3736248633330873e-10
GC_2_241 b_2 NI_2 NS_241 0 -3.1793573529091818e-05
GC_2_242 b_2 NI_2 NS_242 0 3.5424378234236163e-06
GC_2_243 b_2 NI_2 NS_243 0 -1.3247016244259810e-08
GC_2_244 b_2 NI_2 NS_244 0 3.4619122456230193e-10
GC_2_245 b_2 NI_2 NS_245 0 2.0231536468614670e-06
GC_2_246 b_2 NI_2 NS_246 0 2.9210661916247262e-07
GC_2_247 b_2 NI_2 NS_247 0 1.7678880691984389e-06
GC_2_248 b_2 NI_2 NS_248 0 -1.7931419403378394e-06
GC_2_249 b_2 NI_2 NS_249 0 2.2220719255206669e-06
GC_2_250 b_2 NI_2 NS_250 0 -1.9594594941982678e-06
GC_2_251 b_2 NI_2 NS_251 0 1.2037175642543786e-06
GC_2_252 b_2 NI_2 NS_252 0 -1.4894341770626221e-06
GC_2_253 b_2 NI_2 NS_253 0 1.6529547174242388e-06
GC_2_254 b_2 NI_2 NS_254 0 -1.3652561397798644e-06
GC_2_255 b_2 NI_2 NS_255 0 1.7719400771501643e-06
GC_2_256 b_2 NI_2 NS_256 0 -3.2630848438480849e-06
GC_2_257 b_2 NI_2 NS_257 0 1.9918528084035700e-06
GC_2_258 b_2 NI_2 NS_258 0 -3.6175779313296203e-06
GC_2_259 b_2 NI_2 NS_259 0 7.3162851047263495e-07
GC_2_260 b_2 NI_2 NS_260 0 -3.2936016375505469e-06
GC_2_261 b_2 NI_2 NS_261 0 3.3990069601850210e-06
GC_2_262 b_2 NI_2 NS_262 0 -1.4915449350852330e-06
GC_2_263 b_2 NI_2 NS_263 0 2.6897948219837712e-07
GC_2_264 b_2 NI_2 NS_264 0 3.2033132458016121e-08
GC_2_265 b_2 NI_2 NS_265 0 1.3100791047908568e-08
GC_2_266 b_2 NI_2 NS_266 0 1.2281189687862081e-07
GC_2_267 b_2 NI_2 NS_267 0 2.5320003958778054e-11
GC_2_268 b_2 NI_2 NS_268 0 1.2029520784905085e-10
GC_2_269 b_2 NI_2 NS_269 0 3.7619860952150127e-11
GC_2_270 b_2 NI_2 NS_270 0 1.6471739417392505e-10
GC_2_271 b_2 NI_2 NS_271 0 1.7965861797371931e-05
GC_2_272 b_2 NI_2 NS_272 0 -2.5639519500940998e-06
GC_2_273 b_2 NI_2 NS_273 0 1.0272994988560639e-08
GC_2_274 b_2 NI_2 NS_274 0 -2.6568078946026766e-10
GC_2_275 b_2 NI_2 NS_275 0 -1.2437459975973932e-06
GC_2_276 b_2 NI_2 NS_276 0 -1.1106323162281758e-06
GC_2_277 b_2 NI_2 NS_277 0 -2.4819748656303872e-06
GC_2_278 b_2 NI_2 NS_278 0 5.4032062050823426e-07
GC_2_279 b_2 NI_2 NS_279 0 -1.2563619757899755e-06
GC_2_280 b_2 NI_2 NS_280 0 2.6678121234005862e-06
GC_2_281 b_2 NI_2 NS_281 0 1.8212420090990724e-06
GC_2_282 b_2 NI_2 NS_282 0 7.7843852075432266e-07
GC_2_283 b_2 NI_2 NS_283 0 -2.7681914998404720e-06
GC_2_284 b_2 NI_2 NS_284 0 -1.3641178129456397e-06
GC_2_285 b_2 NI_2 NS_285 0 -2.1614706859116978e-06
GC_2_286 b_2 NI_2 NS_286 0 3.4589233062556999e-06
GC_2_287 b_2 NI_2 NS_287 0 1.2662035953028954e-06
GC_2_288 b_2 NI_2 NS_288 0 2.3623979147263239e-06
GC_2_289 b_2 NI_2 NS_289 0 -9.1304848062052170e-07
GC_2_290 b_2 NI_2 NS_290 0 -3.9147086914891022e-07
GC_2_291 b_2 NI_2 NS_291 0 -3.3032133222126457e-06
GC_2_292 b_2 NI_2 NS_292 0 6.2694718191815283e-07
GC_2_293 b_2 NI_2 NS_293 0 -1.4109287200359197e-07
GC_2_294 b_2 NI_2 NS_294 0 -7.7483885978549345e-08
GC_2_295 b_2 NI_2 NS_295 0 2.3769447646566807e-08
GC_2_296 b_2 NI_2 NS_296 0 -5.0980976241574899e-08
GC_2_297 b_2 NI_2 NS_297 0 -1.7923333291363817e-11
GC_2_298 b_2 NI_2 NS_298 0 -1.0091409175816505e-10
GC_2_299 b_2 NI_2 NS_299 0 -3.8139225202536526e-11
GC_2_300 b_2 NI_2 NS_300 0 -1.6276483846663709e-10
GC_2_301 b_2 NI_2 NS_301 0 -1.5512838963412092e-05
GC_2_302 b_2 NI_2 NS_302 0 5.0657948591386815e-07
GC_2_303 b_2 NI_2 NS_303 0 9.6809805599882063e-09
GC_2_304 b_2 NI_2 NS_304 0 -7.2853267454243433e-11
GC_2_305 b_2 NI_2 NS_305 0 1.1250117505983639e-06
GC_2_306 b_2 NI_2 NS_306 0 2.1547633630149899e-07
GC_2_307 b_2 NI_2 NS_307 0 1.1958320984711174e-06
GC_2_308 b_2 NI_2 NS_308 0 -1.3674766167420031e-07
GC_2_309 b_2 NI_2 NS_309 0 9.0974009160248183e-07
GC_2_310 b_2 NI_2 NS_310 0 -1.0540137489237922e-06
GC_2_311 b_2 NI_2 NS_311 0 8.4885470350700835e-07
GC_2_312 b_2 NI_2 NS_312 0 -4.8307583523757187e-07
GC_2_313 b_2 NI_2 NS_313 0 1.5466602851058459e-06
GC_2_314 b_2 NI_2 NS_314 0 -9.6833602555422640e-07
GC_2_315 b_2 NI_2 NS_315 0 1.0931328100884654e-06
GC_2_316 b_2 NI_2 NS_316 0 -1.7311313532477137e-06
GC_2_317 b_2 NI_2 NS_317 0 1.0586181103382640e-06
GC_2_318 b_2 NI_2 NS_318 0 -2.2535260994625728e-06
GC_2_319 b_2 NI_2 NS_319 0 6.5143340144887638e-07
GC_2_320 b_2 NI_2 NS_320 0 -1.7389301313369657e-06
GC_2_321 b_2 NI_2 NS_321 0 1.7338385641467393e-06
GC_2_322 b_2 NI_2 NS_322 0 -2.0387001201420721e-06
GC_2_323 b_2 NI_2 NS_323 0 1.4316551614484683e-09
GC_2_324 b_2 NI_2 NS_324 0 -2.3457319693319715e-07
GC_2_325 b_2 NI_2 NS_325 0 1.1736229159126305e-07
GC_2_326 b_2 NI_2 NS_326 0 2.0439108621049986e-08
GC_2_327 b_2 NI_2 NS_327 0 -7.0685152823505588e-11
GC_2_328 b_2 NI_2 NS_328 0 5.3530547790474028e-11
GC_2_329 b_2 NI_2 NS_329 0 3.3461061496168521e-11
GC_2_330 b_2 NI_2 NS_330 0 1.2644062363800532e-10
GC_2_331 b_2 NI_2 NS_331 0 -3.0823726913123485e-05
GC_2_332 b_2 NI_2 NS_332 0 4.3670088130998961e-06
GC_2_333 b_2 NI_2 NS_333 0 -1.9330853593359727e-08
GC_2_334 b_2 NI_2 NS_334 0 3.1701889080545857e-10
GC_2_335 b_2 NI_2 NS_335 0 1.4873613528276718e-06
GC_2_336 b_2 NI_2 NS_336 0 4.2934781911002894e-07
GC_2_337 b_2 NI_2 NS_337 0 1.3519114405975383e-06
GC_2_338 b_2 NI_2 NS_338 0 -4.6262466542331226e-07
GC_2_339 b_2 NI_2 NS_339 0 2.0703115455988080e-06
GC_2_340 b_2 NI_2 NS_340 0 -5.7999535522853430e-07
GC_2_341 b_2 NI_2 NS_341 0 2.2940195668170827e-06
GC_2_342 b_2 NI_2 NS_342 0 -9.4237083997098930e-07
GC_2_343 b_2 NI_2 NS_343 0 1.8336243360095074e-06
GC_2_344 b_2 NI_2 NS_344 0 -2.7427284313265883e-06
GC_2_345 b_2 NI_2 NS_345 0 9.1064040817943276e-07
GC_2_346 b_2 NI_2 NS_346 0 -2.2464260729603807e-06
GC_2_347 b_2 NI_2 NS_347 0 1.6377248763060868e-06
GC_2_348 b_2 NI_2 NS_348 0 -2.1621584658267294e-06
GC_2_349 b_2 NI_2 NS_349 0 1.5040333640258170e-06
GC_2_350 b_2 NI_2 NS_350 0 -1.7689261022890319e-06
GC_2_351 b_2 NI_2 NS_351 0 5.2308081919982187e-06
GC_2_352 b_2 NI_2 NS_352 0 -4.1145695548180041e-07
GC_2_353 b_2 NI_2 NS_353 0 3.8002143867841813e-07
GC_2_354 b_2 NI_2 NS_354 0 -1.9138288237275258e-08
GC_2_355 b_2 NI_2 NS_355 0 3.5325231967939288e-08
GC_2_356 b_2 NI_2 NS_356 0 1.6834529642056422e-07
GC_2_357 b_2 NI_2 NS_357 0 8.1397299508614123e-11
GC_2_358 b_2 NI_2 NS_358 0 -1.5430842811938193e-12
GC_2_359 b_2 NI_2 NS_359 0 -4.0249872354478894e-11
GC_2_360 b_2 NI_2 NS_360 0 -1.3801720844569949e-10
GD_2_1 b_2 NI_2 NA_1 0 -1.0827123500652965e-02
GD_2_2 b_2 NI_2 NA_2 0 -4.0049975508414104e-02
GD_2_3 b_2 NI_2 NA_3 0 -9.1324786502561072e-05
GD_2_4 b_2 NI_2 NA_4 0 1.6053745417191796e-02
GD_2_5 b_2 NI_2 NA_5 0 -6.0795871331765681e-05
GD_2_6 b_2 NI_2 NA_6 0 1.7077821718938373e-04
GD_2_7 b_2 NI_2 NA_7 0 8.6020242704384235e-06
GD_2_8 b_2 NI_2 NA_8 0 2.0740546162087024e-06
GD_2_9 b_2 NI_2 NA_9 0 7.7100767523544134e-06
GD_2_10 b_2 NI_2 NA_10 0 -1.7050921443983463e-06
GD_2_11 b_2 NI_2 NA_11 0 2.7280703225996946e-06
GD_2_12 b_2 NI_2 NA_12 0 5.1396599975742974e-06
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 -5.4930026805734234e-04
GC_3_2 b_3 NI_3 NS_2 0 -2.9018693022415851e-03
GC_3_3 b_3 NI_3 NS_3 0 -6.1489190989435889e-06
GC_3_4 b_3 NI_3 NS_4 0 -3.8642013610519308e-07
GC_3_5 b_3 NI_3 NS_5 0 2.6865571608067490e-03
GC_3_6 b_3 NI_3 NS_6 0 -1.9871345790794513e-03
GC_3_7 b_3 NI_3 NS_7 0 -6.1989446682094041e-03
GC_3_8 b_3 NI_3 NS_8 0 1.7530826878390260e-03
GC_3_9 b_3 NI_3 NS_9 0 4.7648950909667601e-03
GC_3_10 b_3 NI_3 NS_10 0 -5.5284542855493111e-03
GC_3_11 b_3 NI_3 NS_11 0 -2.4813945917556501e-04
GC_3_12 b_3 NI_3 NS_12 0 7.2493802967724544e-03
GC_3_13 b_3 NI_3 NS_13 0 -6.3155980978114139e-03
GC_3_14 b_3 NI_3 NS_14 0 -5.0550518692203681e-03
GC_3_15 b_3 NI_3 NS_15 0 4.5025743711785120e-03
GC_3_16 b_3 NI_3 NS_16 0 -1.7116291151872309e-03
GC_3_17 b_3 NI_3 NS_17 0 -5.9124273565081442e-04
GC_3_18 b_3 NI_3 NS_18 0 6.9477768462132394e-03
GC_3_19 b_3 NI_3 NS_19 0 -3.4362381852350975e-03
GC_3_20 b_3 NI_3 NS_20 0 -3.6821939951054016e-03
GC_3_21 b_3 NI_3 NS_21 0 5.9242818960603561e-03
GC_3_22 b_3 NI_3 NS_22 0 3.9701299788724893e-04
GC_3_23 b_3 NI_3 NS_23 0 6.3747582452010977e-05
GC_3_24 b_3 NI_3 NS_24 0 8.4790923774613675e-06
GC_3_25 b_3 NI_3 NS_25 0 1.5085785272715415e-05
GC_3_26 b_3 NI_3 NS_26 0 3.9927089988351425e-05
GC_3_27 b_3 NI_3 NS_27 0 7.1121045721107145e-09
GC_3_28 b_3 NI_3 NS_28 0 -2.9352073930732085e-08
GC_3_29 b_3 NI_3 NS_29 0 -1.8854152519888644e-09
GC_3_30 b_3 NI_3 NS_30 0 -5.6020820707857826e-10
GC_3_31 b_3 NI_3 NS_31 0 1.3560956931443606e-03
GC_3_32 b_3 NI_3 NS_32 0 -1.2038969097071814e-03
GC_3_33 b_3 NI_3 NS_33 0 3.7358057956577209e-06
GC_3_34 b_3 NI_3 NS_34 0 2.8902002799590245e-07
GC_3_35 b_3 NI_3 NS_35 0 1.2295927369714905e-04
GC_3_36 b_3 NI_3 NS_36 0 8.9417218286711321e-04
GC_3_37 b_3 NI_3 NS_37 0 1.8425109571019210e-03
GC_3_38 b_3 NI_3 NS_38 0 -8.6745731531467213e-04
GC_3_39 b_3 NI_3 NS_39 0 -2.9666009059735538e-03
GC_3_40 b_3 NI_3 NS_40 0 -1.6486043781858617e-03
GC_3_41 b_3 NI_3 NS_41 0 2.2194918497218863e-03
GC_3_42 b_3 NI_3 NS_42 0 2.6689302766800711e-03
GC_3_43 b_3 NI_3 NS_43 0 -1.4401401008550009e-03
GC_3_44 b_3 NI_3 NS_44 0 -2.9129078564214127e-03
GC_3_45 b_3 NI_3 NS_45 0 1.0698830025113227e-03
GC_3_46 b_3 NI_3 NS_46 0 2.2566979248096405e-03
GC_3_47 b_3 NI_3 NS_47 0 -1.6275461966845928e-03
GC_3_48 b_3 NI_3 NS_48 0 -2.1363605764622719e-03
GC_3_49 b_3 NI_3 NS_49 0 4.2046424896205876e-04
GC_3_50 b_3 NI_3 NS_50 0 2.0118561391834450e-03
GC_3_51 b_3 NI_3 NS_51 0 2.1506914840130199e-04
GC_3_52 b_3 NI_3 NS_52 0 -2.1102665001296950e-03
GC_3_53 b_3 NI_3 NS_53 0 -4.3297295367409808e-06
GC_3_54 b_3 NI_3 NS_54 0 4.3533505059811302e-06
GC_3_55 b_3 NI_3 NS_55 0 -7.8987709029423220e-07
GC_3_56 b_3 NI_3 NS_56 0 -3.5253651605178683e-06
GC_3_57 b_3 NI_3 NS_57 0 -7.5480235291728289e-09
GC_3_58 b_3 NI_3 NS_58 0 2.2567513572473928e-08
GC_3_59 b_3 NI_3 NS_59 0 2.3359255152441992e-09
GC_3_60 b_3 NI_3 NS_60 0 1.5101863938417655e-09
GC_3_61 b_3 NI_3 NS_61 0 1.2659768848160130e-01
GC_3_62 b_3 NI_3 NS_62 0 -9.9682227254338038e-03
GC_3_63 b_3 NI_3 NS_63 0 -2.0418483468456343e-05
GC_3_64 b_3 NI_3 NS_64 0 -3.8273614983901576e-06
GC_3_65 b_3 NI_3 NS_65 0 -8.0908262368300562e-03
GC_3_66 b_3 NI_3 NS_66 0 6.4296865047940141e-04
GC_3_67 b_3 NI_3 NS_67 0 -1.9909408466115956e-03
GC_3_68 b_3 NI_3 NS_68 0 6.7356143800925632e-05
GC_3_69 b_3 NI_3 NS_69 0 -1.2598719640679382e-02
GC_3_70 b_3 NI_3 NS_70 0 8.2477800777836872e-03
GC_3_71 b_3 NI_3 NS_71 0 -1.0271311615499384e-02
GC_3_72 b_3 NI_3 NS_72 0 -6.2357295410833452e-04
GC_3_73 b_3 NI_3 NS_73 0 -3.5565617083853258e-03
GC_3_74 b_3 NI_3 NS_74 0 1.6966131517386275e-02
GC_3_75 b_3 NI_3 NS_75 0 -7.7825903588609972e-03
GC_3_76 b_3 NI_3 NS_76 0 1.3370076548945831e-02
GC_3_77 b_3 NI_3 NS_77 0 -3.9902897788398799e-03
GC_3_78 b_3 NI_3 NS_78 0 6.9628713158745156e-03
GC_3_79 b_3 NI_3 NS_79 0 -2.7633627349993558e-03
GC_3_80 b_3 NI_3 NS_80 0 1.2313497559275612e-02
GC_3_81 b_3 NI_3 NS_81 0 -2.2964005253819374e-02
GC_3_82 b_3 NI_3 NS_82 0 5.9629952375129733e-03
GC_3_83 b_3 NI_3 NS_83 0 -8.6294474345638601e-04
GC_3_84 b_3 NI_3 NS_84 0 8.0344033683356624e-04
GC_3_85 b_3 NI_3 NS_85 0 -5.1358560300163571e-04
GC_3_86 b_3 NI_3 NS_86 0 -4.3937271563943101e-04
GC_3_87 b_3 NI_3 NS_87 0 -6.4174241182784420e-08
GC_3_88 b_3 NI_3 NS_88 0 -1.9155149919510570e-07
GC_3_89 b_3 NI_3 NS_89 0 -3.0939598424255364e-09
GC_3_90 b_3 NI_3 NS_90 0 5.6381472190732542e-09
GC_3_91 b_3 NI_3 NS_91 0 -7.5349163815256998e-02
GC_3_92 b_3 NI_3 NS_92 0 2.4900079417694981e-02
GC_3_93 b_3 NI_3 NS_93 0 1.9200031946918058e-05
GC_3_94 b_3 NI_3 NS_94 0 5.3863145950413912e-06
GC_3_95 b_3 NI_3 NS_95 0 1.8353491281154828e-02
GC_3_96 b_3 NI_3 NS_96 0 2.7965422967468477e-02
GC_3_97 b_3 NI_3 NS_97 0 -1.9176288461739178e-02
GC_3_98 b_3 NI_3 NS_98 0 8.3761626446775973e-03
GC_3_99 b_3 NI_3 NS_99 0 -5.5264497699069413e-03
GC_3_100 b_3 NI_3 NS_100 0 -2.3054181826065476e-02
GC_3_101 b_3 NI_3 NS_101 0 2.6687341783097281e-02
GC_3_102 b_3 NI_3 NS_102 0 -1.4576068776458622e-02
GC_3_103 b_3 NI_3 NS_103 0 3.4517374059684892e-02
GC_3_104 b_3 NI_3 NS_104 0 4.8628324173480217e-03
GC_3_105 b_3 NI_3 NS_105 0 9.6719524326555634e-03
GC_3_106 b_3 NI_3 NS_106 0 1.3692459401495893e-02
GC_3_107 b_3 NI_3 NS_107 0 -1.2370833783429231e-02
GC_3_108 b_3 NI_3 NS_108 0 1.1007973578273853e-02
GC_3_109 b_3 NI_3 NS_109 0 -1.1774494690440420e-02
GC_3_110 b_3 NI_3 NS_110 0 -1.2014107182198362e-02
GC_3_111 b_3 NI_3 NS_111 0 1.9794036474421774e-02
GC_3_112 b_3 NI_3 NS_112 0 -2.6023915309449790e-02
GC_3_113 b_3 NI_3 NS_113 0 9.6721712997440215e-04
GC_3_114 b_3 NI_3 NS_114 0 -1.0822083477013040e-03
GC_3_115 b_3 NI_3 NS_115 0 6.3094709279558445e-04
GC_3_116 b_3 NI_3 NS_116 0 3.4914543307700794e-04
GC_3_117 b_3 NI_3 NS_117 0 9.7107606131496305e-08
GC_3_118 b_3 NI_3 NS_118 0 4.1868728972869690e-07
GC_3_119 b_3 NI_3 NS_119 0 -1.0314548937310278e-08
GC_3_120 b_3 NI_3 NS_120 0 -1.9789285278344030e-08
GC_3_121 b_3 NI_3 NS_121 0 2.2651865886728025e-03
GC_3_122 b_3 NI_3 NS_122 0 -7.3251972011387765e-04
GC_3_123 b_3 NI_3 NS_123 0 -1.8149120175332799e-06
GC_3_124 b_3 NI_3 NS_124 0 -1.2099866005212076e-07
GC_3_125 b_3 NI_3 NS_125 0 3.5975567735478827e-04
GC_3_126 b_3 NI_3 NS_126 0 -3.7511051392757764e-04
GC_3_127 b_3 NI_3 NS_127 0 -1.2775980892526990e-03
GC_3_128 b_3 NI_3 NS_128 0 3.4322578639535661e-04
GC_3_129 b_3 NI_3 NS_129 0 7.1263690545177421e-04
GC_3_130 b_3 NI_3 NS_130 0 -8.2807530089469930e-04
GC_3_131 b_3 NI_3 NS_131 0 -1.5003852361326436e-04
GC_3_132 b_3 NI_3 NS_132 0 1.3910695890866915e-03
GC_3_133 b_3 NI_3 NS_133 0 -1.3010597841858007e-03
GC_3_134 b_3 NI_3 NS_134 0 -7.6485404590085119e-04
GC_3_135 b_3 NI_3 NS_135 0 6.8667001039798977e-04
GC_3_136 b_3 NI_3 NS_136 0 -2.8752446521080150e-05
GC_3_137 b_3 NI_3 NS_137 0 -1.3686847991479029e-04
GC_3_138 b_3 NI_3 NS_138 0 1.4680977678805170e-03
GC_3_139 b_3 NI_3 NS_139 0 -7.1828111558766485e-04
GC_3_140 b_3 NI_3 NS_140 0 -5.4315200812502548e-04
GC_3_141 b_3 NI_3 NS_141 0 6.5114860902977848e-04
GC_3_142 b_3 NI_3 NS_142 0 1.9303369668886660e-04
GC_3_143 b_3 NI_3 NS_143 0 -3.0047597070758387e-06
GC_3_144 b_3 NI_3 NS_144 0 2.6001120928764995e-05
GC_3_145 b_3 NI_3 NS_145 0 -9.9139321315056861e-06
GC_3_146 b_3 NI_3 NS_146 0 -1.4183971022526131e-06
GC_3_147 b_3 NI_3 NS_147 0 7.0603582380030274e-09
GC_3_148 b_3 NI_3 NS_148 0 -1.0479502326700760e-08
GC_3_149 b_3 NI_3 NS_149 0 -6.2226005295801224e-10
GC_3_150 b_3 NI_3 NS_150 0 -2.1194094617202473e-09
GC_3_151 b_3 NI_3 NS_151 0 9.8221998051327181e-04
GC_3_152 b_3 NI_3 NS_152 0 -3.4568850905820241e-04
GC_3_153 b_3 NI_3 NS_153 0 2.1363463108302340e-06
GC_3_154 b_3 NI_3 NS_154 0 8.2059870942344138e-08
GC_3_155 b_3 NI_3 NS_155 0 1.1716130537776617e-05
GC_3_156 b_3 NI_3 NS_156 0 8.7365700679801738e-05
GC_3_157 b_3 NI_3 NS_157 0 3.1568141578055251e-04
GC_3_158 b_3 NI_3 NS_158 0 -1.1545538121775877e-04
GC_3_159 b_3 NI_3 NS_159 0 -5.1920690098359332e-04
GC_3_160 b_3 NI_3 NS_160 0 -2.4290506669826195e-04
GC_3_161 b_3 NI_3 NS_161 0 3.2786513421190693e-04
GC_3_162 b_3 NI_3 NS_162 0 3.8890657171528395e-04
GC_3_163 b_3 NI_3 NS_163 0 -3.2493457998835143e-04
GC_3_164 b_3 NI_3 NS_164 0 -5.5994745677548363e-04
GC_3_165 b_3 NI_3 NS_165 0 7.3914987846073466e-05
GC_3_166 b_3 NI_3 NS_166 0 3.8468218659057780e-04
GC_3_167 b_3 NI_3 NS_167 0 -3.5604590653043355e-04
GC_3_168 b_3 NI_3 NS_168 0 -2.6839971511717886e-04
GC_3_169 b_3 NI_3 NS_169 0 5.3171183721004391e-06
GC_3_170 b_3 NI_3 NS_170 0 4.0801918374313564e-04
GC_3_171 b_3 NI_3 NS_171 0 -9.5155443024379693e-05
GC_3_172 b_3 NI_3 NS_172 0 -3.4082770314449937e-04
GC_3_173 b_3 NI_3 NS_173 0 -1.4814525093495929e-05
GC_3_174 b_3 NI_3 NS_174 0 -8.4884339744399655e-06
GC_3_175 b_3 NI_3 NS_175 0 2.7375555553973949e-06
GC_3_176 b_3 NI_3 NS_176 0 -6.6722604982037556e-06
GC_3_177 b_3 NI_3 NS_177 0 -7.7198142249859095e-09
GC_3_178 b_3 NI_3 NS_178 0 4.8069215178103958e-09
GC_3_179 b_3 NI_3 NS_179 0 1.1496323391478625e-09
GC_3_180 b_3 NI_3 NS_180 0 2.7805482816878410e-09
GC_3_181 b_3 NI_3 NS_181 0 1.2346779190605095e-04
GC_3_182 b_3 NI_3 NS_182 0 3.0700836473075641e-06
GC_3_183 b_3 NI_3 NS_183 0 -2.0465933414965203e-07
GC_3_184 b_3 NI_3 NS_184 0 -9.2708994522849683e-09
GC_3_185 b_3 NI_3 NS_185 0 5.0562971753782661e-05
GC_3_186 b_3 NI_3 NS_186 0 -1.7974655073981246e-06
GC_3_187 b_3 NI_3 NS_187 0 2.6615715036229555e-05
GC_3_188 b_3 NI_3 NS_188 0 -7.4108933215336073e-06
GC_3_189 b_3 NI_3 NS_189 0 2.3162181185390882e-05
GC_3_190 b_3 NI_3 NS_190 0 -2.6930191863051270e-04
GC_3_191 b_3 NI_3 NS_191 0 -2.9060536158607281e-04
GC_3_192 b_3 NI_3 NS_192 0 4.0320326539138950e-05
GC_3_193 b_3 NI_3 NS_193 0 -5.3916150546226429e-05
GC_3_194 b_3 NI_3 NS_194 0 2.2026889071697335e-04
GC_3_195 b_3 NI_3 NS_195 0 1.6852299406448234e-04
GC_3_196 b_3 NI_3 NS_196 0 -1.0673931075432540e-04
GC_3_197 b_3 NI_3 NS_197 0 -1.8008568489094343e-04
GC_3_198 b_3 NI_3 NS_198 0 6.0276502310352042e-05
GC_3_199 b_3 NI_3 NS_199 0 -4.9794891956701930e-05
GC_3_200 b_3 NI_3 NS_200 0 1.1982017633548768e-04
GC_3_201 b_3 NI_3 NS_201 0 1.3938970307412801e-04
GC_3_202 b_3 NI_3 NS_202 0 7.0034128345583809e-05
GC_3_203 b_3 NI_3 NS_203 0 3.3249792773291863e-08
GC_3_204 b_3 NI_3 NS_204 0 4.2541382642850515e-06
GC_3_205 b_3 NI_3 NS_205 0 -1.9651708590014324e-06
GC_3_206 b_3 NI_3 NS_206 0 8.5734784682591364e-08
GC_3_207 b_3 NI_3 NS_207 0 6.1371543351702125e-10
GC_3_208 b_3 NI_3 NS_208 0 -6.3978986292656802e-10
GC_3_209 b_3 NI_3 NS_209 0 -1.4671798310330668e-10
GC_3_210 b_3 NI_3 NS_210 0 -1.2237848164274736e-09
GC_3_211 b_3 NI_3 NS_211 0 5.4738142254738950e-05
GC_3_212 b_3 NI_3 NS_212 0 9.2112454947429774e-05
GC_3_213 b_3 NI_3 NS_213 0 2.8701181671316087e-07
GC_3_214 b_3 NI_3 NS_214 0 8.4903205062482310e-09
GC_3_215 b_3 NI_3 NS_215 0 -4.0119214570263636e-05
GC_3_216 b_3 NI_3 NS_216 0 -8.6005710790264226e-05
GC_3_217 b_3 NI_3 NS_217 0 -2.2672226251827820e-04
GC_3_218 b_3 NI_3 NS_218 0 9.6554307080355472e-05
GC_3_219 b_3 NI_3 NS_219 0 2.8122318367176512e-04
GC_3_220 b_3 NI_3 NS_220 0 1.5448269687313356e-04
GC_3_221 b_3 NI_3 NS_221 0 -3.0715716472208066e-04
GC_3_222 b_3 NI_3 NS_222 0 -2.0845982562297770e-04
GC_3_223 b_3 NI_3 NS_223 0 1.8399114315724541e-04
GC_3_224 b_3 NI_3 NS_224 0 3.9106493892931331e-04
GC_3_225 b_3 NI_3 NS_225 0 -9.4953716186659820e-05
GC_3_226 b_3 NI_3 NS_226 0 -1.5522812341873580e-04
GC_3_227 b_3 NI_3 NS_227 0 2.3741515441041042e-04
GC_3_228 b_3 NI_3 NS_228 0 2.1644233246770407e-04
GC_3_229 b_3 NI_3 NS_229 0 -5.9512661747001294e-05
GC_3_230 b_3 NI_3 NS_230 0 -2.0712465687151645e-04
GC_3_231 b_3 NI_3 NS_231 0 -2.1944906459053293e-06
GC_3_232 b_3 NI_3 NS_232 0 2.1430415344084327e-04
GC_3_233 b_3 NI_3 NS_233 0 -2.2385951198962805e-06
GC_3_234 b_3 NI_3 NS_234 0 6.4696319832445258e-08
GC_3_235 b_3 NI_3 NS_235 0 -4.6490700168098333e-07
GC_3_236 b_3 NI_3 NS_236 0 -4.5323122638434135e-07
GC_3_237 b_3 NI_3 NS_237 0 -7.2776868068408527e-10
GC_3_238 b_3 NI_3 NS_238 0 5.1680379588721952e-10
GC_3_239 b_3 NI_3 NS_239 0 1.4749278244528328e-10
GC_3_240 b_3 NI_3 NS_240 0 1.2209615790827941e-09
GC_3_241 b_3 NI_3 NS_241 0 -1.2017602622377574e-05
GC_3_242 b_3 NI_3 NS_242 0 4.3917202626908535e-07
GC_3_243 b_3 NI_3 NS_243 0 -2.5636464384690413e-08
GC_3_244 b_3 NI_3 NS_244 0 4.9337581068022287e-11
GC_3_245 b_3 NI_3 NS_245 0 -1.4663206633840265e-06
GC_3_246 b_3 NI_3 NS_246 0 -5.4509487118505087e-07
GC_3_247 b_3 NI_3 NS_247 0 -5.9487633602346990e-06
GC_3_248 b_3 NI_3 NS_248 0 2.4734450213973576e-06
GC_3_249 b_3 NI_3 NS_249 0 3.5848772826826232e-06
GC_3_250 b_3 NI_3 NS_250 0 1.3123316781799856e-05
GC_3_251 b_3 NI_3 NS_251 0 1.7633552096752774e-05
GC_3_252 b_3 NI_3 NS_252 0 1.5693730819128222e-06
GC_3_253 b_3 NI_3 NS_253 0 -1.8870594741350989e-06
GC_3_254 b_3 NI_3 NS_254 0 -1.5992004065328842e-05
GC_3_255 b_3 NI_3 NS_255 0 -4.9788853158623889e-06
GC_3_256 b_3 NI_3 NS_256 0 6.1974140408280859e-06
GC_3_257 b_3 NI_3 NS_257 0 1.1466516882034917e-05
GC_3_258 b_3 NI_3 NS_258 0 -6.6423527527889808e-07
GC_3_259 b_3 NI_3 NS_259 0 -3.8491871955770115e-07
GC_3_260 b_3 NI_3 NS_260 0 -1.0150638830138417e-05
GC_3_261 b_3 NI_3 NS_261 0 -3.8412894907652661e-06
GC_3_262 b_3 NI_3 NS_262 0 -1.7054666366948979e-06
GC_3_263 b_3 NI_3 NS_263 0 2.6625126058609800e-07
GC_3_264 b_3 NI_3 NS_264 0 9.8849098098793554e-08
GC_3_265 b_3 NI_3 NS_265 0 -1.4789729520445455e-08
GC_3_266 b_3 NI_3 NS_266 0 7.1362538897597923e-08
GC_3_267 b_3 NI_3 NS_267 0 1.4820035755027780e-10
GC_3_268 b_3 NI_3 NS_268 0 -3.5112421499616157e-11
GC_3_269 b_3 NI_3 NS_269 0 -6.6614191008634860e-11
GC_3_270 b_3 NI_3 NS_270 0 -2.6888833407031348e-10
GC_3_271 b_3 NI_3 NS_271 0 6.5825891513705958e-05
GC_3_272 b_3 NI_3 NS_272 0 -5.5593684677632027e-06
GC_3_273 b_3 NI_3 NS_273 0 3.0838598031295373e-08
GC_3_274 b_3 NI_3 NS_274 0 -1.4027711099414041e-10
GC_3_275 b_3 NI_3 NS_275 0 -2.7028171348269357e-06
GC_3_276 b_3 NI_3 NS_276 0 -1.1672689865501828e-06
GC_3_277 b_3 NI_3 NS_277 0 -4.9273589081516935e-06
GC_3_278 b_3 NI_3 NS_278 0 5.6497627019122873e-06
GC_3_279 b_3 NI_3 NS_279 0 9.6714840220185317e-06
GC_3_280 b_3 NI_3 NS_280 0 3.4362363515155606e-06
GC_3_281 b_3 NI_3 NS_281 0 -3.2948860225927133e-06
GC_3_282 b_3 NI_3 NS_282 0 -1.0812297997235533e-05
GC_3_283 b_3 NI_3 NS_283 0 -3.1204246287508559e-06
GC_3_284 b_3 NI_3 NS_284 0 -1.6758468453126991e-06
GC_3_285 b_3 NI_3 NS_285 0 -1.7488156366597079e-05
GC_3_286 b_3 NI_3 NS_286 0 -3.8613093728828136e-06
GC_3_287 b_3 NI_3 NS_287 0 -8.5222345623995185e-06
GC_3_288 b_3 NI_3 NS_288 0 1.4169312521207763e-05
GC_3_289 b_3 NI_3 NS_289 0 -7.0349684868613688e-06
GC_3_290 b_3 NI_3 NS_290 0 5.2061725462638876e-06
GC_3_291 b_3 NI_3 NS_291 0 -8.8717702006538550e-06
GC_3_292 b_3 NI_3 NS_292 0 1.0862361563844579e-05
GC_3_293 b_3 NI_3 NS_293 0 -5.7880790918862616e-07
GC_3_294 b_3 NI_3 NS_294 0 -6.3442370187768608e-08
GC_3_295 b_3 NI_3 NS_295 0 -3.7786182905142634e-08
GC_3_296 b_3 NI_3 NS_296 0 -2.6268891035065533e-07
GC_3_297 b_3 NI_3 NS_297 0 -1.5841789011023595e-10
GC_3_298 b_3 NI_3 NS_298 0 2.0132313187787053e-11
GC_3_299 b_3 NI_3 NS_299 0 6.8079753641076832e-11
GC_3_300 b_3 NI_3 NS_300 0 2.7024522741836943e-10
GC_3_301 b_3 NI_3 NS_301 0 1.7901683391939836e-05
GC_3_302 b_3 NI_3 NS_302 0 -2.5568014595303126e-06
GC_3_303 b_3 NI_3 NS_303 0 1.0257139039559033e-08
GC_3_304 b_3 NI_3 NS_304 0 -2.6532696844572411e-10
GC_3_305 b_3 NI_3 NS_305 0 -1.2423327534459854e-06
GC_3_306 b_3 NI_3 NS_306 0 -1.1108574190715826e-06
GC_3_307 b_3 NI_3 NS_307 0 -2.4790778225795314e-06
GC_3_308 b_3 NI_3 NS_308 0 5.4356147900346171e-07
GC_3_309 b_3 NI_3 NS_309 0 -1.2528111218071501e-06
GC_3_310 b_3 NI_3 NS_310 0 2.6650236151270064e-06
GC_3_311 b_3 NI_3 NS_311 0 1.8273669405964116e-06
GC_3_312 b_3 NI_3 NS_312 0 7.7991587334217560e-07
GC_3_313 b_3 NI_3 NS_313 0 -2.7635942949232997e-06
GC_3_314 b_3 NI_3 NS_314 0 -1.3704503509517564e-06
GC_3_315 b_3 NI_3 NS_315 0 -2.1566728526465934e-06
GC_3_316 b_3 NI_3 NS_316 0 3.4557465886562390e-06
GC_3_317 b_3 NI_3 NS_317 0 1.2689233611965959e-06
GC_3_318 b_3 NI_3 NS_318 0 2.3550489396651073e-06
GC_3_319 b_3 NI_3 NS_319 0 -9.0819751829936203e-07
GC_3_320 b_3 NI_3 NS_320 0 -3.9371809741033430e-07
GC_3_321 b_3 NI_3 NS_321 0 -3.2916088792914510e-06
GC_3_322 b_3 NI_3 NS_322 0 6.2256363987555933e-07
GC_3_323 b_3 NI_3 NS_323 0 -1.4055846380776007e-07
GC_3_324 b_3 NI_3 NS_324 0 -7.7795693281227011e-08
GC_3_325 b_3 NI_3 NS_325 0 2.3942272708108484e-08
GC_3_326 b_3 NI_3 NS_326 0 -5.0742625325521971e-08
GC_3_327 b_3 NI_3 NS_327 0 -1.7904003408457901e-11
GC_3_328 b_3 NI_3 NS_328 0 -1.0084237457694805e-10
GC_3_329 b_3 NI_3 NS_329 0 -3.8149508300604012e-11
GC_3_330 b_3 NI_3 NS_330 0 -1.6277829009824855e-10
GC_3_331 b_3 NI_3 NS_331 0 -3.1942315072336629e-05
GC_3_332 b_3 NI_3 NS_332 0 3.5545369002805564e-06
GC_3_333 b_3 NI_3 NS_333 0 -1.3272797153789374e-08
GC_3_334 b_3 NI_3 NS_334 0 3.4691757974356507e-10
GC_3_335 b_3 NI_3 NS_335 0 2.0364670298846815e-06
GC_3_336 b_3 NI_3 NS_336 0 2.9512198655430224e-07
GC_3_337 b_3 NI_3 NS_337 0 1.7829865509264036e-06
GC_3_338 b_3 NI_3 NS_338 0 -1.7976012084968925e-06
GC_3_339 b_3 NI_3 NS_339 0 2.2339251346981760e-06
GC_3_340 b_3 NI_3 NS_340 0 -1.9710652533886366e-06
GC_3_341 b_3 NI_3 NS_341 0 1.2218455895156565e-06
GC_3_342 b_3 NI_3 NS_342 0 -1.5034943224834136e-06
GC_3_343 b_3 NI_3 NS_343 0 1.6567993256610509e-06
GC_3_344 b_3 NI_3 NS_344 0 -1.3902509339825437e-06
GC_3_345 b_3 NI_3 NS_345 0 1.7716180769555136e-06
GC_3_346 b_3 NI_3 NS_346 0 -3.2805698815984926e-06
GC_3_347 b_3 NI_3 NS_347 0 1.9903680886095316e-06
GC_3_348 b_3 NI_3 NS_348 0 -3.6368214863882628e-06
GC_3_349 b_3 NI_3 NS_349 0 7.3352828664693958e-07
GC_3_350 b_3 NI_3 NS_350 0 -3.3032757435453469e-06
GC_3_351 b_3 NI_3 NS_351 0 3.4149821357894885e-06
GC_3_352 b_3 NI_3 NS_352 0 -1.5015847156298875e-06
GC_3_353 b_3 NI_3 NS_353 0 2.6974185792305801e-07
GC_3_354 b_3 NI_3 NS_354 0 3.1441944318786620e-08
GC_3_355 b_3 NI_3 NS_355 0 1.3484806677803301e-08
GC_3_356 b_3 NI_3 NS_356 0 1.2312561565015122e-07
GC_3_357 b_3 NI_3 NS_357 0 2.5347160353453281e-11
GC_3_358 b_3 NI_3 NS_358 0 1.2044965500239512e-10
GC_3_359 b_3 NI_3 NS_359 0 3.7594583543093844e-11
GC_3_360 b_3 NI_3 NS_360 0 1.6468103053449742e-10
GD_3_1 b_3 NI_3 NA_1 0 1.6053745417191803e-02
GD_3_2 b_3 NI_3 NA_2 0 -9.1340177342169774e-05
GD_3_3 b_3 NI_3 NA_3 0 -4.0270206208655776e-02
GD_3_4 b_3 NI_3 NA_4 0 -9.9682735972884962e-03
GD_3_5 b_3 NI_3 NA_5 0 2.3300350421506378e-03
GD_3_6 b_3 NI_3 NA_6 0 -4.6783139508794080e-05
GD_3_7 b_3 NI_3 NA_7 0 1.7128697648621010e-04
GD_3_8 b_3 NI_3 NA_8 0 -6.2842245982104374e-05
GD_3_9 b_3 NI_3 NA_9 0 -1.1548347624455805e-06
GD_3_10 b_3 NI_3 NA_10 0 -9.0627077179041734e-06
GD_3_11 b_3 NI_3 NA_11 0 -1.6971830497440935e-06
GD_3_12 b_3 NI_3 NA_12 0 7.7454572573918705e-06
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 1.3559977266702022e-03
GC_4_2 b_4 NI_4 NS_2 0 -1.2038876436080150e-03
GC_4_3 b_4 NI_4 NS_3 0 3.7357899062390004e-06
GC_4_4 b_4 NI_4 NS_4 0 2.8902025643847683e-07
GC_4_5 b_4 NI_4 NS_5 0 1.2297103897685650e-04
GC_4_6 b_4 NI_4 NS_6 0 8.9417681564551163e-04
GC_4_7 b_4 NI_4 NS_7 0 1.8425181613924266e-03
GC_4_8 b_4 NI_4 NS_8 0 -8.6745204795826193e-04
GC_4_9 b_4 NI_4 NS_9 0 -2.9665984448669185e-03
GC_4_10 b_4 NI_4 NS_10 0 -1.6486215866960755e-03
GC_4_11 b_4 NI_4 NS_11 0 2.2194995090952458e-03
GC_4_12 b_4 NI_4 NS_12 0 2.6689300497430980e-03
GC_4_13 b_4 NI_4 NS_13 0 -1.4401272077439915e-03
GC_4_14 b_4 NI_4 NS_14 0 -2.9129239481868485e-03
GC_4_15 b_4 NI_4 NS_15 0 1.0698835745811112e-03
GC_4_16 b_4 NI_4 NS_16 0 2.2566924764740206e-03
GC_4_17 b_4 NI_4 NS_17 0 -1.6275425023295667e-03
GC_4_18 b_4 NI_4 NS_18 0 -2.1363730378474630e-03
GC_4_19 b_4 NI_4 NS_19 0 4.2046566768488711e-04
GC_4_20 b_4 NI_4 NS_20 0 2.0118498158381028e-03
GC_4_21 b_4 NI_4 NS_21 0 2.1508326771051717e-04
GC_4_22 b_4 NI_4 NS_22 0 -2.1102726803271040e-03
GC_4_23 b_4 NI_4 NS_23 0 -4.3290758021995981e-06
GC_4_24 b_4 NI_4 NS_24 0 4.3528691030463468e-06
GC_4_25 b_4 NI_4 NS_25 0 -7.8953772070042473e-07
GC_4_26 b_4 NI_4 NS_26 0 -3.5250190153895121e-06
GC_4_27 b_4 NI_4 NS_27 0 -7.5479910794354111e-09
GC_4_28 b_4 NI_4 NS_28 0 2.2567545206178911e-08
GC_4_29 b_4 NI_4 NS_29 0 2.3359230281106339e-09
GC_4_30 b_4 NI_4 NS_30 0 1.5101849077686995e-09
GC_4_31 b_4 NI_4 NS_31 0 -5.5801074599777880e-04
GC_4_32 b_4 NI_4 NS_32 0 -2.9007616243612875e-03
GC_4_33 b_4 NI_4 NS_33 0 -6.1510250246002188e-06
GC_4_34 b_4 NI_4 NS_34 0 -3.8641528467944275e-07
GC_4_35 b_4 NI_4 NS_35 0 2.6869528711998660e-03
GC_4_36 b_4 NI_4 NS_36 0 -1.9871035345229893e-03
GC_4_37 b_4 NI_4 NS_37 0 -6.1985251461633053e-03
GC_4_38 b_4 NI_4 NS_38 0 1.7528631976828446e-03
GC_4_39 b_4 NI_4 NS_39 0 4.7654008991423269e-03
GC_4_40 b_4 NI_4 NS_40 0 -5.5287242487402121e-03
GC_4_41 b_4 NI_4 NS_41 0 -2.4763103516912976e-04
GC_4_42 b_4 NI_4 NS_42 0 7.2490216894870972e-03
GC_4_43 b_4 NI_4 NS_43 0 -6.3151021330279441e-03
GC_4_44 b_4 NI_4 NS_44 0 -5.0558253063733658e-03
GC_4_45 b_4 NI_4 NS_45 0 4.5028162175496898e-03
GC_4_46 b_4 NI_4 NS_46 0 -1.7122915625266630e-03
GC_4_47 b_4 NI_4 NS_47 0 -5.9096753127079653e-04
GC_4_48 b_4 NI_4 NS_48 0 6.9470776364957331e-03
GC_4_49 b_4 NI_4 NS_49 0 -3.4358105681654414e-03
GC_4_50 b_4 NI_4 NS_50 0 -3.6826697955017469e-03
GC_4_51 b_4 NI_4 NS_51 0 5.9256580380445600e-03
GC_4_52 b_4 NI_4 NS_52 0 3.9686148945753216e-04
GC_4_53 b_4 NI_4 NS_53 0 6.3856041306214559e-05
GC_4_54 b_4 NI_4 NS_54 0 8.4381967260811374e-06
GC_4_55 b_4 NI_4 NS_55 0 1.5113680856155398e-05
GC_4_56 b_4 NI_4 NS_56 0 3.9976674193447948e-05
GC_4_57 b_4 NI_4 NS_57 0 7.1156028022573029e-09
GC_4_58 b_4 NI_4 NS_58 0 -2.9351516618504965e-08
GC_4_59 b_4 NI_4 NS_59 0 -1.8855648137956497e-09
GC_4_60 b_4 NI_4 NS_60 0 -5.6002683984500131e-10
GC_4_61 b_4 NI_4 NS_61 0 -7.5349046462616531e-02
GC_4_62 b_4 NI_4 NS_62 0 2.4900050708905077e-02
GC_4_63 b_4 NI_4 NS_63 0 1.9199962318260712e-05
GC_4_64 b_4 NI_4 NS_64 0 5.3863163438985055e-06
GC_4_65 b_4 NI_4 NS_65 0 1.8353498951985608e-02
GC_4_66 b_4 NI_4 NS_66 0 2.7965358958527108e-02
GC_4_67 b_4 NI_4 NS_67 0 -1.9176261647186877e-02
GC_4_68 b_4 NI_4 NS_68 0 8.3761042118018231e-03
GC_4_69 b_4 NI_4 NS_69 0 -5.5264909658227172e-03
GC_4_70 b_4 NI_4 NS_70 0 -2.3054144747732746e-02
GC_4_71 b_4 NI_4 NS_71 0 2.6687341735551758e-02
GC_4_72 b_4 NI_4 NS_72 0 -1.4576107326727759e-02
GC_4_73 b_4 NI_4 NS_73 0 3.4517302312567943e-02
GC_4_74 b_4 NI_4 NS_74 0 4.8628324083679958e-03
GC_4_75 b_4 NI_4 NS_75 0 9.6719812426988173e-03
GC_4_76 b_4 NI_4 NS_76 0 1.3692421813373457e-02
GC_4_77 b_4 NI_4 NS_77 0 -1.2370876643545995e-02
GC_4_78 b_4 NI_4 NS_78 0 1.1007946209698851e-02
GC_4_79 b_4 NI_4 NS_79 0 -1.1774521606281275e-02
GC_4_80 b_4 NI_4 NS_80 0 -1.2014122209594739e-02
GC_4_81 b_4 NI_4 NS_81 0 1.9793935530302727e-02
GC_4_82 b_4 NI_4 NS_82 0 -2.6023932276003539e-02
GC_4_83 b_4 NI_4 NS_83 0 9.6721681928538489e-04
GC_4_84 b_4 NI_4 NS_84 0 -1.0822028982411520e-03
GC_4_85 b_4 NI_4 NS_85 0 6.3094412014810504e-04
GC_4_86 b_4 NI_4 NS_86 0 3.4914596489023247e-04
GC_4_87 b_4 NI_4 NS_87 0 9.7107874919784162e-08
GC_4_88 b_4 NI_4 NS_88 0 4.1868767422817641e-07
GC_4_89 b_4 NI_4 NS_89 0 -1.0314558722745683e-08
GC_4_90 b_4 NI_4 NS_90 0 -1.9789138220718205e-08
GC_4_91 b_4 NI_4 NS_91 0 1.2659768848160127e-01
GC_4_92 b_4 NI_4 NS_92 0 -9.9682227254338108e-03
GC_4_93 b_4 NI_4 NS_93 0 -2.0418483468457034e-05
GC_4_94 b_4 NI_4 NS_94 0 -3.8273614983901288e-06
GC_4_95 b_4 NI_4 NS_95 0 -8.0908262368300562e-03
GC_4_96 b_4 NI_4 NS_96 0 6.4296865047940542e-04
GC_4_97 b_4 NI_4 NS_97 0 -1.9909408466115626e-03
GC_4_98 b_4 NI_4 NS_98 0 6.7356143800919777e-05
GC_4_99 b_4 NI_4 NS_99 0 -1.2598719640679377e-02
GC_4_100 b_4 NI_4 NS_100 0 8.2477800777836716e-03
GC_4_101 b_4 NI_4 NS_101 0 -1.0271311615499336e-02
GC_4_102 b_4 NI_4 NS_102 0 -6.2357295410835653e-04
GC_4_103 b_4 NI_4 NS_103 0 -3.5565617083853415e-03
GC_4_104 b_4 NI_4 NS_104 0 1.6966131517386220e-02
GC_4_105 b_4 NI_4 NS_105 0 -7.7825903588610371e-03
GC_4_106 b_4 NI_4 NS_106 0 1.3370076548945802e-02
GC_4_107 b_4 NI_4 NS_107 0 -3.9902897788399094e-03
GC_4_108 b_4 NI_4 NS_108 0 6.9628713158745156e-03
GC_4_109 b_4 NI_4 NS_109 0 -2.7633627349993679e-03
GC_4_110 b_4 NI_4 NS_110 0 1.2313497559275613e-02
GC_4_111 b_4 NI_4 NS_111 0 -2.2964005253819381e-02
GC_4_112 b_4 NI_4 NS_112 0 5.9629952375129681e-03
GC_4_113 b_4 NI_4 NS_113 0 -8.6294474345638720e-04
GC_4_114 b_4 NI_4 NS_114 0 8.0344033683356440e-04
GC_4_115 b_4 NI_4 NS_115 0 -5.1358560300163484e-04
GC_4_116 b_4 NI_4 NS_116 0 -4.3937271563943139e-04
GC_4_117 b_4 NI_4 NS_117 0 -6.4174241182781336e-08
GC_4_118 b_4 NI_4 NS_118 0 -1.9155149919510674e-07
GC_4_119 b_4 NI_4 NS_119 0 -3.0939598424237513e-09
GC_4_120 b_4 NI_4 NS_120 0 5.6381472190783786e-09
GC_4_121 b_4 NI_4 NS_121 0 9.8190999365470170e-04
GC_4_122 b_4 NI_4 NS_122 0 -3.4563276797592874e-04
GC_4_123 b_4 NI_4 NS_123 0 2.1362724149492189e-06
GC_4_124 b_4 NI_4 NS_124 0 8.2060295954657066e-08
GC_4_125 b_4 NI_4 NS_125 0 1.1626324618156408e-05
GC_4_126 b_4 NI_4 NS_126 0 8.7329047514957603e-05
GC_4_127 b_4 NI_4 NS_127 0 3.1565129829292375e-04
GC_4_128 b_4 NI_4 NS_128 0 -1.1550920442199955e-04
GC_4_129 b_4 NI_4 NS_129 0 -5.1916494373669493e-04
GC_4_130 b_4 NI_4 NS_130 0 -2.4271238347770273e-04
GC_4_131 b_4 NI_4 NS_131 0 3.2788951534158656e-04
GC_4_132 b_4 NI_4 NS_132 0 3.8892142575564474e-04
GC_4_133 b_4 NI_4 NS_133 0 -3.2494336485631618e-04
GC_4_134 b_4 NI_4 NS_134 0 -5.5985364423068835e-04
GC_4_135 b_4 NI_4 NS_135 0 7.3996224834266643e-05
GC_4_136 b_4 NI_4 NS_136 0 3.8462470602018640e-04
GC_4_137 b_4 NI_4 NS_137 0 -3.5599393315827453e-04
GC_4_138 b_4 NI_4 NS_138 0 -2.6837281393180456e-04
GC_4_139 b_4 NI_4 NS_139 0 5.3984170047230257e-06
GC_4_140 b_4 NI_4 NS_140 0 4.0799729102666197e-04
GC_4_141 b_4 NI_4 NS_141 0 -9.5062216868778028e-05
GC_4_142 b_4 NI_4 NS_142 0 -3.4082775221454031e-04
GC_4_143 b_4 NI_4 NS_143 0 -1.4810484611842172e-05
GC_4_144 b_4 NI_4 NS_144 0 -8.4933391475198244e-06
GC_4_145 b_4 NI_4 NS_145 0 2.7402888364563581e-06
GC_4_146 b_4 NI_4 NS_146 0 -6.6705469041913801e-06
GC_4_147 b_4 NI_4 NS_147 0 -7.7197156531262780e-09
GC_4_148 b_4 NI_4 NS_148 0 4.8070271996862157e-09
GC_4_149 b_4 NI_4 NS_149 0 1.1496194839768802e-09
GC_4_150 b_4 NI_4 NS_150 0 2.7805417329037762e-09
GC_4_151 b_4 NI_4 NS_151 0 2.2663492400766209e-03
GC_4_152 b_4 NI_4 NS_152 0 -7.3264017963937142e-04
GC_4_153 b_4 NI_4 NS_153 0 -1.8147155500414763e-06
GC_4_154 b_4 NI_4 NS_154 0 -1.2100169703973776e-07
GC_4_155 b_4 NI_4 NS_155 0 3.5969873324481088e-04
GC_4_156 b_4 NI_4 NS_156 0 -3.7511994252593044e-04
GC_4_157 b_4 NI_4 NS_157 0 -1.2776615397505217e-03
GC_4_158 b_4 NI_4 NS_158 0 3.4323472019691842e-04
GC_4_159 b_4 NI_4 NS_159 0 7.1255517818764197e-04
GC_4_160 b_4 NI_4 NS_160 0 -8.2803185444848117e-04
GC_4_161 b_4 NI_4 NS_161 0 -1.5013266752816177e-04
GC_4_162 b_4 NI_4 NS_162 0 1.3911134446684878e-03
GC_4_163 b_4 NI_4 NS_163 0 -1.3011316374249946e-03
GC_4_164 b_4 NI_4 NS_164 0 -7.6474272164763640e-04
GC_4_165 b_4 NI_4 NS_165 0 6.8662633234903097e-04
GC_4_166 b_4 NI_4 NS_166 0 -2.8643590712986572e-05
GC_4_167 b_4 NI_4 NS_167 0 -1.3691314138972424e-04
GC_4_168 b_4 NI_4 NS_168 0 1.4682073596504041e-03
GC_4_169 b_4 NI_4 NS_169 0 -7.1833247192052709e-04
GC_4_170 b_4 NI_4 NS_170 0 -5.4307221124773016e-04
GC_4_171 b_4 NI_4 NS_171 0 6.5097302056588743e-04
GC_4_172 b_4 NI_4 NS_172 0 1.9308955012913460e-04
GC_4_173 b_4 NI_4 NS_173 0 -3.0134567075054201e-06
GC_4_174 b_4 NI_4 NS_174 0 2.6008719631690913e-05
GC_4_175 b_4 NI_4 NS_175 0 -9.9186048049613420e-06
GC_4_176 b_4 NI_4 NS_176 0 -1.4227993878084345e-06
GC_4_177 b_4 NI_4 NS_177 0 7.0599521133360487e-09
GC_4_178 b_4 NI_4 NS_178 0 -1.0479962193339793e-08
GC_4_179 b_4 NI_4 NS_179 0 -6.2224207883282683e-10
GC_4_180 b_4 NI_4 NS_180 0 -2.1193958533872466e-09
GC_4_181 b_4 NI_4 NS_181 0 5.4748275500487317e-05
GC_4_182 b_4 NI_4 NS_182 0 9.2111712053107042e-05
GC_4_183 b_4 NI_4 NS_183 0 2.8701248701860402e-07
GC_4_184 b_4 NI_4 NS_184 0 8.4903050297255276e-09
GC_4_185 b_4 NI_4 NS_185 0 -4.0119717034990485e-05
GC_4_186 b_4 NI_4 NS_186 0 -8.6005427386109292e-05
GC_4_187 b_4 NI_4 NS_187 0 -2.2672225796667981e-04
GC_4_188 b_4 NI_4 NS_188 0 9.6553933990898492e-05
GC_4_189 b_4 NI_4 NS_189 0 2.8122159853187804e-04
GC_4_190 b_4 NI_4 NS_190 0 1.5448308138105325e-04
GC_4_191 b_4 NI_4 NS_191 0 -3.0715791441192336e-04
GC_4_192 b_4 NI_4 NS_192 0 -2.0845896043177292e-04
GC_4_193 b_4 NI_4 NS_193 0 1.8399026107378242e-04
GC_4_194 b_4 NI_4 NS_194 0 3.9106521815177861e-04
GC_4_195 b_4 NI_4 NS_195 0 -9.4954356384519686e-05
GC_4_196 b_4 NI_4 NS_196 0 -1.5522559155525109e-04
GC_4_197 b_4 NI_4 NS_197 0 2.3741529674039684e-04
GC_4_198 b_4 NI_4 NS_198 0 2.1644331571273046e-04
GC_4_199 b_4 NI_4 NS_199 0 -5.9513295464940577e-05
GC_4_200 b_4 NI_4 NS_200 0 -2.0712363327951932e-04
GC_4_201 b_4 NI_4 NS_201 0 -2.1951623178621124e-06
GC_4_202 b_4 NI_4 NS_202 0 2.1430507822037460e-04
GC_4_203 b_4 NI_4 NS_203 0 -2.2386607227584789e-06
GC_4_204 b_4 NI_4 NS_204 0 6.4753763987386544e-08
GC_4_205 b_4 NI_4 NS_205 0 -4.6493723018620398e-07
GC_4_206 b_4 NI_4 NS_206 0 -4.5326362444998958e-07
GC_4_207 b_4 NI_4 NS_207 0 -7.2777010751582435e-10
GC_4_208 b_4 NI_4 NS_208 0 5.1680156730104860e-10
GC_4_209 b_4 NI_4 NS_209 0 1.4749280946134943e-10
GC_4_210 b_4 NI_4 NS_210 0 1.2209615416459595e-09
GC_4_211 b_4 NI_4 NS_211 0 1.3848393088197942e-04
GC_4_212 b_4 NI_4 NS_212 0 1.3826450016982999e-06
GC_4_213 b_4 NI_4 NS_213 0 -2.0149254752494797e-07
GC_4_214 b_4 NI_4 NS_214 0 -9.3083372698525652e-09
GC_4_215 b_4 NI_4 NS_215 0 4.9978472404074885e-05
GC_4_216 b_4 NI_4 NS_216 0 -1.9598857449514031e-06
GC_4_217 b_4 NI_4 NS_217 0 2.5680848674533730e-05
GC_4_218 b_4 NI_4 NS_218 0 -7.5195352630806116e-06
GC_4_219 b_4 NI_4 NS_219 0 2.2272049107698274e-05
GC_4_220 b_4 NI_4 NS_220 0 -2.6882874601804365e-04
GC_4_221 b_4 NI_4 NS_221 0 -2.9200588247558758e-04
GC_4_222 b_4 NI_4 NS_222 0 4.0810790293972405e-05
GC_4_223 b_4 NI_4 NS_223 0 -5.4965812311936194e-05
GC_4_224 b_4 NI_4 NS_224 0 2.2142104820023655e-04
GC_4_225 b_4 NI_4 NS_225 0 1.6790676995051836e-04
GC_4_226 b_4 NI_4 NS_226 0 -1.0526825956219975e-04
GC_4_227 b_4 NI_4 NS_227 0 -1.8088182198440516e-04
GC_4_228 b_4 NI_4 NS_228 0 6.1686549046416708e-05
GC_4_229 b_4 NI_4 NS_229 0 -5.0481355937145995e-05
GC_4_230 b_4 NI_4 NS_230 0 1.2078608421046147e-04
GC_4_231 b_4 NI_4 NS_231 0 1.3701556669134230e-04
GC_4_232 b_4 NI_4 NS_232 0 7.0686012430378389e-05
GC_4_233 b_4 NI_4 NS_233 0 -1.0585899887850897e-07
GC_4_234 b_4 NI_4 NS_234 0 4.3444543621580961e-06
GC_4_235 b_4 NI_4 NS_235 0 -2.0219892617724642e-06
GC_4_236 b_4 NI_4 NS_236 0 1.8441426281312162e-08
GC_4_237 b_4 NI_4 NS_237 0 6.0917257188967162e-10
GC_4_238 b_4 NI_4 NS_238 0 -6.4486073250166914e-10
GC_4_239 b_4 NI_4 NS_239 0 -1.4660653939035876e-10
GC_4_240 b_4 NI_4 NS_240 0 -1.2238416602021871e-09
GC_4_241 b_4 NI_4 NS_241 0 6.6256704782338525e-05
GC_4_242 b_4 NI_4 NS_242 0 -5.6124273705929551e-06
GC_4_243 b_4 NI_4 NS_243 0 3.0931090795227231e-08
GC_4_244 b_4 NI_4 NS_244 0 -1.4166221354264636e-10
GC_4_245 b_4 NI_4 NS_245 0 -2.7183688476798192e-06
GC_4_246 b_4 NI_4 NS_246 0 -1.1809898579077868e-06
GC_4_247 b_4 NI_4 NS_247 0 -4.9372986987460440e-06
GC_4_248 b_4 NI_4 NS_248 0 5.6220223569934645e-06
GC_4_249 b_4 NI_4 NS_249 0 9.6526166152277768e-06
GC_4_250 b_4 NI_4 NS_250 0 3.4537878604461652e-06
GC_4_251 b_4 NI_4 NS_251 0 -3.3260945440092885e-06
GC_4_252 b_4 NI_4 NS_252 0 -1.0830891410264642e-05
GC_4_253 b_4 NI_4 NS_253 0 -3.1844543716836622e-06
GC_4_254 b_4 NI_4 NS_254 0 -1.6471618457476845e-06
GC_4_255 b_4 NI_4 NS_255 0 -1.7516679419389536e-05
GC_4_256 b_4 NI_4 NS_256 0 -3.8364715831123949e-06
GC_4_257 b_4 NI_4 NS_257 0 -8.5579003325221651e-06
GC_4_258 b_4 NI_4 NS_258 0 1.4206941889774643e-05
GC_4_259 b_4 NI_4 NS_259 0 -7.0646554803662881e-06
GC_4_260 b_4 NI_4 NS_260 0 5.2325198035238452e-06
GC_4_261 b_4 NI_4 NS_261 0 -8.9556861729502751e-06
GC_4_262 b_4 NI_4 NS_262 0 1.0881313074297142e-05
GC_4_263 b_4 NI_4 NS_263 0 -5.8293540085292760e-07
GC_4_264 b_4 NI_4 NS_264 0 -6.0298293263903377e-08
GC_4_265 b_4 NI_4 NS_265 0 -3.9873529413292808e-08
GC_4_266 b_4 NI_4 NS_266 0 -2.6482637929326490e-07
GC_4_267 b_4 NI_4 NS_267 0 -1.5857049041594667e-10
GC_4_268 b_4 NI_4 NS_268 0 1.9903933077555555e-11
GC_4_269 b_4 NI_4 NS_269 0 6.8097742761519369e-11
GC_4_270 b_4 NI_4 NS_270 0 2.7026123815119156e-10
GC_4_271 b_4 NI_4 NS_271 0 -1.2017262780358764e-05
GC_4_272 b_4 NI_4 NS_272 0 4.3913093417956436e-07
GC_4_273 b_4 NI_4 NS_273 0 -2.5636372905260088e-08
GC_4_274 b_4 NI_4 NS_274 0 4.9336614949738579e-11
GC_4_275 b_4 NI_4 NS_275 0 -1.4663436336132777e-06
GC_4_276 b_4 NI_4 NS_276 0 -5.4508427484617660e-07
GC_4_277 b_4 NI_4 NS_277 0 -5.9487779151976121e-06
GC_4_278 b_4 NI_4 NS_278 0 2.4734516617288765e-06
GC_4_279 b_4 NI_4 NS_279 0 3.5848581235509793e-06
GC_4_280 b_4 NI_4 NS_280 0 1.3123341739084130e-05
GC_4_281 b_4 NI_4 NS_281 0 1.7633528732675042e-05
GC_4_282 b_4 NI_4 NS_282 0 1.5693913643780166e-06
GC_4_283 b_4 NI_4 NS_283 0 -1.8870706510097454e-06
GC_4_284 b_4 NI_4 NS_284 0 -1.5991965655372383e-05
GC_4_285 b_4 NI_4 NS_285 0 -4.9788798257646478e-06
GC_4_286 b_4 NI_4 NS_286 0 6.1974437392069866e-06
GC_4_287 b_4 NI_4 NS_287 0 1.1466512972220433e-05
GC_4_288 b_4 NI_4 NS_288 0 -6.6421532169824602e-07
GC_4_289 b_4 NI_4 NS_289 0 -3.8493444823072789e-07
GC_4_290 b_4 NI_4 NS_290 0 -1.0150630316590273e-05
GC_4_291 b_4 NI_4 NS_291 0 -3.8413498438681415e-06
GC_4_292 b_4 NI_4 NS_292 0 -1.7054593190541120e-06
GC_4_293 b_4 NI_4 NS_293 0 2.6624763081564505e-07
GC_4_294 b_4 NI_4 NS_294 0 9.8851575228242991e-08
GC_4_295 b_4 NI_4 NS_295 0 -1.4791292705375124e-08
GC_4_296 b_4 NI_4 NS_296 0 7.1360551376685940e-08
GC_4_297 b_4 NI_4 NS_297 0 1.4820020789333931e-10
GC_4_298 b_4 NI_4 NS_298 0 -3.5112530526918983e-11
GC_4_299 b_4 NI_4 NS_299 0 -6.6614212516923096e-11
GC_4_300 b_4 NI_4 NS_300 0 -2.6888835790607818e-10
GC_4_301 b_4 NI_4 NS_301 0 -3.1941709615194003e-05
GC_4_302 b_4 NI_4 NS_302 0 3.5544762558064761e-06
GC_4_303 b_4 NI_4 NS_303 0 -1.3272659813696286e-08
GC_4_304 b_4 NI_4 NS_304 0 3.4691406679945140e-10
GC_4_305 b_4 NI_4 NS_305 0 2.0364022761505049e-06
GC_4_306 b_4 NI_4 NS_306 0 2.9506704211061977e-07
GC_4_307 b_4 NI_4 NS_307 0 1.7829378320922602e-06
GC_4_308 b_4 NI_4 NS_308 0 -1.7976020546785272e-06
GC_4_309 b_4 NI_4 NS_309 0 2.2338177776627805e-06
GC_4_310 b_4 NI_4 NS_310 0 -1.9709266593095548e-06
GC_4_311 b_4 NI_4 NS_311 0 1.2218262728179620e-06
GC_4_312 b_4 NI_4 NS_312 0 -1.5034225397465892e-06
GC_4_313 b_4 NI_4 NS_313 0 1.6567931372790353e-06
GC_4_314 b_4 NI_4 NS_314 0 -1.3901781948702357e-06
GC_4_315 b_4 NI_4 NS_315 0 1.7716545670443709e-06
GC_4_316 b_4 NI_4 NS_316 0 -3.2805214595957028e-06
GC_4_317 b_4 NI_4 NS_317 0 1.9903583895526049e-06
GC_4_318 b_4 NI_4 NS_318 0 -3.6367828456687892e-06
GC_4_319 b_4 NI_4 NS_319 0 7.3350442361600154e-07
GC_4_320 b_4 NI_4 NS_320 0 -3.3032497007314505e-06
GC_4_321 b_4 NI_4 NS_321 0 3.4148903294441744e-06
GC_4_322 b_4 NI_4 NS_322 0 -1.5015526483621118e-06
GC_4_323 b_4 NI_4 NS_323 0 2.6973770729350292e-07
GC_4_324 b_4 NI_4 NS_324 0 3.1444604385075089e-08
GC_4_325 b_4 NI_4 NS_325 0 1.3483178619824344e-08
GC_4_326 b_4 NI_4 NS_326 0 1.2312365042139022e-07
GC_4_327 b_4 NI_4 NS_327 0 2.5346957051249125e-11
GC_4_328 b_4 NI_4 NS_328 0 1.2044891685038952e-10
GC_4_329 b_4 NI_4 NS_329 0 3.7594671267634705e-11
GC_4_330 b_4 NI_4 NS_330 0 1.6468111637915960e-10
GC_4_331 b_4 NI_4 NS_331 0 1.8113430302228979e-05
GC_4_332 b_4 NI_4 NS_332 0 -2.5825692430325210e-06
GC_4_333 b_4 NI_4 NS_333 0 1.0317756114455756e-08
GC_4_334 b_4 NI_4 NS_334 0 -2.6663560478129995e-10
GC_4_335 b_4 NI_4 NS_335 0 -1.2543602284430799e-06
GC_4_336 b_4 NI_4 NS_336 0 -1.1114241245212727e-06
GC_4_337 b_4 NI_4 NS_337 0 -2.4906503821511758e-06
GC_4_338 b_4 NI_4 NS_338 0 5.3778958607147823e-07
GC_4_339 b_4 NI_4 NS_339 0 -1.2738987908451755e-06
GC_4_340 b_4 NI_4 NS_340 0 2.6842757648173644e-06
GC_4_341 b_4 NI_4 NS_341 0 1.8130844990356743e-06
GC_4_342 b_4 NI_4 NS_342 0 7.9201541686079354e-07
GC_4_343 b_4 NI_4 NS_343 0 -2.7645306722504840e-06
GC_4_344 b_4 NI_4 NS_344 0 -1.3551197428563171e-06
GC_4_345 b_4 NI_4 NS_345 0 -2.1678155432626801e-06
GC_4_346 b_4 NI_4 NS_346 0 3.4714091903030629e-06
GC_4_347 b_4 NI_4 NS_347 0 1.2584624740127084e-06
GC_4_348 b_4 NI_4 NS_348 0 2.3719290211840732e-06
GC_4_349 b_4 NI_4 NS_349 0 -9.1723703482140815e-07
GC_4_350 b_4 NI_4 NS_350 0 -3.8008705975106569e-07
GC_4_351 b_4 NI_4 NS_351 0 -3.3257346719917357e-06
GC_4_352 b_4 NI_4 NS_352 0 6.2805334174153310e-07
GC_4_353 b_4 NI_4 NS_353 0 -1.4282103217836559e-07
GC_4_354 b_4 NI_4 NS_354 0 -7.6712430003939633e-08
GC_4_355 b_4 NI_4 NS_355 0 2.3256076133010276e-08
GC_4_356 b_4 NI_4 NS_356 0 -5.1807329263716241e-08
GC_4_357 b_4 NI_4 NS_357 0 -1.7982957075372901e-11
GC_4_358 b_4 NI_4 NS_358 0 -1.0110893089282082e-10
GC_4_359 b_4 NI_4 NS_359 0 -3.8114121570143458e-11
GC_4_360 b_4 NI_4 NS_360 0 -1.6273680829229972e-10
GD_4_1 b_4 NI_4 NA_1 0 -9.1324786499264325e-05
GD_4_2 b_4 NI_4 NA_2 0 1.6056004849540367e-02
GD_4_3 b_4 NI_4 NA_3 0 -9.9681698811546673e-03
GD_4_4 b_4 NI_4 NA_4 0 -4.0270206208655887e-02
GD_4_5 b_4 NI_4 NA_5 0 -4.6772755112167041e-05
GD_4_6 b_4 NI_4 NA_6 0 2.3298014152276958e-03
GD_4_7 b_4 NI_4 NA_7 0 -6.2844767913684731e-05
GD_4_8 b_4 NI_4 NA_8 0 1.6924455739742713e-04
GD_4_9 b_4 NI_4 NA_9 0 -9.0925705668893068e-06
GD_4_10 b_4 NI_4 NA_10 0 -1.1549172007867563e-06
GD_4_11 b_4 NI_4 NA_11 0 7.7453325151464186e-06
GD_4_12 b_4 NI_4 NA_12 0 -1.7302922205302330e-06
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 1.2794855363909669e-04
GC_5_2 b_5 NI_5 NS_2 0 2.8895180758200148e-06
GC_5_3 b_5 NI_5 NS_3 0 -2.0789759302606578e-07
GC_5_4 b_5 NI_5 NS_4 0 -9.2148620618220835e-09
GC_5_5 b_5 NI_5 NS_5 0 5.0391238670461804e-05
GC_5_6 b_5 NI_5 NS_6 0 -1.8561640353577073e-06
GC_5_7 b_5 NI_5 NS_7 0 2.6276469901156174e-05
GC_5_8 b_5 NI_5 NS_8 0 -7.5099482509492870e-06
GC_5_9 b_5 NI_5 NS_9 0 2.3050776556802502e-05
GC_5_10 b_5 NI_5 NS_10 0 -2.6914133545999992e-04
GC_5_11 b_5 NI_5 NS_11 0 -2.9117457354196398e-04
GC_5_12 b_5 NI_5 NS_12 0 4.0238017546484322e-05
GC_5_13 b_5 NI_5 NS_13 0 -5.4545162114372599e-05
GC_5_14 b_5 NI_5 NS_14 0 2.2062130341976441e-04
GC_5_15 b_5 NI_5 NS_15 0 1.6841453138073120e-04
GC_5_16 b_5 NI_5 NS_16 0 -1.0598925855322593e-04
GC_5_17 b_5 NI_5 NS_17 0 -1.8032968846687958e-04
GC_5_18 b_5 NI_5 NS_18 0 6.0705395883476211e-05
GC_5_19 b_5 NI_5 NS_19 0 -5.0071063583628667e-05
GC_5_20 b_5 NI_5 NS_20 0 1.2013387940195742e-04
GC_5_21 b_5 NI_5 NS_21 0 1.3866115923107195e-04
GC_5_22 b_5 NI_5 NS_22 0 7.0602025256552369e-05
GC_5_23 b_5 NI_5 NS_23 0 4.2957798923436088e-08
GC_5_24 b_5 NI_5 NS_24 0 4.3451731471030420e-06
GC_5_25 b_5 NI_5 NS_25 0 -2.0150898786427323e-06
GC_5_26 b_5 NI_5 NS_26 0 7.7203150116131309e-08
GC_5_27 b_5 NI_5 NS_27 0 6.2847950070478097e-10
GC_5_28 b_5 NI_5 NS_28 0 -6.3035850343910785e-10
GC_5_29 b_5 NI_5 NS_29 0 -1.5189614196007946e-10
GC_5_30 b_5 NI_5 NS_30 0 -1.2381203670678952e-09
GC_5_31 b_5 NI_5 NS_31 0 4.7532271596050444e-05
GC_5_32 b_5 NI_5 NS_32 0 9.2489064230913301e-05
GC_5_33 b_5 NI_5 NS_33 0 2.8963097943998230e-07
GC_5_34 b_5 NI_5 NS_34 0 8.4382805071568453e-09
GC_5_35 b_5 NI_5 NS_35 0 -3.9637599879923364e-05
GC_5_36 b_5 NI_5 NS_36 0 -8.5805859504887221e-05
GC_5_37 b_5 NI_5 NS_37 0 -2.2607906816322812e-04
GC_5_38 b_5 NI_5 NS_38 0 9.6527611055115015e-05
GC_5_39 b_5 NI_5 NS_39 0 2.8256934672354472e-04
GC_5_40 b_5 NI_5 NS_40 0 1.5421120020302117e-04
GC_5_41 b_5 NI_5 NS_41 0 -3.0587235591508636e-04
GC_5_42 b_5 NI_5 NS_42 0 -2.0977069140036444e-04
GC_5_43 b_5 NI_5 NS_43 0 1.8405493487707466e-04
GC_5_44 b_5 NI_5 NS_44 0 3.8935394446277003e-04
GC_5_45 b_5 NI_5 NS_45 0 -9.5573094897882603e-05
GC_5_46 b_5 NI_5 NS_46 0 -1.5669758067639837e-04
GC_5_47 b_5 NI_5 NS_47 0 2.3688406440780253e-04
GC_5_48 b_5 NI_5 NS_48 0 2.1604672656049765e-04
GC_5_49 b_5 NI_5 NS_49 0 -5.9367849581231100e-05
GC_5_50 b_5 NI_5 NS_50 0 -2.0749584543929898e-04
GC_5_51 b_5 NI_5 NS_51 0 -1.3067184353581168e-06
GC_5_52 b_5 NI_5 NS_52 0 2.1379961139234038e-04
GC_5_53 b_5 NI_5 NS_53 0 -2.2338729205544724e-06
GC_5_54 b_5 NI_5 NS_54 0 -4.4289049168842147e-08
GC_5_55 b_5 NI_5 NS_55 0 -4.0520391191200959e-07
GC_5_56 b_5 NI_5 NS_56 0 -4.3742199189929629e-07
GC_5_57 b_5 NI_5 NS_57 0 -7.4128424070471881e-10
GC_5_58 b_5 NI_5 NS_58 0 5.0839396958302212e-10
GC_5_59 b_5 NI_5 NS_59 0 1.5218546103283184e-10
GC_5_60 b_5 NI_5 NS_60 0 1.2347107454218802e-09
GC_5_61 b_5 NI_5 NS_61 0 2.2663492400739412e-03
GC_5_62 b_5 NI_5 NS_62 0 -7.3264017964000578e-04
GC_5_63 b_5 NI_5 NS_63 0 -1.8147155500376210e-06
GC_5_64 b_5 NI_5 NS_64 0 -1.2100169703979443e-07
GC_5_65 b_5 NI_5 NS_65 0 3.5969873324490092e-04
GC_5_66 b_5 NI_5 NS_66 0 -3.7511994252585683e-04
GC_5_67 b_5 NI_5 NS_67 0 -1.2776615397503814e-03
GC_5_68 b_5 NI_5 NS_68 0 3.4323472019698374e-04
GC_5_69 b_5 NI_5 NS_69 0 7.1255517818788038e-04
GC_5_70 b_5 NI_5 NS_70 0 -8.2803185444845211e-04
GC_5_71 b_5 NI_5 NS_71 0 -1.5013266752782648e-04
GC_5_72 b_5 NI_5 NS_72 0 1.3911134446685433e-03
GC_5_73 b_5 NI_5 NS_73 0 -1.3011316374245403e-03
GC_5_74 b_5 NI_5 NS_74 0 -7.6474272164783752e-04
GC_5_75 b_5 NI_5 NS_75 0 6.8662633234941586e-04
GC_5_76 b_5 NI_5 NS_76 0 -2.8643590713356133e-05
GC_5_77 b_5 NI_5 NS_77 0 -1.3691314138931173e-04
GC_5_78 b_5 NI_5 NS_78 0 1.4682073596498950e-03
GC_5_79 b_5 NI_5 NS_79 0 -7.1833247192018969e-04
GC_5_80 b_5 NI_5 NS_80 0 -5.4307221124832853e-04
GC_5_81 b_5 NI_5 NS_81 0 6.5097302056624663e-04
GC_5_82 b_5 NI_5 NS_82 0 1.9308955012773335e-04
GC_5_83 b_5 NI_5 NS_83 0 -3.0134567077198736e-06
GC_5_84 b_5 NI_5 NS_84 0 2.6008719631645675e-05
GC_5_85 b_5 NI_5 NS_85 0 -9.9186048049076909e-06
GC_5_86 b_5 NI_5 NS_86 0 -1.4227993879476176e-06
GC_5_87 b_5 NI_5 NS_87 0 7.0599521133265253e-09
GC_5_88 b_5 NI_5 NS_88 0 -1.0479962193349236e-08
GC_5_89 b_5 NI_5 NS_89 0 -6.2224207883245853e-10
GC_5_90 b_5 NI_5 NS_90 0 -2.1193958533875435e-09
GC_5_91 b_5 NI_5 NS_91 0 9.8221998845326054e-04
GC_5_92 b_5 NI_5 NS_92 0 -3.4568851057396112e-04
GC_5_93 b_5 NI_5 NS_93 0 2.1363463180268923e-06
GC_5_94 b_5 NI_5 NS_94 0 8.2059870812672897e-08
GC_5_95 b_5 NI_5 NS_95 0 1.1716130561782913e-05
GC_5_96 b_5 NI_5 NS_96 0 8.7365700629615686e-05
GC_5_97 b_5 NI_5 NS_97 0 3.1568141584907583e-04
GC_5_98 b_5 NI_5 NS_98 0 -1.1545538138936188e-04
GC_5_99 b_5 NI_5 NS_99 0 -5.1920690108400096e-04
GC_5_100 b_5 NI_5 NS_100 0 -2.4290506716328645e-04
GC_5_101 b_5 NI_5 NS_101 0 3.2786513367049784e-04
GC_5_102 b_5 NI_5 NS_102 0 3.8890657095702190e-04
GC_5_103 b_5 NI_5 NS_103 0 -3.2493458129559144e-04
GC_5_104 b_5 NI_5 NS_104 0 -5.5994745674540396e-04
GC_5_105 b_5 NI_5 NS_105 0 7.3914986946115204e-05
GC_5_106 b_5 NI_5 NS_106 0 3.8468218724308813e-04
GC_5_107 b_5 NI_5 NS_107 0 -3.5604590721878852e-04
GC_5_108 b_5 NI_5 NS_108 0 -2.6839971444927204e-04
GC_5_109 b_5 NI_5 NS_109 0 5.3171178191500111e-06
GC_5_110 b_5 NI_5 NS_110 0 4.0801918413498213e-04
GC_5_111 b_5 NI_5 NS_111 0 -9.5155444612180412e-05
GC_5_112 b_5 NI_5 NS_112 0 -3.4082770335301985e-04
GC_5_113 b_5 NI_5 NS_113 0 -1.4814525261919984e-05
GC_5_114 b_5 NI_5 NS_114 0 -8.4884339860686031e-06
GC_5_115 b_5 NI_5 NS_115 0 2.7375555611239975e-06
GC_5_116 b_5 NI_5 NS_116 0 -6.6722605757409203e-06
GC_5_117 b_5 NI_5 NS_117 0 -7.7198142445263988e-09
GC_5_118 b_5 NI_5 NS_118 0 4.8069214989750035e-09
GC_5_119 b_5 NI_5 NS_119 0 1.1496323406989099e-09
GC_5_120 b_5 NI_5 NS_120 0 2.7805482828933964e-09
GC_5_121 b_5 NI_5 NS_121 0 1.2599073411321338e-01
GC_5_122 b_5 NI_5 NS_122 0 -9.9112046575705205e-03
GC_5_123 b_5 NI_5 NS_123 0 -2.0441620544481966e-05
GC_5_124 b_5 NI_5 NS_124 0 -3.8242974047395100e-06
GC_5_125 b_5 NI_5 NS_125 0 -8.0690521573809418e-03
GC_5_126 b_5 NI_5 NS_126 0 6.6387660765239670e-04
GC_5_127 b_5 NI_5 NS_127 0 -1.9547018341130773e-03
GC_5_128 b_5 NI_5 NS_128 0 7.9835925108020080e-05
GC_5_129 b_5 NI_5 NS_129 0 -1.2548140616111760e-02
GC_5_130 b_5 NI_5 NS_130 0 8.2410841278418214e-03
GC_5_131 b_5 NI_5 NS_131 0 -1.0211192193654756e-02
GC_5_132 b_5 NI_5 NS_132 0 -6.2935718798827305e-04
GC_5_133 b_5 NI_5 NS_133 0 -3.4910900895131435e-03
GC_5_134 b_5 NI_5 NS_134 0 1.6912355268116880e-02
GC_5_135 b_5 NI_5 NS_135 0 -7.7475177972904418e-03
GC_5_136 b_5 NI_5 NS_136 0 1.3307965400227450e-02
GC_5_137 b_5 NI_5 NS_137 0 -3.9569349728180219e-03
GC_5_138 b_5 NI_5 NS_138 0 6.8929693074706406e-03
GC_5_139 b_5 NI_5 NS_139 0 -2.7322523917513073e-03
GC_5_140 b_5 NI_5 NS_140 0 1.2270495815720282e-02
GC_5_141 b_5 NI_5 NS_141 0 -2.2866218902057801e-02
GC_5_142 b_5 NI_5 NS_142 0 5.9252171672498780e-03
GC_5_143 b_5 NI_5 NS_143 0 -8.5896972971984673e-04
GC_5_144 b_5 NI_5 NS_144 0 7.9678382317308213e-04
GC_5_145 b_5 NI_5 NS_145 0 -5.1011835263954164e-04
GC_5_146 b_5 NI_5 NS_146 0 -4.3700565859872435e-04
GC_5_147 b_5 NI_5 NS_147 0 -6.4199781599864623e-08
GC_5_148 b_5 NI_5 NS_148 0 -1.9083794022158586e-07
GC_5_149 b_5 NI_5 NS_149 0 -3.1376277601997439e-09
GC_5_150 b_5 NI_5 NS_150 0 5.5114951277711807e-09
GC_5_151 b_5 NI_5 NS_151 0 -7.5339287960270285e-02
GC_5_152 b_5 NI_5 NS_152 0 2.4883719958362357e-02
GC_5_153 b_5 NI_5 NS_153 0 1.9330117856678718e-05
GC_5_154 b_5 NI_5 NS_154 0 5.3843329167051454e-06
GC_5_155 b_5 NI_5 NS_155 0 1.8356557396898576e-02
GC_5_156 b_5 NI_5 NS_156 0 2.7965826876807414e-02
GC_5_157 b_5 NI_5 NS_157 0 -1.9176395669313090e-02
GC_5_158 b_5 NI_5 NS_158 0 8.3763404895768750e-03
GC_5_159 b_5 NI_5 NS_159 0 -5.5267126897673262e-03
GC_5_160 b_5 NI_5 NS_160 0 -2.3054644493507179e-02
GC_5_161 b_5 NI_5 NS_161 0 2.6686336640670615e-02
GC_5_162 b_5 NI_5 NS_162 0 -1.4570101276776361e-02
GC_5_163 b_5 NI_5 NS_163 0 3.4524049652831075e-02
GC_5_164 b_5 NI_5 NS_164 0 4.8600737671339912e-03
GC_5_165 b_5 NI_5 NS_165 0 9.6777166167375684e-03
GC_5_166 b_5 NI_5 NS_166 0 1.3687348593047830e-02
GC_5_167 b_5 NI_5 NS_167 0 -1.2366663074878274e-02
GC_5_168 b_5 NI_5 NS_168 0 1.1002978815462425e-02
GC_5_169 b_5 NI_5 NS_169 0 -1.1776695103622958e-02
GC_5_170 b_5 NI_5 NS_170 0 -1.2018476729940423e-02
GC_5_171 b_5 NI_5 NS_171 0 1.9787646023365330e-02
GC_5_172 b_5 NI_5 NS_172 0 -2.6040607983496011e-02
GC_5_173 b_5 NI_5 NS_173 0 9.6541124240875215e-04
GC_5_174 b_5 NI_5 NS_174 0 -1.0850257884336776e-03
GC_5_175 b_5 NI_5 NS_175 0 6.3206443218429996e-04
GC_5_176 b_5 NI_5 NS_176 0 3.4856855840376859e-04
GC_5_177 b_5 NI_5 NS_177 0 9.6067328075935982e-08
GC_5_178 b_5 NI_5 NS_178 0 4.1718991135252917e-07
GC_5_179 b_5 NI_5 NS_179 0 -1.0291304675965502e-08
GC_5_180 b_5 NI_5 NS_180 0 -1.9939744778825817e-08
GC_5_181 b_5 NI_5 NS_181 0 -4.2988330634103863e-04
GC_5_182 b_5 NI_5 NS_182 0 -2.9336419347796099e-03
GC_5_183 b_5 NI_5 NS_183 0 -5.9839363530273596e-06
GC_5_184 b_5 NI_5 NS_184 0 -3.8844120751574824e-07
GC_5_185 b_5 NI_5 NS_185 0 2.6783420245401453e-03
GC_5_186 b_5 NI_5 NS_186 0 -1.9922212538343257e-03
GC_5_187 b_5 NI_5 NS_187 0 -6.2097779188802545e-03
GC_5_188 b_5 NI_5 NS_188 0 1.7605677112088223e-03
GC_5_189 b_5 NI_5 NS_189 0 4.7592134835835838e-03
GC_5_190 b_5 NI_5 NS_190 0 -5.5072000653056752e-03
GC_5_191 b_5 NI_5 NS_191 0 -2.2146105042580277e-04
GC_5_192 b_5 NI_5 NS_192 0 7.2473058667639739e-03
GC_5_193 b_5 NI_5 NS_193 0 -6.3292949808905199e-03
GC_5_194 b_5 NI_5 NS_194 0 -5.0696862845352767e-03
GC_5_195 b_5 NI_5 NS_195 0 4.4823184746202293e-03
GC_5_196 b_5 NI_5 NS_196 0 -1.6976964447727319e-03
GC_5_197 b_5 NI_5 NS_197 0 -5.7700526280905784e-04
GC_5_198 b_5 NI_5 NS_198 0 6.9526872290205308e-03
GC_5_199 b_5 NI_5 NS_199 0 -3.4461625867765583e-03
GC_5_200 b_5 NI_5 NS_200 0 -3.6908762062469193e-03
GC_5_201 b_5 NI_5 NS_201 0 5.8924903735889760e-03
GC_5_202 b_5 NI_5 NS_202 0 3.8135561389996976e-04
GC_5_203 b_5 NI_5 NS_203 0 6.0575586239378041e-05
GC_5_204 b_5 NI_5 NS_204 0 6.7951232327458209e-06
GC_5_205 b_5 NI_5 NS_205 0 1.5523892175816139e-05
GC_5_206 b_5 NI_5 NS_206 0 3.8659076368952927e-05
GC_5_207 b_5 NI_5 NS_207 0 6.7893114148684876e-09
GC_5_208 b_5 NI_5 NS_208 0 -2.9476097763899797e-08
GC_5_209 b_5 NI_5 NS_209 0 -1.8905813639732721e-09
GC_5_210 b_5 NI_5 NS_210 0 -5.6443499378434953e-10
GC_5_211 b_5 NI_5 NS_211 0 1.0840922670246537e-03
GC_5_212 b_5 NI_5 NS_212 0 -1.1636889249524048e-03
GC_5_213 b_5 NI_5 NS_213 0 3.5431778317845473e-06
GC_5_214 b_5 NI_5 NS_214 0 2.9212403421921495e-07
GC_5_215 b_5 NI_5 NS_215 0 1.4064404222740798e-04
GC_5_216 b_5 NI_5 NS_216 0 8.9896530515383433e-04
GC_5_217 b_5 NI_5 NS_217 0 1.8646089535908404e-03
GC_5_218 b_5 NI_5 NS_218 0 -8.6916670552580834e-04
GC_5_219 b_5 NI_5 NS_219 0 -2.9480987198010214e-03
GC_5_220 b_5 NI_5 NS_220 0 -1.6595206254428928e-03
GC_5_221 b_5 NI_5 NS_221 0 2.2564581467825525e-03
GC_5_222 b_5 NI_5 NS_222 0 2.6488456344150326e-03
GC_5_223 b_5 NI_5 NS_223 0 -1.4346094264205717e-03
GC_5_224 b_5 NI_5 NS_224 0 -2.9589610827340752e-03
GC_5_225 b_5 NI_5 NS_225 0 1.0713443603436201e-03
GC_5_226 b_5 NI_5 NS_226 0 2.2277942478627082e-03
GC_5_227 b_5 NI_5 NS_227 0 -1.6363481363665196e-03
GC_5_228 b_5 NI_5 NS_228 0 -2.1584332926056944e-03
GC_5_229 b_5 NI_5 NS_229 0 4.3014456973562395e-04
GC_5_230 b_5 NI_5 NS_230 0 2.0082070964713167e-03
GC_5_231 b_5 NI_5 NS_231 0 2.5563233020226136e-04
GC_5_232 b_5 NI_5 NS_232 0 -2.1120365753270086e-03
GC_5_233 b_5 NI_5 NS_233 0 -8.3367111622941104e-08
GC_5_234 b_5 NI_5 NS_234 0 5.0560805793950593e-06
GC_5_235 b_5 NI_5 NS_235 0 -7.2970510681857430e-07
GC_5_236 b_5 NI_5 NS_236 0 -1.7733987878528091e-06
GC_5_237 b_5 NI_5 NS_237 0 -6.9274348772880443e-09
GC_5_238 b_5 NI_5 NS_238 0 2.2849910037722338e-08
GC_5_239 b_5 NI_5 NS_239 0 2.3580829732977999e-09
GC_5_240 b_5 NI_5 NS_240 0 1.5278538684477850e-09
GC_5_241 b_5 NI_5 NS_241 0 1.3866250998233166e-04
GC_5_242 b_5 NI_5 NS_242 0 1.3581110085285046e-06
GC_5_243 b_5 NI_5 NS_243 0 -2.0145404758696825e-07
GC_5_244 b_5 NI_5 NS_244 0 -9.3088469343320933e-09
GC_5_245 b_5 NI_5 NS_245 0 4.9967109803108552e-05
GC_5_246 b_5 NI_5 NS_246 0 -1.9693983487925595e-06
GC_5_247 b_5 NI_5 NS_247 0 2.5673319972904892e-05
GC_5_248 b_5 NI_5 NS_248 0 -7.4987205064210960e-06
GC_5_249 b_5 NI_5 NS_249 0 2.2259867693761837e-05
GC_5_250 b_5 NI_5 NS_250 0 -2.6884224295157757e-04
GC_5_251 b_5 NI_5 NS_251 0 -2.9200887642031817e-04
GC_5_252 b_5 NI_5 NS_252 0 4.0827743177611885e-05
GC_5_253 b_5 NI_5 NS_253 0 -5.4990127725812295e-05
GC_5_254 b_5 NI_5 NS_254 0 2.2142040487331522e-04
GC_5_255 b_5 NI_5 NS_255 0 1.6790480567854780e-04
GC_5_256 b_5 NI_5 NS_256 0 -1.0524497964760553e-04
GC_5_257 b_5 NI_5 NS_257 0 -1.8089903864450030e-04
GC_5_258 b_5 NI_5 NS_258 0 6.1698513663450497e-05
GC_5_259 b_5 NI_5 NS_259 0 -5.0485828620764860e-05
GC_5_260 b_5 NI_5 NS_260 0 1.2080567342422545e-04
GC_5_261 b_5 NI_5 NS_261 0 1.3699039547090055e-04
GC_5_262 b_5 NI_5 NS_262 0 7.0683380379048139e-05
GC_5_263 b_5 NI_5 NS_263 0 -1.0789922691433554e-07
GC_5_264 b_5 NI_5 NS_264 0 4.3458261472479927e-06
GC_5_265 b_5 NI_5 NS_265 0 -2.0228967171568218e-06
GC_5_266 b_5 NI_5 NS_266 0 1.7344805700208079e-08
GC_5_267 b_5 NI_5 NS_267 0 6.0908628667259715e-10
GC_5_268 b_5 NI_5 NS_268 0 -6.4494215331581564e-10
GC_5_269 b_5 NI_5 NS_269 0 -1.4660392294238869e-10
GC_5_270 b_5 NI_5 NS_270 0 -1.2238406329097938e-09
GC_5_271 b_5 NI_5 NS_271 0 5.4736157365917097e-05
GC_5_272 b_5 NI_5 NS_272 0 9.2111711913235570e-05
GC_5_273 b_5 NI_5 NS_273 0 2.8700364147984924e-07
GC_5_274 b_5 NI_5 NS_274 0 8.4904567927957700e-09
GC_5_275 b_5 NI_5 NS_275 0 -4.0121829155476122e-05
GC_5_276 b_5 NI_5 NS_276 0 -8.6000256087875925e-05
GC_5_277 b_5 NI_5 NS_277 0 -2.2672035668295568e-04
GC_5_278 b_5 NI_5 NS_278 0 9.6541664979615991e-05
GC_5_279 b_5 NI_5 NS_279 0 2.8121763860729010e-04
GC_5_280 b_5 NI_5 NS_280 0 1.5448808038517854e-04
GC_5_281 b_5 NI_5 NS_281 0 -3.0713745717624383e-04
GC_5_282 b_5 NI_5 NS_282 0 -2.0845289344767454e-04
GC_5_283 b_5 NI_5 NS_283 0 1.8397833612047101e-04
GC_5_284 b_5 NI_5 NS_284 0 3.9105516817663735e-04
GC_5_285 b_5 NI_5 NS_285 0 -9.4946752798195046e-05
GC_5_286 b_5 NI_5 NS_286 0 -1.5522233052538625e-04
GC_5_287 b_5 NI_5 NS_287 0 2.3740762421901201e-04
GC_5_288 b_5 NI_5 NS_288 0 2.1642595954322622e-04
GC_5_289 b_5 NI_5 NS_289 0 -5.9516953202888661e-05
GC_5_290 b_5 NI_5 NS_290 0 -2.0711938485895175e-04
GC_5_291 b_5 NI_5 NS_291 0 -2.1936488950665667e-06
GC_5_292 b_5 NI_5 NS_292 0 2.1430580406028437e-04
GC_5_293 b_5 NI_5 NS_293 0 -2.2383105557292624e-06
GC_5_294 b_5 NI_5 NS_294 0 6.4589087905182799e-08
GC_5_295 b_5 NI_5 NS_295 0 -4.6477950398045753e-07
GC_5_296 b_5 NI_5 NS_296 0 -4.5309975196156832e-07
GC_5_297 b_5 NI_5 NS_297 0 -7.2775450551601326e-10
GC_5_298 b_5 NI_5 NS_298 0 5.1682454624757206e-10
GC_5_299 b_5 NI_5 NS_299 0 1.4748960385655192e-10
GC_5_300 b_5 NI_5 NS_300 0 1.2209581969797276e-09
GC_5_301 b_5 NI_5 NS_301 0 -5.9716322557720316e-05
GC_5_302 b_5 NI_5 NS_302 0 -4.9579621579383842e-06
GC_5_303 b_5 NI_5 NS_303 0 -5.3052465503349670e-08
GC_5_304 b_5 NI_5 NS_304 0 -5.8065271579881540e-10
GC_5_305 b_5 NI_5 NS_305 0 -6.6914496789007247e-06
GC_5_306 b_5 NI_5 NS_306 0 -5.1560606394719605e-06
GC_5_307 b_5 NI_5 NS_307 0 -3.1757005693071985e-05
GC_5_308 b_5 NI_5 NS_308 0 1.3388490798042759e-05
GC_5_309 b_5 NI_5 NS_309 0 2.0727018835374842e-05
GC_5_310 b_5 NI_5 NS_310 0 6.7059935058316850e-05
GC_5_311 b_5 NI_5 NS_311 0 9.6715112075965111e-05
GC_5_312 b_5 NI_5 NS_312 0 4.8803892988421818e-06
GC_5_313 b_5 NI_5 NS_313 0 -1.5545038749323558e-05
GC_5_314 b_5 NI_5 NS_314 0 -9.0322206993421651e-05
GC_5_315 b_5 NI_5 NS_315 0 -2.8410494895256944e-05
GC_5_316 b_5 NI_5 NS_316 0 3.3441985403512281e-05
GC_5_317 b_5 NI_5 NS_317 0 5.9984035844904709e-05
GC_5_318 b_5 NI_5 NS_318 0 -4.9318773355950769e-06
GC_5_319 b_5 NI_5 NS_319 0 -4.5492025202810974e-06
GC_5_320 b_5 NI_5 NS_320 0 -5.6348575872755769e-05
GC_5_321 b_5 NI_5 NS_321 0 -2.2571981502333436e-05
GC_5_322 b_5 NI_5 NS_322 0 -1.3235097030034714e-05
GC_5_323 b_5 NI_5 NS_323 0 6.7403410032988561e-07
GC_5_324 b_5 NI_5 NS_324 0 -6.8468780766671817e-07
GC_5_325 b_5 NI_5 NS_325 0 3.8201624646954823e-07
GC_5_326 b_5 NI_5 NS_326 0 1.4911380177891462e-07
GC_5_327 b_5 NI_5 NS_327 0 1.7058242704298835e-10
GC_5_328 b_5 NI_5 NS_328 0 -7.6198339762411669e-11
GC_5_329 b_5 NI_5 NS_329 0 -7.2508425668359924e-11
GC_5_330 b_5 NI_5 NS_330 0 -4.3770158798917940e-10
GC_5_331 b_5 NI_5 NS_331 0 9.7557392191026631e-05
GC_5_332 b_5 NI_5 NS_332 0 -6.3842772047081272e-08
GC_5_333 b_5 NI_5 NS_333 0 3.9237401502712176e-08
GC_5_334 b_5 NI_5 NS_334 0 7.0029800210339005e-10
GC_5_335 b_5 NI_5 NS_335 0 3.8317144813175806e-07
GC_5_336 b_5 NI_5 NS_336 0 -1.4093022637636299e-06
GC_5_337 b_5 NI_5 NS_337 0 -9.1557182083264747e-06
GC_5_338 b_5 NI_5 NS_338 0 2.4452150564102485e-05
GC_5_339 b_5 NI_5 NS_339 0 7.9465466162662940e-05
GC_5_340 b_5 NI_5 NS_340 0 8.7690498026679645e-06
GC_5_341 b_5 NI_5 NS_341 0 1.1469116865467569e-05
GC_5_342 b_5 NI_5 NS_342 0 -7.9811145215118493e-05
GC_5_343 b_5 NI_5 NS_343 0 -6.7934157587539218e-06
GC_5_344 b_5 NI_5 NS_344 0 -4.3503399520720265e-05
GC_5_345 b_5 NI_5 NS_345 0 -9.4941652747991832e-05
GC_5_346 b_5 NI_5 NS_346 0 -5.4391210426731962e-05
GC_5_347 b_5 NI_5 NS_347 0 -4.5788268805694557e-05
GC_5_348 b_5 NI_5 NS_348 0 5.2625383147314133e-05
GC_5_349 b_5 NI_5 NS_349 0 -3.1146648000068158e-05
GC_5_350 b_5 NI_5 NS_350 0 1.2605040995304574e-05
GC_5_351 b_5 NI_5 NS_351 0 -1.5816706532082337e-05
GC_5_352 b_5 NI_5 NS_352 0 4.9605030885793370e-05
GC_5_353 b_5 NI_5 NS_353 0 -7.3647506731346872e-07
GC_5_354 b_5 NI_5 NS_354 0 -4.4503384430488927e-07
GC_5_355 b_5 NI_5 NS_355 0 1.3570641549335845e-07
GC_5_356 b_5 NI_5 NS_356 0 -3.6538833814225624e-07
GC_5_357 b_5 NI_5 NS_357 0 -1.5129395351170996e-10
GC_5_358 b_5 NI_5 NS_358 0 9.3552987448571220e-11
GC_5_359 b_5 NI_5 NS_359 0 7.1163721531462728e-11
GC_5_360 b_5 NI_5 NS_360 0 4.3626480470848610e-10
GD_5_1 b_5 NI_5 NA_1 0 1.7077821725073578e-04
GD_5_2 b_5 NI_5 NA_2 0 -6.0788958049236536e-05
GD_5_3 b_5 NI_5 NA_3 0 2.3298014152281260e-03
GD_5_4 b_5 NI_5 NA_4 0 -4.6783139904390105e-05
GD_5_5 b_5 NI_5 NA_5 0 -4.0224699724402471e-02
GD_5_6 b_5 NI_5 NA_6 0 -9.9740445305878528e-03
GD_5_7 b_5 NI_5 NA_7 0 1.6033810802924379e-02
GD_5_8 b_5 NI_5 NA_8 0 -3.7759943577884097e-05
GD_5_9 b_5 NI_5 NA_9 0 1.6921919722808469e-04
GD_5_10 b_5 NI_5 NA_10 0 -6.2836548667596917e-05
GD_5_11 b_5 NI_5 NA_11 0 3.8174511259994853e-06
GD_5_12 b_5 NI_5 NA_12 0 8.3909789437812144e-06
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 4.7529404043407935e-05
GC_6_2 b_6 NI_6 NS_2 0 9.2489246294779400e-05
GC_6_3 b_6 NI_6 NS_3 0 2.8963833700943906e-07
GC_6_4 b_6 NI_6 NS_4 0 8.4383177632276242e-09
GC_6_5 b_6 NI_6 NS_5 0 -3.9637640095678359e-05
GC_6_6 b_6 NI_6 NS_6 0 -8.5800994712951072e-05
GC_6_7 b_6 NI_6 NS_7 0 -2.2608169022328715e-04
GC_6_8 b_6 NI_6 NS_8 0 9.6531803615791670e-05
GC_6_9 b_6 NI_6 NS_9 0 2.8257314199459045e-04
GC_6_10 b_6 NI_6 NS_10 0 1.5420735143575182e-04
GC_6_11 b_6 NI_6 NS_11 0 -3.0587341594500686e-04
GC_6_12 b_6 NI_6 NS_12 0 -2.0976792639094632e-04
GC_6_13 b_6 NI_6 NS_13 0 1.8406147744641260e-04
GC_6_14 b_6 NI_6 NS_14 0 3.8935567182311860e-04
GC_6_15 b_6 NI_6 NS_15 0 -9.5573710850402739e-05
GC_6_16 b_6 NI_6 NS_16 0 -1.5669664151134820e-04
GC_6_17 b_6 NI_6 NS_17 0 2.3688714669774244e-04
GC_6_18 b_6 NI_6 NS_18 0 2.1604584814134955e-04
GC_6_19 b_6 NI_6 NS_19 0 -5.9368011261115722e-05
GC_6_20 b_6 NI_6 NS_20 0 -2.0749699671023439e-04
GC_6_21 b_6 NI_6 NS_21 0 -1.3040362945613148e-06
GC_6_22 b_6 NI_6 NS_22 0 2.1379953049746638e-04
GC_6_23 b_6 NI_6 NS_23 0 -2.2339328122456738e-06
GC_6_24 b_6 NI_6 NS_24 0 -4.4443761451502109e-08
GC_6_25 b_6 NI_6 NS_25 0 -4.0519950343567944e-07
GC_6_26 b_6 NI_6 NS_26 0 -4.3752051445754023e-07
GC_6_27 b_6 NI_6 NS_27 0 -7.4130870403326556e-10
GC_6_28 b_6 NI_6 NS_28 0 5.0839026590189672e-10
GC_6_29 b_6 NI_6 NS_29 0 1.5218849885232036e-10
GC_6_30 b_6 NI_6 NS_30 0 1.2347152130959892e-09
GC_6_31 b_6 NI_6 NS_31 0 1.4263880614678263e-04
GC_6_32 b_6 NI_6 NS_32 0 1.2397282086845646e-06
GC_6_33 b_6 NI_6 NS_33 0 -2.0479871770124067e-07
GC_6_34 b_6 NI_6 NS_34 0 -9.2517560415118182e-09
GC_6_35 b_6 NI_6 NS_35 0 4.9822047756304829e-05
GC_6_36 b_6 NI_6 NS_36 0 -2.0166476431603002e-06
GC_6_37 b_6 NI_6 NS_37 0 2.5357888587942720e-05
GC_6_38 b_6 NI_6 NS_38 0 -7.6229365303167256e-06
GC_6_39 b_6 NI_6 NS_39 0 2.2183853277334241e-05
GC_6_40 b_6 NI_6 NS_40 0 -2.6867991399770041e-04
GC_6_41 b_6 NI_6 NS_41 0 -2.9255258097777529e-04
GC_6_42 b_6 NI_6 NS_42 0 4.0714051658204878e-05
GC_6_43 b_6 NI_6 NS_43 0 -5.5577241348226784e-05
GC_6_44 b_6 NI_6 NS_44 0 2.2174315920000116e-04
GC_6_45 b_6 NI_6 NS_45 0 1.6780985302961121e-04
GC_6_46 b_6 NI_6 NS_46 0 -1.0454530626151895e-04
GC_6_47 b_6 NI_6 NS_47 0 -1.8111484377603969e-04
GC_6_48 b_6 NI_6 NS_48 0 6.2085961479670158e-05
GC_6_49 b_6 NI_6 NS_49 0 -5.0743165088658386e-05
GC_6_50 b_6 NI_6 NS_50 0 1.2107951040554659e-04
GC_6_51 b_6 NI_6 NS_51 0 1.3633682334685782e-04
GC_6_52 b_6 NI_6 NS_52 0 7.1243819744348325e-05
GC_6_53 b_6 NI_6 NS_53 0 -9.2884404553346596e-08
GC_6_54 b_6 NI_6 NS_54 0 4.4336494120841090e-06
GC_6_55 b_6 NI_6 NS_55 0 -2.0707155175282032e-06
GC_6_56 b_6 NI_6 NS_56 0 1.1473729833120061e-08
GC_6_57 b_6 NI_6 NS_57 0 6.2405872942276581e-10
GC_6_58 b_6 NI_6 NS_58 0 -6.3535515236878582e-10
GC_6_59 b_6 NI_6 NS_59 0 -1.5179186304188703e-10
GC_6_60 b_6 NI_6 NS_60 0 -1.2381860264181437e-09
GC_6_61 b_6 NI_6 NS_61 0 9.8191000710233641e-04
GC_6_62 b_6 NI_6 NS_62 0 -3.4563276908159953e-04
GC_6_63 b_6 NI_6 NS_63 0 2.1362724158167818e-06
GC_6_64 b_6 NI_6 NS_64 0 8.2060295943127796e-08
GC_6_65 b_6 NI_6 NS_65 0 1.1626324372703267e-05
GC_6_66 b_6 NI_6 NS_66 0 8.7329047216630932e-05
GC_6_67 b_6 NI_6 NS_67 0 3.1565129779423623e-04
GC_6_68 b_6 NI_6 NS_68 0 -1.1550920472581685e-04
GC_6_69 b_6 NI_6 NS_69 0 -5.1916494456237538e-04
GC_6_70 b_6 NI_6 NS_70 0 -2.4271238356379294e-04
GC_6_71 b_6 NI_6 NS_71 0 3.2788951433130291e-04
GC_6_72 b_6 NI_6 NS_72 0 3.8892142555885570e-04
GC_6_73 b_6 NI_6 NS_73 0 -3.2494336627801769e-04
GC_6_74 b_6 NI_6 NS_74 0 -5.5985364379252539e-04
GC_6_75 b_6 NI_6 NS_75 0 7.3996223445681162e-05
GC_6_76 b_6 NI_6 NS_76 0 3.8462470696021809e-04
GC_6_77 b_6 NI_6 NS_77 0 -3.5599393468439670e-04
GC_6_78 b_6 NI_6 NS_78 0 -2.6837281247813150e-04
GC_6_79 b_6 NI_6 NS_79 0 5.3984160093501751e-06
GC_6_80 b_6 NI_6 NS_80 0 4.0799729250003358e-04
GC_6_81 b_6 NI_6 NS_81 0 -9.5062218967622577e-05
GC_6_82 b_6 NI_6 NS_82 0 -3.4082775084778302e-04
GC_6_83 b_6 NI_6 NS_83 0 -1.4810484634238721e-05
GC_6_84 b_6 NI_6 NS_84 0 -8.4933390569874658e-06
GC_6_85 b_6 NI_6 NS_85 0 2.7402887748044267e-06
GC_6_86 b_6 NI_6 NS_86 0 -6.6705469056713432e-06
GC_6_87 b_6 NI_6 NS_87 0 -7.7197156543075300e-09
GC_6_88 b_6 NI_6 NS_88 0 4.8070271978097383e-09
GC_6_89 b_6 NI_6 NS_89 0 1.1496194840926708e-09
GC_6_90 b_6 NI_6 NS_90 0 2.7805417329395022e-09
GC_6_91 b_6 NI_6 NS_91 0 2.2651865886702265e-03
GC_6_92 b_6 NI_6 NS_92 0 -7.3251972011469774e-04
GC_6_93 b_6 NI_6 NS_93 0 -1.8149120175278200e-06
GC_6_94 b_6 NI_6 NS_94 0 -1.2099866005222807e-07
GC_6_95 b_6 NI_6 NS_95 0 3.5975567735494065e-04
GC_6_96 b_6 NI_6 NS_96 0 -3.7511051392748846e-04
GC_6_97 b_6 NI_6 NS_97 0 -1.2775980892524533e-03
GC_6_98 b_6 NI_6 NS_98 0 3.4322578639538160e-04
GC_6_99 b_6 NI_6 NS_99 0 7.1263690545207280e-04
GC_6_100 b_6 NI_6 NS_100 0 -8.2807530089480457e-04
GC_6_101 b_6 NI_6 NS_101 0 -1.5003852361291151e-04
GC_6_102 b_6 NI_6 NS_102 0 1.3910695890865991e-03
GC_6_103 b_6 NI_6 NS_103 0 -1.3010597841854343e-03
GC_6_104 b_6 NI_6 NS_104 0 -7.6485404590117536e-04
GC_6_105 b_6 NI_6 NS_105 0 6.8667001039827849e-04
GC_6_106 b_6 NI_6 NS_106 0 -2.8752446521507342e-05
GC_6_107 b_6 NI_6 NS_107 0 -1.3686847991445145e-04
GC_6_108 b_6 NI_6 NS_108 0 1.4680977678799656e-03
GC_6_109 b_6 NI_6 NS_109 0 -7.1828111558737699e-04
GC_6_110 b_6 NI_6 NS_110 0 -5.4315200812566256e-04
GC_6_111 b_6 NI_6 NS_111 0 6.5114860903004162e-04
GC_6_112 b_6 NI_6 NS_112 0 1.9303369668727900e-04
GC_6_113 b_6 NI_6 NS_113 0 -3.0047597073234193e-06
GC_6_114 b_6 NI_6 NS_114 0 2.6001120928722230e-05
GC_6_115 b_6 NI_6 NS_115 0 -9.9139321314521452e-06
GC_6_116 b_6 NI_6 NS_116 0 -1.4183971024163971e-06
GC_6_117 b_6 NI_6 NS_117 0 7.0603582379898926e-09
GC_6_118 b_6 NI_6 NS_118 0 -1.0479502326724456e-08
GC_6_119 b_6 NI_6 NS_119 0 -6.2226005295884097e-10
GC_6_120 b_6 NI_6 NS_120 0 -2.1194094617205798e-09
GC_6_121 b_6 NI_6 NS_121 0 -7.5339607420133514e-02
GC_6_122 b_6 NI_6 NS_122 0 2.4883759867721199e-02
GC_6_123 b_6 NI_6 NS_123 0 1.9330040494682609e-05
GC_6_124 b_6 NI_6 NS_124 0 5.3843347150347869e-06
GC_6_125 b_6 NI_6 NS_125 0 1.8356559574355742e-02
GC_6_126 b_6 NI_6 NS_126 0 2.7965832958539282e-02
GC_6_127 b_6 NI_6 NS_127 0 -1.9176389900470495e-02
GC_6_128 b_6 NI_6 NS_128 0 8.3763509093365222e-03
GC_6_129 b_6 NI_6 NS_129 0 -5.5266929072144812e-03
GC_6_130 b_6 NI_6 NS_130 0 -2.3054635236206183e-02
GC_6_131 b_6 NI_6 NS_131 0 2.6686362654414701e-02
GC_6_132 b_6 NI_6 NS_132 0 -1.4570094127759631e-02
GC_6_133 b_6 NI_6 NS_133 0 3.4524082293192114e-02
GC_6_134 b_6 NI_6 NS_134 0 4.8600630401891640e-03
GC_6_135 b_6 NI_6 NS_135 0 9.6777441253077853e-03
GC_6_136 b_6 NI_6 NS_136 0 1.3687329180206211e-02
GC_6_137 b_6 NI_6 NS_137 0 -1.2366631894203018e-02
GC_6_138 b_6 NI_6 NS_138 0 1.1002955997739376e-02
GC_6_139 b_6 NI_6 NS_139 0 -1.1776667060433298e-02
GC_6_140 b_6 NI_6 NS_140 0 -1.2018498437579350e-02
GC_6_141 b_6 NI_6 NS_141 0 1.9787709408560897e-02
GC_6_142 b_6 NI_6 NS_142 0 -2.6040623008703984e-02
GC_6_143 b_6 NI_6 NS_143 0 9.6541417395488234e-04
GC_6_144 b_6 NI_6 NS_144 0 -1.0850280594338689e-03
GC_6_145 b_6 NI_6 NS_145 0 6.3206587651109527e-04
GC_6_146 b_6 NI_6 NS_146 0 3.4856993383115521e-04
GC_6_147 b_6 NI_6 NS_147 0 9.6067446224714915e-08
GC_6_148 b_6 NI_6 NS_148 0 4.1719029748693908e-07
GC_6_149 b_6 NI_6 NS_149 0 -1.0291342080483950e-08
GC_6_150 b_6 NI_6 NS_150 0 -1.9939776031229145e-08
GC_6_151 b_6 NI_6 NS_151 0 1.2599073411321318e-01
GC_6_152 b_6 NI_6 NS_152 0 -9.9112046575704875e-03
GC_6_153 b_6 NI_6 NS_153 0 -2.0441620544482329e-05
GC_6_154 b_6 NI_6 NS_154 0 -3.8242974047395007e-06
GC_6_155 b_6 NI_6 NS_155 0 -8.0690521573809470e-03
GC_6_156 b_6 NI_6 NS_156 0 6.6387660765240050e-04
GC_6_157 b_6 NI_6 NS_157 0 -1.9547018341130634e-03
GC_6_158 b_6 NI_6 NS_158 0 7.9835925108028848e-05
GC_6_159 b_6 NI_6 NS_159 0 -1.2548140616111755e-02
GC_6_160 b_6 NI_6 NS_160 0 8.2410841278418266e-03
GC_6_161 b_6 NI_6 NS_161 0 -1.0211192193654725e-02
GC_6_162 b_6 NI_6 NS_162 0 -6.2935718798827305e-04
GC_6_163 b_6 NI_6 NS_163 0 -3.4910900895131262e-03
GC_6_164 b_6 NI_6 NS_164 0 1.6912355268116862e-02
GC_6_165 b_6 NI_6 NS_165 0 -7.7475177972904452e-03
GC_6_166 b_6 NI_6 NS_166 0 1.3307965400227439e-02
GC_6_167 b_6 NI_6 NS_167 0 -3.9569349728180115e-03
GC_6_168 b_6 NI_6 NS_168 0 6.8929693074706328e-03
GC_6_169 b_6 NI_6 NS_169 0 -2.7322523917512991e-03
GC_6_170 b_6 NI_6 NS_170 0 1.2270495815720281e-02
GC_6_171 b_6 NI_6 NS_171 0 -2.2866218902057773e-02
GC_6_172 b_6 NI_6 NS_172 0 5.9252171672498841e-03
GC_6_173 b_6 NI_6 NS_173 0 -8.5896972971984337e-04
GC_6_174 b_6 NI_6 NS_174 0 7.9678382317308462e-04
GC_6_175 b_6 NI_6 NS_175 0 -5.1011835263954294e-04
GC_6_176 b_6 NI_6 NS_176 0 -4.3700565859872321e-04
GC_6_177 b_6 NI_6 NS_177 0 -6.4199781599866701e-08
GC_6_178 b_6 NI_6 NS_178 0 -1.9083794022158308e-07
GC_6_179 b_6 NI_6 NS_179 0 -3.1376277602029876e-09
GC_6_180 b_6 NI_6 NS_180 0 5.5114951277674799e-09
GC_6_181 b_6 NI_6 NS_181 0 1.0838823714819001e-03
GC_6_182 b_6 NI_6 NS_182 0 -1.1636685271583383e-03
GC_6_183 b_6 NI_6 NS_183 0 3.5431451647806048e-06
GC_6_184 b_6 NI_6 NS_184 0 2.9212450531121249e-07
GC_6_185 b_6 NI_6 NS_185 0 1.4066769082717007e-04
GC_6_186 b_6 NI_6 NS_186 0 8.9897478263251617e-04
GC_6_187 b_6 NI_6 NS_187 0 1.8646238121185926e-03
GC_6_188 b_6 NI_6 NS_188 0 -8.6915567389506294e-04
GC_6_189 b_6 NI_6 NS_189 0 -2.9480926598205465e-03
GC_6_190 b_6 NI_6 NS_190 0 -1.6595552023057878e-03
GC_6_191 b_6 NI_6 NS_191 0 2.2564741451611024e-03
GC_6_192 b_6 NI_6 NS_192 0 2.6488447170502087e-03
GC_6_193 b_6 NI_6 NS_193 0 -1.4345831403094888e-03
GC_6_194 b_6 NI_6 NS_194 0 -2.9589936278453526e-03
GC_6_195 b_6 NI_6 NS_195 0 1.0713461029232478e-03
GC_6_196 b_6 NI_6 NS_196 0 2.2277830754690326e-03
GC_6_197 b_6 NI_6 NS_197 0 -1.6363393827163884e-03
GC_6_198 b_6 NI_6 NS_198 0 -2.1584583419812578e-03
GC_6_199 b_6 NI_6 NS_199 0 4.3014902104061966e-04
GC_6_200 b_6 NI_6 NS_200 0 2.0081938847509003e-03
GC_6_201 b_6 NI_6 NS_201 0 2.5566390069106572e-04
GC_6_202 b_6 NI_6 NS_202 0 -2.1120493070928030e-03
GC_6_203 b_6 NI_6 NS_203 0 -8.1917109482818723e-08
GC_6_204 b_6 NI_6 NS_204 0 5.0549397308268994e-06
GC_6_205 b_6 NI_6 NS_205 0 -7.2891361720862673e-07
GC_6_206 b_6 NI_6 NS_206 0 -1.7726258484745412e-06
GC_6_207 b_6 NI_6 NS_207 0 -6.9273595010498190e-09
GC_6_208 b_6 NI_6 NS_208 0 2.2849982943392392e-08
GC_6_209 b_6 NI_6 NS_209 0 2.3580775129936354e-09
GC_6_210 b_6 NI_6 NS_210 0 1.5278505482418853e-09
GC_6_211 b_6 NI_6 NS_211 0 -4.2988052038240470e-04
GC_6_212 b_6 NI_6 NS_212 0 -2.9336422244617454e-03
GC_6_213 b_6 NI_6 NS_213 0 -5.9839359493122031e-06
GC_6_214 b_6 NI_6 NS_214 0 -3.8844121115236810e-07
GC_6_215 b_6 NI_6 NS_215 0 2.6783419208677587e-03
GC_6_216 b_6 NI_6 NS_216 0 -1.9922212938142236e-03
GC_6_217 b_6 NI_6 NS_217 0 -6.2097780491404044e-03
GC_6_218 b_6 NI_6 NS_218 0 1.7605677202605975e-03
GC_6_219 b_6 NI_6 NS_219 0 4.7592133388197231e-03
GC_6_220 b_6 NI_6 NS_220 0 -5.5072000178070088e-03
GC_6_221 b_6 NI_6 NS_221 0 -2.2146125338751835e-04
GC_6_222 b_6 NI_6 NS_222 0 7.2473058856116594e-03
GC_6_223 b_6 NI_6 NS_223 0 -6.3292952035544966e-03
GC_6_224 b_6 NI_6 NS_224 0 -5.0696861088136294e-03
GC_6_225 b_6 NI_6 NS_225 0 4.4823182983335314e-03
GC_6_226 b_6 NI_6 NS_226 0 -1.6976962329513855e-03
GC_6_227 b_6 NI_6 NS_227 0 -5.7700545307214741e-04
GC_6_228 b_6 NI_6 NS_228 0 6.9526874784096799e-03
GC_6_229 b_6 NI_6 NS_229 0 -3.4461627633188552e-03
GC_6_230 b_6 NI_6 NS_230 0 -3.6908760057206657e-03
GC_6_231 b_6 NI_6 NS_231 0 5.8924899006940123e-03
GC_6_232 b_6 NI_6 NS_232 0 3.8135578020032313e-04
GC_6_233 b_6 NI_6 NS_233 0 6.0575568528386798e-05
GC_6_234 b_6 NI_6 NS_234 0 6.7951427454913578e-06
GC_6_235 b_6 NI_6 NS_235 0 1.5523879572242515e-05
GC_6_236 b_6 NI_6 NS_236 0 3.8659068401755665e-05
GC_6_237 b_6 NI_6 NS_237 0 6.7893105569913257e-09
GC_6_238 b_6 NI_6 NS_238 0 -2.9476098365486250e-08
GC_6_239 b_6 NI_6 NS_239 0 -1.8905813247337954e-09
GC_6_240 b_6 NI_6 NS_240 0 -5.6443499855355768e-10
GC_6_241 b_6 NI_6 NS_241 0 5.4752154018401094e-05
GC_6_242 b_6 NI_6 NS_242 0 9.2110310902821118e-05
GC_6_243 b_6 NI_6 NS_243 0 2.8700554578277191e-07
GC_6_244 b_6 NI_6 NS_244 0 8.4904237329906508e-09
GC_6_245 b_6 NI_6 NS_245 0 -4.0122562833061902e-05
GC_6_246 b_6 NI_6 NS_246 0 -8.5999951812822177e-05
GC_6_247 b_6 NI_6 NS_247 0 -2.2672065800386594e-04
GC_6_248 b_6 NI_6 NS_248 0 9.6541364452455353e-05
GC_6_249 b_6 NI_6 NS_249 0 2.8121580720593515e-04
GC_6_250 b_6 NI_6 NS_250 0 1.5448853371768229e-04
GC_6_251 b_6 NI_6 NS_251 0 -3.0713872740714514e-04
GC_6_252 b_6 NI_6 NS_252 0 -2.0845193557348331e-04
GC_6_253 b_6 NI_6 NS_253 0 1.8397692249118327e-04
GC_6_254 b_6 NI_6 NS_254 0 3.9105606887090245e-04
GC_6_255 b_6 NI_6 NS_255 0 -9.4947559103984109e-05
GC_6_256 b_6 NI_6 NS_256 0 -1.5521933874865012e-04
GC_6_257 b_6 NI_6 NS_257 0 2.3740745873390717e-04
GC_6_258 b_6 NI_6 NS_258 0 2.1642751423899185e-04
GC_6_259 b_6 NI_6 NS_259 0 -5.9517836592164968e-05
GC_6_260 b_6 NI_6 NS_260 0 -2.0711790671541942e-04
GC_6_261 b_6 NI_6 NS_261 0 -2.1951773753940714e-06
GC_6_262 b_6 NI_6 NS_262 0 2.1430694893296009e-04
GC_6_263 b_6 NI_6 NS_263 0 -2.2384337330811990e-06
GC_6_264 b_6 NI_6 NS_264 0 6.4681908962421275e-08
GC_6_265 b_6 NI_6 NS_265 0 -4.6483139812305991e-07
GC_6_266 b_6 NI_6 NS_266 0 -4.5316246825355049e-07
GC_6_267 b_6 NI_6 NS_267 0 -7.2775863886637205e-10
GC_6_268 b_6 NI_6 NS_268 0 5.1681952777835940e-10
GC_6_269 b_6 NI_6 NS_269 0 1.4748977677629137e-10
GC_6_270 b_6 NI_6 NS_270 0 1.2209582719587393e-09
GC_6_271 b_6 NI_6 NS_271 0 1.2368801880826365e-04
GC_6_272 b_6 NI_6 NS_272 0 3.0410909185759357e-06
GC_6_273 b_6 NI_6 NS_273 0 -2.0461318705688850e-07
GC_6_274 b_6 NI_6 NS_274 0 -9.2714568243557466e-09
GC_6_275 b_6 NI_6 NS_275 0 5.0549171103322381e-05
GC_6_276 b_6 NI_6 NS_276 0 -1.8064784689245983e-06
GC_6_277 b_6 NI_6 NS_277 0 2.6605830004787285e-05
GC_6_278 b_6 NI_6 NS_278 0 -7.3891975037747517e-06
GC_6_279 b_6 NI_6 NS_279 0 2.3147543089910568e-05
GC_6_280 b_6 NI_6 NS_280 0 -2.6931280935142086e-04
GC_6_281 b_6 NI_6 NS_281 0 -2.9061129598189223e-04
GC_6_282 b_6 NI_6 NS_282 0 4.0339509825974434e-05
GC_6_283 b_6 NI_6 NS_283 0 -5.3941966830330908e-05
GC_6_284 b_6 NI_6 NS_284 0 2.2027267087789797e-04
GC_6_285 b_6 NI_6 NS_285 0 1.6852043013720373e-04
GC_6_286 b_6 NI_6 NS_286 0 -1.0671238681479294e-04
GC_6_287 b_6 NI_6 NS_287 0 -1.8010365291132869e-04
GC_6_288 b_6 NI_6 NS_288 0 6.0291836817617495e-05
GC_6_289 b_6 NI_6 NS_289 0 -4.9801218002541373e-05
GC_6_290 b_6 NI_6 NS_290 0 1.1984178022802449e-04
GC_6_291 b_6 NI_6 NS_291 0 1.3935796540507175e-04
GC_6_292 b_6 NI_6 NS_292 0 7.0033210100102394e-05
GC_6_293 b_6 NI_6 NS_293 0 3.0857760248737267e-08
GC_6_294 b_6 NI_6 NS_294 0 4.2557785679217513e-06
GC_6_295 b_6 NI_6 NS_295 0 -1.9662424748091160e-06
GC_6_296 b_6 NI_6 NS_296 0 8.4457542172029461e-08
GC_6_297 b_6 NI_6 NS_297 0 6.1361185702443315e-10
GC_6_298 b_6 NI_6 NS_298 0 -6.3988311696128989e-10
GC_6_299 b_6 NI_6 NS_299 0 -1.4671369787257862e-10
GC_6_300 b_6 NI_6 NS_300 0 -1.2237817828820434e-09
GC_6_301 b_6 NI_6 NS_301 0 9.6421903142094074e-05
GC_6_302 b_6 NI_6 NS_302 0 2.8798942808375614e-08
GC_6_303 b_6 NI_6 NS_303 0 3.9109900084154727e-08
GC_6_304 b_6 NI_6 NS_304 0 7.0175518736752990e-10
GC_6_305 b_6 NI_6 NS_305 0 5.3823017471570829e-07
GC_6_306 b_6 NI_6 NS_306 0 -1.3492803942277510e-06
GC_6_307 b_6 NI_6 NS_307 0 -9.0392074173722785e-06
GC_6_308 b_6 NI_6 NS_308 0 2.4491118510374457e-05
GC_6_309 b_6 NI_6 NS_309 0 7.9496248941772387e-05
GC_6_310 b_6 NI_6 NS_310 0 8.5223802660384004e-06
GC_6_311 b_6 NI_6 NS_311 0 1.1537152693099601e-05
GC_6_312 b_6 NI_6 NS_312 0 -7.9841300237395502e-05
GC_6_313 b_6 NI_6 NS_313 0 -6.6585356190823244e-06
GC_6_314 b_6 NI_6 NS_314 0 -4.3699588905623617e-05
GC_6_315 b_6 NI_6 NS_315 0 -9.4957032571641096e-05
GC_6_316 b_6 NI_6 NS_316 0 -5.4470338024552317e-05
GC_6_317 b_6 NI_6 NS_317 0 -4.5766854779251573e-05
GC_6_318 b_6 NI_6 NS_318 0 5.2480776904457839e-05
GC_6_319 b_6 NI_6 NS_319 0 -3.1138984358084375e-05
GC_6_320 b_6 NI_6 NS_320 0 1.2530530356615284e-05
GC_6_321 b_6 NI_6 NS_321 0 -1.5669043613081356e-05
GC_6_322 b_6 NI_6 NS_322 0 4.9521444069564177e-05
GC_6_323 b_6 NI_6 NS_323 0 -7.3125483167829450e-07
GC_6_324 b_6 NI_6 NS_324 0 -4.5045374740569141e-07
GC_6_325 b_6 NI_6 NS_325 0 1.3959010129329322e-07
GC_6_326 b_6 NI_6 NS_326 0 -3.6272330391987479e-07
GC_6_327 b_6 NI_6 NS_327 0 -1.5098901171692854e-10
GC_6_328 b_6 NI_6 NS_328 0 9.3782714050161526e-11
GC_6_329 b_6 NI_6 NS_329 0 7.1151105110165018e-11
GC_6_330 b_6 NI_6 NS_330 0 4.3624309285304850e-10
GC_6_331 b_6 NI_6 NS_331 0 -5.9645810639020153e-05
GC_6_332 b_6 NI_6 NS_332 0 -4.9654237923381193e-06
GC_6_333 b_6 NI_6 NS_333 0 -5.3039122392498771e-08
GC_6_334 b_6 NI_6 NS_334 0 -5.8090607943560715e-10
GC_6_335 b_6 NI_6 NS_335 0 -6.6949085763660875e-06
GC_6_336 b_6 NI_6 NS_336 0 -5.1567311069344485e-06
GC_6_337 b_6 NI_6 NS_337 0 -3.1760424633388274e-05
GC_6_338 b_6 NI_6 NS_338 0 1.3387790186596356e-05
GC_6_339 b_6 NI_6 NS_339 0 2.0720936055482408e-05
GC_6_340 b_6 NI_6 NS_340 0 6.7062458822982987e-05
GC_6_341 b_6 NI_6 NS_341 0 9.6708352088478201e-05
GC_6_342 b_6 NI_6 NS_342 0 4.8828677692217225e-06
GC_6_343 b_6 NI_6 NS_343 0 -1.5549097444661938e-05
GC_6_344 b_6 NI_6 NS_344 0 -9.0315249085946522e-05
GC_6_345 b_6 NI_6 NS_345 0 -2.8413734678947043e-05
GC_6_346 b_6 NI_6 NS_346 0 3.3448569770489025e-05
GC_6_347 b_6 NI_6 NS_347 0 5.9980502394869641e-05
GC_6_348 b_6 NI_6 NS_348 0 -4.9248339743263402e-06
GC_6_349 b_6 NI_6 NS_349 0 -4.5519426586499097e-06
GC_6_350 b_6 NI_6 NS_350 0 -5.6343191562886423e-05
GC_6_351 b_6 NI_6 NS_351 0 -2.2582441882314114e-05
GC_6_352 b_6 NI_6 NS_352 0 -1.3231851780265377e-05
GC_6_353 b_6 NI_6 NS_353 0 6.7346331455528897e-07
GC_6_354 b_6 NI_6 NS_354 0 -6.8427533394890893e-07
GC_6_355 b_6 NI_6 NS_355 0 3.8175830392045661e-07
GC_6_356 b_6 NI_6 NS_356 0 1.4884424098441611e-07
GC_6_357 b_6 NI_6 NS_357 0 1.7055251146698510e-10
GC_6_358 b_6 NI_6 NS_358 0 -7.6241216315748699e-11
GC_6_359 b_6 NI_6 NS_359 0 -7.2505238354709801e-11
GC_6_360 b_6 NI_6 NS_360 0 -4.3769883077108661e-10
GD_6_1 b_6 NI_6 NA_1 0 -6.0795871134196025e-05
GD_6_2 b_6 NI_6 NA_2 0 1.6881266759593416e-04
GD_6_3 b_6 NI_6 NA_3 0 -4.6772756379743946e-05
GD_6_4 b_6 NI_6 NA_4 0 2.3300350421512597e-03
GD_6_5 b_6 NI_6 NA_5 0 -9.9740241344489049e-03
GD_6_6 b_6 NI_6 NA_6 0 -4.0224699724402360e-02
GD_6_7 b_6 NI_6 NA_7 0 -3.7727936103095701e-05
GD_6_8 b_6 NI_6 NA_8 0 1.6033810388021666e-02
GD_6_9 b_6 NI_6 NA_9 0 -6.2840282483554412e-05
GD_6_10 b_6 NI_6 NA_10 0 1.7125087286493391e-04
GD_6_11 b_6 NI_6 NA_11 0 8.6158352242780212e-06
GD_6_12 b_6 NI_6 NA_12 0 3.8071666632870531e-06
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 -4.8135716527291533e-05
GC_7_2 b_7 NI_7 NS_2 0 -6.1994505327946950e-06
GC_7_3 b_7 NI_7 NS_3 0 -5.0843105329247058e-08
GC_7_4 b_7 NI_7 NS_4 0 -6.2431948966900872e-10
GC_7_5 b_7 NI_7 NS_5 0 -7.2065667168328169e-06
GC_7_6 b_7 NI_7 NS_6 0 -5.3857708290721351e-06
GC_7_7 b_7 NI_7 NS_7 0 -3.2442024566157802e-05
GC_7_8 b_7 NI_7 NS_8 0 1.3398299576138161e-05
GC_7_9 b_7 NI_7 NS_9 0 1.9876528227259883e-05
GC_7_10 b_7 NI_7 NS_10 0 6.7339623836336457e-05
GC_7_11 b_7 NI_7 NS_11 0 9.5704756306467937e-05
GC_7_12 b_7 NI_7 NS_12 0 5.2308313805063917e-06
GC_7_13 b_7 NI_7 NS_13 0 -1.6517241266969708e-05
GC_7_14 b_7 NI_7 NS_14 0 -8.9259113685169440e-05
GC_7_15 b_7 NI_7 NS_15 0 -2.8888132854508985e-05
GC_7_16 b_7 NI_7 NS_16 0 3.4594520369884967e-05
GC_7_17 b_7 NI_7 NS_17 0 5.9457511427339758e-05
GC_7_18 b_7 NI_7 NS_18 0 -3.7031010492686586e-06
GC_7_19 b_7 NI_7 NS_19 0 -5.0255515141290581e-06
GC_7_20 b_7 NI_7 NS_20 0 -5.5563156270066863e-05
GC_7_21 b_7 NI_7 NS_21 0 -2.4322595081285289e-05
GC_7_22 b_7 NI_7 NS_22 0 -1.2674778812100727e-05
GC_7_23 b_7 NI_7 NS_23 0 5.7935595020851473e-07
GC_7_24 b_7 NI_7 NS_24 0 -6.2107062017573765e-07
GC_7_25 b_7 NI_7 NS_25 0 3.4453227700198468e-07
GC_7_26 b_7 NI_7 NS_26 0 1.0390768773123015e-07
GC_7_27 b_7 NI_7 NS_27 0 1.6608213807425085e-10
GC_7_28 b_7 NI_7 NS_28 0 -8.2866519517203862e-11
GC_7_29 b_7 NI_7 NS_29 0 -7.1942968445088252e-11
GC_7_30 b_7 NI_7 NS_30 0 -4.3736248567944955e-10
GC_7_31 b_7 NI_7 NS_31 0 9.9930229682326503e-05
GC_7_32 b_7 NI_7 NS_32 0 -2.5739261910817974e-07
GC_7_33 b_7 NI_7 NS_33 0 3.9431180019964886e-08
GC_7_34 b_7 NI_7 NS_34 0 6.8131648305051008e-10
GC_7_35 b_7 NI_7 NS_35 0 2.6782844498636717e-07
GC_7_36 b_7 NI_7 NS_36 0 -1.4818921682127701e-06
GC_7_37 b_7 NI_7 NS_37 0 -9.2953821889630012e-06
GC_7_38 b_7 NI_7 NS_38 0 2.4293152316411805e-05
GC_7_39 b_7 NI_7 NS_39 0 7.9303136592429244e-05
GC_7_40 b_7 NI_7 NS_40 0 8.7579687659913919e-06
GC_7_41 b_7 NI_7 NS_41 0 1.1180702426789234e-05
GC_7_42 b_7 NI_7 NS_42 0 -7.9803303970227862e-05
GC_7_43 b_7 NI_7 NS_43 0 -7.1787621358255896e-06
GC_7_44 b_7 NI_7 NS_44 0 -4.3358680079807133e-05
GC_7_45 b_7 NI_7 NS_45 0 -9.5157367919046992e-05
GC_7_46 b_7 NI_7 NS_46 0 -5.4098639092592564e-05
GC_7_47 b_7 NI_7 NS_47 0 -4.5957062077985595e-05
GC_7_48 b_7 NI_7 NS_48 0 5.3040645159368834e-05
GC_7_49 b_7 NI_7 NS_49 0 -3.1272898078277762e-05
GC_7_50 b_7 NI_7 NS_50 0 1.2847064456430015e-05
GC_7_51 b_7 NI_7 NS_51 0 -1.6072318556668330e-05
GC_7_52 b_7 NI_7 NS_52 0 4.9857336992617643e-05
GC_7_53 b_7 NI_7 NS_53 0 -7.4582985130104990e-07
GC_7_54 b_7 NI_7 NS_54 0 -4.3446850349217280e-07
GC_7_55 b_7 NI_7 NS_55 0 1.2918945522139137e-07
GC_7_56 b_7 NI_7 NS_56 0 -3.6965426676560518e-07
GC_7_57 b_7 NI_7 NS_57 0 -1.5102427386712086e-10
GC_7_58 b_7 NI_7 NS_58 0 9.1264380995904376e-11
GC_7_59 b_7 NI_7 NS_59 0 7.1484119795148135e-11
GC_7_60 b_7 NI_7 NS_60 0 4.3623182074164620e-10
GC_7_61 b_7 NI_7 NS_61 0 1.3848393150009489e-04
GC_7_62 b_7 NI_7 NS_62 0 1.3826445703650613e-06
GC_7_63 b_7 NI_7 NS_63 0 -2.0149254429599302e-07
GC_7_64 b_7 NI_7 NS_64 0 -9.3083373162940698e-09
GC_7_65 b_7 NI_7 NS_65 0 4.9978472949828316e-05
GC_7_66 b_7 NI_7 NS_66 0 -1.9598859220419896e-06
GC_7_67 b_7 NI_7 NS_67 0 2.5680848987425014e-05
GC_7_68 b_7 NI_7 NS_68 0 -7.5195360073093233e-06
GC_7_69 b_7 NI_7 NS_69 0 2.2272048670392264e-05
GC_7_70 b_7 NI_7 NS_70 0 -2.6882874683454807e-04
GC_7_71 b_7 NI_7 NS_71 0 -2.9200588313070671e-04
GC_7_72 b_7 NI_7 NS_72 0 4.0810789813992810e-05
GC_7_73 b_7 NI_7 NS_73 0 -5.4965813040212242e-05
GC_7_74 b_7 NI_7 NS_74 0 2.2142104839290133e-04
GC_7_75 b_7 NI_7 NS_75 0 1.6790676971944953e-04
GC_7_76 b_7 NI_7 NS_76 0 -1.0526825919102777e-04
GC_7_77 b_7 NI_7 NS_77 0 -1.8088182197284995e-04
GC_7_78 b_7 NI_7 NS_78 0 6.1686549163056303e-05
GC_7_79 b_7 NI_7 NS_79 0 -5.0481355991807749e-05
GC_7_80 b_7 NI_7 NS_80 0 1.2078608411477899e-04
GC_7_81 b_7 NI_7 NS_81 0 1.3701556639138590e-04
GC_7_82 b_7 NI_7 NS_82 0 7.0686012092327106e-05
GC_7_83 b_7 NI_7 NS_83 0 -1.0585906323335231e-07
GC_7_84 b_7 NI_7 NS_84 0 4.3444543426625791e-06
GC_7_85 b_7 NI_7 NS_85 0 -2.0219892499067320e-06
GC_7_86 b_7 NI_7 NS_86 0 1.8441394708677857e-08
GC_7_87 b_7 NI_7 NS_87 0 6.0917253196313035e-10
GC_7_88 b_7 NI_7 NS_88 0 -6.4486072827060391e-10
GC_7_89 b_7 NI_7 NS_89 0 -1.4660654046829325e-10
GC_7_90 b_7 NI_7 NS_90 0 -1.2238416593714880e-09
GC_7_91 b_7 NI_7 NS_91 0 5.4738142990692918e-05
GC_7_92 b_7 NI_7 NS_92 0 9.2112448095261283e-05
GC_7_93 b_7 NI_7 NS_93 0 2.8701184943729348e-07
GC_7_94 b_7 NI_7 NS_94 0 8.4903194648835753e-09
GC_7_95 b_7 NI_7 NS_95 0 -4.0119214290223885e-05
GC_7_96 b_7 NI_7 NS_96 0 -8.6005710747797653e-05
GC_7_97 b_7 NI_7 NS_97 0 -2.2672226237512087e-04
GC_7_98 b_7 NI_7 NS_98 0 9.6554307186504191e-05
GC_7_99 b_7 NI_7 NS_99 0 2.8122318410562499e-04
GC_7_100 b_7 NI_7 NS_100 0 1.5448269748406074e-04
GC_7_101 b_7 NI_7 NS_101 0 -3.0715716311536015e-04
GC_7_102 b_7 NI_7 NS_102 0 -2.0845982436700156e-04
GC_7_103 b_7 NI_7 NS_103 0 1.8399114651144514e-04
GC_7_104 b_7 NI_7 NS_104 0 3.9106493780154675e-04
GC_7_105 b_7 NI_7 NS_105 0 -9.4953714286868880e-05
GC_7_106 b_7 NI_7 NS_106 0 -1.5522812663418273e-04
GC_7_107 b_7 NI_7 NS_107 0 2.3741515494735480e-04
GC_7_108 b_7 NI_7 NS_108 0 2.1644232841872105e-04
GC_7_109 b_7 NI_7 NS_109 0 -5.9512662437023274e-05
GC_7_110 b_7 NI_7 NS_110 0 -2.0712466055223551e-04
GC_7_111 b_7 NI_7 NS_111 0 -2.1944935212442949e-06
GC_7_112 b_7 NI_7 NS_112 0 2.1430414522613912e-04
GC_7_113 b_7 NI_7 NS_113 0 -2.2385967373590619e-06
GC_7_114 b_7 NI_7 NS_114 0 6.4695993464487365e-08
GC_7_115 b_7 NI_7 NS_115 0 -4.6490657568477761e-07
GC_7_116 b_7 NI_7 NS_116 0 -4.5323208971717019e-07
GC_7_117 b_7 NI_7 NS_117 0 -7.2776886970675795e-10
GC_7_118 b_7 NI_7 NS_118 0 5.1680350425232345e-10
GC_7_119 b_7 NI_7 NS_119 0 1.4749279529941489e-10
GC_7_120 b_7 NI_7 NS_120 0 1.2209615899592015e-09
GC_7_121 b_7 NI_7 NS_121 0 -4.2988052038290566e-04
GC_7_122 b_7 NI_7 NS_122 0 -2.9336422244616292e-03
GC_7_123 b_7 NI_7 NS_123 0 -5.9839359493132102e-06
GC_7_124 b_7 NI_7 NS_124 0 -3.8844121115232374e-07
GC_7_125 b_7 NI_7 NS_125 0 2.6783419208677630e-03
GC_7_126 b_7 NI_7 NS_126 0 -1.9922212938142192e-03
GC_7_127 b_7 NI_7 NS_127 0 -6.2097780491403871e-03
GC_7_128 b_7 NI_7 NS_128 0 1.7605677202605996e-03
GC_7_129 b_7 NI_7 NS_129 0 4.7592133388197439e-03
GC_7_130 b_7 NI_7 NS_130 0 -5.5072000178070105e-03
GC_7_131 b_7 NI_7 NS_131 0 -2.2146125338748989e-04
GC_7_132 b_7 NI_7 NS_132 0 7.2473058856116481e-03
GC_7_133 b_7 NI_7 NS_133 0 -6.3292952035544766e-03
GC_7_134 b_7 NI_7 NS_134 0 -5.0696861088136563e-03
GC_7_135 b_7 NI_7 NS_135 0 4.4823182983335340e-03
GC_7_136 b_7 NI_7 NS_136 0 -1.6976962329514004e-03
GC_7_137 b_7 NI_7 NS_137 0 -5.7700545307211976e-04
GC_7_138 b_7 NI_7 NS_138 0 6.9526874784096790e-03
GC_7_139 b_7 NI_7 NS_139 0 -3.4461627633188170e-03
GC_7_140 b_7 NI_7 NS_140 0 -3.6908760057206614e-03
GC_7_141 b_7 NI_7 NS_141 0 5.8924899006941329e-03
GC_7_142 b_7 NI_7 NS_142 0 3.8135578020036888e-04
GC_7_143 b_7 NI_7 NS_143 0 6.0575568528399606e-05
GC_7_144 b_7 NI_7 NS_144 0 6.7951427454909233e-06
GC_7_145 b_7 NI_7 NS_145 0 1.5523879572243372e-05
GC_7_146 b_7 NI_7 NS_146 0 3.8659068401762116e-05
GC_7_147 b_7 NI_7 NS_147 0 6.7893105569896342e-09
GC_7_148 b_7 NI_7 NS_148 0 -2.9476098365481575e-08
GC_7_149 b_7 NI_7 NS_149 0 -1.8905813247331097e-09
GC_7_150 b_7 NI_7 NS_150 0 -5.6443499855184025e-10
GC_7_151 b_7 NI_7 NS_151 0 1.0840922670246537e-03
GC_7_152 b_7 NI_7 NS_152 0 -1.1636889249524048e-03
GC_7_153 b_7 NI_7 NS_153 0 3.5431778317845473e-06
GC_7_154 b_7 NI_7 NS_154 0 2.9212403421921495e-07
GC_7_155 b_7 NI_7 NS_155 0 1.4064404222740798e-04
GC_7_156 b_7 NI_7 NS_156 0 8.9896530515383433e-04
GC_7_157 b_7 NI_7 NS_157 0 1.8646089535908404e-03
GC_7_158 b_7 NI_7 NS_158 0 -8.6916670552580834e-04
GC_7_159 b_7 NI_7 NS_159 0 -2.9480987198010214e-03
GC_7_160 b_7 NI_7 NS_160 0 -1.6595206254428928e-03
GC_7_161 b_7 NI_7 NS_161 0 2.2564581467825525e-03
GC_7_162 b_7 NI_7 NS_162 0 2.6488456344150326e-03
GC_7_163 b_7 NI_7 NS_163 0 -1.4346094264205717e-03
GC_7_164 b_7 NI_7 NS_164 0 -2.9589610827340752e-03
GC_7_165 b_7 NI_7 NS_165 0 1.0713443603436201e-03
GC_7_166 b_7 NI_7 NS_166 0 2.2277942478627082e-03
GC_7_167 b_7 NI_7 NS_167 0 -1.6363481363665196e-03
GC_7_168 b_7 NI_7 NS_168 0 -2.1584332926056944e-03
GC_7_169 b_7 NI_7 NS_169 0 4.3014456973562395e-04
GC_7_170 b_7 NI_7 NS_170 0 2.0082070964713167e-03
GC_7_171 b_7 NI_7 NS_171 0 2.5563233020226136e-04
GC_7_172 b_7 NI_7 NS_172 0 -2.1120365753270086e-03
GC_7_173 b_7 NI_7 NS_173 0 -8.3367111622941104e-08
GC_7_174 b_7 NI_7 NS_174 0 5.0560805793950593e-06
GC_7_175 b_7 NI_7 NS_175 0 -7.2970510681857430e-07
GC_7_176 b_7 NI_7 NS_176 0 -1.7733987878528091e-06
GC_7_177 b_7 NI_7 NS_177 0 -6.9274348772880443e-09
GC_7_178 b_7 NI_7 NS_178 0 2.2849910037722338e-08
GC_7_179 b_7 NI_7 NS_179 0 2.3580829732977999e-09
GC_7_180 b_7 NI_7 NS_180 0 1.5278538684477850e-09
GC_7_181 b_7 NI_7 NS_181 0 1.2599076361271955e-01
GC_7_182 b_7 NI_7 NS_182 0 -9.9112080127415313e-03
GC_7_183 b_7 NI_7 NS_183 0 -2.0441607351726244e-05
GC_7_184 b_7 NI_7 NS_184 0 -3.8242989525754314e-06
GC_7_185 b_7 NI_7 NS_185 0 -8.0690526843633960e-03
GC_7_186 b_7 NI_7 NS_186 0 6.6387582309224288e-04
GC_7_187 b_7 NI_7 NS_187 0 -1.9547028587339576e-03
GC_7_188 b_7 NI_7 NS_188 0 7.9835083278134968e-05
GC_7_189 b_7 NI_7 NS_189 0 -1.2548143124636722e-02
GC_7_190 b_7 NI_7 NS_190 0 8.2410833341110250e-03
GC_7_191 b_7 NI_7 NS_191 0 -1.0211195942393347e-02
GC_7_192 b_7 NI_7 NS_192 0 -6.2935725908548461e-04
GC_7_193 b_7 NI_7 NS_193 0 -3.4910933020387007e-03
GC_7_194 b_7 NI_7 NS_194 0 1.6912358811950193e-02
GC_7_195 b_7 NI_7 NS_195 0 -7.7475184677850278e-03
GC_7_196 b_7 NI_7 NS_196 0 1.3307968081950096e-02
GC_7_197 b_7 NI_7 NS_197 0 -3.9569371169058641e-03
GC_7_198 b_7 NI_7 NS_198 0 6.8929712631648071e-03
GC_7_199 b_7 NI_7 NS_199 0 -2.7322546574418006e-03
GC_7_200 b_7 NI_7 NS_200 0 1.2270498206423825e-02
GC_7_201 b_7 NI_7 NS_201 0 -2.2866223595561938e-02
GC_7_202 b_7 NI_7 NS_202 0 5.9252190904824425e-03
GC_7_203 b_7 NI_7 NS_203 0 -8.5896996238840530e-04
GC_7_204 b_7 NI_7 NS_204 0 7.9678388920307306e-04
GC_7_205 b_7 NI_7 NS_205 0 -5.1011839415658080e-04
GC_7_206 b_7 NI_7 NS_206 0 -4.3700574101341249e-04
GC_7_207 b_7 NI_7 NS_207 0 -6.4199378436639210e-08
GC_7_208 b_7 NI_7 NS_208 0 -1.9083810202951794e-07
GC_7_209 b_7 NI_7 NS_209 0 -3.1375533761581488e-09
GC_7_210 b_7 NI_7 NS_210 0 5.5115721586700449e-09
GC_7_211 b_7 NI_7 NS_211 0 -7.5339438971634878e-02
GC_7_212 b_7 NI_7 NS_212 0 2.4883735290169115e-02
GC_7_213 b_7 NI_7 NS_213 0 1.9330101656498309e-05
GC_7_214 b_7 NI_7 NS_214 0 5.3843320981045828e-06
GC_7_215 b_7 NI_7 NS_215 0 1.8356559283443815e-02
GC_7_216 b_7 NI_7 NS_216 0 2.7965831409430483e-02
GC_7_217 b_7 NI_7 NS_217 0 -1.9176389408365472e-02
GC_7_218 b_7 NI_7 NS_218 0 8.3763464295342933e-03
GC_7_219 b_7 NI_7 NS_219 0 -5.5266990683682047e-03
GC_7_220 b_7 NI_7 NS_220 0 -2.3054642516386264e-02
GC_7_221 b_7 NI_7 NS_221 0 2.6686352844859890e-02
GC_7_222 b_7 NI_7 NS_222 0 -1.4570102538051653e-02
GC_7_223 b_7 NI_7 NS_223 0 3.4524064253645251e-02
GC_7_224 b_7 NI_7 NS_224 0 4.8600617039194129e-03
GC_7_225 b_7 NI_7 NS_225 0 9.6777250457072833e-03
GC_7_226 b_7 NI_7 NS_226 0 1.3687334236118405e-02
GC_7_227 b_7 NI_7 NS_227 0 -1.2366653928528707e-02
GC_7_228 b_7 NI_7 NS_228 0 1.1002968061165630e-02
GC_7_229 b_7 NI_7 NS_229 0 -1.1776682646439770e-02
GC_7_230 b_7 NI_7 NS_230 0 -1.2018486469441121e-02
GC_7_231 b_7 NI_7 NS_231 0 1.9787674007401265e-02
GC_7_232 b_7 NI_7 NS_232 0 -2.6040618793129522e-02
GC_7_233 b_7 NI_7 NS_233 0 9.6541196834647180e-04
GC_7_234 b_7 NI_7 NS_234 0 -1.0850268989447927e-03
GC_7_235 b_7 NI_7 NS_235 0 6.3206516088480560e-04
GC_7_236 b_7 NI_7 NS_236 0 3.4856881828651965e-04
GC_7_237 b_7 NI_7 NS_237 0 9.6067727322425791e-08
GC_7_238 b_7 NI_7 NS_238 0 4.1718988322608288e-07
GC_7_239 b_7 NI_7 NS_239 0 -1.0291247108829765e-08
GC_7_240 b_7 NI_7 NS_240 0 -1.9939675234813333e-08
GC_7_241 b_7 NI_7 NS_241 0 2.2669800212217731e-03
GC_7_242 b_7 NI_7 NS_242 0 -7.3271184793637653e-04
GC_7_243 b_7 NI_7 NS_243 0 -1.8145925515516780e-06
GC_7_244 b_7 NI_7 NS_244 0 -1.2100366346738890e-07
GC_7_245 b_7 NI_7 NS_245 0 3.5967389933553201e-04
GC_7_246 b_7 NI_7 NS_246 0 -3.7513265312498115e-04
GC_7_247 b_7 NI_7 NS_247 0 -1.2776934268300304e-03
GC_7_248 b_7 NI_7 NS_248 0 3.4323481760049527e-04
GC_7_249 b_7 NI_7 NS_249 0 7.1251046995014224e-04
GC_7_250 b_7 NI_7 NS_250 0 -8.2802878810151197e-04
GC_7_251 b_7 NI_7 NS_251 0 -1.5019445020390099e-04
GC_7_252 b_7 NI_7 NS_252 0 1.3911406003856085e-03
GC_7_253 b_7 NI_7 NS_253 0 -1.3011798115130772e-03
GC_7_254 b_7 NI_7 NS_254 0 -7.6470496628228417e-04
GC_7_255 b_7 NI_7 NS_255 0 6.8660249326417291e-04
GC_7_256 b_7 NI_7 NS_256 0 -2.8573053935910821e-05
GC_7_257 b_7 NI_7 NS_257 0 -1.3696246576587400e-04
GC_7_258 b_7 NI_7 NS_258 0 1.4682625691808586e-03
GC_7_259 b_7 NI_7 NS_259 0 -7.1835131342257933e-04
GC_7_260 b_7 NI_7 NS_260 0 -5.4301922806738979e-04
GC_7_261 b_7 NI_7 NS_261 0 6.5087457235514891e-04
GC_7_262 b_7 NI_7 NS_262 0 1.9310986966556548e-04
GC_7_263 b_7 NI_7 NS_263 0 -3.0193392365254942e-06
GC_7_264 b_7 NI_7 NS_264 0 2.6012932966880591e-05
GC_7_265 b_7 NI_7 NS_265 0 -9.9212370796079498e-06
GC_7_266 b_7 NI_7 NS_266 0 -1.4257832993561649e-06
GC_7_267 b_7 NI_7 NS_267 0 7.0597005966563206e-09
GC_7_268 b_7 NI_7 NS_268 0 -1.0480243407384705e-08
GC_7_269 b_7 NI_7 NS_269 0 -6.2223258839125395e-10
GC_7_270 b_7 NI_7 NS_270 0 -2.1193868104308223e-09
GC_7_271 b_7 NI_7 NS_271 0 9.8222030621349077e-04
GC_7_272 b_7 NI_7 NS_272 0 -3.4568952204080809e-04
GC_7_273 b_7 NI_7 NS_273 0 2.1363494648340069e-06
GC_7_274 b_7 NI_7 NS_274 0 8.2059474661047428e-08
GC_7_275 b_7 NI_7 NS_275 0 1.1718806334637791e-05
GC_7_276 b_7 NI_7 NS_276 0 8.7362348539828964e-05
GC_7_277 b_7 NI_7 NS_277 0 3.1568319952669522e-04
GC_7_278 b_7 NI_7 NS_278 0 -1.1545911805289533e-04
GC_7_279 b_7 NI_7 NS_279 0 -5.1920857260506781e-04
GC_7_280 b_7 NI_7 NS_280 0 -2.4291005045192613e-04
GC_7_281 b_7 NI_7 NS_281 0 3.2786467014177825e-04
GC_7_282 b_7 NI_7 NS_282 0 3.8890649165207729e-04
GC_7_283 b_7 NI_7 NS_283 0 -3.2493968117156729e-04
GC_7_284 b_7 NI_7 NS_284 0 -5.5996074920638332e-04
GC_7_285 b_7 NI_7 NS_285 0 7.3917211881945085e-05
GC_7_286 b_7 NI_7 NS_286 0 3.8468623991006449e-04
GC_7_287 b_7 NI_7 NS_287 0 -3.5604784948680269e-04
GC_7_288 b_7 NI_7 NS_288 0 -2.6841050059363177e-04
GC_7_289 b_7 NI_7 NS_289 0 5.3022462075263313e-06
GC_7_290 b_7 NI_7 NS_290 0 4.0801997346943979e-04
GC_7_291 b_7 NI_7 NS_291 0 -9.5158001109067210e-05
GC_7_292 b_7 NI_7 NS_292 0 -3.4082250144684234e-04
GC_7_293 b_7 NI_7 NS_293 0 -1.4814592615129901e-05
GC_7_294 b_7 NI_7 NS_294 0 -8.4885222527748674e-06
GC_7_295 b_7 NI_7 NS_295 0 2.7376409654283980e-06
GC_7_296 b_7 NI_7 NS_296 0 -6.6723225822819260e-06
GC_7_297 b_7 NI_7 NS_297 0 -7.7197737704248881e-09
GC_7_298 b_7 NI_7 NS_298 0 4.8068825250161712e-09
GC_7_299 b_7 NI_7 NS_299 0 1.1496283846969446e-09
GC_7_300 b_7 NI_7 NS_300 0 2.7805514270402454e-09
GC_7_301 b_7 NI_7 NS_301 0 1.1737144757328107e-04
GC_7_302 b_7 NI_7 NS_302 0 4.0259730818298561e-06
GC_7_303 b_7 NI_7 NS_303 0 -2.0970088800893805e-07
GC_7_304 b_7 NI_7 NS_304 0 -9.1846099447886345e-09
GC_7_305 b_7 NI_7 NS_305 0 5.0822812799751389e-05
GC_7_306 b_7 NI_7 NS_306 0 -1.6606067970578384e-06
GC_7_307 b_7 NI_7 NS_307 0 2.6862077357652854e-05
GC_7_308 b_7 NI_7 NS_308 0 -7.4538578576212163e-06
GC_7_309 b_7 NI_7 NS_309 0 2.3829669918133206e-05
GC_7_310 b_7 NI_7 NS_310 0 -2.6937137615299885e-04
GC_7_311 b_7 NI_7 NS_311 0 -2.9022335991201907e-04
GC_7_312 b_7 NI_7 NS_312 0 3.9958670656614478e-05
GC_7_313 b_7 NI_7 NS_313 0 -5.3672778565882958e-05
GC_7_314 b_7 NI_7 NS_314 0 2.1969145544923889e-04
GC_7_315 b_7 NI_7 NS_315 0 1.6888955693291675e-04
GC_7_316 b_7 NI_7 NS_316 0 -1.0703566531095523e-04
GC_7_317 b_7 NI_7 NS_317 0 -1.7982839593148122e-04
GC_7_318 b_7 NI_7 NS_318 0 5.9624845915312533e-05
GC_7_319 b_7 NI_7 NS_319 0 -4.9612695057050068e-05
GC_7_320 b_7 NI_7 NS_320 0 1.1944079420544327e-04
GC_7_321 b_7 NI_7 NS_321 0 1.4033724948066560e-04
GC_7_322 b_7 NI_7 NS_322 0 7.0104839797677760e-05
GC_7_323 b_7 NI_7 NS_323 0 1.2844109247913522e-07
GC_7_324 b_7 NI_7 NS_324 0 4.2771201675911977e-06
GC_7_325 b_7 NI_7 NS_325 0 -1.9736722875100915e-06
GC_7_326 b_7 NI_7 NS_326 0 1.1969799575953979e-07
GC_7_327 b_7 NI_7 NS_327 0 6.3201777010922842e-10
GC_7_328 b_7 NI_7 NS_328 0 -6.2610964396799064e-10
GC_7_329 b_7 NI_7 NS_329 0 -1.5199178566256865e-10
GC_7_330 b_7 NI_7 NS_330 0 -1.2381057969313265e-09
GC_7_331 b_7 NI_7 NS_331 0 4.6478479905190400e-05
GC_7_332 b_7 NI_7 NS_332 0 9.2529797701376140e-05
GC_7_333 b_7 NI_7 NS_333 0 2.8968373871606788e-07
GC_7_334 b_7 NI_7 NS_334 0 8.4521572703754866e-09
GC_7_335 b_7 NI_7 NS_335 0 -3.9577689814023113e-05
GC_7_336 b_7 NI_7 NS_336 0 -8.5753646966473101e-05
GC_7_337 b_7 NI_7 NS_337 0 -2.2600523007570736e-04
GC_7_338 b_7 NI_7 NS_338 0 9.6583221706585145e-05
GC_7_339 b_7 NI_7 NS_339 0 2.8263681002332869e-04
GC_7_340 b_7 NI_7 NS_340 0 1.5421636275975359e-04
GC_7_341 b_7 NI_7 NS_341 0 -3.0568636052722868e-04
GC_7_342 b_7 NI_7 NS_342 0 -2.0974779162364344e-04
GC_7_343 b_7 NI_7 NS_343 0 1.8427059531911008e-04
GC_7_344 b_7 NI_7 NS_344 0 3.8931159002504286e-04
GC_7_345 b_7 NI_7 NS_345 0 -9.5460094141764287e-05
GC_7_346 b_7 NI_7 NS_346 0 -1.5686561283551089e-04
GC_7_347 b_7 NI_7 NS_347 0 2.3694532129009345e-04
GC_7_348 b_7 NI_7 NS_348 0 2.1575073803471837e-04
GC_7_349 b_7 NI_7 NS_349 0 -5.9308460819697873e-05
GC_7_350 b_7 NI_7 NS_350 0 -2.0763778256266616e-04
GC_7_351 b_7 NI_7 NS_351 0 -1.2638894916257193e-06
GC_7_352 b_7 NI_7 NS_352 0 2.1361782612738488e-04
GC_7_353 b_7 NI_7 NS_353 0 -2.2353357046790214e-06
GC_7_354 b_7 NI_7 NS_354 0 -4.6168220698467330e-08
GC_7_355 b_7 NI_7 NS_355 0 -4.0400834376076010e-07
GC_7_356 b_7 NI_7 NS_356 0 -4.3854113048578428e-07
GC_7_357 b_7 NI_7 NS_357 0 -7.4184943205256972e-10
GC_7_358 b_7 NI_7 NS_358 0 5.0959123194604516e-10
GC_7_359 b_7 NI_7 NS_359 0 1.5238772785782757e-10
GC_7_360 b_7 NI_7 NS_360 0 1.2350645631444497e-09
GD_7_1 b_7 NI_7 NA_1 0 2.0740548355161132e-06
GD_7_2 b_7 NI_7 NA_2 0 8.3717115848551148e-06
GD_7_3 b_7 NI_7 NA_3 0 1.6924455844464866e-04
GD_7_4 b_7 NI_7 NA_4 0 -6.2842244272549432e-05
GD_7_5 b_7 NI_7 NA_5 0 1.6033810388021739e-02
GD_7_6 b_7 NI_7 NA_6 0 -3.7759943577884097e-05
GD_7_7 b_7 NI_7 NA_7 0 -4.0224702549935182e-02
GD_7_8 b_7 NI_7 NA_8 0 -9.9740318182197293e-03
GD_7_9 b_7 NI_7 NA_9 0 2.3297112132932554e-03
GD_7_10 b_7 NI_7 NA_10 0 -4.6762441596145187e-05
GD_7_11 b_7 NI_7 NA_11 0 1.7232177003560184e-04
GD_7_12 b_7 NI_7 NA_12 0 -6.0828850588476980e-05
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 9.8877786572450113e-05
GC_8_2 b_8 NI_8 NS_2 0 -1.7559974497400706e-07
GC_8_3 b_8 NI_8 NS_3 0 3.9323533028354311e-08
GC_8_4 b_8 NI_8 NS_4 0 6.8242734945029720e-10
GC_8_5 b_8 NI_8 NS_5 0 4.2701060512216410e-07
GC_8_6 b_8 NI_8 NS_6 0 -1.4257168160955722e-06
GC_8_7 b_8 NI_8 NS_7 0 -9.1784464471381652e-06
GC_8_8 b_8 NI_8 NS_8 0 2.4322921138164567e-05
GC_8_9 b_8 NI_8 NS_9 0 7.9325301007692787e-05
GC_8_10 b_8 NI_8 NS_10 0 8.5014430489423639e-06
GC_8_11 b_8 NI_8 NS_11 0 1.1235554762359245e-05
GC_8_12 b_8 NI_8 NS_12 0 -7.9840732596104733e-05
GC_8_13 b_8 NI_8 NS_13 0 -7.0607551267935109e-06
GC_8_14 b_8 NI_8 NS_14 0 -4.3550071605079858e-05
GC_8_15 b_8 NI_8 NS_15 0 -9.5183559618506659e-05
GC_8_16 b_8 NI_8 NS_16 0 -5.4168022900665610e-05
GC_8_17 b_8 NI_8 NS_17 0 -4.5943856557457020e-05
GC_8_18 b_8 NI_8 NS_18 0 5.2906451290963879e-05
GC_8_19 b_8 NI_8 NS_19 0 -3.1270743278443057e-05
GC_8_20 b_8 NI_8 NS_20 0 1.2779482423343480e-05
GC_8_21 b_8 NI_8 NS_21 0 -1.5940310585770982e-05
GC_8_22 b_8 NI_8 NS_22 0 4.9776957101643266e-05
GC_8_23 b_8 NI_8 NS_23 0 -7.4154406111243682e-07
GC_8_24 b_8 NI_8 NS_24 0 -4.3929228906798716e-07
GC_8_25 b_8 NI_8 NS_25 0 1.3271423576487225e-07
GC_8_26 b_8 NI_8 NS_26 0 -3.6747224688624590e-07
GC_8_27 b_8 NI_8 NS_27 0 -1.5075737032610264e-10
GC_8_28 b_8 NI_8 NS_28 0 9.1441469323521283e-11
GC_8_29 b_8 NI_8 NS_29 0 7.1476089426826352e-11
GC_8_30 b_8 NI_8 NS_30 0 4.3621313945372260e-10
GC_8_31 b_8 NI_8 NS_31 0 -4.8030176433698773e-05
GC_8_32 b_8 NI_8 NS_32 0 -6.2106734560762067e-06
GC_8_33 b_8 NI_8 NS_33 0 -5.0822347351583310e-08
GC_8_34 b_8 NI_8 NS_34 0 -6.2461126638357417e-10
GC_8_35 b_8 NI_8 NS_35 0 -7.2122565890876776e-06
GC_8_36 b_8 NI_8 NS_36 0 -5.3858958983423357e-06
GC_8_37 b_8 NI_8 NS_37 0 -3.2447467519246173e-05
GC_8_38 b_8 NI_8 NS_38 0 1.3398731295429836e-05
GC_8_39 b_8 NI_8 NS_39 0 1.9868488164544676e-05
GC_8_40 b_8 NI_8 NS_40 0 6.7344523967674368e-05
GC_8_41 b_8 NI_8 NS_41 0 9.5695706517679821e-05
GC_8_42 b_8 NI_8 NS_42 0 5.2354548788194113e-06
GC_8_43 b_8 NI_8 NS_43 0 -1.6522316905091303e-05
GC_8_44 b_8 NI_8 NS_44 0 -8.9248188846275935e-05
GC_8_45 b_8 NI_8 NS_45 0 -2.8891587537652362e-05
GC_8_46 b_8 NI_8 NS_46 0 3.4604100542195937e-05
GC_8_47 b_8 NI_8 NS_47 0 5.9453626652958950e-05
GC_8_48 b_8 NI_8 NS_48 0 -3.6932690027875347e-06
GC_8_49 b_8 NI_8 NS_49 0 -5.0298055173996108e-06
GC_8_50 b_8 NI_8 NS_50 0 -5.5556149421469150e-05
GC_8_51 b_8 NI_8 NS_51 0 -2.4338390153477108e-05
GC_8_52 b_8 NI_8 NS_52 0 -1.2670120704755404e-05
GC_8_53 b_8 NI_8 NS_53 0 5.7847784004585310e-07
GC_8_54 b_8 NI_8 NS_54 0 -6.2045984768338244e-07
GC_8_55 b_8 NI_8 NS_55 0 3.4415512365595091e-07
GC_8_56 b_8 NI_8 NS_56 0 1.0348450793764513e-07
GC_8_57 b_8 NI_8 NS_57 0 1.6603336845254201e-10
GC_8_58 b_8 NI_8 NS_58 0 -8.2919047685956579e-11
GC_8_59 b_8 NI_8 NS_59 0 -7.1939845563505141e-11
GC_8_60 b_8 NI_8 NS_60 0 -4.3735874460077014e-10
GC_8_61 b_8 NI_8 NS_61 0 5.4748184181781756e-05
GC_8_62 b_8 NI_8 NS_62 0 9.2111723374299411e-05
GC_8_63 b_8 NI_8 NS_63 0 2.8701247430131636e-07
GC_8_64 b_8 NI_8 NS_64 0 8.4903048168274525e-09
GC_8_65 b_8 NI_8 NS_65 0 -4.0119715726193095e-05
GC_8_66 b_8 NI_8 NS_66 0 -8.6005424880713377e-05
GC_8_67 b_8 NI_8 NS_67 0 -2.2672225462969778e-04
GC_8_68 b_8 NI_8 NS_68 0 9.6553936958964403e-05
GC_8_69 b_8 NI_8 NS_69 0 2.8122160575699037e-04
GC_8_70 b_8 NI_8 NS_70 0 1.5448308319063498e-04
GC_8_71 b_8 NI_8 NS_71 0 -3.0715790431761202e-04
GC_8_72 b_8 NI_8 NS_72 0 -2.0845896011364203e-04
GC_8_73 b_8 NI_8 NS_73 0 1.8399027048539315e-04
GC_8_74 b_8 NI_8 NS_74 0 3.9106521065542573e-04
GC_8_75 b_8 NI_8 NS_75 0 -9.4954350926528070e-05
GC_8_76 b_8 NI_8 NS_76 0 -1.5522560000865652e-04
GC_8_77 b_8 NI_8 NS_77 0 2.3741530242283657e-04
GC_8_78 b_8 NI_8 NS_78 0 2.1644330777361291e-04
GC_8_79 b_8 NI_8 NS_79 0 -5.9513289841488136e-05
GC_8_80 b_8 NI_8 NS_80 0 -2.0712363904909671e-04
GC_8_81 b_8 NI_8 NS_81 0 -2.1951460559558422e-06
GC_8_82 b_8 NI_8 NS_82 0 2.1430507509019061e-04
GC_8_83 b_8 NI_8 NS_83 0 -2.2386596911463824e-06
GC_8_84 b_8 NI_8 NS_84 0 6.4753172592564529e-08
GC_8_85 b_8 NI_8 NS_85 0 -4.6493689574682810e-07
GC_8_86 b_8 NI_8 NS_86 0 -4.5326311216055111e-07
GC_8_87 b_8 NI_8 NS_87 0 -7.2777013558652311e-10
GC_8_88 b_8 NI_8 NS_88 0 5.1680150851728063e-10
GC_8_89 b_8 NI_8 NS_89 0 1.4749281167501391e-10
GC_8_90 b_8 NI_8 NS_90 0 1.2209615432424778e-09
GC_8_91 b_8 NI_8 NS_91 0 1.2346779882590840e-04
GC_8_92 b_8 NI_8 NS_92 0 3.0700828568269275e-06
GC_8_93 b_8 NI_8 NS_93 0 -2.0465933803461428e-07
GC_8_94 b_8 NI_8 NS_94 0 -9.2708993117117741e-09
GC_8_95 b_8 NI_8 NS_95 0 5.0562971618427196e-05
GC_8_96 b_8 NI_8 NS_96 0 -1.7974656437339510e-06
GC_8_97 b_8 NI_8 NS_97 0 2.6615714796355954e-05
GC_8_98 b_8 NI_8 NS_98 0 -7.4108934580294550e-06
GC_8_99 b_8 NI_8 NS_99 0 2.3162180768712834e-05
GC_8_100 b_8 NI_8 NS_100 0 -2.6930191864011553e-04
GC_8_101 b_8 NI_8 NS_101 0 -2.9060536205790719e-04
GC_8_102 b_8 NI_8 NS_102 0 4.0320326514362795e-05
GC_8_103 b_8 NI_8 NS_103 0 -5.3916151138489314e-05
GC_8_104 b_8 NI_8 NS_104 0 2.2026889096772291e-04
GC_8_105 b_8 NI_8 NS_105 0 1.6852299351769734e-04
GC_8_106 b_8 NI_8 NS_106 0 -1.0673931031527922e-04
GC_8_107 b_8 NI_8 NS_107 0 -1.8008568543910675e-04
GC_8_108 b_8 NI_8 NS_108 0 6.0276502861850281e-05
GC_8_109 b_8 NI_8 NS_109 0 -4.9794892428343184e-05
GC_8_110 b_8 NI_8 NS_110 0 1.1982017671940831e-04
GC_8_111 b_8 NI_8 NS_111 0 1.3938970163785292e-04
GC_8_112 b_8 NI_8 NS_112 0 7.0034128480645909e-05
GC_8_113 b_8 NI_8 NS_113 0 3.3249683710629592e-08
GC_8_114 b_8 NI_8 NS_114 0 4.2541384003551304e-06
GC_8_115 b_8 NI_8 NS_115 0 -1.9651709190248167e-06
GC_8_116 b_8 NI_8 NS_116 0 8.5734706838959041e-08
GC_8_117 b_8 NI_8 NS_117 0 6.1371545072206439e-10
GC_8_118 b_8 NI_8 NS_118 0 -6.3978983669841191e-10
GC_8_119 b_8 NI_8 NS_119 0 -1.4671798609537537e-10
GC_8_120 b_8 NI_8 NS_120 0 -1.2237848149088651e-09
GC_8_121 b_8 NI_8 NS_121 0 1.0838825755828875e-03
GC_8_122 b_8 NI_8 NS_122 0 -1.1636685876998533e-03
GC_8_123 b_8 NI_8 NS_123 0 3.5431453499449500e-06
GC_8_124 b_8 NI_8 NS_124 0 2.9212450276130969e-07
GC_8_125 b_8 NI_8 NS_125 0 1.4066770003435118e-04
GC_8_126 b_8 NI_8 NS_126 0 8.9897477137551194e-04
GC_8_127 b_8 NI_8 NS_127 0 1.8646238070248017e-03
GC_8_128 b_8 NI_8 NS_128 0 -8.6915569569320154e-04
GC_8_129 b_8 NI_8 NS_129 0 -2.9480926838601298e-03
GC_8_130 b_8 NI_8 NS_130 0 -1.6595552138660634e-03
GC_8_131 b_8 NI_8 NS_131 0 2.2564741211461943e-03
GC_8_132 b_8 NI_8 NS_132 0 2.6488447144518610e-03
GC_8_133 b_8 NI_8 NS_133 0 -1.4345831598167121e-03
GC_8_134 b_8 NI_8 NS_134 0 -2.9589936147707326e-03
GC_8_135 b_8 NI_8 NS_135 0 1.0713460933028146e-03
GC_8_136 b_8 NI_8 NS_136 0 2.2277830877607376e-03
GC_8_137 b_8 NI_8 NS_137 0 -1.6363393917880765e-03
GC_8_138 b_8 NI_8 NS_138 0 -2.1584583361198692e-03
GC_8_139 b_8 NI_8 NS_139 0 4.3014900976300036e-04
GC_8_140 b_8 NI_8 NS_140 0 2.0081938809727888e-03
GC_8_141 b_8 NI_8 NS_141 0 2.5566385172536650e-04
GC_8_142 b_8 NI_8 NS_142 0 -2.1120493467362191e-03
GC_8_143 b_8 NI_8 NS_143 0 -8.1927604122682648e-08
GC_8_144 b_8 NI_8 NS_144 0 5.0549410016988348e-06
GC_8_145 b_8 NI_8 NS_145 0 -7.2891355749680300e-07
GC_8_146 b_8 NI_8 NS_146 0 -1.7726323538580892e-06
GC_8_147 b_8 NI_8 NS_147 0 -6.9273598869386547e-09
GC_8_148 b_8 NI_8 NS_148 0 2.2849982543066883e-08
GC_8_149 b_8 NI_8 NS_149 0 2.3580775417406213e-09
GC_8_150 b_8 NI_8 NS_150 0 1.5278505673224266e-09
GC_8_151 b_8 NI_8 NS_151 0 -4.2988330634121763e-04
GC_8_152 b_8 NI_8 NS_152 0 -2.9336419347796060e-03
GC_8_153 b_8 NI_8 NS_153 0 -5.9839363530271233e-06
GC_8_154 b_8 NI_8 NS_154 0 -3.8844120751575242e-07
GC_8_155 b_8 NI_8 NS_155 0 2.6783420245401388e-03
GC_8_156 b_8 NI_8 NS_156 0 -1.9922212538343136e-03
GC_8_157 b_8 NI_8 NS_157 0 -6.2097779188802415e-03
GC_8_158 b_8 NI_8 NS_158 0 1.7605677112088312e-03
GC_8_159 b_8 NI_8 NS_159 0 4.7592134835835881e-03
GC_8_160 b_8 NI_8 NS_160 0 -5.5072000653056691e-03
GC_8_161 b_8 NI_8 NS_161 0 -2.2146105042577938e-04
GC_8_162 b_8 NI_8 NS_162 0 7.2473058667639808e-03
GC_8_163 b_8 NI_8 NS_163 0 -6.3292949808905008e-03
GC_8_164 b_8 NI_8 NS_164 0 -5.0696862845352846e-03
GC_8_165 b_8 NI_8 NS_165 0 4.4823184746202544e-03
GC_8_166 b_8 NI_8 NS_166 0 -1.6976964447727469e-03
GC_8_167 b_8 NI_8 NS_167 0 -5.7700526280904114e-04
GC_8_168 b_8 NI_8 NS_168 0 6.9526872290205134e-03
GC_8_169 b_8 NI_8 NS_169 0 -3.4461625867765414e-03
GC_8_170 b_8 NI_8 NS_170 0 -3.6908762062469336e-03
GC_8_171 b_8 NI_8 NS_171 0 5.8924903735890211e-03
GC_8_172 b_8 NI_8 NS_172 0 3.8135561389994482e-04
GC_8_173 b_8 NI_8 NS_173 0 6.0575586239374924e-05
GC_8_174 b_8 NI_8 NS_174 0 6.7951232327423930e-06
GC_8_175 b_8 NI_8 NS_175 0 1.5523892175819358e-05
GC_8_176 b_8 NI_8 NS_176 0 3.8659076368951002e-05
GC_8_177 b_8 NI_8 NS_177 0 6.7893114148697358e-09
GC_8_178 b_8 NI_8 NS_178 0 -2.9476097763905418e-08
GC_8_179 b_8 NI_8 NS_179 0 -1.8905813639738569e-09
GC_8_180 b_8 NI_8 NS_180 0 -5.6443499378471121e-10
GC_8_181 b_8 NI_8 NS_181 0 -7.5339251406161614e-02
GC_8_182 b_8 NI_8 NS_182 0 2.4883709961722154e-02
GC_8_183 b_8 NI_8 NS_183 0 1.9330156888161319e-05
GC_8_184 b_8 NI_8 NS_184 0 5.3843307724518299e-06
GC_8_185 b_8 NI_8 NS_185 0 1.8356556297536568e-02
GC_8_186 b_8 NI_8 NS_186 0 2.7965825867945611e-02
GC_8_187 b_8 NI_8 NS_187 0 -1.9176397571209421e-02
GC_8_188 b_8 NI_8 NS_188 0 8.3763414589274939e-03
GC_8_189 b_8 NI_8 NS_189 0 -5.5267117168074078e-03
GC_8_190 b_8 NI_8 NS_190 0 -2.3054643020709600e-02
GC_8_191 b_8 NI_8 NS_191 0 2.6686338102362494e-02
GC_8_192 b_8 NI_8 NS_192 0 -1.4570103098377531e-02
GC_8_193 b_8 NI_8 NS_193 0 3.4524047394794415e-02
GC_8_194 b_8 NI_8 NS_194 0 4.8600710812115545e-03
GC_8_195 b_8 NI_8 NS_195 0 9.6777117074828122e-03
GC_8_196 b_8 NI_8 NS_196 0 1.3687347256441185e-02
GC_8_197 b_8 NI_8 NS_197 0 -1.2366667403668654e-02
GC_8_198 b_8 NI_8 NS_198 0 1.1002982427814868e-02
GC_8_199 b_8 NI_8 NS_199 0 -1.1776695604821837e-02
GC_8_200 b_8 NI_8 NS_200 0 -1.2018476843498296e-02
GC_8_201 b_8 NI_8 NS_201 0 1.9787636315845049e-02
GC_8_202 b_8 NI_8 NS_202 0 -2.6040614865922615e-02
GC_8_203 b_8 NI_8 NS_203 0 9.6540988525443136e-04
GC_8_204 b_8 NI_8 NS_204 0 -1.0850255176153222e-03
GC_8_205 b_8 NI_8 NS_205 0 6.3206423816375532e-04
GC_8_206 b_8 NI_8 NS_206 0 3.4856778305341680e-04
GC_8_207 b_8 NI_8 NS_207 0 9.6067639663910073e-08
GC_8_208 b_8 NI_8 NS_208 0 4.1718959648248321e-07
GC_8_209 b_8 NI_8 NS_209 0 -1.0291219725212227e-08
GC_8_210 b_8 NI_8 NS_210 0 -1.9939654620964741e-08
GC_8_211 b_8 NI_8 NS_211 0 1.2599076361271946e-01
GC_8_212 b_8 NI_8 NS_212 0 -9.9112080127415243e-03
GC_8_213 b_8 NI_8 NS_213 0 -2.0441607351726437e-05
GC_8_214 b_8 NI_8 NS_214 0 -3.8242989525754551e-06
GC_8_215 b_8 NI_8 NS_215 0 -8.0690526843633908e-03
GC_8_216 b_8 NI_8 NS_216 0 6.6387582309224429e-04
GC_8_217 b_8 NI_8 NS_217 0 -1.9547028587339702e-03
GC_8_218 b_8 NI_8 NS_218 0 7.9835083278136920e-05
GC_8_219 b_8 NI_8 NS_219 0 -1.2548143124636722e-02
GC_8_220 b_8 NI_8 NS_220 0 8.2410833341110372e-03
GC_8_221 b_8 NI_8 NS_221 0 -1.0211195942393352e-02
GC_8_222 b_8 NI_8 NS_222 0 -6.2935725908546682e-04
GC_8_223 b_8 NI_8 NS_223 0 -3.4910933020386834e-03
GC_8_224 b_8 NI_8 NS_224 0 1.6912358811950207e-02
GC_8_225 b_8 NI_8 NS_225 0 -7.7475184677849984e-03
GC_8_226 b_8 NI_8 NS_226 0 1.3307968081950092e-02
GC_8_227 b_8 NI_8 NS_227 0 -3.9569371169058572e-03
GC_8_228 b_8 NI_8 NS_228 0 6.8929712631647950e-03
GC_8_229 b_8 NI_8 NS_229 0 -2.7322546574417936e-03
GC_8_230 b_8 NI_8 NS_230 0 1.2270498206423824e-02
GC_8_231 b_8 NI_8 NS_231 0 -2.2866223595561921e-02
GC_8_232 b_8 NI_8 NS_232 0 5.9252190904824364e-03
GC_8_233 b_8 NI_8 NS_233 0 -8.5896996238840650e-04
GC_8_234 b_8 NI_8 NS_234 0 7.9678388920307274e-04
GC_8_235 b_8 NI_8 NS_235 0 -5.1011839415657982e-04
GC_8_236 b_8 NI_8 NS_236 0 -4.3700574101341336e-04
GC_8_237 b_8 NI_8 NS_237 0 -6.4199378436638893e-08
GC_8_238 b_8 NI_8 NS_238 0 -1.9083810202951847e-07
GC_8_239 b_8 NI_8 NS_239 0 -3.1375533761577952e-09
GC_8_240 b_8 NI_8 NS_240 0 5.5115721586691292e-09
GC_8_241 b_8 NI_8 NS_241 0 9.8191779966069412e-04
GC_8_242 b_8 NI_8 NS_242 0 -3.4563458345370196e-04
GC_8_243 b_8 NI_8 NS_243 0 2.1362772083741888e-06
GC_8_244 b_8 NI_8 NS_244 0 8.2059868492505990e-08
GC_8_245 b_8 NI_8 NS_245 0 1.1628698289643525e-05
GC_8_246 b_8 NI_8 NS_246 0 8.7325783942707836e-05
GC_8_247 b_8 NI_8 NS_247 0 3.1565263708250918e-04
GC_8_248 b_8 NI_8 NS_248 0 -1.1551278690767940e-04
GC_8_249 b_8 NI_8 NS_249 0 -5.1916689050861406e-04
GC_8_250 b_8 NI_8 NS_250 0 -2.4271731263572128e-04
GC_8_251 b_8 NI_8 NS_251 0 3.2788840301512505e-04
GC_8_252 b_8 NI_8 NS_252 0 3.8892152452892867e-04
GC_8_253 b_8 NI_8 NS_253 0 -3.2494902875157105e-04
GC_8_254 b_8 NI_8 NS_254 0 -5.5986616108802130e-04
GC_8_255 b_8 NI_8 NS_255 0 7.3998216474239906e-05
GC_8_256 b_8 NI_8 NS_256 0 3.8462936641480962e-04
GC_8_257 b_8 NI_8 NS_257 0 -3.5599623989953201e-04
GC_8_258 b_8 NI_8 NS_258 0 -2.6838291499796721e-04
GC_8_259 b_8 NI_8 NS_259 0 5.3831814408468356e-06
GC_8_260 b_8 NI_8 NS_260 0 4.0799864329136757e-04
GC_8_261 b_8 NI_8 NS_261 0 -9.5065871464297913e-05
GC_8_262 b_8 NI_8 NS_262 0 -3.4082220314271495e-04
GC_8_263 b_8 NI_8 NS_263 0 -1.4810614235155547e-05
GC_8_264 b_8 NI_8 NS_264 0 -8.4933832275382277e-06
GC_8_265 b_8 NI_8 NS_265 0 2.7403456806307032e-06
GC_8_266 b_8 NI_8 NS_266 0 -6.6706399607702683e-06
GC_8_267 b_8 NI_8 NS_267 0 -7.7196779497810798e-09
GC_8_268 b_8 NI_8 NS_268 0 4.8069828057303069e-09
GC_8_269 b_8 NI_8 NS_269 0 1.1496159315032387e-09
GC_8_270 b_8 NI_8 NS_270 0 2.7805452068155977e-09
GC_8_271 b_8 NI_8 NS_271 0 2.2658564448318520e-03
GC_8_272 b_8 NI_8 NS_272 0 -7.3259609540744807e-04
GC_8_273 b_8 NI_8 NS_273 0 -1.8147797949500816e-06
GC_8_274 b_8 NI_8 NS_274 0 -1.2100069774820966e-07
GC_8_275 b_8 NI_8 NS_275 0 3.5972857013983803e-04
GC_8_276 b_8 NI_8 NS_276 0 -3.7512259089745508e-04
GC_8_277 b_8 NI_8 NS_277 0 -1.2776319317232246e-03
GC_8_278 b_8 NI_8 NS_278 0 3.4322714293510390e-04
GC_8_279 b_8 NI_8 NS_279 0 7.1259047115004718e-04
GC_8_280 b_8 NI_8 NS_280 0 -8.2806986813786299e-04
GC_8_281 b_8 NI_8 NS_281 0 -1.5010235007434676e-04
GC_8_282 b_8 NI_8 NS_282 0 1.3910986753145926e-03
GC_8_283 b_8 NI_8 NS_283 0 -1.3011090185239187e-03
GC_8_284 b_8 NI_8 NS_284 0 -7.6481278553710576e-04
GC_8_285 b_8 NI_8 NS_285 0 6.8664558429670124e-04
GC_8_286 b_8 NI_8 NS_286 0 -2.8679358344318256e-05
GC_8_287 b_8 NI_8 NS_287 0 -1.3691887213993368e-04
GC_8_288 b_8 NI_8 NS_288 0 1.4681555604078185e-03
GC_8_289 b_8 NI_8 NS_289 0 -7.1830203043518853e-04
GC_8_290 b_8 NI_8 NS_290 0 -5.4309744759253485e-04
GC_8_291 b_8 NI_8 NS_291 0 6.5104338262691032e-04
GC_8_292 b_8 NI_8 NS_292 0 1.9305495674247394e-04
GC_8_293 b_8 NI_8 NS_293 0 -3.0110342850914789e-06
GC_8_294 b_8 NI_8 NS_294 0 2.6005608500362293e-05
GC_8_295 b_8 NI_8 NS_295 0 -9.9167465879538548e-06
GC_8_296 b_8 NI_8 NS_296 0 -1.4215860849892076e-06
GC_8_297 b_8 NI_8 NS_297 0 7.0600819132830297e-09
GC_8_298 b_8 NI_8 NS_298 0 -1.0479797431619891e-08
GC_8_299 b_8 NI_8 NS_299 0 -6.2224917871337336e-10
GC_8_300 b_8 NI_8 NS_300 0 -2.1194002757355828e-09
GC_8_301 b_8 NI_8 NS_301 0 4.6469696800314238e-05
GC_8_302 b_8 NI_8 NS_302 0 9.2530535087370608e-05
GC_8_303 b_8 NI_8 NS_303 0 2.8969073334388427e-07
GC_8_304 b_8 NI_8 NS_304 0 8.4521963972296529e-09
GC_8_305 b_8 NI_8 NS_305 0 -3.9577516123419140e-05
GC_8_306 b_8 NI_8 NS_306 0 -8.5748799005896568e-05
GC_8_307 b_8 NI_8 NS_307 0 -2.2600756427561326e-04
GC_8_308 b_8 NI_8 NS_308 0 9.6587366021181573e-05
GC_8_309 b_8 NI_8 NS_309 0 2.8264086022554419e-04
GC_8_310 b_8 NI_8 NS_310 0 1.5421249329740491e-04
GC_8_311 b_8 NI_8 NS_311 0 -3.0568685860313927e-04
GC_8_312 b_8 NI_8 NS_312 0 -2.0974507171819386e-04
GC_8_313 b_8 NI_8 NS_313 0 1.8427774460842684e-04
GC_8_314 b_8 NI_8 NS_314 0 3.8931269031669893e-04
GC_8_315 b_8 NI_8 NS_315 0 -9.5460495572826859e-05
GC_8_316 b_8 NI_8 NS_316 0 -1.5686517369835316e-04
GC_8_317 b_8 NI_8 NS_317 0 2.3694874016147503e-04
GC_8_318 b_8 NI_8 NS_318 0 2.1574923644893600e-04
GC_8_319 b_8 NI_8 NS_319 0 -5.9308357006091284e-05
GC_8_320 b_8 NI_8 NS_320 0 -2.0763943777584487e-04
GC_8_321 b_8 NI_8 NS_321 0 -1.2603417247180772e-06
GC_8_322 b_8 NI_8 NS_322 0 2.1361740066367410e-04
GC_8_323 b_8 NI_8 NS_323 0 -2.2353604784447700e-06
GC_8_324 b_8 NI_8 NS_324 0 -4.6374166823600213e-08
GC_8_325 b_8 NI_8 NS_325 0 -4.0397125876825967e-07
GC_8_326 b_8 NI_8 NS_326 0 -4.3861915382881299e-07
GC_8_327 b_8 NI_8 NS_327 0 -7.4187305906314540e-10
GC_8_328 b_8 NI_8 NS_328 0 5.0958795454954410e-10
GC_8_329 b_8 NI_8 NS_329 0 1.5239076169513229e-10
GC_8_330 b_8 NI_8 NS_330 0 1.2350690274386145e-09
GC_8_331 b_8 NI_8 NS_331 0 1.3201863525887680e-04
GC_8_332 b_8 NI_8 NS_332 0 2.3805703140939459e-06
GC_8_333 b_8 NI_8 NS_333 0 -2.0660918475835331e-07
GC_8_334 b_8 NI_8 NS_334 0 -9.2214648069959954e-09
GC_8_335 b_8 NI_8 NS_335 0 5.0256255519114230e-05
GC_8_336 b_8 NI_8 NS_336 0 -1.8215604444958026e-06
GC_8_337 b_8 NI_8 NS_337 0 2.5946087031741702e-05
GC_8_338 b_8 NI_8 NS_338 0 -7.5678259914522154e-06
GC_8_339 b_8 NI_8 NS_339 0 2.2965371885432535e-05
GC_8_340 b_8 NI_8 NS_340 0 -2.6891282361119596e-04
GC_8_341 b_8 NI_8 NS_341 0 -2.9159830509612632e-04
GC_8_342 b_8 NI_8 NS_342 0 4.0432224445736778e-05
GC_8_343 b_8 NI_8 NS_343 0 -5.4703353845516494e-05
GC_8_344 b_8 NI_8 NS_344 0 2.2080859855683505e-04
GC_8_345 b_8 NI_8 NS_345 0 1.6828542721788984e-04
GC_8_346 b_8 NI_8 NS_346 0 -1.0559560020126229e-04
GC_8_347 b_8 NI_8 NS_347 0 -1.8061281390630457e-04
GC_8_348 b_8 NI_8 NS_348 0 6.1001806843218892e-05
GC_8_349 b_8 NI_8 NS_349 0 -5.0282957471464693e-05
GC_8_350 b_8 NI_8 NS_350 0 1.2038418620468663e-04
GC_8_351 b_8 NI_8 NS_351 0 1.3801948292061514e-04
GC_8_352 b_8 NI_8 NS_352 0 7.0744592420768758e-05
GC_8_353 b_8 NI_8 NS_353 0 -7.0769554280203108e-09
GC_8_354 b_8 NI_8 NS_354 0 4.3653237249695982e-06
GC_8_355 b_8 NI_8 NS_355 0 -2.0291298626015703e-06
GC_8_356 b_8 NI_8 NS_356 0 5.4131833807096357e-08
GC_8_357 b_8 NI_8 NS_357 0 6.2761202080330391e-10
GC_8_358 b_8 NI_8 NS_358 0 -6.3109557501478250e-10
GC_8_359 b_8 NI_8 NS_359 0 -1.5188948279510850e-10
GC_8_360 b_8 NI_8 NS_360 0 -1.2381737925183406e-09
GD_8_1 b_8 NI_8 NA_1 0 8.6020236710722875e-06
GD_8_2 b_8 NI_8 NA_2 0 2.0534848324926025e-06
GD_8_3 b_8 NI_8 NA_3 0 -6.2844760212509557e-05
GD_8_4 b_8 NI_8 NA_4 0 1.7128697586485863e-04
GD_8_5 b_8 NI_8 NA_5 0 -3.7727923170489692e-05
GD_8_6 b_8 NI_8 NA_6 0 1.6033810802924393e-02
GD_8_7 b_8 NI_8 NA_7 0 -9.9740453537863587e-03
GD_8_8 b_8 NI_8 NA_8 0 -4.0224702549935133e-02
GD_8_9 b_8 NI_8 NA_9 0 -4.6753669872355310e-05
GD_8_10 b_8 NI_8 NA_10 0 2.3299342725127143e-03
GD_8_11 b_8 NI_8 NA_11 0 -6.0834572687309590e-05
GD_8_12 b_8 NI_8 NA_12 0 1.7036754114433696e-04
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 1.7965862534325096e-05
GC_9_2 b_9 NI_9 NS_2 0 -2.5639521233869823e-06
GC_9_3 b_9 NI_9 NS_3 0 1.0272995194283881e-08
GC_9_4 b_9 NI_9 NS_4 0 -2.6568076290986142e-10
GC_9_5 b_9 NI_9 NS_5 0 -1.2437460577103881e-06
GC_9_6 b_9 NI_9 NS_6 0 -1.1106323020428648e-06
GC_9_7 b_9 NI_9 NS_7 0 -2.4819749076115991e-06
GC_9_8 b_9 NI_9 NS_8 0 5.4032068287584329e-07
GC_9_9 b_9 NI_9 NS_9 0 -1.2563619615356070e-06
GC_9_10 b_9 NI_9 NS_10 0 2.6678122058687846e-06
GC_9_11 b_9 NI_9 NS_11 0 1.8212420645204424e-06
GC_9_12 b_9 NI_9 NS_12 0 7.7843856860556934e-07
GC_9_13 b_9 NI_9 NS_13 0 -2.7681914611851447e-06
GC_9_14 b_9 NI_9 NS_14 0 -1.3641178516243669e-06
GC_9_15 b_9 NI_9 NS_15 0 -2.1614707222325172e-06
GC_9_16 b_9 NI_9 NS_16 0 3.4589232704707156e-06
GC_9_17 b_9 NI_9 NS_17 0 1.2662035217219895e-06
GC_9_18 b_9 NI_9 NS_18 0 2.3623979199001294e-06
GC_9_19 b_9 NI_9 NS_19 0 -9.1304853469336822e-07
GC_9_20 b_9 NI_9 NS_20 0 -3.9147084966136301e-07
GC_9_21 b_9 NI_9 NS_21 0 -3.3032134648907243e-06
GC_9_22 b_9 NI_9 NS_22 0 6.2694710403989278e-07
GC_9_23 b_9 NI_9 NS_23 0 -1.4109290578332321e-07
GC_9_24 b_9 NI_9 NS_24 0 -7.7483884113157127e-08
GC_9_25 b_9 NI_9 NS_25 0 2.3769451642188750e-08
GC_9_26 b_9 NI_9 NS_26 0 -5.0980995248401498e-08
GC_9_27 b_9 NI_9 NS_27 0 -1.7923342531526524e-11
GC_9_28 b_9 NI_9 NS_28 0 -1.0091409063182721e-10
GC_9_29 b_9 NI_9 NS_29 0 -3.8139229193087308e-11
GC_9_30 b_9 NI_9 NS_30 0 -1.6276484380667015e-10
GC_9_31 b_9 NI_9 NS_31 0 -3.1794853349395027e-05
GC_9_32 b_9 NI_9 NS_32 0 3.5425563920605988e-06
GC_9_33 b_9 NI_9 NS_33 0 -1.3247270519106439e-08
GC_9_34 b_9 NI_9 NS_34 0 3.4619751891358576e-10
GC_9_35 b_9 NI_9 NS_35 0 2.0232774240098874e-06
GC_9_36 b_9 NI_9 NS_36 0 2.9214617545888664e-07
GC_9_37 b_9 NI_9 NS_37 0 1.7680035689554480e-06
GC_9_38 b_9 NI_9 NS_38 0 -1.7931868137553251e-06
GC_9_39 b_9 NI_9 NS_39 0 2.2222057876235132e-06
GC_9_40 b_9 NI_9 NS_40 0 -1.9596521030794661e-06
GC_9_41 b_9 NI_9 NS_41 0 1.2037877436428755e-06
GC_9_42 b_9 NI_9 NS_42 0 -1.4895731794631647e-06
GC_9_43 b_9 NI_9 NS_43 0 1.6529682573680742e-06
GC_9_44 b_9 NI_9 NS_44 0 -1.3654354008721489e-06
GC_9_45 b_9 NI_9 NS_45 0 1.7718821580779961e-06
GC_9_46 b_9 NI_9 NS_46 0 -3.2631845564199825e-06
GC_9_47 b_9 NI_9 NS_47 0 1.9918743339194487e-06
GC_9_48 b_9 NI_9 NS_48 0 -3.6176771660968299e-06
GC_9_49 b_9 NI_9 NS_49 0 7.3166907068881413e-07
GC_9_50 b_9 NI_9 NS_50 0 -3.2936831498660870e-06
GC_9_51 b_9 NI_9 NS_51 0 3.3991701054777536e-06
GC_9_52 b_9 NI_9 NS_52 0 -1.4916171613632386e-06
GC_9_53 b_9 NI_9 NS_53 0 2.6898777537254595e-07
GC_9_54 b_9 NI_9 NS_54 0 3.2027541649795704e-08
GC_9_55 b_9 NI_9 NS_55 0 1.3104225572732653e-08
GC_9_56 b_9 NI_9 NS_56 0 1.2281585014913009e-07
GC_9_57 b_9 NI_9 NS_57 0 2.5320410122473425e-11
GC_9_58 b_9 NI_9 NS_58 0 1.2029656017908744e-10
GC_9_59 b_9 NI_9 NS_59 0 3.7619720459493197e-11
GC_9_60 b_9 NI_9 NS_60 0 1.6471727625893579e-10
GC_9_61 b_9 NI_9 NS_61 0 -1.2017263142849770e-05
GC_9_62 b_9 NI_9 NS_62 0 4.3913043627566363e-07
GC_9_63 b_9 NI_9 NS_63 0 -2.5636367894331522e-08
GC_9_64 b_9 NI_9 NS_64 0 4.9336463364820488e-11
GC_9_65 b_9 NI_9 NS_65 0 -1.4663435723364255e-06
GC_9_66 b_9 NI_9 NS_66 0 -5.4508423698794246e-07
GC_9_67 b_9 NI_9 NS_67 0 -5.9487778233890154e-06
GC_9_68 b_9 NI_9 NS_68 0 2.4734516874726930e-06
GC_9_69 b_9 NI_9 NS_69 0 3.5848582715789755e-06
GC_9_70 b_9 NI_9 NS_70 0 1.3123341729813182e-05
GC_9_71 b_9 NI_9 NS_71 0 1.7633528953758116e-05
GC_9_72 b_9 NI_9 NS_72 0 1.5693913569878104e-06
GC_9_73 b_9 NI_9 NS_73 0 -1.8870703810707708e-06
GC_9_74 b_9 NI_9 NS_74 0 -1.5991965880253694e-05
GC_9_75 b_9 NI_9 NS_75 0 -4.9788796957794986e-06
GC_9_76 b_9 NI_9 NS_76 0 6.1974433531420502e-06
GC_9_77 b_9 NI_9 NS_77 0 1.1466512911358343e-05
GC_9_78 b_9 NI_9 NS_78 0 -6.6421576205495945e-07
GC_9_79 b_9 NI_9 NS_79 0 -3.8493460031581052e-07
GC_9_80 b_9 NI_9 NS_80 0 -1.0150630604222460e-05
GC_9_81 b_9 NI_9 NS_81 0 -3.8413500580221466e-06
GC_9_82 b_9 NI_9 NS_82 0 -1.7054598505634006e-06
GC_9_83 b_9 NI_9 NS_83 0 2.6624755775860252e-07
GC_9_84 b_9 NI_9 NS_84 0 9.8851510652547883e-08
GC_9_85 b_9 NI_9 NS_85 0 -1.4791259754942896e-08
GC_9_86 b_9 NI_9 NS_86 0 7.1360524537594004e-08
GC_9_87 b_9 NI_9 NS_87 0 1.4820019780720761e-10
GC_9_88 b_9 NI_9 NS_88 0 -3.5112568514766597e-11
GC_9_89 b_9 NI_9 NS_89 0 -6.6614209572715231e-11
GC_9_90 b_9 NI_9 NS_90 0 -2.6888835529788139e-10
GC_9_91 b_9 NI_9 NS_91 0 6.5825889225615018e-05
GC_9_92 b_9 NI_9 NS_92 0 -5.5593679973246308e-06
GC_9_93 b_9 NI_9 NS_93 0 3.0838594547824003e-08
GC_9_94 b_9 NI_9 NS_94 0 -1.4027678957444510e-10
GC_9_95 b_9 NI_9 NS_95 0 -2.7028172792487684e-06
GC_9_96 b_9 NI_9 NS_96 0 -1.1672689884994515e-06
GC_9_97 b_9 NI_9 NS_97 0 -4.9273591119479189e-06
GC_9_98 b_9 NI_9 NS_98 0 5.6497628020823605e-06
GC_9_99 b_9 NI_9 NS_99 0 9.6714838536575655e-06
GC_9_100 b_9 NI_9 NS_100 0 3.4362367337449998e-06
GC_9_101 b_9 NI_9 NS_101 0 -3.2948859741385112e-06
GC_9_102 b_9 NI_9 NS_102 0 -1.0812297424601746e-05
GC_9_103 b_9 NI_9 NS_103 0 -3.1204240488103253e-06
GC_9_104 b_9 NI_9 NS_104 0 -1.6758464889545716e-06
GC_9_105 b_9 NI_9 NS_105 0 -1.7488155820008276e-05
GC_9_106 b_9 NI_9 NS_106 0 -3.8613094108538048e-06
GC_9_107 b_9 NI_9 NS_107 0 -8.5222341166006217e-06
GC_9_108 b_9 NI_9 NS_108 0 1.4169312406542509e-05
GC_9_109 b_9 NI_9 NS_109 0 -7.0349681133197238e-06
GC_9_110 b_9 NI_9 NS_110 0 5.2061724342106046e-06
GC_9_111 b_9 NI_9 NS_111 0 -8.8717695143738834e-06
GC_9_112 b_9 NI_9 NS_112 0 1.0862361534895165e-05
GC_9_113 b_9 NI_9 NS_113 0 -5.7880788183911326e-07
GC_9_114 b_9 NI_9 NS_114 0 -6.3442362931488058e-08
GC_9_115 b_9 NI_9 NS_115 0 -3.7786179315891758e-08
GC_9_116 b_9 NI_9 NS_116 0 -2.6268890772987271e-07
GC_9_117 b_9 NI_9 NS_117 0 -1.5841793705445433e-10
GC_9_118 b_9 NI_9 NS_118 0 2.0132399410059364e-11
GC_9_119 b_9 NI_9 NS_119 0 6.8079745427445194e-11
GC_9_120 b_9 NI_9 NS_120 0 2.7024521902442259e-10
GC_9_121 b_9 NI_9 NS_121 0 1.2368801473949608e-04
GC_9_122 b_9 NI_9 NS_122 0 3.0410920225731186e-06
GC_9_123 b_9 NI_9 NS_123 0 -2.0461318876398280e-07
GC_9_124 b_9 NI_9 NS_124 0 -9.2714568781587583e-09
GC_9_125 b_9 NI_9 NS_125 0 5.0549170996789753e-05
GC_9_126 b_9 NI_9 NS_126 0 -1.8064784730913099e-06
GC_9_127 b_9 NI_9 NS_127 0 2.6605829830742435e-05
GC_9_128 b_9 NI_9 NS_128 0 -7.3891974108727244e-06
GC_9_129 b_9 NI_9 NS_129 0 2.3147543003967054e-05
GC_9_130 b_9 NI_9 NS_130 0 -2.6931280902044803e-04
GC_9_131 b_9 NI_9 NS_131 0 -2.9061129591903653e-04
GC_9_132 b_9 NI_9 NS_132 0 4.0339510218830524e-05
GC_9_133 b_9 NI_9 NS_133 0 -5.3941966477438374e-05
GC_9_134 b_9 NI_9 NS_134 0 2.2027267117522668e-04
GC_9_135 b_9 NI_9 NS_135 0 1.6852043053352343e-04
GC_9_136 b_9 NI_9 NS_136 0 -1.0671238666487607e-04
GC_9_137 b_9 NI_9 NS_137 0 -1.8010365244191693e-04
GC_9_138 b_9 NI_9 NS_138 0 6.0291836990389651e-05
GC_9_139 b_9 NI_9 NS_139 0 -4.9801217461142626e-05
GC_9_140 b_9 NI_9 NS_140 0 1.1984178044380441e-04
GC_9_141 b_9 NI_9 NS_141 0 1.3935796692703779e-04
GC_9_142 b_9 NI_9 NS_142 0 7.0033210780019359e-05
GC_9_143 b_9 NI_9 NS_143 0 3.0857897980873246e-08
GC_9_144 b_9 NI_9 NS_144 0 4.2557784859203764e-06
GC_9_145 b_9 NI_9 NS_145 0 -1.9662424219448834e-06
GC_9_146 b_9 NI_9 NS_146 0 8.4457627824057878e-08
GC_9_147 b_9 NI_9 NS_147 0 6.1361187741076143e-10
GC_9_148 b_9 NI_9 NS_148 0 -6.3988312600160801e-10
GC_9_149 b_9 NI_9 NS_149 0 -1.4671369425863314e-10
GC_9_150 b_9 NI_9 NS_150 0 -1.2237817799299295e-09
GC_9_151 b_9 NI_9 NS_151 0 5.4736180129007222e-05
GC_9_152 b_9 NI_9 NS_152 0 9.2111704618688523e-05
GC_9_153 b_9 NI_9 NS_153 0 2.8700366870423736e-07
GC_9_154 b_9 NI_9 NS_154 0 8.4904563937908963e-09
GC_9_155 b_9 NI_9 NS_155 0 -4.0121829880024276e-05
GC_9_156 b_9 NI_9 NS_156 0 -8.6000256292131930e-05
GC_9_157 b_9 NI_9 NS_157 0 -2.2672035750797583e-04
GC_9_158 b_9 NI_9 NS_158 0 9.6541665037368785e-05
GC_9_159 b_9 NI_9 NS_159 0 2.8121763751696565e-04
GC_9_160 b_9 NI_9 NS_160 0 1.5448808075185785e-04
GC_9_161 b_9 NI_9 NS_161 0 -3.0713745864391210e-04
GC_9_162 b_9 NI_9 NS_162 0 -2.0845289291345525e-04
GC_9_163 b_9 NI_9 NS_163 0 1.8397833523902451e-04
GC_9_164 b_9 NI_9 NS_164 0 3.9105516979648976e-04
GC_9_165 b_9 NI_9 NS_165 0 -9.4946753031781877e-05
GC_9_166 b_9 NI_9 NS_166 0 -1.5522232931490155e-04
GC_9_167 b_9 NI_9 NS_167 0 2.3740762382043097e-04
GC_9_168 b_9 NI_9 NS_168 0 2.1642596031168430e-04
GC_9_169 b_9 NI_9 NS_169 0 -5.9516953681097131e-05
GC_9_170 b_9 NI_9 NS_170 0 -2.0711938507905157e-04
GC_9_171 b_9 NI_9 NS_171 0 -2.1936527619352149e-06
GC_9_172 b_9 NI_9 NS_172 0 2.1430579906381552e-04
GC_9_173 b_9 NI_9 NS_173 0 -2.2383120276810301e-06
GC_9_174 b_9 NI_9 NS_174 0 6.4588990630521810e-08
GC_9_175 b_9 NI_9 NS_175 0 -4.6477925149707233e-07
GC_9_176 b_9 NI_9 NS_176 0 -4.5310063349281602e-07
GC_9_177 b_9 NI_9 NS_177 0 -7.2775456933964774e-10
GC_9_178 b_9 NI_9 NS_178 0 5.1682448181456334e-10
GC_9_179 b_9 NI_9 NS_179 0 1.4748960743037531e-10
GC_9_180 b_9 NI_9 NS_180 0 1.2209581998831445e-09
GC_9_181 b_9 NI_9 NS_181 0 2.2658564431924091e-03
GC_9_182 b_9 NI_9 NS_182 0 -7.3259609460769241e-04
GC_9_183 b_9 NI_9 NS_183 0 -1.8147798015694404e-06
GC_9_184 b_9 NI_9 NS_184 0 -1.2100069733947770e-07
GC_9_185 b_9 NI_9 NS_185 0 3.5972857007827557e-04
GC_9_186 b_9 NI_9 NS_186 0 -3.7512259088591326e-04
GC_9_187 b_9 NI_9 NS_187 0 -1.2776319317895878e-03
GC_9_188 b_9 NI_9 NS_188 0 3.4322714298305843e-04
GC_9_189 b_9 NI_9 NS_189 0 7.1259047109704357e-04
GC_9_190 b_9 NI_9 NS_190 0 -8.2806986803091783e-04
GC_9_191 b_9 NI_9 NS_191 0 -1.5010235012802542e-04
GC_9_192 b_9 NI_9 NS_192 0 1.3910986754601059e-03
GC_9_193 b_9 NI_9 NS_193 0 -1.3011090184595249e-03
GC_9_194 b_9 NI_9 NS_194 0 -7.6481278533339556e-04
GC_9_195 b_9 NI_9 NS_195 0 6.8664558444414320e-04
GC_9_196 b_9 NI_9 NS_196 0 -2.8679358179347108e-05
GC_9_197 b_9 NI_9 NS_197 0 -1.3691887193630219e-04
GC_9_198 b_9 NI_9 NS_198 0 1.4681555605746256e-03
GC_9_199 b_9 NI_9 NS_199 0 -7.1830203020495939e-04
GC_9_200 b_9 NI_9 NS_200 0 -5.4309744743232067e-04
GC_9_201 b_9 NI_9 NS_201 0 6.5104338320360255e-04
GC_9_202 b_9 NI_9 NS_202 0 1.9305495729484822e-04
GC_9_203 b_9 NI_9 NS_203 0 -3.0110341711249124e-06
GC_9_204 b_9 NI_9 NS_204 0 2.6005608542399902e-05
GC_9_205 b_9 NI_9 NS_205 0 -9.9167466130714327e-06
GC_9_206 b_9 NI_9 NS_206 0 -1.4215860318450902e-06
GC_9_207 b_9 NI_9 NS_207 0 7.0600818737195675e-09
GC_9_208 b_9 NI_9 NS_208 0 -1.0479797327162022e-08
GC_9_209 b_9 NI_9 NS_209 0 -6.2224924868716404e-10
GC_9_210 b_9 NI_9 NS_210 0 -2.1194002561654577e-09
GC_9_211 b_9 NI_9 NS_211 0 9.8222022760814935e-04
GC_9_212 b_9 NI_9 NS_212 0 -3.4568950576806918e-04
GC_9_213 b_9 NI_9 NS_213 0 2.1363493972984145e-06
GC_9_214 b_9 NI_9 NS_214 0 8.2059475521024335e-08
GC_9_215 b_9 NI_9 NS_215 0 1.1718806563855454e-05
GC_9_216 b_9 NI_9 NS_216 0 8.7362349435559584e-05
GC_9_217 b_9 NI_9 NS_217 0 3.1568319997713932e-04
GC_9_218 b_9 NI_9 NS_218 0 -1.1545911643438253e-04
GC_9_219 b_9 NI_9 NS_219 0 -5.1920857029678349e-04
GC_9_220 b_9 NI_9 NS_220 0 -2.4291004803810864e-04
GC_9_221 b_9 NI_9 NS_221 0 3.2786467375423820e-04
GC_9_222 b_9 NI_9 NS_222 0 3.8890649503389068e-04
GC_9_223 b_9 NI_9 NS_223 0 -3.2493967352261875e-04
GC_9_224 b_9 NI_9 NS_224 0 -5.5996074854649299e-04
GC_9_225 b_9 NI_9 NS_225 0 7.3917219149957855e-05
GC_9_226 b_9 NI_9 NS_226 0 3.8468623706292915e-04
GC_9_227 b_9 NI_9 NS_227 0 -3.5604784217616866e-04
GC_9_228 b_9 NI_9 NS_228 0 -2.6841050401765168e-04
GC_9_229 b_9 NI_9 NS_229 0 5.3022531504096291e-06
GC_9_230 b_9 NI_9 NS_230 0 4.0801997125193426e-04
GC_9_231 b_9 NI_9 NS_231 0 -9.5157983113976726e-05
GC_9_232 b_9 NI_9 NS_232 0 -3.4082249767297803e-04
GC_9_233 b_9 NI_9 NS_233 0 -1.4814590733117278e-05
GC_9_234 b_9 NI_9 NS_234 0 -8.4885222856912979e-06
GC_9_235 b_9 NI_9 NS_235 0 2.7376409896317390e-06
GC_9_236 b_9 NI_9 NS_236 0 -6.6723216765000272e-06
GC_9_237 b_9 NI_9 NS_237 0 -7.7197736137596098e-09
GC_9_238 b_9 NI_9 NS_238 0 4.8068825892666659e-09
GC_9_239 b_9 NI_9 NS_239 0 1.1496283780445532e-09
GC_9_240 b_9 NI_9 NS_240 0 2.7805514223049851e-09
GC_9_241 b_9 NI_9 NS_241 0 1.2659773860458268e-01
GC_9_242 b_9 NI_9 NS_242 0 -9.9682294588668424e-03
GC_9_243 b_9 NI_9 NS_243 0 -2.0418473141989946e-05
GC_9_244 b_9 NI_9 NS_244 0 -3.8273616432283193e-06
GC_9_245 b_9 NI_9 NS_245 0 -8.0908251645516616e-03
GC_9_246 b_9 NI_9 NS_246 0 6.4296780914414355e-04
GC_9_247 b_9 NI_9 NS_247 0 -1.9909397529217568e-03
GC_9_248 b_9 NI_9 NS_248 0 6.7353868360028852e-05
GC_9_249 b_9 NI_9 NS_249 0 -1.2598721021315521e-02
GC_9_250 b_9 NI_9 NS_250 0 8.2477756362525981e-03
GC_9_251 b_9 NI_9 NS_251 0 -1.0271315651357403e-02
GC_9_252 b_9 NI_9 NS_252 0 -6.2357810582910466e-04
GC_9_253 b_9 NI_9 NS_253 0 -3.5565687463906342e-03
GC_9_254 b_9 NI_9 NS_254 0 1.6966131545998242e-02
GC_9_255 b_9 NI_9 NS_255 0 -7.7825975278901323e-03
GC_9_256 b_9 NI_9 NS_256 0 1.3370077146006586e-02
GC_9_257 b_9 NI_9 NS_257 0 -3.9902969105566352e-03
GC_9_258 b_9 NI_9 NS_258 0 6.9628750442002115e-03
GC_9_259 b_9 NI_9 NS_259 0 -2.7633689428856129e-03
GC_9_260 b_9 NI_9 NS_260 0 1.2313501087860952e-02
GC_9_261 b_9 NI_9 NS_261 0 -2.2964016853188465e-02
GC_9_262 b_9 NI_9 NS_262 0 5.9629979338305114e-03
GC_9_263 b_9 NI_9 NS_263 0 -8.6294521792626444e-04
GC_9_264 b_9 NI_9 NS_264 0 8.0344078006493083e-04
GC_9_265 b_9 NI_9 NS_265 0 -5.1358588480691783e-04
GC_9_266 b_9 NI_9 NS_266 0 -4.3937294384617531e-04
GC_9_267 b_9 NI_9 NS_267 0 -6.4174258942452756e-08
GC_9_268 b_9 NI_9 NS_268 0 -1.9155152348216248e-07
GC_9_269 b_9 NI_9 NS_269 0 -3.0939577975646501e-09
GC_9_270 b_9 NI_9 NS_270 0 5.6381487193437262e-09
GC_9_271 b_9 NI_9 NS_271 0 -7.5348993576201326e-02
GC_9_272 b_9 NI_9 NS_272 0 2.4900053766048813e-02
GC_9_273 b_9 NI_9 NS_273 0 1.9200088562089617e-05
GC_9_274 b_9 NI_9 NS_274 0 5.3863132218958305e-06
GC_9_275 b_9 NI_9 NS_275 0 1.8353490408803595e-02
GC_9_276 b_9 NI_9 NS_276 0 2.7965421093143230e-02
GC_9_277 b_9 NI_9 NS_277 0 -1.9176289837020410e-02
GC_9_278 b_9 NI_9 NS_278 0 8.3761603397304839e-03
GC_9_279 b_9 NI_9 NS_279 0 -5.5264526429188963e-03
GC_9_280 b_9 NI_9 NS_280 0 -2.3054185939361101e-02
GC_9_281 b_9 NI_9 NS_281 0 2.6687335929769802e-02
GC_9_282 b_9 NI_9 NS_282 0 -1.4576077176349195e-02
GC_9_283 b_9 NI_9 NS_283 0 3.4517359662758693e-02
GC_9_284 b_9 NI_9 NS_284 0 4.8628291368667661e-03
GC_9_285 b_9 NI_9 NS_285 0 9.6719352021881217e-03
GC_9_286 b_9 NI_9 NS_286 0 1.3692458946476064e-02
GC_9_287 b_9 NI_9 NS_287 0 -1.2370858371226754e-02
GC_9_288 b_9 NI_9 NS_288 0 1.1007980187933194e-02
GC_9_289 b_9 NI_9 NS_289 0 -1.1774514058568844e-02
GC_9_290 b_9 NI_9 NS_290 0 -1.2014097021479530e-02
GC_9_291 b_9 NI_9 NS_291 0 1.9793996337900681e-02
GC_9_292 b_9 NI_9 NS_292 0 -2.6023911237968479e-02
GC_9_293 b_9 NI_9 NS_293 0 9.6721498585233096e-04
GC_9_294 b_9 NI_9 NS_294 0 -1.0822069829665283e-03
GC_9_295 b_9 NI_9 NS_295 0 6.3094621163340694e-04
GC_9_296 b_9 NI_9 NS_296 0 3.4914437967213170e-04
GC_9_297 b_9 NI_9 NS_297 0 9.7107516730023475e-08
GC_9_298 b_9 NI_9 NS_298 0 4.1868699176562550e-07
GC_9_299 b_9 NI_9 NS_299 0 -1.0314520371142416e-08
GC_9_300 b_9 NI_9 NS_300 0 -1.9789263145178136e-08
GC_9_301 b_9 NI_9 NS_301 0 -5.4915841993808875e-04
GC_9_302 b_9 NI_9 NS_302 0 -2.9018837039708296e-03
GC_9_303 b_9 NI_9 NS_303 0 -6.1488955598811034e-06
GC_9_304 b_9 NI_9 NS_304 0 -3.8642052853340799e-07
GC_9_305 b_9 NI_9 NS_305 0 2.6865516591988749e-03
GC_9_306 b_9 NI_9 NS_306 0 -1.9871372582523921e-03
GC_9_307 b_9 NI_9 NS_307 0 -6.1989513832137275e-03
GC_9_308 b_9 NI_9 NS_308 0 1.7530828200673320e-03
GC_9_309 b_9 NI_9 NS_309 0 4.7648850850489236e-03
GC_9_310 b_9 NI_9 NS_310 0 -5.5284540635730864e-03
GC_9_311 b_9 NI_9 NS_311 0 -2.4815306869972059e-04
GC_9_312 b_9 NI_9 NS_312 0 7.2493849593844575e-03
GC_9_313 b_9 NI_9 NS_313 0 -6.3156107463805443e-03
GC_9_314 b_9 NI_9 NS_314 0 -5.0550429424194524e-03
GC_9_315 b_9 NI_9 NS_315 0 4.5025677458851313e-03
GC_9_316 b_9 NI_9 NS_316 0 -1.7116128853888381e-03
GC_9_317 b_9 NI_9 NS_317 0 -5.9125367198868412e-04
GC_9_318 b_9 NI_9 NS_318 0 6.9477907108374598e-03
GC_9_319 b_9 NI_9 NS_319 0 -3.4362430168487067e-03
GC_9_320 b_9 NI_9 NS_320 0 -3.6821810458767435e-03
GC_9_321 b_9 NI_9 NS_321 0 5.9242608986460410e-03
GC_9_322 b_9 NI_9 NS_322 0 3.9702052908980353e-04
GC_9_323 b_9 NI_9 NS_323 0 6.3746601294586234e-05
GC_9_324 b_9 NI_9 NS_324 0 8.4799176107691170e-06
GC_9_325 b_9 NI_9 NS_325 0 1.5085273241362107e-05
GC_9_326 b_9 NI_9 NS_326 0 3.9926660865903014e-05
GC_9_327 b_9 NI_9 NS_327 0 7.1120485370220176e-09
GC_9_328 b_9 NI_9 NS_328 0 -2.9352136411090104e-08
GC_9_329 b_9 NI_9 NS_329 0 -1.8854126658506922e-09
GC_9_330 b_9 NI_9 NS_330 0 -5.6020611491903549e-10
GC_9_331 b_9 NI_9 NS_331 0 1.3561032718190709e-03
GC_9_332 b_9 NI_9 NS_332 0 -1.2038975406755130e-03
GC_9_333 b_9 NI_9 NS_333 0 3.7358057183382851e-06
GC_9_334 b_9 NI_9 NS_334 0 2.8901996539223217e-07
GC_9_335 b_9 NI_9 NS_335 0 1.2295932909834015e-04
GC_9_336 b_9 NI_9 NS_336 0 8.9417142188338687e-04
GC_9_337 b_9 NI_9 NS_337 0 1.8425106140205765e-03
GC_9_338 b_9 NI_9 NS_338 0 -8.6745792168850218e-04
GC_9_339 b_9 NI_9 NS_339 0 -2.9666020918209190e-03
GC_9_340 b_9 NI_9 NS_340 0 -1.6486044684690816e-03
GC_9_341 b_9 NI_9 NS_341 0 2.2194915709220714e-03
GC_9_342 b_9 NI_9 NS_342 0 2.6689308128691100e-03
GC_9_343 b_9 NI_9 NS_343 0 -1.4401415521705441e-03
GC_9_344 b_9 NI_9 NS_344 0 -2.9129099036704258e-03
GC_9_345 b_9 NI_9 NS_345 0 1.0698831151070159e-03
GC_9_346 b_9 NI_9 NS_346 0 2.2566994843893399e-03
GC_9_347 b_9 NI_9 NS_347 0 -1.6275472028653586e-03
GC_9_348 b_9 NI_9 NS_348 0 -2.1363613895425330e-03
GC_9_349 b_9 NI_9 NS_349 0 4.2046148382028176e-04
GC_9_350 b_9 NI_9 NS_350 0 2.0118573278588596e-03
GC_9_351 b_9 NI_9 NS_351 0 2.1506806916417667e-04
GC_9_352 b_9 NI_9 NS_352 0 -2.1102648323654927e-03
GC_9_353 b_9 NI_9 NS_353 0 -4.3297592914652035e-06
GC_9_354 b_9 NI_9 NS_354 0 4.3533743092581193e-06
GC_9_355 b_9 NI_9 NS_355 0 -7.8987902033922279e-07
GC_9_356 b_9 NI_9 NS_356 0 -3.5253886213821896e-06
GC_9_357 b_9 NI_9 NS_357 0 -7.5480237649974902e-09
GC_9_358 b_9 NI_9 NS_358 0 2.2567511706671412e-08
GC_9_359 b_9 NI_9 NS_359 0 2.3359259828195180e-09
GC_9_360 b_9 NI_9 NS_360 0 1.5101887849105698e-09
GD_9_1 b_9 NI_9 NA_1 0 -1.7050923126667179e-06
GD_9_2 b_9 NI_9 NA_2 0 7.7104334434857245e-06
GD_9_3 b_9 NI_9 NA_3 0 -1.1549169558395701e-06
GD_9_4 b_9 NI_9 NA_4 0 -9.0627079894041708e-06
GD_9_5 b_9 NI_9 NA_5 0 1.7125087270432532e-04
GD_9_6 b_9 NI_9 NA_6 0 -6.2836551426455922e-05
GD_9_7 b_9 NI_9 NA_7 0 2.3299342723291385e-03
GD_9_8 b_9 NI_9 NA_8 0 -4.6762438048733507e-05
GD_9_9 b_9 NI_9 NA_9 0 -4.0270205362664090e-02
GD_9_10 b_9 NI_9 NA_10 0 -9.9682817487122821e-03
GD_9_11 b_9 NI_9 NA_11 0 1.6053724364173561e-02
GD_9_12 b_9 NI_9 NA_12 0 -9.1338169335060580e-05
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 -3.1793575120580654e-05
GC_10_2 b_10 NI_10 NS_2 0 3.5424378043569224e-06
GC_10_3 b_10 NI_10 NS_3 0 -1.3247016182661042e-08
GC_10_4 b_10 NI_10 NS_4 0 3.4619120895328476e-10
GC_10_5 b_10 NI_10 NS_5 0 2.0231536813855486e-06
GC_10_6 b_10 NI_10 NS_6 0 2.9210670963746515e-07
GC_10_7 b_10 NI_10 NS_7 0 1.7678881579961950e-06
GC_10_8 b_10 NI_10 NS_8 0 -1.7931418331852966e-06
GC_10_9 b_10 NI_10 NS_9 0 2.2220721400375270e-06
GC_10_10 b_10 NI_10 NS_10 0 -1.9594593712809157e-06
GC_10_11 b_10 NI_10 NS_11 0 1.2037180123768188e-06
GC_10_12 b_10 NI_10 NS_12 0 -1.4894340290034103e-06
GC_10_13 b_10 NI_10 NS_13 0 1.6529552467767675e-06
GC_10_14 b_10 NI_10 NS_14 0 -1.3652565625220923e-06
GC_10_15 b_10 NI_10 NS_15 0 1.7719402119347430e-06
GC_10_16 b_10 NI_10 NS_16 0 -3.2630854029293619e-06
GC_10_17 b_10 NI_10 NS_17 0 1.9918527508190866e-06
GC_10_18 b_10 NI_10 NS_18 0 -3.6175784220806373e-06
GC_10_19 b_10 NI_10 NS_19 0 7.3162840412348144e-07
GC_10_20 b_10 NI_10 NS_20 0 -3.2936019099166414e-06
GC_10_21 b_10 NI_10 NS_21 0 3.3990069366955819e-06
GC_10_22 b_10 NI_10 NS_22 0 -1.4915452347026693e-06
GC_10_23 b_10 NI_10 NS_23 0 2.6897946638989878e-07
GC_10_24 b_10 NI_10 NS_24 0 3.2033133029752071e-08
GC_10_25 b_10 NI_10 NS_25 0 1.3100790320465231e-08
GC_10_26 b_10 NI_10 NS_26 0 1.2281188663500836e-07
GC_10_27 b_10 NI_10 NS_27 0 2.5320005813120942e-11
GC_10_28 b_10 NI_10 NS_28 0 1.2029519948515463e-10
GC_10_29 b_10 NI_10 NS_29 0 3.7619861964098403e-11
GC_10_30 b_10 NI_10 NS_30 0 1.6471739537554982e-10
GC_10_31 b_10 NI_10 NS_31 0 1.8182627614184791e-05
GC_10_32 b_10 NI_10 NS_32 0 -2.5901341950131765e-06
GC_10_33 b_10 NI_10 NS_33 0 1.0334195313759740e-08
GC_10_34 b_10 NI_10 NS_34 0 -2.6700214895846905e-10
GC_10_35 b_10 NI_10 NS_35 0 -1.2561972240480255e-06
GC_10_36 b_10 NI_10 NS_36 0 -1.1110382747613928e-06
GC_10_37 b_10 NI_10 NS_37 0 -2.4938859600926695e-06
GC_10_38 b_10 NI_10 NS_38 0 5.3481703630228151e-07
GC_10_39 b_10 NI_10 NS_39 0 -1.2776559239347972e-06
GC_10_40 b_10 NI_10 NS_40 0 2.6875757086234610e-06
GC_10_41 b_10 NI_10 NS_41 0 1.8066986446091088e-06
GC_10_42 b_10 NI_10 NS_42 0 7.9089573360123267e-07
GC_10_43 b_10 NI_10 NS_43 0 -2.7692144886105533e-06
GC_10_44 b_10 NI_10 NS_44 0 -1.3482201235263328e-06
GC_10_45 b_10 NI_10 NS_45 0 -2.1726550298531809e-06
GC_10_46 b_10 NI_10 NS_46 0 3.4750576385032522e-06
GC_10_47 b_10 NI_10 NS_47 0 1.2557145191618845e-06
GC_10_48 b_10 NI_10 NS_48 0 2.3797764732273320e-06
GC_10_49 b_10 NI_10 NS_49 0 -9.2223793712865595e-07
GC_10_50 b_10 NI_10 NS_50 0 -3.7752720443769691e-07
GC_10_51 b_10 NI_10 NS_51 0 -3.3379677302476039e-06
GC_10_52 b_10 NI_10 NS_52 0 6.3278216094284929e-07
GC_10_53 b_10 NI_10 NS_53 0 -1.4338076363007125e-07
GC_10_54 b_10 NI_10 NS_54 0 -7.6374244603797899e-08
GC_10_55 b_10 NI_10 NS_55 0 2.3067696263226196e-08
GC_10_56 b_10 NI_10 NS_56 0 -5.2057516728874935e-08
GC_10_57 b_10 NI_10 NS_57 0 -1.8003842956577788e-11
GC_10_58 b_10 NI_10 NS_58 0 -1.0118382916136453e-10
GC_10_59 b_10 NI_10 NS_59 0 -3.8103999483278552e-11
GC_10_60 b_10 NI_10 NS_60 0 -1.6272437015848249e-10
GC_10_61 b_10 NI_10 NS_61 0 6.6256689617543731e-05
GC_10_62 b_10 NI_10 NS_62 0 -5.6124249325245599e-06
GC_10_63 b_10 NI_10 NS_63 0 3.0931084320127369e-08
GC_10_64 b_10 NI_10 NS_64 0 -1.4166196453141024e-10
GC_10_65 b_10 NI_10 NS_65 0 -2.7183688788801816e-06
GC_10_66 b_10 NI_10 NS_66 0 -1.1809895673134519e-06
GC_10_67 b_10 NI_10 NS_67 0 -4.9372985382801448e-06
GC_10_68 b_10 NI_10 NS_68 0 5.6220228218073454e-06
GC_10_69 b_10 NI_10 NS_69 0 9.6526171982338680e-06
GC_10_70 b_10 NI_10 NS_70 0 3.4537884098533883e-06
GC_10_71 b_10 NI_10 NS_71 0 -3.3260936580128930e-06
GC_10_72 b_10 NI_10 NS_72 0 -1.0830890682061186e-05
GC_10_73 b_10 NI_10 NS_73 0 -3.1844527093074772e-06
GC_10_74 b_10 NI_10 NS_74 0 -1.6471617803173969e-06
GC_10_75 b_10 NI_10 NS_75 0 -1.7516677792472084e-05
GC_10_76 b_10 NI_10 NS_76 0 -3.8364721951655624e-06
GC_10_77 b_10 NI_10 NS_77 0 -8.5578986087408962e-06
GC_10_78 b_10 NI_10 NS_78 0 1.4206940937329282e-05
GC_10_79 b_10 NI_10 NS_79 0 -7.0646540710165132e-06
GC_10_80 b_10 NI_10 NS_80 0 5.2325189170539283e-06
GC_10_81 b_10 NI_10 NS_81 0 -8.9556829121472553e-06
GC_10_82 b_10 NI_10 NS_82 0 1.0881312971276958e-05
GC_10_83 b_10 NI_10 NS_83 0 -5.8293515448929081e-07
GC_10_84 b_10 NI_10 NS_84 0 -6.0298377478652792e-08
GC_10_85 b_10 NI_10 NS_85 0 -3.9873479783716724e-08
GC_10_86 b_10 NI_10 NS_86 0 -2.6482625466718598e-07
GC_10_87 b_10 NI_10 NS_87 0 -1.5857053539954890e-10
GC_10_88 b_10 NI_10 NS_88 0 1.9903998835457215e-11
GC_10_89 b_10 NI_10 NS_89 0 6.8097740535777061e-11
GC_10_90 b_10 NI_10 NS_90 0 2.7026123862286742e-10
GC_10_91 b_10 NI_10 NS_91 0 -1.2017600754582061e-05
GC_10_92 b_10 NI_10 NS_92 0 4.3917146397351328e-07
GC_10_93 b_10 NI_10 NS_93 0 -2.5636463744052287e-08
GC_10_94 b_10 NI_10 NS_94 0 4.9337643492046543e-11
GC_10_95 b_10 NI_10 NS_95 0 -1.4663206416779239e-06
GC_10_96 b_10 NI_10 NS_96 0 -5.4509489287444058e-07
GC_10_97 b_10 NI_10 NS_97 0 -5.9487633472919509e-06
GC_10_98 b_10 NI_10 NS_98 0 2.4734449764692922e-06
GC_10_99 b_10 NI_10 NS_99 0 3.5848772641100311e-06
GC_10_100 b_10 NI_10 NS_100 0 1.3123316712635292e-05
GC_10_101 b_10 NI_10 NS_101 0 1.7633552067163037e-05
GC_10_102 b_10 NI_10 NS_102 0 1.5693729928652510e-06
GC_10_103 b_10 NI_10 NS_103 0 -1.8870595810546831e-06
GC_10_104 b_10 NI_10 NS_104 0 -1.5992004150509057e-05
GC_10_105 b_10 NI_10 NS_105 0 -4.9788854600051602e-06
GC_10_106 b_10 NI_10 NS_106 0 6.1974139912781451e-06
GC_10_107 b_10 NI_10 NS_107 0 1.1466516694150449e-05
GC_10_108 b_10 NI_10 NS_108 0 -6.6423532744954216e-07
GC_10_109 b_10 NI_10 NS_109 0 -3.8491893212015234e-07
GC_10_110 b_10 NI_10 NS_110 0 -1.0150638891604437e-05
GC_10_111 b_10 NI_10 NS_111 0 -3.8412900477125309e-06
GC_10_112 b_10 NI_10 NS_112 0 -1.7054669522090318e-06
GC_10_113 b_10 NI_10 NS_113 0 2.6625117038399535e-07
GC_10_114 b_10 NI_10 NS_114 0 9.8849096428814987e-08
GC_10_115 b_10 NI_10 NS_115 0 -1.4789722842684261e-08
GC_10_116 b_10 NI_10 NS_116 0 7.1362494094801019e-08
GC_10_117 b_10 NI_10 NS_117 0 1.4820036648792503e-10
GC_10_118 b_10 NI_10 NS_118 0 -3.5112405867222798e-11
GC_10_119 b_10 NI_10 NS_119 0 -6.6614192287498829e-11
GC_10_120 b_10 NI_10 NS_120 0 -2.6888833528515993e-10
GC_10_121 b_10 NI_10 NS_121 0 5.4752131756256967e-05
GC_10_122 b_10 NI_10 NS_122 0 9.2110312088026982e-05
GC_10_123 b_10 NI_10 NS_123 0 2.8700555372227213e-07
GC_10_124 b_10 NI_10 NS_124 0 8.4904230633084132e-09
GC_10_125 b_10 NI_10 NS_125 0 -4.0122562585976387e-05
GC_10_126 b_10 NI_10 NS_126 0 -8.5999951195783530e-05
GC_10_127 b_10 NI_10 NS_127 0 -2.2672065736546956e-04
GC_10_128 b_10 NI_10 NS_128 0 9.6541365297674294e-05
GC_10_129 b_10 NI_10 NS_129 0 2.8121580880630234e-04
GC_10_130 b_10 NI_10 NS_130 0 1.5448853467131304e-04
GC_10_131 b_10 NI_10 NS_131 0 -3.0713872454817074e-04
GC_10_132 b_10 NI_10 NS_132 0 -2.0845193420367182e-04
GC_10_133 b_10 NI_10 NS_133 0 1.8397692698793509e-04
GC_10_134 b_10 NI_10 NS_134 0 3.9105606697686696e-04
GC_10_135 b_10 NI_10 NS_135 0 -9.4947556848771762e-05
GC_10_136 b_10 NI_10 NS_136 0 -1.5521934250054722e-04
GC_10_137 b_10 NI_10 NS_137 0 2.3740746001518276e-04
GC_10_138 b_10 NI_10 NS_138 0 2.1642751075658291e-04
GC_10_139 b_10 NI_10 NS_139 0 -5.9517835685953021e-05
GC_10_140 b_10 NI_10 NS_140 0 -2.0711790913539890e-04
GC_10_141 b_10 NI_10 NS_141 0 -2.1951743490265657e-06
GC_10_142 b_10 NI_10 NS_142 0 2.1430694636684892e-04
GC_10_143 b_10 NI_10 NS_143 0 -2.2384337647571552e-06
GC_10_144 b_10 NI_10 NS_144 0 6.4681666266890886e-08
GC_10_145 b_10 NI_10 NS_145 0 -4.6483124857781362e-07
GC_10_146 b_10 NI_10 NS_146 0 -4.5316248144194348e-07
GC_10_147 b_10 NI_10 NS_147 0 -7.2775856801077230e-10
GC_10_148 b_10 NI_10 NS_148 0 5.1681931366362099e-10
GC_10_149 b_10 NI_10 NS_149 0 1.4748978102905751e-10
GC_10_150 b_10 NI_10 NS_150 0 1.2209582720388090e-09
GC_10_151 b_10 NI_10 NS_151 0 1.3866248409621836e-04
GC_10_152 b_10 NI_10 NS_152 0 1.3581155374805223e-06
GC_10_153 b_10 NI_10 NS_153 0 -2.0145405486085696e-07
GC_10_154 b_10 NI_10 NS_154 0 -9.3088468483846660e-09
GC_10_155 b_10 NI_10 NS_155 0 4.9967109856868900e-05
GC_10_156 b_10 NI_10 NS_156 0 -1.9693981016066081e-06
GC_10_157 b_10 NI_10 NS_157 0 2.5673320102397615e-05
GC_10_158 b_10 NI_10 NS_158 0 -7.4987201559846379e-06
GC_10_159 b_10 NI_10 NS_159 0 2.2259868070879740e-05
GC_10_160 b_10 NI_10 NS_160 0 -2.6884224242147974e-04
GC_10_161 b_10 NI_10 NS_161 0 -2.9200887591968158e-04
GC_10_162 b_10 NI_10 NS_162 0 4.0827744081241385e-05
GC_10_163 b_10 NI_10 NS_163 0 -5.4990126274054561e-05
GC_10_164 b_10 NI_10 NS_164 0 2.2142040575059247e-04
GC_10_165 b_10 NI_10 NS_165 0 1.6790480777281489e-04
GC_10_166 b_10 NI_10 NS_166 0 -1.0524497912790598e-04
GC_10_167 b_10 NI_10 NS_167 0 -1.8089903548837942e-04
GC_10_168 b_10 NI_10 NS_168 0 6.1698514030793155e-05
GC_10_169 b_10 NI_10 NS_169 0 -5.0485824938456516e-05
GC_10_170 b_10 NI_10 NS_170 0 1.2080567320384622e-04
GC_10_171 b_10 NI_10 NS_171 0 1.3699040315422108e-04
GC_10_172 b_10 NI_10 NS_172 0 7.0683380697144531e-05
GC_10_173 b_10 NI_10 NS_173 0 -1.0789883801949112e-07
GC_10_174 b_10 NI_10 NS_174 0 4.3458258228282219e-06
GC_10_175 b_10 NI_10 NS_175 0 -2.0228965017355681e-06
GC_10_176 b_10 NI_10 NS_176 0 1.7345012944490243e-08
GC_10_177 b_10 NI_10 NS_177 0 6.0908630078237221e-10
GC_10_178 b_10 NI_10 NS_178 0 -6.4494214291664770e-10
GC_10_179 b_10 NI_10 NS_179 0 -1.4660392980888061e-10
GC_10_180 b_10 NI_10 NS_180 0 -1.2238406444678684e-09
GC_10_181 b_10 NI_10 NS_181 0 9.8191781229332734e-04
GC_10_182 b_10 NI_10 NS_182 0 -3.4563458490509652e-04
GC_10_183 b_10 NI_10 NS_183 0 2.1362772100010917e-06
GC_10_184 b_10 NI_10 NS_184 0 8.2059868472045922e-08
GC_10_185 b_10 NI_10 NS_185 0 1.1628698311457659e-05
GC_10_186 b_10 NI_10 NS_186 0 8.7325783699856456e-05
GC_10_187 b_10 NI_10 NS_187 0 3.1565263696006052e-04
GC_10_188 b_10 NI_10 NS_188 0 -1.1551278727261860e-04
GC_10_189 b_10 NI_10 NS_189 0 -5.1916689092184600e-04
GC_10_190 b_10 NI_10 NS_190 0 -2.4271731305418399e-04
GC_10_191 b_10 NI_10 NS_191 0 3.2788840250700264e-04
GC_10_192 b_10 NI_10 NS_192 0 3.8892152388608710e-04
GC_10_193 b_10 NI_10 NS_193 0 -3.2494903009044576e-04
GC_10_194 b_10 NI_10 NS_194 0 -5.5986616154216117e-04
GC_10_195 b_10 NI_10 NS_195 0 7.3998214808362197e-05
GC_10_196 b_10 NI_10 NS_196 0 3.8462936667805402e-04
GC_10_197 b_10 NI_10 NS_197 0 -3.5599624180046970e-04
GC_10_198 b_10 NI_10 NS_198 0 -2.6838291423287816e-04
GC_10_199 b_10 NI_10 NS_199 0 5.3831799127637378e-06
GC_10_200 b_10 NI_10 NS_200 0 4.0799864439013480e-04
GC_10_201 b_10 NI_10 NS_201 0 -9.5065874195527665e-05
GC_10_202 b_10 NI_10 NS_202 0 -3.4082220217833295e-04
GC_10_203 b_10 NI_10 NS_203 0 -1.4810614307717058e-05
GC_10_204 b_10 NI_10 NS_204 0 -8.4933831161579369e-06
GC_10_205 b_10 NI_10 NS_205 0 2.7403456071686013e-06
GC_10_206 b_10 NI_10 NS_206 0 -6.6706399905351272e-06
GC_10_207 b_10 NI_10 NS_207 0 -7.7196779521421328e-09
GC_10_208 b_10 NI_10 NS_208 0 4.8069828023510631e-09
GC_10_209 b_10 NI_10 NS_209 0 1.1496159317838916e-09
GC_10_210 b_10 NI_10 NS_210 0 2.7805452070943426e-09
GC_10_211 b_10 NI_10 NS_211 0 2.2669800208487182e-03
GC_10_212 b_10 NI_10 NS_212 0 -7.3271184797746086e-04
GC_10_213 b_10 NI_10 NS_213 0 -1.8145925512065822e-06
GC_10_214 b_10 NI_10 NS_214 0 -1.2100366347261348e-07
GC_10_215 b_10 NI_10 NS_215 0 3.5967389934464771e-04
GC_10_216 b_10 NI_10 NS_216 0 -3.7513265311666104e-04
GC_10_217 b_10 NI_10 NS_217 0 -1.2776934268155008e-03
GC_10_218 b_10 NI_10 NS_218 0 3.4323481760863866e-04
GC_10_219 b_10 NI_10 NS_219 0 7.1251046997574004e-04
GC_10_220 b_10 NI_10 NS_220 0 -8.2802878809652410e-04
GC_10_221 b_10 NI_10 NS_221 0 -1.5019445016822380e-04
GC_10_222 b_10 NI_10 NS_222 0 1.3911406003945406e-03
GC_10_223 b_10 NI_10 NS_223 0 -1.3011798114619636e-03
GC_10_224 b_10 NI_10 NS_224 0 -7.6470496629918406e-04
GC_10_225 b_10 NI_10 NS_225 0 6.8660249331077170e-04
GC_10_226 b_10 NI_10 NS_226 0 -2.8573053971484439e-05
GC_10_227 b_10 NI_10 NS_227 0 -1.3696246571377591e-04
GC_10_228 b_10 NI_10 NS_228 0 1.4682625691307702e-03
GC_10_229 b_10 NI_10 NS_229 0 -7.1835131337681277e-04
GC_10_230 b_10 NI_10 NS_230 0 -5.4301922812627194e-04
GC_10_231 b_10 NI_10 NS_231 0 6.5087457242265373e-04
GC_10_232 b_10 NI_10 NS_232 0 1.9310986953437130e-04
GC_10_233 b_10 NI_10 NS_233 0 -3.0193392553707872e-06
GC_10_234 b_10 NI_10 NS_234 0 2.6012932960704071e-05
GC_10_235 b_10 NI_10 NS_235 0 -9.9212370732036759e-06
GC_10_236 b_10 NI_10 NS_236 0 -1.4257833116477586e-06
GC_10_237 b_10 NI_10 NS_237 0 7.0597005958012905e-09
GC_10_238 b_10 NI_10 NS_238 0 -1.0480243408264042e-08
GC_10_239 b_10 NI_10 NS_239 0 -6.2223258833533499e-10
GC_10_240 b_10 NI_10 NS_240 0 -2.1193868103984828e-09
GC_10_241 b_10 NI_10 NS_241 0 -7.5349025098013139e-02
GC_10_242 b_10 NI_10 NS_242 0 2.4900038185669118e-02
GC_10_243 b_10 NI_10 NS_243 0 1.9200001151674604e-05
GC_10_244 b_10 NI_10 NS_244 0 5.3863153288023733e-06
GC_10_245 b_10 NI_10 NS_245 0 1.8353501457195189e-02
GC_10_246 b_10 NI_10 NS_246 0 2.7965362161056183e-02
GC_10_247 b_10 NI_10 NS_247 0 -1.9176254794619312e-02
GC_10_248 b_10 NI_10 NS_248 0 8.3761062563849527e-03
GC_10_249 b_10 NI_10 NS_249 0 -5.5264811615611462e-03
GC_10_250 b_10 NI_10 NS_250 0 -2.3054149389419763e-02
GC_10_251 b_10 NI_10 NS_251 0 2.6687350720135401e-02
GC_10_252 b_10 NI_10 NS_252 0 -1.4576116513831968e-02
GC_10_253 b_10 NI_10 NS_253 0 3.4517304099459363e-02
GC_10_254 b_10 NI_10 NS_254 0 4.8628185950539042e-03
GC_10_255 b_10 NI_10 NS_255 0 9.6719768518995723e-03
GC_10_256 b_10 NI_10 NS_256 0 1.3692405563896538e-02
GC_10_257 b_10 NI_10 NS_257 0 -1.2370890739813352e-02
GC_10_258 b_10 NI_10 NS_258 0 1.1007933557513816e-02
GC_10_259 b_10 NI_10 NS_259 0 -1.1774534279057692e-02
GC_10_260 b_10 NI_10 NS_260 0 -1.2014125921970464e-02
GC_10_261 b_10 NI_10 NS_261 0 1.9793916906631927e-02
GC_10_262 b_10 NI_10 NS_262 0 -2.6023940213583004e-02
GC_10_263 b_10 NI_10 NS_263 0 9.6721527689412536e-04
GC_10_264 b_10 NI_10 NS_264 0 -1.0822023848425894e-03
GC_10_265 b_10 NI_10 NS_265 0 6.3094378459886691e-04
GC_10_266 b_10 NI_10 NS_266 0 3.4914512290628783e-04
GC_10_267 b_10 NI_10 NS_267 0 9.7107810517780465e-08
GC_10_268 b_10 NI_10 NS_268 0 4.1868745006954798e-07
GC_10_269 b_10 NI_10 NS_269 0 -1.0314537484996732e-08
GC_10_270 b_10 NI_10 NS_270 0 -1.9789123308592280e-08
GC_10_271 b_10 NI_10 NS_271 0 1.2659773860458307e-01
GC_10_272 b_10 NI_10 NS_272 0 -9.9682294588669361e-03
GC_10_273 b_10 NI_10 NS_273 0 -2.0418473141989621e-05
GC_10_274 b_10 NI_10 NS_274 0 -3.8273616432282964e-06
GC_10_275 b_10 NI_10 NS_275 0 -8.0908251645516703e-03
GC_10_276 b_10 NI_10 NS_276 0 6.4296780914413975e-04
GC_10_277 b_10 NI_10 NS_277 0 -1.9909397529217711e-03
GC_10_278 b_10 NI_10 NS_278 0 6.7353868360024935e-05
GC_10_279 b_10 NI_10 NS_279 0 -1.2598721021315526e-02
GC_10_280 b_10 NI_10 NS_280 0 8.2477756362525981e-03
GC_10_281 b_10 NI_10 NS_281 0 -1.0271315651357435e-02
GC_10_282 b_10 NI_10 NS_282 0 -6.2357810582910022e-04
GC_10_283 b_10 NI_10 NS_283 0 -3.5565687463906446e-03
GC_10_284 b_10 NI_10 NS_284 0 1.6966131545998259e-02
GC_10_285 b_10 NI_10 NS_285 0 -7.7825975278901357e-03
GC_10_286 b_10 NI_10 NS_286 0 1.3370077146006588e-02
GC_10_287 b_10 NI_10 NS_287 0 -3.9902969105566535e-03
GC_10_288 b_10 NI_10 NS_288 0 6.9628750442002054e-03
GC_10_289 b_10 NI_10 NS_289 0 -2.7633689428856480e-03
GC_10_290 b_10 NI_10 NS_290 0 1.2313501087860945e-02
GC_10_291 b_10 NI_10 NS_291 0 -2.2964016853188558e-02
GC_10_292 b_10 NI_10 NS_292 0 5.9629979338304768e-03
GC_10_293 b_10 NI_10 NS_293 0 -8.6294521792627408e-04
GC_10_294 b_10 NI_10 NS_294 0 8.0344078006492963e-04
GC_10_295 b_10 NI_10 NS_295 0 -5.1358588480691773e-04
GC_10_296 b_10 NI_10 NS_296 0 -4.3937294384617975e-04
GC_10_297 b_10 NI_10 NS_297 0 -6.4174258942450096e-08
GC_10_298 b_10 NI_10 NS_298 0 -1.9155152348216894e-07
GC_10_299 b_10 NI_10 NS_299 0 -3.0939577975637042e-09
GC_10_300 b_10 NI_10 NS_300 0 5.6381487193444053e-09
GC_10_301 b_10 NI_10 NS_301 0 1.3559941333469981e-03
GC_10_302 b_10 NI_10 NS_302 0 -1.2038862725508366e-03
GC_10_303 b_10 NI_10 NS_303 0 3.7357854959704748e-06
GC_10_304 b_10 NI_10 NS_304 0 2.8902026035869836e-07
GC_10_305 b_10 NI_10 NS_305 0 1.2297142344565206e-04
GC_10_306 b_10 NI_10 NS_306 0 8.9417630350379339e-04
GC_10_307 b_10 NI_10 NS_307 0 1.8425184633426490e-03
GC_10_308 b_10 NI_10 NS_308 0 -8.6745250025173847e-04
GC_10_309 b_10 NI_10 NS_309 0 -2.9665987272878436e-03
GC_10_310 b_10 NI_10 NS_310 0 -1.6486220358267413e-03
GC_10_311 b_10 NI_10 NS_311 0 2.2195000405747464e-03
GC_10_312 b_10 NI_10 NS_312 0 2.6689299046905438e-03
GC_10_313 b_10 NI_10 NS_313 0 -1.4401285736990593e-03
GC_10_314 b_10 NI_10 NS_314 0 -2.9129269897473424e-03
GC_10_315 b_10 NI_10 NS_315 0 1.0698835469290962e-03
GC_10_316 b_10 NI_10 NS_316 0 2.2566937004190159e-03
GC_10_317 b_10 NI_10 NS_317 0 -1.6275429696302858e-03
GC_10_318 b_10 NI_10 NS_318 0 -2.1363737894757092e-03
GC_10_319 b_10 NI_10 NS_319 0 4.2046390500930262e-04
GC_10_320 b_10 NI_10 NS_320 0 2.0118509055250845e-03
GC_10_321 b_10 NI_10 NS_321 0 2.1508474918553440e-04
GC_10_322 b_10 NI_10 NS_322 0 -2.1102705443109587e-03
GC_10_323 b_10 NI_10 NS_323 0 -4.3288629883400822e-06
GC_10_324 b_10 NI_10 NS_324 0 4.3527946950789731e-06
GC_10_325 b_10 NI_10 NS_325 0 -7.8948787043224797e-07
GC_10_326 b_10 NI_10 NS_326 0 -3.5249024235589959e-06
GC_10_327 b_10 NI_10 NS_327 0 -7.5479782475711162e-09
GC_10_328 b_10 NI_10 NS_328 0 2.2567554930169281e-08
GC_10_329 b_10 NI_10 NS_329 0 2.3359227883048457e-09
GC_10_330 b_10 NI_10 NS_330 0 1.5101868391132197e-09
GC_10_331 b_10 NI_10 NS_331 0 -5.5793667744484434e-04
GC_10_332 b_10 NI_10 NS_332 0 -2.9007725959459378e-03
GC_10_333 b_10 NI_10 NS_333 0 -6.1510036392310192e-06
GC_10_334 b_10 NI_10 NS_334 0 -3.8641563261376772e-07
GC_10_335 b_10 NI_10 NS_335 0 2.6869490494028630e-03
GC_10_336 b_10 NI_10 NS_336 0 -1.9871038099452520e-03
GC_10_337 b_10 NI_10 NS_337 0 -6.1985279242058227e-03
GC_10_338 b_10 NI_10 NS_338 0 1.7528661756157470e-03
GC_10_339 b_10 NI_10 NS_339 0 4.7653988676771859e-03
GC_10_340 b_10 NI_10 NS_340 0 -5.5287233157844951e-03
GC_10_341 b_10 NI_10 NS_341 0 -2.4763410507989937e-04
GC_10_342 b_10 NI_10 NS_342 0 7.2490256057337905e-03
GC_10_343 b_10 NI_10 NS_343 0 -6.3151048482298694e-03
GC_10_344 b_10 NI_10 NS_344 0 -5.0558262301611014e-03
GC_10_345 b_10 NI_10 NS_345 0 4.5028131999799671e-03
GC_10_346 b_10 NI_10 NS_346 0 -1.7122871003182898e-03
GC_10_347 b_10 NI_10 NS_347 0 -5.9097652360970085e-04
GC_10_348 b_10 NI_10 NS_348 0 6.9470812017020222e-03
GC_10_349 b_10 NI_10 NS_349 0 -3.4358134815053493e-03
GC_10_350 b_10 NI_10 NS_350 0 -3.6826642571445014e-03
GC_10_351 b_10 NI_10 NS_351 0 5.9256440462513420e-03
GC_10_352 b_10 NI_10 NS_352 0 3.9686043464200513e-04
GC_10_353 b_10 NI_10 NS_353 0 6.3854894322719412e-05
GC_10_354 b_10 NI_10 NS_354 0 8.4387918009252830e-06
GC_10_355 b_10 NI_10 NS_355 0 1.5113326183366396e-05
GC_10_356 b_10 NI_10 NS_356 0 3.9976048949888710e-05
GC_10_357 b_10 NI_10 NS_357 0 7.1155597467534361e-09
GC_10_358 b_10 NI_10 NS_358 0 -2.9351570048651540e-08
GC_10_359 b_10 NI_10 NS_359 0 -1.8855630146795669e-09
GC_10_360 b_10 NI_10 NS_360 0 -5.6002472516809174e-10
GD_10_1 b_10 NI_10 NA_1 0 7.7100769182345930e-06
GD_10_2 b_10 NI_10 NA_2 0 -1.7399465855375127e-06
GD_10_3 b_10 NI_10 NA_3 0 -9.0925700446016019e-06
GD_10_4 b_10 NI_10 NA_4 0 -1.1548347358558561e-06
GD_10_5 b_10 NI_10 NA_5 0 -6.2840280532848594e-05
GD_10_6 b_10 NI_10 NA_6 0 1.6921919802865686e-04
GD_10_7 b_10 NI_10 NA_7 0 -4.6753670194391321e-05
GD_10_8 b_10 NI_10 NA_8 0 2.3297112133392230e-03
GD_10_9 b_10 NI_10 NA_9 0 -9.9681628022031711e-03
GD_10_10 b_10 NI_10 NA_10 0 -4.0270205362663979e-02
GD_10_11 b_10 NI_10 NA_11 0 -9.1321497460458625e-05
GD_10_12 b_10 NI_10 NA_12 0 1.6055992846919956e-02
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 -3.0823727631184004e-05
GC_11_2 b_11 NI_11 NS_2 0 4.3670089324541465e-06
GC_11_3 b_11 NI_11 NS_3 0 -1.9330853974161223e-08
GC_11_4 b_11 NI_11 NS_4 0 3.1701890685135231e-10
GC_11_5 b_11 NI_11 NS_5 0 1.4873613175647958e-06
GC_11_6 b_11 NI_11 NS_6 0 4.2934783312556167e-07
GC_11_7 b_11 NI_11 NS_7 0 1.3519114160366522e-06
GC_11_8 b_11 NI_11 NS_8 0 -4.6262462874732642e-07
GC_11_9 b_11 NI_11 NS_9 0 2.0703115333573366e-06
GC_11_10 b_11 NI_11 NS_10 0 -5.7999530492363719e-07
GC_11_11 b_11 NI_11 NS_11 0 2.2940195380625270e-06
GC_11_12 b_11 NI_11 NS_12 0 -9.4237075984345602e-07
GC_11_13 b_11 NI_11 NS_13 0 1.8336243914951854e-06
GC_11_14 b_11 NI_11 NS_14 0 -2.7427283120849237e-06
GC_11_15 b_11 NI_11 NS_15 0 9.1064052578015001e-07
GC_11_16 b_11 NI_11 NS_16 0 -2.2464259863473185e-06
GC_11_17 b_11 NI_11 NS_17 0 1.6377250559358612e-06
GC_11_18 b_11 NI_11 NS_18 0 -2.1621584168854685e-06
GC_11_19 b_11 NI_11 NS_19 0 1.5040335360500440e-06
GC_11_20 b_11 NI_11 NS_20 0 -1.7689261237386512e-06
GC_11_21 b_11 NI_11 NS_21 0 5.2308084643623338e-06
GC_11_22 b_11 NI_11 NS_22 0 -4.1145699078184788e-07
GC_11_23 b_11 NI_11 NS_23 0 3.8002143715184491e-07
GC_11_24 b_11 NI_11 NS_24 0 -1.9138298657502977e-08
GC_11_25 b_11 NI_11 NS_25 0 3.5325243304420956e-08
GC_11_26 b_11 NI_11 NS_26 0 1.6834529456802702e-07
GC_11_27 b_11 NI_11 NS_27 0 8.1397291643913634e-11
GC_11_28 b_11 NI_11 NS_28 0 -1.5430950235420870e-12
GC_11_29 b_11 NI_11 NS_29 0 -4.0249872941911430e-11
GC_11_30 b_11 NI_11 NS_30 0 -1.3801720832448385e-10
GC_11_31 b_11 NI_11 NS_31 0 -1.5473889988650606e-05
GC_11_32 b_11 NI_11 NS_32 0 5.0273892886776762e-07
GC_11_33 b_11 NI_11 NS_33 0 9.6893771470450580e-09
GC_11_34 b_11 NI_11 NS_34 0 -7.3056664862293245e-11
GC_11_35 b_11 NI_11 NS_35 0 1.1231108643043090e-06
GC_11_36 b_11 NI_11 NS_36 0 2.1488802086211543e-07
GC_11_37 b_11 NI_11 NS_37 0 1.1947568429386556e-06
GC_11_38 b_11 NI_11 NS_38 0 -1.3852140496333040e-07
GC_11_39 b_11 NI_11 NS_39 0 9.0379855897045188e-07
GC_11_40 b_11 NI_11 NS_40 0 -1.0516120417753235e-06
GC_11_41 b_11 NI_11 NS_41 0 8.4623794634136026e-07
GC_11_42 b_11 NI_11 NS_42 0 -4.8065447231958376e-07
GC_11_43 b_11 NI_11 NS_43 0 1.5417938605430643e-06
GC_11_44 b_11 NI_11 NS_44 0 -9.6405365084387797e-07
GC_11_45 b_11 NI_11 NS_45 0 1.0933705349972386e-06
GC_11_46 b_11 NI_11 NS_46 0 -1.7255577280143064e-06
GC_11_47 b_11 NI_11 NS_47 0 1.0576544219613491e-06
GC_11_48 b_11 NI_11 NS_48 0 -2.2497661937693762e-06
GC_11_49 b_11 NI_11 NS_49 0 6.5021012309269962e-07
GC_11_50 b_11 NI_11 NS_50 0 -1.7357121787071843e-06
GC_11_51 b_11 NI_11 NS_51 0 1.7290798398709556e-06
GC_11_52 b_11 NI_11 NS_52 0 -2.0366571645801701e-06
GC_11_53 b_11 NI_11 NS_53 0 1.1291027791057958e-09
GC_11_54 b_11 NI_11 NS_54 0 -2.3439243766772798e-07
GC_11_55 b_11 NI_11 NS_55 0 1.1724055836403782e-07
GC_11_56 b_11 NI_11 NS_56 0 2.0287765950960443e-08
GC_11_57 b_11 NI_11 NS_57 0 -7.0700056815783025e-11
GC_11_58 b_11 NI_11 NS_58 0 5.3485839817208973e-11
GC_11_59 b_11 NI_11 NS_59 0 3.3464772892254874e-11
GC_11_60 b_11 NI_11 NS_60 0 1.2644123404053072e-10
GC_11_61 b_11 NI_11 NS_61 0 1.8113431637388908e-05
GC_11_62 b_11 NI_11 NS_62 0 -2.5825694303074572e-06
GC_11_63 b_11 NI_11 NS_63 0 1.0317757766121547e-08
GC_11_64 b_11 NI_11 NS_64 0 -2.6663569641060849e-10
GC_11_65 b_11 NI_11 NS_65 0 -1.2543602180116303e-06
GC_11_66 b_11 NI_11 NS_66 0 -1.1114242070879598e-06
GC_11_67 b_11 NI_11 NS_67 0 -2.4906504724769173e-06
GC_11_68 b_11 NI_11 NS_68 0 5.3778947066627186e-07
GC_11_69 b_11 NI_11 NS_69 0 -1.2738989980249836e-06
GC_11_70 b_11 NI_11 NS_70 0 2.6842757357846372e-06
GC_11_71 b_11 NI_11 NS_71 0 1.8130842781738599e-06
GC_11_72 b_11 NI_11 NS_72 0 7.9201546304975120e-07
GC_11_73 b_11 NI_11 NS_73 0 -2.7645308213271354e-06
GC_11_74 b_11 NI_11 NS_74 0 -1.3551195624953273e-06
GC_11_75 b_11 NI_11 NS_75 0 -2.1678156199766106e-06
GC_11_76 b_11 NI_11 NS_76 0 3.4714093661015785e-06
GC_11_77 b_11 NI_11 NS_77 0 1.2584624010284561e-06
GC_11_78 b_11 NI_11 NS_78 0 2.3719291982769907e-06
GC_11_79 b_11 NI_11 NS_79 0 -9.1723707796371916e-07
GC_11_80 b_11 NI_11 NS_80 0 -3.8008691972654707e-07
GC_11_81 b_11 NI_11 NS_81 0 -3.3257347950062878e-06
GC_11_82 b_11 NI_11 NS_82 0 6.2805342374894917e-07
GC_11_83 b_11 NI_11 NS_83 0 -1.4282104756105754e-07
GC_11_84 b_11 NI_11 NS_84 0 -7.6712456164825457e-08
GC_11_85 b_11 NI_11 NS_85 0 2.3256090064681787e-08
GC_11_86 b_11 NI_11 NS_86 0 -5.1807327356946550e-08
GC_11_87 b_11 NI_11 NS_87 0 -1.7982955237986058e-11
GC_11_88 b_11 NI_11 NS_88 0 -1.0110897146739927e-10
GC_11_89 b_11 NI_11 NS_89 0 -3.8114116637051826e-11
GC_11_90 b_11 NI_11 NS_90 0 -1.6273682434605962e-10
GC_11_91 b_11 NI_11 NS_91 0 -3.1942314572016432e-05
GC_11_92 b_11 NI_11 NS_92 0 3.5545366105807008e-06
GC_11_93 b_11 NI_11 NS_93 0 -1.3272793485770076e-08
GC_11_94 b_11 NI_11 NS_94 0 3.4691728173365932e-10
GC_11_95 b_11 NI_11 NS_95 0 2.0364670001880829e-06
GC_11_96 b_11 NI_11 NS_96 0 2.9512191742107880e-07
GC_11_97 b_11 NI_11 NS_97 0 1.7829864226807915e-06
GC_11_98 b_11 NI_11 NS_98 0 -1.7976013084453299e-06
GC_11_99 b_11 NI_11 NS_99 0 2.2339248333473268e-06
GC_11_100 b_11 NI_11 NS_100 0 -1.9710652114333812e-06
GC_11_101 b_11 NI_11 NS_101 0 1.2218452513452848e-06
GC_11_102 b_11 NI_11 NS_102 0 -1.5034940598631287e-06
GC_11_103 b_11 NI_11 NS_103 0 1.6567993701168351e-06
GC_11_104 b_11 NI_11 NS_104 0 -1.3902503954709503e-06
GC_11_105 b_11 NI_11 NS_105 0 1.7716184557332945e-06
GC_11_106 b_11 NI_11 NS_106 0 -3.2805696111864899e-06
GC_11_107 b_11 NI_11 NS_107 0 1.9903684318866199e-06
GC_11_108 b_11 NI_11 NS_108 0 -3.6368215152100026e-06
GC_11_109 b_11 NI_11 NS_109 0 7.3352842286435871e-07
GC_11_110 b_11 NI_11 NS_110 0 -3.3032759000963517e-06
GC_11_111 b_11 NI_11 NS_111 0 3.4149821290816017e-06
GC_11_112 b_11 NI_11 NS_112 0 -1.5015850174776164e-06
GC_11_113 b_11 NI_11 NS_113 0 2.6974181392513493e-07
GC_11_114 b_11 NI_11 NS_114 0 3.1441902922022971e-08
GC_11_115 b_11 NI_11 NS_115 0 1.3484828492346425e-08
GC_11_116 b_11 NI_11 NS_116 0 1.2312559914878238e-07
GC_11_117 b_11 NI_11 NS_117 0 2.5347194597801394e-11
GC_11_118 b_11 NI_11 NS_118 0 1.2044959952356605e-10
GC_11_119 b_11 NI_11 NS_119 0 3.7594593042667965e-11
GC_11_120 b_11 NI_11 NS_120 0 1.6468105670542902e-10
GC_11_121 b_11 NI_11 NS_121 0 -5.9645814179589012e-05
GC_11_122 b_11 NI_11 NS_122 0 -4.9654226832329376e-06
GC_11_123 b_11 NI_11 NS_123 0 -5.3039127016581464e-08
GC_11_124 b_11 NI_11 NS_124 0 -5.8090600318894306e-10
GC_11_125 b_11 NI_11 NS_125 0 -6.6949085803085650e-06
GC_11_126 b_11 NI_11 NS_126 0 -5.1567310813506849e-06
GC_11_127 b_11 NI_11 NS_127 0 -3.1760424629077256e-05
GC_11_128 b_11 NI_11 NS_128 0 1.3387790232780343e-05
GC_11_129 b_11 NI_11 NS_129 0 2.0720936087136196e-05
GC_11_130 b_11 NI_11 NS_130 0 6.7062458897435015e-05
GC_11_131 b_11 NI_11 NS_131 0 9.6708352137577259e-05
GC_11_132 b_11 NI_11 NS_132 0 4.8828679046986395e-06
GC_11_133 b_11 NI_11 NS_133 0 -1.5549097244462126e-05
GC_11_134 b_11 NI_11 NS_134 0 -9.0315248961858160e-05
GC_11_135 b_11 NI_11 NS_135 0 -2.8413734419844103e-05
GC_11_136 b_11 NI_11 NS_136 0 3.3448569808901569e-05
GC_11_137 b_11 NI_11 NS_137 0 5.9980502701859169e-05
GC_11_138 b_11 NI_11 NS_138 0 -4.9248339402518150e-06
GC_11_139 b_11 NI_11 NS_139 0 -4.5519423252404368e-06
GC_11_140 b_11 NI_11 NS_140 0 -5.6343191474996116e-05
GC_11_141 b_11 NI_11 NS_141 0 -2.2582440948652834e-05
GC_11_142 b_11 NI_11 NS_142 0 -1.3231851167627702e-05
GC_11_143 b_11 NI_11 NS_143 0 6.7346349071930674e-07
GC_11_144 b_11 NI_11 NS_144 0 -6.8427530532769317e-07
GC_11_145 b_11 NI_11 NS_145 0 3.8175827499149662e-07
GC_11_146 b_11 NI_11 NS_146 0 1.4884432558861510e-07
GC_11_147 b_11 NI_11 NS_147 0 1.7055251482896459e-10
GC_11_148 b_11 NI_11 NS_148 0 -7.6241219073555975e-11
GC_11_149 b_11 NI_11 NS_149 0 -7.2505239526567230e-11
GC_11_150 b_11 NI_11 NS_150 0 -4.3769883131512950e-10
GC_11_151 b_11 NI_11 NS_151 0 9.7557395329886029e-05
GC_11_152 b_11 NI_11 NS_152 0 -6.3843707189847951e-08
GC_11_153 b_11 NI_11 NS_153 0 3.9237402772074103e-08
GC_11_154 b_11 NI_11 NS_154 0 7.0029793324240431e-10
GC_11_155 b_11 NI_11 NS_155 0 3.8317168032099586e-07
GC_11_156 b_11 NI_11 NS_156 0 -1.4093022854415997e-06
GC_11_157 b_11 NI_11 NS_157 0 -9.1557179410113740e-06
GC_11_158 b_11 NI_11 NS_158 0 2.4452150415078876e-05
GC_11_159 b_11 NI_11 NS_159 0 7.9465466458638817e-05
GC_11_160 b_11 NI_11 NS_160 0 8.7690493634677645e-06
GC_11_161 b_11 NI_11 NS_161 0 1.1469116997558431e-05
GC_11_162 b_11 NI_11 NS_162 0 -7.9811146028748811e-05
GC_11_163 b_11 NI_11 NS_163 0 -6.7934164376543840e-06
GC_11_164 b_11 NI_11 NS_164 0 -4.3503400171874512e-05
GC_11_165 b_11 NI_11 NS_165 0 -9.4941653448967731e-05
GC_11_166 b_11 NI_11 NS_166 0 -5.4391210605067479e-05
GC_11_167 b_11 NI_11 NS_167 0 -4.5788269463091457e-05
GC_11_168 b_11 NI_11 NS_168 0 5.2625383098840877e-05
GC_11_169 b_11 NI_11 NS_169 0 -3.1146648530543229e-05
GC_11_170 b_11 NI_11 NS_170 0 1.2605040941722188e-05
GC_11_171 b_11 NI_11 NS_171 0 -1.5816707738013603e-05
GC_11_172 b_11 NI_11 NS_172 0 4.9605030382544310e-05
GC_11_173 b_11 NI_11 NS_173 0 -7.3647521127344567e-07
GC_11_174 b_11 NI_11 NS_174 0 -4.4503378163759115e-07
GC_11_175 b_11 NI_11 NS_175 0 1.3570639180348460e-07
GC_11_176 b_11 NI_11 NS_176 0 -3.6538842981793888e-07
GC_11_177 b_11 NI_11 NS_177 0 -1.5129394464217304e-10
GC_11_178 b_11 NI_11 NS_178 0 9.3552939172471939e-11
GC_11_179 b_11 NI_11 NS_179 0 7.1163720541317350e-11
GC_11_180 b_11 NI_11 NS_180 0 4.3626480307279723e-10
GC_11_181 b_11 NI_11 NS_181 0 1.3201864306430165e-04
GC_11_182 b_11 NI_11 NS_182 0 2.3805681736583100e-06
GC_11_183 b_11 NI_11 NS_183 0 -2.0660917225322691e-07
GC_11_184 b_11 NI_11 NS_184 0 -9.2214651690512373e-09
GC_11_185 b_11 NI_11 NS_185 0 5.0256255547160094e-05
GC_11_186 b_11 NI_11 NS_186 0 -1.8215604839286691e-06
GC_11_187 b_11 NI_11 NS_187 0 2.5946087105737084e-05
GC_11_188 b_11 NI_11 NS_188 0 -7.5678260738690886e-06
GC_11_189 b_11 NI_11 NS_189 0 2.2965371940241984e-05
GC_11_190 b_11 NI_11 NS_190 0 -2.6891282391372506e-04
GC_11_191 b_11 NI_11 NS_191 0 -2.9159830523542391e-04
GC_11_192 b_11 NI_11 NS_192 0 4.0432223915224275e-05
GC_11_193 b_11 NI_11 NS_193 0 -5.4703354488949928e-05
GC_11_194 b_11 NI_11 NS_194 0 2.2080859819961370e-04
GC_11_195 b_11 NI_11 NS_195 0 1.6828542649852067e-04
GC_11_196 b_11 NI_11 NS_196 0 -1.0559560027124265e-04
GC_11_197 b_11 NI_11 NS_197 0 -1.8061281475558486e-04
GC_11_198 b_11 NI_11 NS_198 0 6.1001806811667681e-05
GC_11_199 b_11 NI_11 NS_199 0 -5.0282958352480020e-05
GC_11_200 b_11 NI_11 NS_200 0 1.2038418616110363e-04
GC_11_201 b_11 NI_11 NS_201 0 1.3801948080609372e-04
GC_11_202 b_11 NI_11 NS_202 0 7.0744591543147879e-05
GC_11_203 b_11 NI_11 NS_203 0 -7.0772161959050636e-09
GC_11_204 b_11 NI_11 NS_204 0 4.3653236796635033e-06
GC_11_205 b_11 NI_11 NS_205 0 -2.0291298390963895e-06
GC_11_206 b_11 NI_11 NS_206 0 5.4131714189655765e-08
GC_11_207 b_11 NI_11 NS_207 0 6.2761200539424835e-10
GC_11_208 b_11 NI_11 NS_208 0 -6.3109571132238463e-10
GC_11_209 b_11 NI_11 NS_209 0 -1.5188949591625093e-10
GC_11_210 b_11 NI_11 NS_210 0 -1.2381738205099187e-09
GC_11_211 b_11 NI_11 NS_211 0 4.6478457846633833e-05
GC_11_212 b_11 NI_11 NS_212 0 9.2529799983019737e-05
GC_11_213 b_11 NI_11 NS_213 0 2.8968373521672612e-07
GC_11_214 b_11 NI_11 NS_214 0 8.4521573109726061e-09
GC_11_215 b_11 NI_11 NS_215 0 -3.9577689407224088e-05
GC_11_216 b_11 NI_11 NS_216 0 -8.5753646500502374e-05
GC_11_217 b_11 NI_11 NS_217 0 -2.2600522934228568e-04
GC_11_218 b_11 NI_11 NS_218 0 9.6583222237372243e-05
GC_11_219 b_11 NI_11 NS_219 0 2.8263681148531732e-04
GC_11_220 b_11 NI_11 NS_220 0 1.5421636311087781e-04
GC_11_221 b_11 NI_11 NS_221 0 -3.0568635839092669e-04
GC_11_222 b_11 NI_11 NS_222 0 -2.0974779126653104e-04
GC_11_223 b_11 NI_11 NS_223 0 1.8427059781613069e-04
GC_11_224 b_11 NI_11 NS_224 0 3.8931158859503625e-04
GC_11_225 b_11 NI_11 NS_225 0 -9.5460092402372318e-05
GC_11_226 b_11 NI_11 NS_226 0 -1.5686561480074757e-04
GC_11_227 b_11 NI_11 NS_227 0 2.3694532313688323e-04
GC_11_228 b_11 NI_11 NS_228 0 2.1575073577385638e-04
GC_11_229 b_11 NI_11 NS_229 0 -5.9308459434402274e-05
GC_11_230 b_11 NI_11 NS_230 0 -2.0763778450584754e-04
GC_11_231 b_11 NI_11 NS_231 0 -1.2638859607301856e-06
GC_11_232 b_11 NI_11 NS_232 0 2.1361782465272820e-04
GC_11_233 b_11 NI_11 NS_233 0 -2.2353355517798852e-06
GC_11_234 b_11 NI_11 NS_234 0 -4.6168357245215342e-08
GC_11_235 b_11 NI_11 NS_235 0 -4.0400826112504691e-07
GC_11_236 b_11 NI_11 NS_236 0 -4.3854105858847051e-07
GC_11_237 b_11 NI_11 NS_237 0 -7.4184942470670140e-10
GC_11_238 b_11 NI_11 NS_238 0 5.0959123862200379e-10
GC_11_239 b_11 NI_11 NS_239 0 1.5238772740126830e-10
GC_11_240 b_11 NI_11 NS_240 0 1.2350645627168486e-09
GC_11_241 b_11 NI_11 NS_241 0 -5.5793667744495872e-04
GC_11_242 b_11 NI_11 NS_242 0 -2.9007725959458949e-03
GC_11_243 b_11 NI_11 NS_243 0 -6.1510036392317366e-06
GC_11_244 b_11 NI_11 NS_244 0 -3.8641563261374454e-07
GC_11_245 b_11 NI_11 NS_245 0 2.6869490494028573e-03
GC_11_246 b_11 NI_11 NS_246 0 -1.9871038099452572e-03
GC_11_247 b_11 NI_11 NS_247 0 -6.1985279242058348e-03
GC_11_248 b_11 NI_11 NS_248 0 1.7528661756157518e-03
GC_11_249 b_11 NI_11 NS_249 0 4.7653988676771824e-03
GC_11_250 b_11 NI_11 NS_250 0 -5.5287233157844768e-03
GC_11_251 b_11 NI_11 NS_251 0 -2.4763410507990137e-04
GC_11_252 b_11 NI_11 NS_252 0 7.2490256057338156e-03
GC_11_253 b_11 NI_11 NS_253 0 -6.3151048482298373e-03
GC_11_254 b_11 NI_11 NS_254 0 -5.0558262301610866e-03
GC_11_255 b_11 NI_11 NS_255 0 4.5028131999799818e-03
GC_11_256 b_11 NI_11 NS_256 0 -1.7122871003182926e-03
GC_11_257 b_11 NI_11 NS_257 0 -5.9097652360967623e-04
GC_11_258 b_11 NI_11 NS_258 0 6.9470812017020135e-03
GC_11_259 b_11 NI_11 NS_259 0 -3.4358134815053419e-03
GC_11_260 b_11 NI_11 NS_260 0 -3.6826642571445062e-03
GC_11_261 b_11 NI_11 NS_261 0 5.9256440462513681e-03
GC_11_262 b_11 NI_11 NS_262 0 3.9686043464202503e-04
GC_11_263 b_11 NI_11 NS_263 0 6.3854894322724209e-05
GC_11_264 b_11 NI_11 NS_264 0 8.4387918009285204e-06
GC_11_265 b_11 NI_11 NS_265 0 1.5113326183364838e-05
GC_11_266 b_11 NI_11 NS_266 0 3.9976048949890865e-05
GC_11_267 b_11 NI_11 NS_267 0 7.1155597467522541e-09
GC_11_268 b_11 NI_11 NS_268 0 -2.9351570048644324e-08
GC_11_269 b_11 NI_11 NS_269 0 -1.8855630146804706e-09
GC_11_270 b_11 NI_11 NS_270 0 -5.6002472516841082e-10
GC_11_271 b_11 NI_11 NS_271 0 1.3561032718190709e-03
GC_11_272 b_11 NI_11 NS_272 0 -1.2038975406755130e-03
GC_11_273 b_11 NI_11 NS_273 0 3.7358057183382851e-06
GC_11_274 b_11 NI_11 NS_274 0 2.8901996539223217e-07
GC_11_275 b_11 NI_11 NS_275 0 1.2295932909834015e-04
GC_11_276 b_11 NI_11 NS_276 0 8.9417142188338687e-04
GC_11_277 b_11 NI_11 NS_277 0 1.8425106140205765e-03
GC_11_278 b_11 NI_11 NS_278 0 -8.6745792168850218e-04
GC_11_279 b_11 NI_11 NS_279 0 -2.9666020918209190e-03
GC_11_280 b_11 NI_11 NS_280 0 -1.6486044684690816e-03
GC_11_281 b_11 NI_11 NS_281 0 2.2194915709220714e-03
GC_11_282 b_11 NI_11 NS_282 0 2.6689308128691100e-03
GC_11_283 b_11 NI_11 NS_283 0 -1.4401415521705441e-03
GC_11_284 b_11 NI_11 NS_284 0 -2.9129099036704258e-03
GC_11_285 b_11 NI_11 NS_285 0 1.0698831151070159e-03
GC_11_286 b_11 NI_11 NS_286 0 2.2566994843893399e-03
GC_11_287 b_11 NI_11 NS_287 0 -1.6275472028653586e-03
GC_11_288 b_11 NI_11 NS_288 0 -2.1363613895425330e-03
GC_11_289 b_11 NI_11 NS_289 0 4.2046148382028176e-04
GC_11_290 b_11 NI_11 NS_290 0 2.0118573278588596e-03
GC_11_291 b_11 NI_11 NS_291 0 2.1506806916417667e-04
GC_11_292 b_11 NI_11 NS_292 0 -2.1102648323654927e-03
GC_11_293 b_11 NI_11 NS_293 0 -4.3297592914652035e-06
GC_11_294 b_11 NI_11 NS_294 0 4.3533743092581193e-06
GC_11_295 b_11 NI_11 NS_295 0 -7.8987902033922279e-07
GC_11_296 b_11 NI_11 NS_296 0 -3.5253886213821896e-06
GC_11_297 b_11 NI_11 NS_297 0 -7.5480237649974902e-09
GC_11_298 b_11 NI_11 NS_298 0 2.2567511706671412e-08
GC_11_299 b_11 NI_11 NS_299 0 2.3359259828195180e-09
GC_11_300 b_11 NI_11 NS_300 0 1.5101887849105698e-09
GC_11_301 b_11 NI_11 NS_301 0 1.2526109539007568e-01
GC_11_302 b_11 NI_11 NS_302 0 -9.7551767127498357e-03
GC_11_303 b_11 NI_11 NS_303 0 -2.1879130952244503e-05
GC_11_304 b_11 NI_11 NS_304 0 -3.7984595388708525e-06
GC_11_305 b_11 NI_11 NS_305 0 -8.0420617900947549e-03
GC_11_306 b_11 NI_11 NS_306 0 6.5371441387693588e-04
GC_11_307 b_11 NI_11 NS_307 0 -1.9771768576952735e-03
GC_11_308 b_11 NI_11 NS_308 0 1.0157035349987814e-04
GC_11_309 b_11 NI_11 NS_309 0 -1.2487318678050897e-02
GC_11_310 b_11 NI_11 NS_310 0 8.2382561606138393e-03
GC_11_311 b_11 NI_11 NS_311 0 -1.0111831129700351e-02
GC_11_312 b_11 NI_11 NS_312 0 -5.9611104333092530e-04
GC_11_313 b_11 NI_11 NS_313 0 -3.4891067426213330e-03
GC_11_314 b_11 NI_11 NS_314 0 1.6807114589681565e-02
GC_11_315 b_11 NI_11 NS_315 0 -7.7156937405831729e-03
GC_11_316 b_11 NI_11 NS_316 0 1.3269795962382869e-02
GC_11_317 b_11 NI_11 NS_317 0 -3.8876506552716931e-03
GC_11_318 b_11 NI_11 NS_318 0 6.8943368294903272e-03
GC_11_319 b_11 NI_11 NS_319 0 -2.7117305920497554e-03
GC_11_320 b_11 NI_11 NS_320 0 1.2199574043009039e-02
GC_11_321 b_11 NI_11 NS_321 0 -2.2742235751446072e-02
GC_11_322 b_11 NI_11 NS_322 0 5.9617076729824381e-03
GC_11_323 b_11 NI_11 NS_323 0 -8.4148616670018915e-04
GC_11_324 b_11 NI_11 NS_324 0 8.1300281436196540e-04
GC_11_325 b_11 NI_11 NS_325 0 -5.1564586368886708e-04
GC_11_326 b_11 NI_11 NS_326 0 -4.3052022749988660e-04
GC_11_327 b_11 NI_11 NS_327 0 -5.9275351095747621e-08
GC_11_328 b_11 NI_11 NS_328 0 -1.8756503205183451e-07
GC_11_329 b_11 NI_11 NS_329 0 -3.3579624240941055e-09
GC_11_330 b_11 NI_11 NS_330 0 5.3365700592452756e-09
GC_11_331 b_11 NI_11 NS_331 0 -7.0424905809883628e-02
GC_11_332 b_11 NI_11 NS_332 0 2.4192876081987787e-02
GC_11_333 b_11 NI_11 NS_333 0 2.2092718039702866e-05
GC_11_334 b_11 NI_11 NS_334 0 5.3186649768010776e-06
GC_11_335 b_11 NI_11 NS_335 0 1.8108336157749056e-02
GC_11_336 b_11 NI_11 NS_336 0 2.7946288701311325e-02
GC_11_337 b_11 NI_11 NS_337 0 -1.9395014030018094e-02
GC_11_338 b_11 NI_11 NS_338 0 8.3724650245715019e-03
GC_11_339 b_11 NI_11 NS_339 0 -5.8925725876615162e-03
GC_11_340 b_11 NI_11 NS_340 0 -2.2930858204175047e-02
GC_11_341 b_11 NI_11 NS_341 0 2.6387227054613955e-02
GC_11_342 b_11 NI_11 NS_342 0 -1.4337546293758328e-02
GC_11_343 b_11 NI_11 NS_343 0 3.4164774325802713e-02
GC_11_344 b_11 NI_11 NS_344 0 5.2157308909303946e-03
GC_11_345 b_11 NI_11 NS_345 0 9.5147656217769820e-03
GC_11_346 b_11 NI_11 NS_346 0 1.4168167210601887e-02
GC_11_347 b_11 NI_11 NS_347 0 -1.2626472890820509e-02
GC_11_348 b_11 NI_11 NS_348 0 1.1356489359880114e-02
GC_11_349 b_11 NI_11 NS_349 0 -1.1978296501839885e-02
GC_11_350 b_11 NI_11 NS_350 0 -1.1686204064082792e-02
GC_11_351 b_11 NI_11 NS_351 0 1.9051213307178776e-02
GC_11_352 b_11 NI_11 NS_352 0 -2.5965268695815308e-02
GC_11_353 b_11 NI_11 NS_353 0 9.0695156094665645e-04
GC_11_354 b_11 NI_11 NS_354 0 -1.0849123617883360e-03
GC_11_355 b_11 NI_11 NS_355 0 6.2679895063856366e-04
GC_11_356 b_11 NI_11 NS_356 0 3.2176415380547621e-04
GC_11_357 b_11 NI_11 NS_357 0 9.0179859031587707e-08
GC_11_358 b_11 NI_11 NS_358 0 4.0615052475847408e-07
GC_11_359 b_11 NI_11 NS_359 0 -9.1806540327368541e-09
GC_11_360 b_11 NI_11 NS_360 0 -1.8630948815939443e-08
GD_11_1 b_11 NI_11 NA_1 0 5.1396599105486145e-06
GD_11_2 b_11 NI_11 NA_2 0 2.7202905211608921e-06
GD_11_3 b_11 NI_11 NA_3 0 -1.7302922944589438e-06
GD_11_4 b_11 NI_11 NA_4 0 7.7454570899349087e-06
GD_11_5 b_11 NI_11 NA_5 0 3.8071667517034134e-06
GD_11_6 b_11 NI_11 NA_6 0 8.3909795482100851e-06
GD_11_7 b_11 NI_11 NA_7 0 1.7036754106096778e-04
GD_11_8 b_11 NI_11 NA_8 0 -6.0828848395370701e-05
GD_11_9 b_11 NI_11 NA_9 0 1.6055992846919932e-02
GD_11_10 b_11 NI_11 NA_10 0 -9.1338169335060580e-05
GD_11_11 b_11 NI_11 NA_11 0 -4.0049979026644353e-02
GD_11_12 b_11 NI_11 NA_12 0 -1.0827019600119886e-02
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -1.5512843760828022e-05
GC_12_2 b_12 NI_12 NS_2 0 5.0658018986112194e-07
GC_12_3 b_12 NI_12 NS_3 0 9.6809792669585177e-09
GC_12_4 b_12 NI_12 NS_4 0 -7.2853288082770494e-11
GC_12_5 b_12 NI_12 NS_5 0 1.1250117987776328e-06
GC_12_6 b_12 NI_12 NS_6 0 2.1547643929355221e-07
GC_12_7 b_12 NI_12 NS_7 0 1.1958322134559715e-06
GC_12_8 b_12 NI_12 NS_8 0 -1.3674754819125972e-07
GC_12_9 b_12 NI_12 NS_9 0 9.0974032144358162e-07
GC_12_10 b_12 NI_12 NS_10 0 -1.0540136594587366e-06
GC_12_11 b_12 NI_12 NS_11 0 8.4885502123982175e-07
GC_12_12 b_12 NI_12 NS_12 0 -4.8307570308525316e-07
GC_12_13 b_12 NI_12 NS_13 0 1.5466607638577416e-06
GC_12_14 b_12 NI_12 NS_14 0 -9.6833614703877404e-07
GC_12_15 b_12 NI_12 NS_15 0 1.0931331871668815e-06
GC_12_16 b_12 NI_12 NS_16 0 -1.7311316268459843e-06
GC_12_17 b_12 NI_12 NS_17 0 1.0586185021998440e-06
GC_12_18 b_12 NI_12 NS_18 0 -2.2535263696143644e-06
GC_12_19 b_12 NI_12 NS_19 0 6.5143382120372656e-07
GC_12_20 b_12 NI_12 NS_20 0 -1.7389303147955882e-06
GC_12_21 b_12 NI_12 NS_21 0 1.7338396595740194e-06
GC_12_22 b_12 NI_12 NS_22 0 -2.0387001691510138e-06
GC_12_23 b_12 NI_12 NS_23 0 1.4317140788886278e-09
GC_12_24 b_12 NI_12 NS_24 0 -2.3457323863841308e-07
GC_12_25 b_12 NI_12 NS_25 0 1.1736231963715717e-07
GC_12_26 b_12 NI_12 NS_26 0 2.0439137536823832e-08
GC_12_27 b_12 NI_12 NS_27 0 -7.0685136076094723e-11
GC_12_28 b_12 NI_12 NS_28 0 5.3530541519299656e-11
GC_12_29 b_12 NI_12 NS_29 0 3.3461059845730853e-11
GC_12_30 b_12 NI_12 NS_30 0 1.2644061918167438e-10
GC_12_31 b_12 NI_12 NS_31 0 -3.0823040270804093e-05
GC_12_32 b_12 NI_12 NS_32 0 4.3669468422745775e-06
GC_12_33 b_12 NI_12 NS_33 0 -1.9330742519410010e-08
GC_12_34 b_12 NI_12 NS_34 0 3.1701658828735141e-10
GC_12_35 b_12 NI_12 NS_35 0 1.4873081199441756e-06
GC_12_36 b_12 NI_12 NS_36 0 4.2936619309321078e-07
GC_12_37 b_12 NI_12 NS_37 0 1.3518704852220470e-06
GC_12_38 b_12 NI_12 NS_38 0 -4.6259409435668413e-07
GC_12_39 b_12 NI_12 NS_39 0 2.0702781927689712e-06
GC_12_40 b_12 NI_12 NS_40 0 -5.7993619335547945e-07
GC_12_41 b_12 NI_12 NS_41 0 2.2939800063288094e-06
GC_12_42 b_12 NI_12 NS_42 0 -9.4232592610279051e-07
GC_12_43 b_12 NI_12 NS_43 0 1.8336065615527967e-06
GC_12_44 b_12 NI_12 NS_44 0 -2.7426509024983493e-06
GC_12_45 b_12 NI_12 NS_45 0 9.1063614964674604e-07
GC_12_46 b_12 NI_12 NS_46 0 -2.2463637348424066e-06
GC_12_47 b_12 NI_12 NS_47 0 1.6377156315622485e-06
GC_12_48 b_12 NI_12 NS_48 0 -2.1620950251060020e-06
GC_12_49 b_12 NI_12 NS_49 0 1.5040099976795839e-06
GC_12_50 b_12 NI_12 NS_50 0 -1.7688845946332439e-06
GC_12_51 b_12 NI_12 NS_51 0 5.2307159666934484e-06
GC_12_52 b_12 NI_12 NS_52 0 -4.1141520671373536e-07
GC_12_53 b_12 NI_12 NS_53 0 3.8001754464708846e-07
GC_12_54 b_12 NI_12 NS_54 0 -1.9134695060663915e-08
GC_12_55 b_12 NI_12 NS_55 0 3.5322959308730633e-08
GC_12_56 b_12 NI_12 NS_56 0 1.6834348662888756e-07
GC_12_57 b_12 NI_12 NS_57 0 8.1397041713145483e-11
GC_12_58 b_12 NI_12 NS_58 0 -1.5436030597837432e-12
GC_12_59 b_12 NI_12 NS_59 0 -4.0249851024499831e-11
GC_12_60 b_12 NI_12 NS_60 0 -1.3801730174680396e-10
GC_12_61 b_12 NI_12 NS_61 0 -3.1941706375645535e-05
GC_12_62 b_12 NI_12 NS_62 0 3.5544757236791198e-06
GC_12_63 b_12 NI_12 NS_63 0 -1.3272658508133015e-08
GC_12_64 b_12 NI_12 NS_64 0 3.4691405420875378e-10
GC_12_65 b_12 NI_12 NS_65 0 2.0364022194153890e-06
GC_12_66 b_12 NI_12 NS_66 0 2.9506699234426061e-07
GC_12_67 b_12 NI_12 NS_67 0 1.7829377447696838e-06
GC_12_68 b_12 NI_12 NS_68 0 -1.7976020737886732e-06
GC_12_69 b_12 NI_12 NS_69 0 2.2338176821819135e-06
GC_12_70 b_12 NI_12 NS_70 0 -1.9709266439781780e-06
GC_12_71 b_12 NI_12 NS_71 0 1.2218261976768591e-06
GC_12_72 b_12 NI_12 NS_72 0 -1.5034225728942779e-06
GC_12_73 b_12 NI_12 NS_73 0 1.6567929693176164e-06
GC_12_74 b_12 NI_12 NS_74 0 -1.3901782539703927e-06
GC_12_75 b_12 NI_12 NS_75 0 1.7716542854877118e-06
GC_12_76 b_12 NI_12 NS_76 0 -3.2805214525178879e-06
GC_12_77 b_12 NI_12 NS_77 0 1.9903580165892476e-06
GC_12_78 b_12 NI_12 NS_78 0 -3.6367827527663803e-06
GC_12_79 b_12 NI_12 NS_79 0 7.3350407191061473e-07
GC_12_80 b_12 NI_12 NS_80 0 -3.3032495696950245e-06
GC_12_81 b_12 NI_12 NS_81 0 3.4148895591534180e-06
GC_12_82 b_12 NI_12 NS_82 0 -1.5015526489099124e-06
GC_12_83 b_12 NI_12 NS_83 0 2.6973765497490347e-07
GC_12_84 b_12 NI_12 NS_84 0 3.1444630836105894e-08
GC_12_85 b_12 NI_12 NS_85 0 1.3483163339089980e-08
GC_12_86 b_12 NI_12 NS_86 0 1.2312362219403316e-07
GC_12_87 b_12 NI_12 NS_87 0 2.5346960573812517e-11
GC_12_88 b_12 NI_12 NS_88 0 1.2044891910472609e-10
GC_12_89 b_12 NI_12 NS_89 0 3.7594669849561823e-11
GC_12_90 b_12 NI_12 NS_90 0 1.6468111867277255e-10
GC_12_91 b_12 NI_12 NS_91 0 1.7901684647746171e-05
GC_12_92 b_12 NI_12 NS_92 0 -2.5568017853157559e-06
GC_12_93 b_12 NI_12 NS_93 0 1.0257140711448923e-08
GC_12_94 b_12 NI_12 NS_94 0 -2.6532702970004855e-10
GC_12_95 b_12 NI_12 NS_95 0 -1.2423327627163728e-06
GC_12_96 b_12 NI_12 NS_96 0 -1.1108574310229257e-06
GC_12_97 b_12 NI_12 NS_97 0 -2.4790778399937317e-06
GC_12_98 b_12 NI_12 NS_98 0 5.4356146833372395e-07
GC_12_99 b_12 NI_12 NS_99 0 -1.2528111426180260e-06
GC_12_100 b_12 NI_12 NS_100 0 2.6650236111097218e-06
GC_12_101 b_12 NI_12 NS_101 0 1.8273669267196241e-06
GC_12_102 b_12 NI_12 NS_102 0 7.7991584884606525e-07
GC_12_103 b_12 NI_12 NS_103 0 -2.7635943481990548e-06
GC_12_104 b_12 NI_12 NS_104 0 -1.3704503864577437e-06
GC_12_105 b_12 NI_12 NS_105 0 -2.1566729364974156e-06
GC_12_106 b_12 NI_12 NS_106 0 3.4557465709135474e-06
GC_12_107 b_12 NI_12 NS_107 0 1.2689232433253989e-06
GC_12_108 b_12 NI_12 NS_108 0 2.3550489266337866e-06
GC_12_109 b_12 NI_12 NS_109 0 -9.0819764939830378e-07
GC_12_110 b_12 NI_12 NS_110 0 -3.9371811200275470e-07
GC_12_111 b_12 NI_12 NS_111 0 -3.2916092198901868e-06
GC_12_112 b_12 NI_12 NS_112 0 6.2256349070727039e-07
GC_12_113 b_12 NI_12 NS_113 0 -1.4055850688761744e-07
GC_12_114 b_12 NI_12 NS_114 0 -7.7795688800129355e-08
GC_12_115 b_12 NI_12 NS_115 0 2.3942271505905175e-08
GC_12_116 b_12 NI_12 NS_116 0 -5.0742649535358238e-08
GC_12_117 b_12 NI_12 NS_117 0 -1.7904008864596788e-11
GC_12_118 b_12 NI_12 NS_118 0 -1.0084239029427359e-10
GC_12_119 b_12 NI_12 NS_119 0 -3.8149507100741912e-11
GC_12_120 b_12 NI_12 NS_120 0 -1.6277828897252798e-10
GC_12_121 b_12 NI_12 NS_121 0 9.6421904204612596e-05
GC_12_122 b_12 NI_12 NS_122 0 2.8798298722863413e-08
GC_12_123 b_12 NI_12 NS_123 0 3.9109902994842181e-08
GC_12_124 b_12 NI_12 NS_124 0 7.0175516133725524e-10
GC_12_125 b_12 NI_12 NS_125 0 5.3823009377278277e-07
GC_12_126 b_12 NI_12 NS_126 0 -1.3492803774882851e-06
GC_12_127 b_12 NI_12 NS_127 0 -9.0392075218832134e-06
GC_12_128 b_12 NI_12 NS_128 0 2.4491118610467673e-05
GC_12_129 b_12 NI_12 NS_129 0 7.9496249003478073e-05
GC_12_130 b_12 NI_12 NS_130 0 8.5223804813320087e-06
GC_12_131 b_12 NI_12 NS_131 0 1.1537152841624553e-05
GC_12_132 b_12 NI_12 NS_132 0 -7.9841300146477330e-05
GC_12_133 b_12 NI_12 NS_133 0 -6.6585354713700961e-06
GC_12_134 b_12 NI_12 NS_134 0 -4.3699588921316881e-05
GC_12_135 b_12 NI_12 NS_135 0 -9.4957032436552500e-05
GC_12_136 b_12 NI_12 NS_136 0 -5.4470338132393808e-05
GC_12_137 b_12 NI_12 NS_137 0 -4.5766854754057635e-05
GC_12_138 b_12 NI_12 NS_138 0 5.2480776703023897e-05
GC_12_139 b_12 NI_12 NS_139 0 -3.1138984417523489e-05
GC_12_140 b_12 NI_12 NS_140 0 1.2530530165198239e-05
GC_12_141 b_12 NI_12 NS_141 0 -1.5669043915097225e-05
GC_12_142 b_12 NI_12 NS_142 0 4.9521443465887577e-05
GC_12_143 b_12 NI_12 NS_143 0 -7.3125496211270450e-07
GC_12_144 b_12 NI_12 NS_144 0 -4.5045377139180121e-07
GC_12_145 b_12 NI_12 NS_145 0 1.3959012716351077e-07
GC_12_146 b_12 NI_12 NS_146 0 -3.6272337742469160e-07
GC_12_147 b_12 NI_12 NS_147 0 -1.5098902260456545e-10
GC_12_148 b_12 NI_12 NS_148 0 9.3782710567231788e-11
GC_12_149 b_12 NI_12 NS_149 0 7.1151103642492952e-11
GC_12_150 b_12 NI_12 NS_150 0 4.3624309224129565e-10
GC_12_151 b_12 NI_12 NS_151 0 -5.9716322203039303e-05
GC_12_152 b_12 NI_12 NS_152 0 -4.9579622987011849e-06
GC_12_153 b_12 NI_12 NS_153 0 -5.3052463737390226e-08
GC_12_154 b_12 NI_12 NS_154 0 -5.8065267811040298e-10
GC_12_155 b_12 NI_12 NS_155 0 -6.6914496936773381e-06
GC_12_156 b_12 NI_12 NS_156 0 -5.1560606179414791e-06
GC_12_157 b_12 NI_12 NS_157 0 -3.1757005679094240e-05
GC_12_158 b_12 NI_12 NS_158 0 1.3388490836460287e-05
GC_12_159 b_12 NI_12 NS_159 0 2.0727018897852640e-05
GC_12_160 b_12 NI_12 NS_160 0 6.7059935066892239e-05
GC_12_161 b_12 NI_12 NS_161 0 9.6715112128875017e-05
GC_12_162 b_12 NI_12 NS_162 0 4.8803892469505836e-06
GC_12_163 b_12 NI_12 NS_163 0 -1.5545038770787305e-05
GC_12_164 b_12 NI_12 NS_164 0 -9.0322207065075258e-05
GC_12_165 b_12 NI_12 NS_165 0 -2.8410494947319909e-05
GC_12_166 b_12 NI_12 NS_166 0 3.3441985365011286e-05
GC_12_167 b_12 NI_12 NS_167 0 5.9984035779289078e-05
GC_12_168 b_12 NI_12 NS_168 0 -4.9318773507814958e-06
GC_12_169 b_12 NI_12 NS_169 0 -4.5492025749072695e-06
GC_12_170 b_12 NI_12 NS_170 0 -5.6348575872212258e-05
GC_12_171 b_12 NI_12 NS_171 0 -2.2571981593789796e-05
GC_12_172 b_12 NI_12 NS_172 0 -1.3235097065899173e-05
GC_12_173 b_12 NI_12 NS_173 0 6.7403410075434685e-07
GC_12_174 b_12 NI_12 NS_174 0 -6.8468783604265267e-07
GC_12_175 b_12 NI_12 NS_175 0 3.8201625269177735e-07
GC_12_176 b_12 NI_12 NS_176 0 1.4911381095379559e-07
GC_12_177 b_12 NI_12 NS_177 0 1.7058240256611561e-10
GC_12_178 b_12 NI_12 NS_178 0 -7.6198341570427871e-11
GC_12_179 b_12 NI_12 NS_179 0 -7.2508428255258335e-11
GC_12_180 b_12 NI_12 NS_180 0 -4.3770158933499988e-10
GC_12_181 b_12 NI_12 NS_181 0 4.6469696041164896e-05
GC_12_182 b_12 NI_12 NS_182 0 9.2530535115958892e-05
GC_12_183 b_12 NI_12 NS_183 0 2.8969073342025043e-07
GC_12_184 b_12 NI_12 NS_184 0 8.4521963959025608e-09
GC_12_185 b_12 NI_12 NS_185 0 -3.9577516136166932e-05
GC_12_186 b_12 NI_12 NS_186 0 -8.5748798994784674e-05
GC_12_187 b_12 NI_12 NS_187 0 -2.2600756429827870e-04
GC_12_188 b_12 NI_12 NS_188 0 9.6587366064429083e-05
GC_12_189 b_12 NI_12 NS_189 0 2.8264086026050385e-04
GC_12_190 b_12 NI_12 NS_190 0 1.5421249338276957e-04
GC_12_191 b_12 NI_12 NS_191 0 -3.0568685852019504e-04
GC_12_192 b_12 NI_12 NS_192 0 -2.0974507162560186e-04
GC_12_193 b_12 NI_12 NS_193 0 1.8427774477804238e-04
GC_12_194 b_12 NI_12 NS_194 0 3.8931269033130184e-04
GC_12_195 b_12 NI_12 NS_195 0 -9.5460495411135669e-05
GC_12_196 b_12 NI_12 NS_196 0 -1.5686517377382306e-04
GC_12_197 b_12 NI_12 NS_197 0 2.3694874029948687e-04
GC_12_198 b_12 NI_12 NS_198 0 2.1574923630679989e-04
GC_12_199 b_12 NI_12 NS_199 0 -5.9308356948110699e-05
GC_12_200 b_12 NI_12 NS_200 0 -2.0763943791568499e-04
GC_12_201 b_12 NI_12 NS_201 0 -1.2603416363086593e-06
GC_12_202 b_12 NI_12 NS_202 0 2.1361740052453635e-04
GC_12_203 b_12 NI_12 NS_203 0 -2.2353604834155045e-06
GC_12_204 b_12 NI_12 NS_204 0 -4.6374170759594547e-08
GC_12_205 b_12 NI_12 NS_205 0 -4.0397125609299340e-07
GC_12_206 b_12 NI_12 NS_206 0 -4.3861915759674144e-07
GC_12_207 b_12 NI_12 NS_207 0 -7.4187305930108949e-10
GC_12_208 b_12 NI_12 NS_208 0 5.0958795430332655e-10
GC_12_209 b_12 NI_12 NS_209 0 1.5239076171078585e-10
GC_12_210 b_12 NI_12 NS_210 0 1.2350690274531419e-09
GC_12_211 b_12 NI_12 NS_211 0 1.1737144650656131e-04
GC_12_212 b_12 NI_12 NS_212 0 4.0259732652204767e-06
GC_12_213 b_12 NI_12 NS_213 0 -2.0970088888442288e-07
GC_12_214 b_12 NI_12 NS_214 0 -9.1846098791167391e-09
GC_12_215 b_12 NI_12 NS_215 0 5.0822812797729352e-05
GC_12_216 b_12 NI_12 NS_216 0 -1.6606067783781579e-06
GC_12_217 b_12 NI_12 NS_217 0 2.6862077367222788e-05
GC_12_218 b_12 NI_12 NS_218 0 -7.4538578238148812e-06
GC_12_219 b_12 NI_12 NS_219 0 2.3829669966672697e-05
GC_12_220 b_12 NI_12 NS_220 0 -2.6937137611487792e-04
GC_12_221 b_12 NI_12 NS_221 0 -2.9022335984535034e-04
GC_12_222 b_12 NI_12 NS_222 0 3.9958670689197653e-05
GC_12_223 b_12 NI_12 NS_223 0 -5.3672778474664171e-05
GC_12_224 b_12 NI_12 NS_224 0 2.1969145544024270e-04
GC_12_225 b_12 NI_12 NS_225 0 1.6888955702016226e-04
GC_12_226 b_12 NI_12 NS_226 0 -1.0703566534036999e-04
GC_12_227 b_12 NI_12 NS_227 0 -1.7982839582278640e-04
GC_12_228 b_12 NI_12 NS_228 0 5.9624845880933247e-05
GC_12_229 b_12 NI_12 NS_229 0 -4.9612694943604356e-05
GC_12_230 b_12 NI_12 NS_230 0 1.1944079417101660e-04
GC_12_231 b_12 NI_12 NS_231 0 1.4033724974236035e-04
GC_12_232 b_12 NI_12 NS_232 0 7.0104839800339260e-05
GC_12_233 b_12 NI_12 NS_233 0 1.2844110657407729e-07
GC_12_234 b_12 NI_12 NS_234 0 4.2771201635959814e-06
GC_12_235 b_12 NI_12 NS_235 0 -1.9736722833413943e-06
GC_12_236 b_12 NI_12 NS_236 0 1.1969800118007441e-07
GC_12_237 b_12 NI_12 NS_237 0 6.3201776309029797e-10
GC_12_238 b_12 NI_12 NS_238 0 -6.2610963007046651e-10
GC_12_239 b_12 NI_12 NS_239 0 -1.5199179183207162e-10
GC_12_240 b_12 NI_12 NS_240 0 -1.2381058098565530e-09
GC_12_241 b_12 NI_12 NS_241 0 1.3559941509461802e-03
GC_12_242 b_12 NI_12 NS_242 0 -1.2038862729302643e-03
GC_12_243 b_12 NI_12 NS_243 0 3.7357854952783150e-06
GC_12_244 b_12 NI_12 NS_244 0 2.8902026037361699e-07
GC_12_245 b_12 NI_12 NS_245 0 1.2297142232693784e-04
GC_12_246 b_12 NI_12 NS_246 0 8.9417630272397913e-04
GC_12_247 b_12 NI_12 NS_247 0 1.8425184615281983e-03
GC_12_248 b_12 NI_12 NS_248 0 -8.6745250080809834e-04
GC_12_249 b_12 NI_12 NS_249 0 -2.9665987303382200e-03
GC_12_250 b_12 NI_12 NS_250 0 -1.6486220355325187e-03
GC_12_251 b_12 NI_12 NS_251 0 2.2195000359709416e-03
GC_12_252 b_12 NI_12 NS_252 0 2.6689299056709128e-03
GC_12_253 b_12 NI_12 NS_253 0 -1.4401285771273558e-03
GC_12_254 b_12 NI_12 NS_254 0 -2.9129269837821986e-03
GC_12_255 b_12 NI_12 NS_255 0 1.0698835480941820e-03
GC_12_256 b_12 NI_12 NS_256 0 2.2566937062412601e-03
GC_12_257 b_12 NI_12 NS_257 0 -1.6275429676173799e-03
GC_12_258 b_12 NI_12 NS_258 0 -2.1363737859431508e-03
GC_12_259 b_12 NI_12 NS_259 0 4.2046390607123452e-04
GC_12_260 b_12 NI_12 NS_260 0 2.0118509072884392e-03
GC_12_261 b_12 NI_12 NS_261 0 2.1508474886420222e-04
GC_12_262 b_12 NI_12 NS_262 0 -2.1102705422550018e-03
GC_12_263 b_12 NI_12 NS_263 0 -4.3288629333587221e-06
GC_12_264 b_12 NI_12 NS_264 0 4.3527947280600229e-06
GC_12_265 b_12 NI_12 NS_265 0 -7.8948788982549123e-07
GC_12_266 b_12 NI_12 NS_266 0 -3.5249023825901023e-06
GC_12_267 b_12 NI_12 NS_267 0 -7.5479782457011023e-09
GC_12_268 b_12 NI_12 NS_268 0 2.2567554932532060e-08
GC_12_269 b_12 NI_12 NS_269 0 2.3359227881260581e-09
GC_12_270 b_12 NI_12 NS_270 0 1.5101868389263613e-09
GC_12_271 b_12 NI_12 NS_271 0 -5.4915841993804029e-04
GC_12_272 b_12 NI_12 NS_272 0 -2.9018837039708405e-03
GC_12_273 b_12 NI_12 NS_273 0 -6.1488955598807146e-06
GC_12_274 b_12 NI_12 NS_274 0 -3.8642052853342371e-07
GC_12_275 b_12 NI_12 NS_275 0 2.6865516591988749e-03
GC_12_276 b_12 NI_12 NS_276 0 -1.9871372582523960e-03
GC_12_277 b_12 NI_12 NS_277 0 -6.1989513832137371e-03
GC_12_278 b_12 NI_12 NS_278 0 1.7530828200673354e-03
GC_12_279 b_12 NI_12 NS_279 0 4.7648850850489262e-03
GC_12_280 b_12 NI_12 NS_280 0 -5.5284540635730838e-03
GC_12_281 b_12 NI_12 NS_281 0 -2.4815306869973078e-04
GC_12_282 b_12 NI_12 NS_282 0 7.2493849593844549e-03
GC_12_283 b_12 NI_12 NS_283 0 -6.3156107463805539e-03
GC_12_284 b_12 NI_12 NS_284 0 -5.0550429424194368e-03
GC_12_285 b_12 NI_12 NS_285 0 4.5025677458851365e-03
GC_12_286 b_12 NI_12 NS_286 0 -1.7116128853888251e-03
GC_12_287 b_12 NI_12 NS_287 0 -5.9125367198867740e-04
GC_12_288 b_12 NI_12 NS_288 0 6.9477907108374632e-03
GC_12_289 b_12 NI_12 NS_289 0 -3.4362430168487028e-03
GC_12_290 b_12 NI_12 NS_290 0 -3.6821810458767443e-03
GC_12_291 b_12 NI_12 NS_291 0 5.9242608986460384e-03
GC_12_292 b_12 NI_12 NS_292 0 3.9702052908979681e-04
GC_12_293 b_12 NI_12 NS_293 0 6.3746601294584852e-05
GC_12_294 b_12 NI_12 NS_294 0 8.4799176107691746e-06
GC_12_295 b_12 NI_12 NS_295 0 1.5085273241361649e-05
GC_12_296 b_12 NI_12 NS_296 0 3.9926660865902120e-05
GC_12_297 b_12 NI_12 NS_297 0 7.1120485370228101e-09
GC_12_298 b_12 NI_12 NS_298 0 -2.9352136411090670e-08
GC_12_299 b_12 NI_12 NS_299 0 -1.8854126658502616e-09
GC_12_300 b_12 NI_12 NS_300 0 -5.6020611491900840e-10
GC_12_301 b_12 NI_12 NS_301 0 -7.0424740245504505e-02
GC_12_302 b_12 NI_12 NS_302 0 2.4192835920643783e-02
GC_12_303 b_12 NI_12 NS_303 0 2.2092931687196073e-05
GC_12_304 b_12 NI_12 NS_304 0 5.3186599719384585e-06
GC_12_305 b_12 NI_12 NS_305 0 1.8108339189770336e-02
GC_12_306 b_12 NI_12 NS_306 0 2.7946335780839403e-02
GC_12_307 b_12 NI_12 NS_307 0 -1.9395057785608683e-02
GC_12_308 b_12 NI_12 NS_308 0 8.3724957898510428e-03
GC_12_309 b_12 NI_12 NS_309 0 -5.8925703625201447e-03
GC_12_310 b_12 NI_12 NS_310 0 -2.2930898492341471e-02
GC_12_311 b_12 NI_12 NS_311 0 2.6387190153252135e-02
GC_12_312 b_12 NI_12 NS_312 0 -1.4337491690516305e-02
GC_12_313 b_12 NI_12 NS_313 0 3.4164840552752068e-02
GC_12_314 b_12 NI_12 NS_314 0 5.2157738563536398e-03
GC_12_315 b_12 NI_12 NS_315 0 9.5147656313803106e-03
GC_12_316 b_12 NI_12 NS_316 0 1.4168220973352096e-02
GC_12_317 b_12 NI_12 NS_317 0 -1.2626417658053848e-02
GC_12_318 b_12 NI_12 NS_318 0 1.1356480837531208e-02
GC_12_319 b_12 NI_12 NS_319 0 -1.1978307887057942e-02
GC_12_320 b_12 NI_12 NS_320 0 -1.1686227988655791e-02
GC_12_321 b_12 NI_12 NS_321 0 1.9051200236770264e-02
GC_12_322 b_12 NI_12 NS_322 0 -2.5965294868455769e-02
GC_12_323 b_12 NI_12 NS_323 0 9.0694550458851652e-04
GC_12_324 b_12 NI_12 NS_324 0 -1.0849120016173143e-03
GC_12_325 b_12 NI_12 NS_325 0 6.2679752285026992e-04
GC_12_326 b_12 NI_12 NS_326 0 3.2175985677567327e-04
GC_12_327 b_12 NI_12 NS_327 0 9.0179353486724931e-08
GC_12_328 b_12 NI_12 NS_328 0 4.0614945231655674e-07
GC_12_329 b_12 NI_12 NS_329 0 -9.1805828425955902e-09
GC_12_330 b_12 NI_12 NS_330 0 -1.8631084947918697e-08
GC_12_331 b_12 NI_12 NS_331 0 1.2526109539007602e-01
GC_12_332 b_12 NI_12 NS_332 0 -9.7551767127499293e-03
GC_12_333 b_12 NI_12 NS_333 0 -2.1879130952243561e-05
GC_12_334 b_12 NI_12 NS_334 0 -3.7984595388708944e-06
GC_12_335 b_12 NI_12 NS_335 0 -8.0420617900947566e-03
GC_12_336 b_12 NI_12 NS_336 0 6.5371441387692883e-04
GC_12_337 b_12 NI_12 NS_337 0 -1.9771768576952735e-03
GC_12_338 b_12 NI_12 NS_338 0 1.0157035349988105e-04
GC_12_339 b_12 NI_12 NS_339 0 -1.2487318678050911e-02
GC_12_340 b_12 NI_12 NS_340 0 8.2382561606138445e-03
GC_12_341 b_12 NI_12 NS_341 0 -1.0111831129700337e-02
GC_12_342 b_12 NI_12 NS_342 0 -5.9611104333092974e-04
GC_12_343 b_12 NI_12 NS_343 0 -3.4891067426213356e-03
GC_12_344 b_12 NI_12 NS_344 0 1.6807114589681548e-02
GC_12_345 b_12 NI_12 NS_345 0 -7.7156937405831972e-03
GC_12_346 b_12 NI_12 NS_346 0 1.3269795962382851e-02
GC_12_347 b_12 NI_12 NS_347 0 -3.8876506552717300e-03
GC_12_348 b_12 NI_12 NS_348 0 6.8943368294903124e-03
GC_12_349 b_12 NI_12 NS_349 0 -2.7117305920497966e-03
GC_12_350 b_12 NI_12 NS_350 0 1.2199574043009030e-02
GC_12_351 b_12 NI_12 NS_351 0 -2.2742235751446176e-02
GC_12_352 b_12 NI_12 NS_352 0 5.9617076729823922e-03
GC_12_353 b_12 NI_12 NS_353 0 -8.4148616670020053e-04
GC_12_354 b_12 NI_12 NS_354 0 8.1300281436196377e-04
GC_12_355 b_12 NI_12 NS_355 0 -5.1564586368886675e-04
GC_12_356 b_12 NI_12 NS_356 0 -4.3052022749989180e-04
GC_12_357 b_12 NI_12 NS_357 0 -5.9275351095744286e-08
GC_12_358 b_12 NI_12 NS_358 0 -1.8756503205184261e-07
GC_12_359 b_12 NI_12 NS_359 0 -3.3579624240905614e-09
GC_12_360 b_12 NI_12 NS_360 0 5.3365700592516714e-09
GD_12_1 b_12 NI_12 NA_1 0 2.7280705906702623e-06
GD_12_2 b_12 NI_12 NA_2 0 5.1394394510151648e-06
GD_12_3 b_12 NI_12 NA_3 0 7.7453323057923730e-06
GD_12_4 b_12 NI_12 NA_4 0 -1.6971831044382806e-06
GD_12_5 b_12 NI_12 NA_5 0 8.6158350037034962e-06
GD_12_6 b_12 NI_12 NA_6 0 3.8174510754971888e-06
GD_12_7 b_12 NI_12 NA_7 0 -6.0834572685209361e-05
GD_12_8 b_12 NI_12 NA_8 0 1.7232177007331942e-04
GD_12_9 b_12 NI_12 NA_9 0 -9.1321501767997800e-05
GD_12_10 b_12 NI_12 NA_10 0 1.6053724364173544e-02
GD_12_11 b_12 NI_12 NA_11 0 -1.0827121564889004e-02
GD_12_12 b_12 NI_12 NA_12 0 -4.0049979026644353e-02
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 7.8204801849513412e+00
GS_1_1 0 NS_1 NA_1 0 7.3338024411935532e-01
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 2.1257837644909412e+01
GS_2_1 0 NS_2 NA_1 0 7.3338024411935532e-01
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 8.8189725508130692e+01
GS_3_1 0 NS_3 NA_1 0 7.3338024411935532e-01
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 4.7583942880173470e+02
GS_4_1 0 NS_4 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 2.4147519902582747e+01
RS_6 NS_6 0 2.4147519902582744e+01
GL_5 0 NS_5 NS_6 0 3.6063062163307147e-01
GL_6 0 NS_6 NS_5 0 -3.6063062163307147e-01
GS_5_1 0 NS_5 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 1.8217846373726687e+01
RS_8 NS_8 0 1.8217846373726687e+01
GL_7 0 NS_7 NS_8 0 3.0904106785287211e-01
GL_8 0 NS_8 NS_7 0 -3.0904106785287211e-01
GS_7_1 0 NS_7 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 1.6355478720039709e+01
RS_10 NS_10 0 1.6355478720039706e+01
GL_9 0 NS_9 NS_10 0 2.6900015870612737e-01
GL_10 0 NS_10 NS_9 0 -2.6900015870612737e-01
GS_9_1 0 NS_9 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 1.6509546628040873e+01
RS_12 NS_12 0 1.6509546628040873e+01
GL_11 0 NS_11 NS_12 0 2.2664475020429389e-01
GL_12 0 NS_12 NS_11 0 -2.2664475020429389e-01
GS_11_1 0 NS_11 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 1.6536240554804539e+01
RS_14 NS_14 0 1.6536240554804539e+01
GL_13 0 NS_13 NS_14 0 1.9441023356946371e-01
GL_14 0 NS_14 NS_13 0 -1.9441023356946371e-01
GS_13_1 0 NS_13 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 1.7105682444637345e+01
RS_16 NS_16 0 1.7105682444637345e+01
GL_15 0 NS_15 NS_16 0 1.6030676643748842e-01
GL_16 0 NS_16 NS_15 0 -1.6030676643748842e-01
GS_15_1 0 NS_15 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 1.7548692376233411e+01
RS_18 NS_18 0 1.7548692376233408e+01
GL_17 0 NS_17 NS_18 0 1.2418335580210092e-01
GL_18 0 NS_18 NS_17 0 -1.2418335580210092e-01
GS_17_1 0 NS_17 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 1.9080711385242900e+01
RS_20 NS_20 0 1.9080711385242903e+01
GL_19 0 NS_19 NS_20 0 9.0245963773871965e-02
GL_20 0 NS_20 NS_19 0 -9.0245963773871965e-02
GS_19_1 0 NS_19 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 1.9398886873467703e+01
RS_22 NS_22 0 1.9398886873467703e+01
GL_21 0 NS_21 NS_22 0 5.0255945091433295e-02
GL_22 0 NS_22 NS_21 0 -5.0255945091433295e-02
GS_21_1 0 NS_21 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 4.6104523042200498e+01
RS_24 NS_24 0 4.6104523042200498e+01
GL_23 0 NS_23 NS_24 0 2.6612229878385272e-02
GL_24 0 NS_24 NS_23 0 -2.6612229878385272e-02
GS_23_1 0 NS_23 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 5.0459916965113045e+01
RS_26 NS_26 0 5.0459916965113038e+01
GL_25 0 NS_25 NS_26 0 3.3991465082001564e-02
GL_26 0 NS_26 NS_25 0 -3.3991465082001564e-02
GS_25_1 0 NS_25 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 1.4140189915393535e+03
RS_28 NS_28 0 1.4140189915393535e+03
GL_27 0 NS_27 NS_28 0 1.8736958636705965e-03
GL_28 0 NS_28 NS_27 0 -1.8736958636705965e-03
GS_27_1 0 NS_27 NA_1 0 7.3338024411935532e-01
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 9.6884954140421924e+03
RS_30 NS_30 0 9.6884954140421905e+03
GL_29 0 NS_29 NS_30 0 7.9053621147275857e-05
GL_30 0 NS_30 NS_29 0 -7.9053621147275857e-05
GS_29_1 0 NS_29 NA_1 0 7.3338024411935532e-01
*
* Real pole n. 31
CS_31 NS_31 0 9.9999999999999998e-13
RS_31 NS_31 0 7.8204801849513412e+00
GS_31_2 0 NS_31 NA_2 0 7.3338024411935532e-01
*
* Real pole n. 32
CS_32 NS_32 0 9.9999999999999998e-13
RS_32 NS_32 0 2.1257837644909412e+01
GS_32_2 0 NS_32 NA_2 0 7.3338024411935532e-01
*
* Real pole n. 33
CS_33 NS_33 0 9.9999999999999998e-13
RS_33 NS_33 0 8.8189725508130692e+01
GS_33_2 0 NS_33 NA_2 0 7.3338024411935532e-01
*
* Real pole n. 34
CS_34 NS_34 0 9.9999999999999998e-13
RS_34 NS_34 0 4.7583942880173470e+02
GS_34_2 0 NS_34 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 2.4147519902582747e+01
RS_36 NS_36 0 2.4147519902582744e+01
GL_35 0 NS_35 NS_36 0 3.6063062163307147e-01
GL_36 0 NS_36 NS_35 0 -3.6063062163307147e-01
GS_35_2 0 NS_35 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 1.8217846373726687e+01
RS_38 NS_38 0 1.8217846373726687e+01
GL_37 0 NS_37 NS_38 0 3.0904106785287211e-01
GL_38 0 NS_38 NS_37 0 -3.0904106785287211e-01
GS_37_2 0 NS_37 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 1.6355478720039709e+01
RS_40 NS_40 0 1.6355478720039706e+01
GL_39 0 NS_39 NS_40 0 2.6900015870612737e-01
GL_40 0 NS_40 NS_39 0 -2.6900015870612737e-01
GS_39_2 0 NS_39 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 1.6509546628040873e+01
RS_42 NS_42 0 1.6509546628040873e+01
GL_41 0 NS_41 NS_42 0 2.2664475020429389e-01
GL_42 0 NS_42 NS_41 0 -2.2664475020429389e-01
GS_41_2 0 NS_41 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 1.6536240554804539e+01
RS_44 NS_44 0 1.6536240554804539e+01
GL_43 0 NS_43 NS_44 0 1.9441023356946371e-01
GL_44 0 NS_44 NS_43 0 -1.9441023356946371e-01
GS_43_2 0 NS_43 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 1.7105682444637345e+01
RS_46 NS_46 0 1.7105682444637345e+01
GL_45 0 NS_45 NS_46 0 1.6030676643748842e-01
GL_46 0 NS_46 NS_45 0 -1.6030676643748842e-01
GS_45_2 0 NS_45 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 1.7548692376233411e+01
RS_48 NS_48 0 1.7548692376233408e+01
GL_47 0 NS_47 NS_48 0 1.2418335580210092e-01
GL_48 0 NS_48 NS_47 0 -1.2418335580210092e-01
GS_47_2 0 NS_47 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 1.9080711385242900e+01
RS_50 NS_50 0 1.9080711385242903e+01
GL_49 0 NS_49 NS_50 0 9.0245963773871965e-02
GL_50 0 NS_50 NS_49 0 -9.0245963773871965e-02
GS_49_2 0 NS_49 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 1.9398886873467703e+01
RS_52 NS_52 0 1.9398886873467703e+01
GL_51 0 NS_51 NS_52 0 5.0255945091433295e-02
GL_52 0 NS_52 NS_51 0 -5.0255945091433295e-02
GS_51_2 0 NS_51 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 4.6104523042200498e+01
RS_54 NS_54 0 4.6104523042200498e+01
GL_53 0 NS_53 NS_54 0 2.6612229878385272e-02
GL_54 0 NS_54 NS_53 0 -2.6612229878385272e-02
GS_53_2 0 NS_53 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 5.0459916965113045e+01
RS_56 NS_56 0 5.0459916965113038e+01
GL_55 0 NS_55 NS_56 0 3.3991465082001564e-02
GL_56 0 NS_56 NS_55 0 -3.3991465082001564e-02
GS_55_2 0 NS_55 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 1.4140189915393535e+03
RS_58 NS_58 0 1.4140189915393535e+03
GL_57 0 NS_57 NS_58 0 1.8736958636705965e-03
GL_58 0 NS_58 NS_57 0 -1.8736958636705965e-03
GS_57_2 0 NS_57 NA_2 0 7.3338024411935532e-01
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 9.6884954140421924e+03
RS_60 NS_60 0 9.6884954140421905e+03
GL_59 0 NS_59 NS_60 0 7.9053621147275857e-05
GL_60 0 NS_60 NS_59 0 -7.9053621147275857e-05
GS_59_2 0 NS_59 NA_2 0 7.3338024411935532e-01
*
* Real pole n. 61
CS_61 NS_61 0 9.9999999999999998e-13
RS_61 NS_61 0 7.8204801849513412e+00
GS_61_3 0 NS_61 NA_3 0 7.3338024411935532e-01
*
* Real pole n. 62
CS_62 NS_62 0 9.9999999999999998e-13
RS_62 NS_62 0 2.1257837644909412e+01
GS_62_3 0 NS_62 NA_3 0 7.3338024411935532e-01
*
* Real pole n. 63
CS_63 NS_63 0 9.9999999999999998e-13
RS_63 NS_63 0 8.8189725508130692e+01
GS_63_3 0 NS_63 NA_3 0 7.3338024411935532e-01
*
* Real pole n. 64
CS_64 NS_64 0 9.9999999999999998e-13
RS_64 NS_64 0 4.7583942880173470e+02
GS_64_3 0 NS_64 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 2.4147519902582747e+01
RS_66 NS_66 0 2.4147519902582744e+01
GL_65 0 NS_65 NS_66 0 3.6063062163307147e-01
GL_66 0 NS_66 NS_65 0 -3.6063062163307147e-01
GS_65_3 0 NS_65 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 1.8217846373726687e+01
RS_68 NS_68 0 1.8217846373726687e+01
GL_67 0 NS_67 NS_68 0 3.0904106785287211e-01
GL_68 0 NS_68 NS_67 0 -3.0904106785287211e-01
GS_67_3 0 NS_67 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 1.6355478720039709e+01
RS_70 NS_70 0 1.6355478720039706e+01
GL_69 0 NS_69 NS_70 0 2.6900015870612737e-01
GL_70 0 NS_70 NS_69 0 -2.6900015870612737e-01
GS_69_3 0 NS_69 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 1.6509546628040873e+01
RS_72 NS_72 0 1.6509546628040873e+01
GL_71 0 NS_71 NS_72 0 2.2664475020429389e-01
GL_72 0 NS_72 NS_71 0 -2.2664475020429389e-01
GS_71_3 0 NS_71 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 1.6536240554804539e+01
RS_74 NS_74 0 1.6536240554804539e+01
GL_73 0 NS_73 NS_74 0 1.9441023356946371e-01
GL_74 0 NS_74 NS_73 0 -1.9441023356946371e-01
GS_73_3 0 NS_73 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 1.7105682444637345e+01
RS_76 NS_76 0 1.7105682444637345e+01
GL_75 0 NS_75 NS_76 0 1.6030676643748842e-01
GL_76 0 NS_76 NS_75 0 -1.6030676643748842e-01
GS_75_3 0 NS_75 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 1.7548692376233411e+01
RS_78 NS_78 0 1.7548692376233408e+01
GL_77 0 NS_77 NS_78 0 1.2418335580210092e-01
GL_78 0 NS_78 NS_77 0 -1.2418335580210092e-01
GS_77_3 0 NS_77 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 1.9080711385242900e+01
RS_80 NS_80 0 1.9080711385242903e+01
GL_79 0 NS_79 NS_80 0 9.0245963773871965e-02
GL_80 0 NS_80 NS_79 0 -9.0245963773871965e-02
GS_79_3 0 NS_79 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 1.9398886873467703e+01
RS_82 NS_82 0 1.9398886873467703e+01
GL_81 0 NS_81 NS_82 0 5.0255945091433295e-02
GL_82 0 NS_82 NS_81 0 -5.0255945091433295e-02
GS_81_3 0 NS_81 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 4.6104523042200498e+01
RS_84 NS_84 0 4.6104523042200498e+01
GL_83 0 NS_83 NS_84 0 2.6612229878385272e-02
GL_84 0 NS_84 NS_83 0 -2.6612229878385272e-02
GS_83_3 0 NS_83 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 5.0459916965113045e+01
RS_86 NS_86 0 5.0459916965113038e+01
GL_85 0 NS_85 NS_86 0 3.3991465082001564e-02
GL_86 0 NS_86 NS_85 0 -3.3991465082001564e-02
GS_85_3 0 NS_85 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 1.4140189915393535e+03
RS_88 NS_88 0 1.4140189915393535e+03
GL_87 0 NS_87 NS_88 0 1.8736958636705965e-03
GL_88 0 NS_88 NS_87 0 -1.8736958636705965e-03
GS_87_3 0 NS_87 NA_3 0 7.3338024411935532e-01
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 9.6884954140421924e+03
RS_90 NS_90 0 9.6884954140421905e+03
GL_89 0 NS_89 NS_90 0 7.9053621147275857e-05
GL_90 0 NS_90 NS_89 0 -7.9053621147275857e-05
GS_89_3 0 NS_89 NA_3 0 7.3338024411935532e-01
*
* Real pole n. 91
CS_91 NS_91 0 9.9999999999999998e-13
RS_91 NS_91 0 7.8204801849513412e+00
GS_91_4 0 NS_91 NA_4 0 7.3338024411935532e-01
*
* Real pole n. 92
CS_92 NS_92 0 9.9999999999999998e-13
RS_92 NS_92 0 2.1257837644909412e+01
GS_92_4 0 NS_92 NA_4 0 7.3338024411935532e-01
*
* Real pole n. 93
CS_93 NS_93 0 9.9999999999999998e-13
RS_93 NS_93 0 8.8189725508130692e+01
GS_93_4 0 NS_93 NA_4 0 7.3338024411935532e-01
*
* Real pole n. 94
CS_94 NS_94 0 9.9999999999999998e-13
RS_94 NS_94 0 4.7583942880173470e+02
GS_94_4 0 NS_94 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 2.4147519902582747e+01
RS_96 NS_96 0 2.4147519902582744e+01
GL_95 0 NS_95 NS_96 0 3.6063062163307147e-01
GL_96 0 NS_96 NS_95 0 -3.6063062163307147e-01
GS_95_4 0 NS_95 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 1.8217846373726687e+01
RS_98 NS_98 0 1.8217846373726687e+01
GL_97 0 NS_97 NS_98 0 3.0904106785287211e-01
GL_98 0 NS_98 NS_97 0 -3.0904106785287211e-01
GS_97_4 0 NS_97 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 1.6355478720039709e+01
RS_100 NS_100 0 1.6355478720039706e+01
GL_99 0 NS_99 NS_100 0 2.6900015870612737e-01
GL_100 0 NS_100 NS_99 0 -2.6900015870612737e-01
GS_99_4 0 NS_99 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 1.6509546628040873e+01
RS_102 NS_102 0 1.6509546628040873e+01
GL_101 0 NS_101 NS_102 0 2.2664475020429389e-01
GL_102 0 NS_102 NS_101 0 -2.2664475020429389e-01
GS_101_4 0 NS_101 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 1.6536240554804539e+01
RS_104 NS_104 0 1.6536240554804539e+01
GL_103 0 NS_103 NS_104 0 1.9441023356946371e-01
GL_104 0 NS_104 NS_103 0 -1.9441023356946371e-01
GS_103_4 0 NS_103 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 1.7105682444637345e+01
RS_106 NS_106 0 1.7105682444637345e+01
GL_105 0 NS_105 NS_106 0 1.6030676643748842e-01
GL_106 0 NS_106 NS_105 0 -1.6030676643748842e-01
GS_105_4 0 NS_105 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 1.7548692376233411e+01
RS_108 NS_108 0 1.7548692376233408e+01
GL_107 0 NS_107 NS_108 0 1.2418335580210092e-01
GL_108 0 NS_108 NS_107 0 -1.2418335580210092e-01
GS_107_4 0 NS_107 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 1.9080711385242900e+01
RS_110 NS_110 0 1.9080711385242903e+01
GL_109 0 NS_109 NS_110 0 9.0245963773871965e-02
GL_110 0 NS_110 NS_109 0 -9.0245963773871965e-02
GS_109_4 0 NS_109 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 1.9398886873467703e+01
RS_112 NS_112 0 1.9398886873467703e+01
GL_111 0 NS_111 NS_112 0 5.0255945091433295e-02
GL_112 0 NS_112 NS_111 0 -5.0255945091433295e-02
GS_111_4 0 NS_111 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 4.6104523042200498e+01
RS_114 NS_114 0 4.6104523042200498e+01
GL_113 0 NS_113 NS_114 0 2.6612229878385272e-02
GL_114 0 NS_114 NS_113 0 -2.6612229878385272e-02
GS_113_4 0 NS_113 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 5.0459916965113045e+01
RS_116 NS_116 0 5.0459916965113038e+01
GL_115 0 NS_115 NS_116 0 3.3991465082001564e-02
GL_116 0 NS_116 NS_115 0 -3.3991465082001564e-02
GS_115_4 0 NS_115 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 1.4140189915393535e+03
RS_118 NS_118 0 1.4140189915393535e+03
GL_117 0 NS_117 NS_118 0 1.8736958636705965e-03
GL_118 0 NS_118 NS_117 0 -1.8736958636705965e-03
GS_117_4 0 NS_117 NA_4 0 7.3338024411935532e-01
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 9.6884954140421924e+03
RS_120 NS_120 0 9.6884954140421905e+03
GL_119 0 NS_119 NS_120 0 7.9053621147275857e-05
GL_120 0 NS_120 NS_119 0 -7.9053621147275857e-05
GS_119_4 0 NS_119 NA_4 0 7.3338024411935532e-01
*
* Real pole n. 121
CS_121 NS_121 0 9.9999999999999998e-13
RS_121 NS_121 0 7.8204801849513412e+00
GS_121_5 0 NS_121 NA_5 0 7.3338024411935532e-01
*
* Real pole n. 122
CS_122 NS_122 0 9.9999999999999998e-13
RS_122 NS_122 0 2.1257837644909412e+01
GS_122_5 0 NS_122 NA_5 0 7.3338024411935532e-01
*
* Real pole n. 123
CS_123 NS_123 0 9.9999999999999998e-13
RS_123 NS_123 0 8.8189725508130692e+01
GS_123_5 0 NS_123 NA_5 0 7.3338024411935532e-01
*
* Real pole n. 124
CS_124 NS_124 0 9.9999999999999998e-13
RS_124 NS_124 0 4.7583942880173470e+02
GS_124_5 0 NS_124 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 2.4147519902582747e+01
RS_126 NS_126 0 2.4147519902582744e+01
GL_125 0 NS_125 NS_126 0 3.6063062163307147e-01
GL_126 0 NS_126 NS_125 0 -3.6063062163307147e-01
GS_125_5 0 NS_125 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 1.8217846373726687e+01
RS_128 NS_128 0 1.8217846373726687e+01
GL_127 0 NS_127 NS_128 0 3.0904106785287211e-01
GL_128 0 NS_128 NS_127 0 -3.0904106785287211e-01
GS_127_5 0 NS_127 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 1.6355478720039709e+01
RS_130 NS_130 0 1.6355478720039706e+01
GL_129 0 NS_129 NS_130 0 2.6900015870612737e-01
GL_130 0 NS_130 NS_129 0 -2.6900015870612737e-01
GS_129_5 0 NS_129 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 1.6509546628040873e+01
RS_132 NS_132 0 1.6509546628040873e+01
GL_131 0 NS_131 NS_132 0 2.2664475020429389e-01
GL_132 0 NS_132 NS_131 0 -2.2664475020429389e-01
GS_131_5 0 NS_131 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 133/134
CS_133 NS_133 0 9.9999999999999998e-13
CS_134 NS_134 0 9.9999999999999998e-13
RS_133 NS_133 0 1.6536240554804539e+01
RS_134 NS_134 0 1.6536240554804539e+01
GL_133 0 NS_133 NS_134 0 1.9441023356946371e-01
GL_134 0 NS_134 NS_133 0 -1.9441023356946371e-01
GS_133_5 0 NS_133 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 1.7105682444637345e+01
RS_136 NS_136 0 1.7105682444637345e+01
GL_135 0 NS_135 NS_136 0 1.6030676643748842e-01
GL_136 0 NS_136 NS_135 0 -1.6030676643748842e-01
GS_135_5 0 NS_135 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 1.7548692376233411e+01
RS_138 NS_138 0 1.7548692376233408e+01
GL_137 0 NS_137 NS_138 0 1.2418335580210092e-01
GL_138 0 NS_138 NS_137 0 -1.2418335580210092e-01
GS_137_5 0 NS_137 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 1.9080711385242900e+01
RS_140 NS_140 0 1.9080711385242903e+01
GL_139 0 NS_139 NS_140 0 9.0245963773871965e-02
GL_140 0 NS_140 NS_139 0 -9.0245963773871965e-02
GS_139_5 0 NS_139 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 1.9398886873467703e+01
RS_142 NS_142 0 1.9398886873467703e+01
GL_141 0 NS_141 NS_142 0 5.0255945091433295e-02
GL_142 0 NS_142 NS_141 0 -5.0255945091433295e-02
GS_141_5 0 NS_141 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 4.6104523042200498e+01
RS_144 NS_144 0 4.6104523042200498e+01
GL_143 0 NS_143 NS_144 0 2.6612229878385272e-02
GL_144 0 NS_144 NS_143 0 -2.6612229878385272e-02
GS_143_5 0 NS_143 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 5.0459916965113045e+01
RS_146 NS_146 0 5.0459916965113038e+01
GL_145 0 NS_145 NS_146 0 3.3991465082001564e-02
GL_146 0 NS_146 NS_145 0 -3.3991465082001564e-02
GS_145_5 0 NS_145 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 1.4140189915393535e+03
RS_148 NS_148 0 1.4140189915393535e+03
GL_147 0 NS_147 NS_148 0 1.8736958636705965e-03
GL_148 0 NS_148 NS_147 0 -1.8736958636705965e-03
GS_147_5 0 NS_147 NA_5 0 7.3338024411935532e-01
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 9.6884954140421924e+03
RS_150 NS_150 0 9.6884954140421905e+03
GL_149 0 NS_149 NS_150 0 7.9053621147275857e-05
GL_150 0 NS_150 NS_149 0 -7.9053621147275857e-05
GS_149_5 0 NS_149 NA_5 0 7.3338024411935532e-01
*
* Real pole n. 151
CS_151 NS_151 0 9.9999999999999998e-13
RS_151 NS_151 0 7.8204801849513412e+00
GS_151_6 0 NS_151 NA_6 0 7.3338024411935532e-01
*
* Real pole n. 152
CS_152 NS_152 0 9.9999999999999998e-13
RS_152 NS_152 0 2.1257837644909412e+01
GS_152_6 0 NS_152 NA_6 0 7.3338024411935532e-01
*
* Real pole n. 153
CS_153 NS_153 0 9.9999999999999998e-13
RS_153 NS_153 0 8.8189725508130692e+01
GS_153_6 0 NS_153 NA_6 0 7.3338024411935532e-01
*
* Real pole n. 154
CS_154 NS_154 0 9.9999999999999998e-13
RS_154 NS_154 0 4.7583942880173470e+02
GS_154_6 0 NS_154 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 2.4147519902582747e+01
RS_156 NS_156 0 2.4147519902582744e+01
GL_155 0 NS_155 NS_156 0 3.6063062163307147e-01
GL_156 0 NS_156 NS_155 0 -3.6063062163307147e-01
GS_155_6 0 NS_155 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 1.8217846373726687e+01
RS_158 NS_158 0 1.8217846373726687e+01
GL_157 0 NS_157 NS_158 0 3.0904106785287211e-01
GL_158 0 NS_158 NS_157 0 -3.0904106785287211e-01
GS_157_6 0 NS_157 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 1.6355478720039709e+01
RS_160 NS_160 0 1.6355478720039706e+01
GL_159 0 NS_159 NS_160 0 2.6900015870612737e-01
GL_160 0 NS_160 NS_159 0 -2.6900015870612737e-01
GS_159_6 0 NS_159 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 1.6509546628040873e+01
RS_162 NS_162 0 1.6509546628040873e+01
GL_161 0 NS_161 NS_162 0 2.2664475020429389e-01
GL_162 0 NS_162 NS_161 0 -2.2664475020429389e-01
GS_161_6 0 NS_161 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 163/164
CS_163 NS_163 0 9.9999999999999998e-13
CS_164 NS_164 0 9.9999999999999998e-13
RS_163 NS_163 0 1.6536240554804539e+01
RS_164 NS_164 0 1.6536240554804539e+01
GL_163 0 NS_163 NS_164 0 1.9441023356946371e-01
GL_164 0 NS_164 NS_163 0 -1.9441023356946371e-01
GS_163_6 0 NS_163 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 1.7105682444637345e+01
RS_166 NS_166 0 1.7105682444637345e+01
GL_165 0 NS_165 NS_166 0 1.6030676643748842e-01
GL_166 0 NS_166 NS_165 0 -1.6030676643748842e-01
GS_165_6 0 NS_165 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 1.7548692376233411e+01
RS_168 NS_168 0 1.7548692376233408e+01
GL_167 0 NS_167 NS_168 0 1.2418335580210092e-01
GL_168 0 NS_168 NS_167 0 -1.2418335580210092e-01
GS_167_6 0 NS_167 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 1.9080711385242900e+01
RS_170 NS_170 0 1.9080711385242903e+01
GL_169 0 NS_169 NS_170 0 9.0245963773871965e-02
GL_170 0 NS_170 NS_169 0 -9.0245963773871965e-02
GS_169_6 0 NS_169 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 1.9398886873467703e+01
RS_172 NS_172 0 1.9398886873467703e+01
GL_171 0 NS_171 NS_172 0 5.0255945091433295e-02
GL_172 0 NS_172 NS_171 0 -5.0255945091433295e-02
GS_171_6 0 NS_171 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 4.6104523042200498e+01
RS_174 NS_174 0 4.6104523042200498e+01
GL_173 0 NS_173 NS_174 0 2.6612229878385272e-02
GL_174 0 NS_174 NS_173 0 -2.6612229878385272e-02
GS_173_6 0 NS_173 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 5.0459916965113045e+01
RS_176 NS_176 0 5.0459916965113038e+01
GL_175 0 NS_175 NS_176 0 3.3991465082001564e-02
GL_176 0 NS_176 NS_175 0 -3.3991465082001564e-02
GS_175_6 0 NS_175 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 1.4140189915393535e+03
RS_178 NS_178 0 1.4140189915393535e+03
GL_177 0 NS_177 NS_178 0 1.8736958636705965e-03
GL_178 0 NS_178 NS_177 0 -1.8736958636705965e-03
GS_177_6 0 NS_177 NA_6 0 7.3338024411935532e-01
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 9.6884954140421924e+03
RS_180 NS_180 0 9.6884954140421905e+03
GL_179 0 NS_179 NS_180 0 7.9053621147275857e-05
GL_180 0 NS_180 NS_179 0 -7.9053621147275857e-05
GS_179_6 0 NS_179 NA_6 0 7.3338024411935532e-01
*
* Real pole n. 181
CS_181 NS_181 0 9.9999999999999998e-13
RS_181 NS_181 0 7.8204801849513412e+00
GS_181_7 0 NS_181 NA_7 0 7.3338024411935532e-01
*
* Real pole n. 182
CS_182 NS_182 0 9.9999999999999998e-13
RS_182 NS_182 0 2.1257837644909412e+01
GS_182_7 0 NS_182 NA_7 0 7.3338024411935532e-01
*
* Real pole n. 183
CS_183 NS_183 0 9.9999999999999998e-13
RS_183 NS_183 0 8.8189725508130692e+01
GS_183_7 0 NS_183 NA_7 0 7.3338024411935532e-01
*
* Real pole n. 184
CS_184 NS_184 0 9.9999999999999998e-13
RS_184 NS_184 0 4.7583942880173470e+02
GS_184_7 0 NS_184 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 2.4147519902582747e+01
RS_186 NS_186 0 2.4147519902582744e+01
GL_185 0 NS_185 NS_186 0 3.6063062163307147e-01
GL_186 0 NS_186 NS_185 0 -3.6063062163307147e-01
GS_185_7 0 NS_185 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 1.8217846373726687e+01
RS_188 NS_188 0 1.8217846373726687e+01
GL_187 0 NS_187 NS_188 0 3.0904106785287211e-01
GL_188 0 NS_188 NS_187 0 -3.0904106785287211e-01
GS_187_7 0 NS_187 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 1.6355478720039709e+01
RS_190 NS_190 0 1.6355478720039706e+01
GL_189 0 NS_189 NS_190 0 2.6900015870612737e-01
GL_190 0 NS_190 NS_189 0 -2.6900015870612737e-01
GS_189_7 0 NS_189 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 1.6509546628040873e+01
RS_192 NS_192 0 1.6509546628040873e+01
GL_191 0 NS_191 NS_192 0 2.2664475020429389e-01
GL_192 0 NS_192 NS_191 0 -2.2664475020429389e-01
GS_191_7 0 NS_191 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 1.6536240554804539e+01
RS_194 NS_194 0 1.6536240554804539e+01
GL_193 0 NS_193 NS_194 0 1.9441023356946371e-01
GL_194 0 NS_194 NS_193 0 -1.9441023356946371e-01
GS_193_7 0 NS_193 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 1.7105682444637345e+01
RS_196 NS_196 0 1.7105682444637345e+01
GL_195 0 NS_195 NS_196 0 1.6030676643748842e-01
GL_196 0 NS_196 NS_195 0 -1.6030676643748842e-01
GS_195_7 0 NS_195 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 1.7548692376233411e+01
RS_198 NS_198 0 1.7548692376233408e+01
GL_197 0 NS_197 NS_198 0 1.2418335580210092e-01
GL_198 0 NS_198 NS_197 0 -1.2418335580210092e-01
GS_197_7 0 NS_197 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 1.9080711385242900e+01
RS_200 NS_200 0 1.9080711385242903e+01
GL_199 0 NS_199 NS_200 0 9.0245963773871965e-02
GL_200 0 NS_200 NS_199 0 -9.0245963773871965e-02
GS_199_7 0 NS_199 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 201/202
CS_201 NS_201 0 9.9999999999999998e-13
CS_202 NS_202 0 9.9999999999999998e-13
RS_201 NS_201 0 1.9398886873467703e+01
RS_202 NS_202 0 1.9398886873467703e+01
GL_201 0 NS_201 NS_202 0 5.0255945091433295e-02
GL_202 0 NS_202 NS_201 0 -5.0255945091433295e-02
GS_201_7 0 NS_201 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 203/204
CS_203 NS_203 0 9.9999999999999998e-13
CS_204 NS_204 0 9.9999999999999998e-13
RS_203 NS_203 0 4.6104523042200498e+01
RS_204 NS_204 0 4.6104523042200498e+01
GL_203 0 NS_203 NS_204 0 2.6612229878385272e-02
GL_204 0 NS_204 NS_203 0 -2.6612229878385272e-02
GS_203_7 0 NS_203 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 5.0459916965113045e+01
RS_206 NS_206 0 5.0459916965113038e+01
GL_205 0 NS_205 NS_206 0 3.3991465082001564e-02
GL_206 0 NS_206 NS_205 0 -3.3991465082001564e-02
GS_205_7 0 NS_205 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 1.4140189915393535e+03
RS_208 NS_208 0 1.4140189915393535e+03
GL_207 0 NS_207 NS_208 0 1.8736958636705965e-03
GL_208 0 NS_208 NS_207 0 -1.8736958636705965e-03
GS_207_7 0 NS_207 NA_7 0 7.3338024411935532e-01
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 9.6884954140421924e+03
RS_210 NS_210 0 9.6884954140421905e+03
GL_209 0 NS_209 NS_210 0 7.9053621147275857e-05
GL_210 0 NS_210 NS_209 0 -7.9053621147275857e-05
GS_209_7 0 NS_209 NA_7 0 7.3338024411935532e-01
*
* Real pole n. 211
CS_211 NS_211 0 9.9999999999999998e-13
RS_211 NS_211 0 7.8204801849513412e+00
GS_211_8 0 NS_211 NA_8 0 7.3338024411935532e-01
*
* Real pole n. 212
CS_212 NS_212 0 9.9999999999999998e-13
RS_212 NS_212 0 2.1257837644909412e+01
GS_212_8 0 NS_212 NA_8 0 7.3338024411935532e-01
*
* Real pole n. 213
CS_213 NS_213 0 9.9999999999999998e-13
RS_213 NS_213 0 8.8189725508130692e+01
GS_213_8 0 NS_213 NA_8 0 7.3338024411935532e-01
*
* Real pole n. 214
CS_214 NS_214 0 9.9999999999999998e-13
RS_214 NS_214 0 4.7583942880173470e+02
GS_214_8 0 NS_214 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 2.4147519902582747e+01
RS_216 NS_216 0 2.4147519902582744e+01
GL_215 0 NS_215 NS_216 0 3.6063062163307147e-01
GL_216 0 NS_216 NS_215 0 -3.6063062163307147e-01
GS_215_8 0 NS_215 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 1.8217846373726687e+01
RS_218 NS_218 0 1.8217846373726687e+01
GL_217 0 NS_217 NS_218 0 3.0904106785287211e-01
GL_218 0 NS_218 NS_217 0 -3.0904106785287211e-01
GS_217_8 0 NS_217 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 1.6355478720039709e+01
RS_220 NS_220 0 1.6355478720039706e+01
GL_219 0 NS_219 NS_220 0 2.6900015870612737e-01
GL_220 0 NS_220 NS_219 0 -2.6900015870612737e-01
GS_219_8 0 NS_219 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 221/222
CS_221 NS_221 0 9.9999999999999998e-13
CS_222 NS_222 0 9.9999999999999998e-13
RS_221 NS_221 0 1.6509546628040873e+01
RS_222 NS_222 0 1.6509546628040873e+01
GL_221 0 NS_221 NS_222 0 2.2664475020429389e-01
GL_222 0 NS_222 NS_221 0 -2.2664475020429389e-01
GS_221_8 0 NS_221 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 223/224
CS_223 NS_223 0 9.9999999999999998e-13
CS_224 NS_224 0 9.9999999999999998e-13
RS_223 NS_223 0 1.6536240554804539e+01
RS_224 NS_224 0 1.6536240554804539e+01
GL_223 0 NS_223 NS_224 0 1.9441023356946371e-01
GL_224 0 NS_224 NS_223 0 -1.9441023356946371e-01
GS_223_8 0 NS_223 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 225/226
CS_225 NS_225 0 9.9999999999999998e-13
CS_226 NS_226 0 9.9999999999999998e-13
RS_225 NS_225 0 1.7105682444637345e+01
RS_226 NS_226 0 1.7105682444637345e+01
GL_225 0 NS_225 NS_226 0 1.6030676643748842e-01
GL_226 0 NS_226 NS_225 0 -1.6030676643748842e-01
GS_225_8 0 NS_225 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 1.7548692376233411e+01
RS_228 NS_228 0 1.7548692376233408e+01
GL_227 0 NS_227 NS_228 0 1.2418335580210092e-01
GL_228 0 NS_228 NS_227 0 -1.2418335580210092e-01
GS_227_8 0 NS_227 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 229/230
CS_229 NS_229 0 9.9999999999999998e-13
CS_230 NS_230 0 9.9999999999999998e-13
RS_229 NS_229 0 1.9080711385242900e+01
RS_230 NS_230 0 1.9080711385242903e+01
GL_229 0 NS_229 NS_230 0 9.0245963773871965e-02
GL_230 0 NS_230 NS_229 0 -9.0245963773871965e-02
GS_229_8 0 NS_229 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 1.9398886873467703e+01
RS_232 NS_232 0 1.9398886873467703e+01
GL_231 0 NS_231 NS_232 0 5.0255945091433295e-02
GL_232 0 NS_232 NS_231 0 -5.0255945091433295e-02
GS_231_8 0 NS_231 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 4.6104523042200498e+01
RS_234 NS_234 0 4.6104523042200498e+01
GL_233 0 NS_233 NS_234 0 2.6612229878385272e-02
GL_234 0 NS_234 NS_233 0 -2.6612229878385272e-02
GS_233_8 0 NS_233 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 5.0459916965113045e+01
RS_236 NS_236 0 5.0459916965113038e+01
GL_235 0 NS_235 NS_236 0 3.3991465082001564e-02
GL_236 0 NS_236 NS_235 0 -3.3991465082001564e-02
GS_235_8 0 NS_235 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 1.4140189915393535e+03
RS_238 NS_238 0 1.4140189915393535e+03
GL_237 0 NS_237 NS_238 0 1.8736958636705965e-03
GL_238 0 NS_238 NS_237 0 -1.8736958636705965e-03
GS_237_8 0 NS_237 NA_8 0 7.3338024411935532e-01
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 9.6884954140421924e+03
RS_240 NS_240 0 9.6884954140421905e+03
GL_239 0 NS_239 NS_240 0 7.9053621147275857e-05
GL_240 0 NS_240 NS_239 0 -7.9053621147275857e-05
GS_239_8 0 NS_239 NA_8 0 7.3338024411935532e-01
*
* Real pole n. 241
CS_241 NS_241 0 9.9999999999999998e-13
RS_241 NS_241 0 7.8204801849513412e+00
GS_241_9 0 NS_241 NA_9 0 7.3338024411935532e-01
*
* Real pole n. 242
CS_242 NS_242 0 9.9999999999999998e-13
RS_242 NS_242 0 2.1257837644909412e+01
GS_242_9 0 NS_242 NA_9 0 7.3338024411935532e-01
*
* Real pole n. 243
CS_243 NS_243 0 9.9999999999999998e-13
RS_243 NS_243 0 8.8189725508130692e+01
GS_243_9 0 NS_243 NA_9 0 7.3338024411935532e-01
*
* Real pole n. 244
CS_244 NS_244 0 9.9999999999999998e-13
RS_244 NS_244 0 4.7583942880173470e+02
GS_244_9 0 NS_244 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 245/246
CS_245 NS_245 0 9.9999999999999998e-13
CS_246 NS_246 0 9.9999999999999998e-13
RS_245 NS_245 0 2.4147519902582747e+01
RS_246 NS_246 0 2.4147519902582744e+01
GL_245 0 NS_245 NS_246 0 3.6063062163307147e-01
GL_246 0 NS_246 NS_245 0 -3.6063062163307147e-01
GS_245_9 0 NS_245 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 247/248
CS_247 NS_247 0 9.9999999999999998e-13
CS_248 NS_248 0 9.9999999999999998e-13
RS_247 NS_247 0 1.8217846373726687e+01
RS_248 NS_248 0 1.8217846373726687e+01
GL_247 0 NS_247 NS_248 0 3.0904106785287211e-01
GL_248 0 NS_248 NS_247 0 -3.0904106785287211e-01
GS_247_9 0 NS_247 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 249/250
CS_249 NS_249 0 9.9999999999999998e-13
CS_250 NS_250 0 9.9999999999999998e-13
RS_249 NS_249 0 1.6355478720039709e+01
RS_250 NS_250 0 1.6355478720039706e+01
GL_249 0 NS_249 NS_250 0 2.6900015870612737e-01
GL_250 0 NS_250 NS_249 0 -2.6900015870612737e-01
GS_249_9 0 NS_249 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 251/252
CS_251 NS_251 0 9.9999999999999998e-13
CS_252 NS_252 0 9.9999999999999998e-13
RS_251 NS_251 0 1.6509546628040873e+01
RS_252 NS_252 0 1.6509546628040873e+01
GL_251 0 NS_251 NS_252 0 2.2664475020429389e-01
GL_252 0 NS_252 NS_251 0 -2.2664475020429389e-01
GS_251_9 0 NS_251 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 253/254
CS_253 NS_253 0 9.9999999999999998e-13
CS_254 NS_254 0 9.9999999999999998e-13
RS_253 NS_253 0 1.6536240554804539e+01
RS_254 NS_254 0 1.6536240554804539e+01
GL_253 0 NS_253 NS_254 0 1.9441023356946371e-01
GL_254 0 NS_254 NS_253 0 -1.9441023356946371e-01
GS_253_9 0 NS_253 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 255/256
CS_255 NS_255 0 9.9999999999999998e-13
CS_256 NS_256 0 9.9999999999999998e-13
RS_255 NS_255 0 1.7105682444637345e+01
RS_256 NS_256 0 1.7105682444637345e+01
GL_255 0 NS_255 NS_256 0 1.6030676643748842e-01
GL_256 0 NS_256 NS_255 0 -1.6030676643748842e-01
GS_255_9 0 NS_255 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 257/258
CS_257 NS_257 0 9.9999999999999998e-13
CS_258 NS_258 0 9.9999999999999998e-13
RS_257 NS_257 0 1.7548692376233411e+01
RS_258 NS_258 0 1.7548692376233408e+01
GL_257 0 NS_257 NS_258 0 1.2418335580210092e-01
GL_258 0 NS_258 NS_257 0 -1.2418335580210092e-01
GS_257_9 0 NS_257 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 259/260
CS_259 NS_259 0 9.9999999999999998e-13
CS_260 NS_260 0 9.9999999999999998e-13
RS_259 NS_259 0 1.9080711385242900e+01
RS_260 NS_260 0 1.9080711385242903e+01
GL_259 0 NS_259 NS_260 0 9.0245963773871965e-02
GL_260 0 NS_260 NS_259 0 -9.0245963773871965e-02
GS_259_9 0 NS_259 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 261/262
CS_261 NS_261 0 9.9999999999999998e-13
CS_262 NS_262 0 9.9999999999999998e-13
RS_261 NS_261 0 1.9398886873467703e+01
RS_262 NS_262 0 1.9398886873467703e+01
GL_261 0 NS_261 NS_262 0 5.0255945091433295e-02
GL_262 0 NS_262 NS_261 0 -5.0255945091433295e-02
GS_261_9 0 NS_261 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 263/264
CS_263 NS_263 0 9.9999999999999998e-13
CS_264 NS_264 0 9.9999999999999998e-13
RS_263 NS_263 0 4.6104523042200498e+01
RS_264 NS_264 0 4.6104523042200498e+01
GL_263 0 NS_263 NS_264 0 2.6612229878385272e-02
GL_264 0 NS_264 NS_263 0 -2.6612229878385272e-02
GS_263_9 0 NS_263 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 265/266
CS_265 NS_265 0 9.9999999999999998e-13
CS_266 NS_266 0 9.9999999999999998e-13
RS_265 NS_265 0 5.0459916965113045e+01
RS_266 NS_266 0 5.0459916965113038e+01
GL_265 0 NS_265 NS_266 0 3.3991465082001564e-02
GL_266 0 NS_266 NS_265 0 -3.3991465082001564e-02
GS_265_9 0 NS_265 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 267/268
CS_267 NS_267 0 9.9999999999999998e-13
CS_268 NS_268 0 9.9999999999999998e-13
RS_267 NS_267 0 1.4140189915393535e+03
RS_268 NS_268 0 1.4140189915393535e+03
GL_267 0 NS_267 NS_268 0 1.8736958636705965e-03
GL_268 0 NS_268 NS_267 0 -1.8736958636705965e-03
GS_267_9 0 NS_267 NA_9 0 7.3338024411935532e-01
*
* Complex pair n. 269/270
CS_269 NS_269 0 9.9999999999999998e-13
CS_270 NS_270 0 9.9999999999999998e-13
RS_269 NS_269 0 9.6884954140421924e+03
RS_270 NS_270 0 9.6884954140421905e+03
GL_269 0 NS_269 NS_270 0 7.9053621147275857e-05
GL_270 0 NS_270 NS_269 0 -7.9053621147275857e-05
GS_269_9 0 NS_269 NA_9 0 7.3338024411935532e-01
*
* Real pole n. 271
CS_271 NS_271 0 9.9999999999999998e-13
RS_271 NS_271 0 7.8204801849513412e+00
GS_271_10 0 NS_271 NA_10 0 7.3338024411935532e-01
*
* Real pole n. 272
CS_272 NS_272 0 9.9999999999999998e-13
RS_272 NS_272 0 2.1257837644909412e+01
GS_272_10 0 NS_272 NA_10 0 7.3338024411935532e-01
*
* Real pole n. 273
CS_273 NS_273 0 9.9999999999999998e-13
RS_273 NS_273 0 8.8189725508130692e+01
GS_273_10 0 NS_273 NA_10 0 7.3338024411935532e-01
*
* Real pole n. 274
CS_274 NS_274 0 9.9999999999999998e-13
RS_274 NS_274 0 4.7583942880173470e+02
GS_274_10 0 NS_274 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 275/276
CS_275 NS_275 0 9.9999999999999998e-13
CS_276 NS_276 0 9.9999999999999998e-13
RS_275 NS_275 0 2.4147519902582747e+01
RS_276 NS_276 0 2.4147519902582744e+01
GL_275 0 NS_275 NS_276 0 3.6063062163307147e-01
GL_276 0 NS_276 NS_275 0 -3.6063062163307147e-01
GS_275_10 0 NS_275 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 277/278
CS_277 NS_277 0 9.9999999999999998e-13
CS_278 NS_278 0 9.9999999999999998e-13
RS_277 NS_277 0 1.8217846373726687e+01
RS_278 NS_278 0 1.8217846373726687e+01
GL_277 0 NS_277 NS_278 0 3.0904106785287211e-01
GL_278 0 NS_278 NS_277 0 -3.0904106785287211e-01
GS_277_10 0 NS_277 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 279/280
CS_279 NS_279 0 9.9999999999999998e-13
CS_280 NS_280 0 9.9999999999999998e-13
RS_279 NS_279 0 1.6355478720039709e+01
RS_280 NS_280 0 1.6355478720039706e+01
GL_279 0 NS_279 NS_280 0 2.6900015870612737e-01
GL_280 0 NS_280 NS_279 0 -2.6900015870612737e-01
GS_279_10 0 NS_279 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 281/282
CS_281 NS_281 0 9.9999999999999998e-13
CS_282 NS_282 0 9.9999999999999998e-13
RS_281 NS_281 0 1.6509546628040873e+01
RS_282 NS_282 0 1.6509546628040873e+01
GL_281 0 NS_281 NS_282 0 2.2664475020429389e-01
GL_282 0 NS_282 NS_281 0 -2.2664475020429389e-01
GS_281_10 0 NS_281 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 283/284
CS_283 NS_283 0 9.9999999999999998e-13
CS_284 NS_284 0 9.9999999999999998e-13
RS_283 NS_283 0 1.6536240554804539e+01
RS_284 NS_284 0 1.6536240554804539e+01
GL_283 0 NS_283 NS_284 0 1.9441023356946371e-01
GL_284 0 NS_284 NS_283 0 -1.9441023356946371e-01
GS_283_10 0 NS_283 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 285/286
CS_285 NS_285 0 9.9999999999999998e-13
CS_286 NS_286 0 9.9999999999999998e-13
RS_285 NS_285 0 1.7105682444637345e+01
RS_286 NS_286 0 1.7105682444637345e+01
GL_285 0 NS_285 NS_286 0 1.6030676643748842e-01
GL_286 0 NS_286 NS_285 0 -1.6030676643748842e-01
GS_285_10 0 NS_285 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 287/288
CS_287 NS_287 0 9.9999999999999998e-13
CS_288 NS_288 0 9.9999999999999998e-13
RS_287 NS_287 0 1.7548692376233411e+01
RS_288 NS_288 0 1.7548692376233408e+01
GL_287 0 NS_287 NS_288 0 1.2418335580210092e-01
GL_288 0 NS_288 NS_287 0 -1.2418335580210092e-01
GS_287_10 0 NS_287 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 289/290
CS_289 NS_289 0 9.9999999999999998e-13
CS_290 NS_290 0 9.9999999999999998e-13
RS_289 NS_289 0 1.9080711385242900e+01
RS_290 NS_290 0 1.9080711385242903e+01
GL_289 0 NS_289 NS_290 0 9.0245963773871965e-02
GL_290 0 NS_290 NS_289 0 -9.0245963773871965e-02
GS_289_10 0 NS_289 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 291/292
CS_291 NS_291 0 9.9999999999999998e-13
CS_292 NS_292 0 9.9999999999999998e-13
RS_291 NS_291 0 1.9398886873467703e+01
RS_292 NS_292 0 1.9398886873467703e+01
GL_291 0 NS_291 NS_292 0 5.0255945091433295e-02
GL_292 0 NS_292 NS_291 0 -5.0255945091433295e-02
GS_291_10 0 NS_291 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 293/294
CS_293 NS_293 0 9.9999999999999998e-13
CS_294 NS_294 0 9.9999999999999998e-13
RS_293 NS_293 0 4.6104523042200498e+01
RS_294 NS_294 0 4.6104523042200498e+01
GL_293 0 NS_293 NS_294 0 2.6612229878385272e-02
GL_294 0 NS_294 NS_293 0 -2.6612229878385272e-02
GS_293_10 0 NS_293 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 295/296
CS_295 NS_295 0 9.9999999999999998e-13
CS_296 NS_296 0 9.9999999999999998e-13
RS_295 NS_295 0 5.0459916965113045e+01
RS_296 NS_296 0 5.0459916965113038e+01
GL_295 0 NS_295 NS_296 0 3.3991465082001564e-02
GL_296 0 NS_296 NS_295 0 -3.3991465082001564e-02
GS_295_10 0 NS_295 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 297/298
CS_297 NS_297 0 9.9999999999999998e-13
CS_298 NS_298 0 9.9999999999999998e-13
RS_297 NS_297 0 1.4140189915393535e+03
RS_298 NS_298 0 1.4140189915393535e+03
GL_297 0 NS_297 NS_298 0 1.8736958636705965e-03
GL_298 0 NS_298 NS_297 0 -1.8736958636705965e-03
GS_297_10 0 NS_297 NA_10 0 7.3338024411935532e-01
*
* Complex pair n. 299/300
CS_299 NS_299 0 9.9999999999999998e-13
CS_300 NS_300 0 9.9999999999999998e-13
RS_299 NS_299 0 9.6884954140421924e+03
RS_300 NS_300 0 9.6884954140421905e+03
GL_299 0 NS_299 NS_300 0 7.9053621147275857e-05
GL_300 0 NS_300 NS_299 0 -7.9053621147275857e-05
GS_299_10 0 NS_299 NA_10 0 7.3338024411935532e-01
*
* Real pole n. 301
CS_301 NS_301 0 9.9999999999999998e-13
RS_301 NS_301 0 7.8204801849513412e+00
GS_301_11 0 NS_301 NA_11 0 7.3338024411935532e-01
*
* Real pole n. 302
CS_302 NS_302 0 9.9999999999999998e-13
RS_302 NS_302 0 2.1257837644909412e+01
GS_302_11 0 NS_302 NA_11 0 7.3338024411935532e-01
*
* Real pole n. 303
CS_303 NS_303 0 9.9999999999999998e-13
RS_303 NS_303 0 8.8189725508130692e+01
GS_303_11 0 NS_303 NA_11 0 7.3338024411935532e-01
*
* Real pole n. 304
CS_304 NS_304 0 9.9999999999999998e-13
RS_304 NS_304 0 4.7583942880173470e+02
GS_304_11 0 NS_304 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 305/306
CS_305 NS_305 0 9.9999999999999998e-13
CS_306 NS_306 0 9.9999999999999998e-13
RS_305 NS_305 0 2.4147519902582747e+01
RS_306 NS_306 0 2.4147519902582744e+01
GL_305 0 NS_305 NS_306 0 3.6063062163307147e-01
GL_306 0 NS_306 NS_305 0 -3.6063062163307147e-01
GS_305_11 0 NS_305 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 307/308
CS_307 NS_307 0 9.9999999999999998e-13
CS_308 NS_308 0 9.9999999999999998e-13
RS_307 NS_307 0 1.8217846373726687e+01
RS_308 NS_308 0 1.8217846373726687e+01
GL_307 0 NS_307 NS_308 0 3.0904106785287211e-01
GL_308 0 NS_308 NS_307 0 -3.0904106785287211e-01
GS_307_11 0 NS_307 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 309/310
CS_309 NS_309 0 9.9999999999999998e-13
CS_310 NS_310 0 9.9999999999999998e-13
RS_309 NS_309 0 1.6355478720039709e+01
RS_310 NS_310 0 1.6355478720039706e+01
GL_309 0 NS_309 NS_310 0 2.6900015870612737e-01
GL_310 0 NS_310 NS_309 0 -2.6900015870612737e-01
GS_309_11 0 NS_309 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 311/312
CS_311 NS_311 0 9.9999999999999998e-13
CS_312 NS_312 0 9.9999999999999998e-13
RS_311 NS_311 0 1.6509546628040873e+01
RS_312 NS_312 0 1.6509546628040873e+01
GL_311 0 NS_311 NS_312 0 2.2664475020429389e-01
GL_312 0 NS_312 NS_311 0 -2.2664475020429389e-01
GS_311_11 0 NS_311 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 313/314
CS_313 NS_313 0 9.9999999999999998e-13
CS_314 NS_314 0 9.9999999999999998e-13
RS_313 NS_313 0 1.6536240554804539e+01
RS_314 NS_314 0 1.6536240554804539e+01
GL_313 0 NS_313 NS_314 0 1.9441023356946371e-01
GL_314 0 NS_314 NS_313 0 -1.9441023356946371e-01
GS_313_11 0 NS_313 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 315/316
CS_315 NS_315 0 9.9999999999999998e-13
CS_316 NS_316 0 9.9999999999999998e-13
RS_315 NS_315 0 1.7105682444637345e+01
RS_316 NS_316 0 1.7105682444637345e+01
GL_315 0 NS_315 NS_316 0 1.6030676643748842e-01
GL_316 0 NS_316 NS_315 0 -1.6030676643748842e-01
GS_315_11 0 NS_315 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 317/318
CS_317 NS_317 0 9.9999999999999998e-13
CS_318 NS_318 0 9.9999999999999998e-13
RS_317 NS_317 0 1.7548692376233411e+01
RS_318 NS_318 0 1.7548692376233408e+01
GL_317 0 NS_317 NS_318 0 1.2418335580210092e-01
GL_318 0 NS_318 NS_317 0 -1.2418335580210092e-01
GS_317_11 0 NS_317 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 319/320
CS_319 NS_319 0 9.9999999999999998e-13
CS_320 NS_320 0 9.9999999999999998e-13
RS_319 NS_319 0 1.9080711385242900e+01
RS_320 NS_320 0 1.9080711385242903e+01
GL_319 0 NS_319 NS_320 0 9.0245963773871965e-02
GL_320 0 NS_320 NS_319 0 -9.0245963773871965e-02
GS_319_11 0 NS_319 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 321/322
CS_321 NS_321 0 9.9999999999999998e-13
CS_322 NS_322 0 9.9999999999999998e-13
RS_321 NS_321 0 1.9398886873467703e+01
RS_322 NS_322 0 1.9398886873467703e+01
GL_321 0 NS_321 NS_322 0 5.0255945091433295e-02
GL_322 0 NS_322 NS_321 0 -5.0255945091433295e-02
GS_321_11 0 NS_321 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 323/324
CS_323 NS_323 0 9.9999999999999998e-13
CS_324 NS_324 0 9.9999999999999998e-13
RS_323 NS_323 0 4.6104523042200498e+01
RS_324 NS_324 0 4.6104523042200498e+01
GL_323 0 NS_323 NS_324 0 2.6612229878385272e-02
GL_324 0 NS_324 NS_323 0 -2.6612229878385272e-02
GS_323_11 0 NS_323 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 325/326
CS_325 NS_325 0 9.9999999999999998e-13
CS_326 NS_326 0 9.9999999999999998e-13
RS_325 NS_325 0 5.0459916965113045e+01
RS_326 NS_326 0 5.0459916965113038e+01
GL_325 0 NS_325 NS_326 0 3.3991465082001564e-02
GL_326 0 NS_326 NS_325 0 -3.3991465082001564e-02
GS_325_11 0 NS_325 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 327/328
CS_327 NS_327 0 9.9999999999999998e-13
CS_328 NS_328 0 9.9999999999999998e-13
RS_327 NS_327 0 1.4140189915393535e+03
RS_328 NS_328 0 1.4140189915393535e+03
GL_327 0 NS_327 NS_328 0 1.8736958636705965e-03
GL_328 0 NS_328 NS_327 0 -1.8736958636705965e-03
GS_327_11 0 NS_327 NA_11 0 7.3338024411935532e-01
*
* Complex pair n. 329/330
CS_329 NS_329 0 9.9999999999999998e-13
CS_330 NS_330 0 9.9999999999999998e-13
RS_329 NS_329 0 9.6884954140421924e+03
RS_330 NS_330 0 9.6884954140421905e+03
GL_329 0 NS_329 NS_330 0 7.9053621147275857e-05
GL_330 0 NS_330 NS_329 0 -7.9053621147275857e-05
GS_329_11 0 NS_329 NA_11 0 7.3338024411935532e-01
*
* Real pole n. 331
CS_331 NS_331 0 9.9999999999999998e-13
RS_331 NS_331 0 7.8204801849513412e+00
GS_331_12 0 NS_331 NA_12 0 7.3338024411935532e-01
*
* Real pole n. 332
CS_332 NS_332 0 9.9999999999999998e-13
RS_332 NS_332 0 2.1257837644909412e+01
GS_332_12 0 NS_332 NA_12 0 7.3338024411935532e-01
*
* Real pole n. 333
CS_333 NS_333 0 9.9999999999999998e-13
RS_333 NS_333 0 8.8189725508130692e+01
GS_333_12 0 NS_333 NA_12 0 7.3338024411935532e-01
*
* Real pole n. 334
CS_334 NS_334 0 9.9999999999999998e-13
RS_334 NS_334 0 4.7583942880173470e+02
GS_334_12 0 NS_334 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 335/336
CS_335 NS_335 0 9.9999999999999998e-13
CS_336 NS_336 0 9.9999999999999998e-13
RS_335 NS_335 0 2.4147519902582747e+01
RS_336 NS_336 0 2.4147519902582744e+01
GL_335 0 NS_335 NS_336 0 3.6063062163307147e-01
GL_336 0 NS_336 NS_335 0 -3.6063062163307147e-01
GS_335_12 0 NS_335 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 337/338
CS_337 NS_337 0 9.9999999999999998e-13
CS_338 NS_338 0 9.9999999999999998e-13
RS_337 NS_337 0 1.8217846373726687e+01
RS_338 NS_338 0 1.8217846373726687e+01
GL_337 0 NS_337 NS_338 0 3.0904106785287211e-01
GL_338 0 NS_338 NS_337 0 -3.0904106785287211e-01
GS_337_12 0 NS_337 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 339/340
CS_339 NS_339 0 9.9999999999999998e-13
CS_340 NS_340 0 9.9999999999999998e-13
RS_339 NS_339 0 1.6355478720039709e+01
RS_340 NS_340 0 1.6355478720039706e+01
GL_339 0 NS_339 NS_340 0 2.6900015870612737e-01
GL_340 0 NS_340 NS_339 0 -2.6900015870612737e-01
GS_339_12 0 NS_339 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 341/342
CS_341 NS_341 0 9.9999999999999998e-13
CS_342 NS_342 0 9.9999999999999998e-13
RS_341 NS_341 0 1.6509546628040873e+01
RS_342 NS_342 0 1.6509546628040873e+01
GL_341 0 NS_341 NS_342 0 2.2664475020429389e-01
GL_342 0 NS_342 NS_341 0 -2.2664475020429389e-01
GS_341_12 0 NS_341 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 343/344
CS_343 NS_343 0 9.9999999999999998e-13
CS_344 NS_344 0 9.9999999999999998e-13
RS_343 NS_343 0 1.6536240554804539e+01
RS_344 NS_344 0 1.6536240554804539e+01
GL_343 0 NS_343 NS_344 0 1.9441023356946371e-01
GL_344 0 NS_344 NS_343 0 -1.9441023356946371e-01
GS_343_12 0 NS_343 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 345/346
CS_345 NS_345 0 9.9999999999999998e-13
CS_346 NS_346 0 9.9999999999999998e-13
RS_345 NS_345 0 1.7105682444637345e+01
RS_346 NS_346 0 1.7105682444637345e+01
GL_345 0 NS_345 NS_346 0 1.6030676643748842e-01
GL_346 0 NS_346 NS_345 0 -1.6030676643748842e-01
GS_345_12 0 NS_345 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 347/348
CS_347 NS_347 0 9.9999999999999998e-13
CS_348 NS_348 0 9.9999999999999998e-13
RS_347 NS_347 0 1.7548692376233411e+01
RS_348 NS_348 0 1.7548692376233408e+01
GL_347 0 NS_347 NS_348 0 1.2418335580210092e-01
GL_348 0 NS_348 NS_347 0 -1.2418335580210092e-01
GS_347_12 0 NS_347 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 349/350
CS_349 NS_349 0 9.9999999999999998e-13
CS_350 NS_350 0 9.9999999999999998e-13
RS_349 NS_349 0 1.9080711385242900e+01
RS_350 NS_350 0 1.9080711385242903e+01
GL_349 0 NS_349 NS_350 0 9.0245963773871965e-02
GL_350 0 NS_350 NS_349 0 -9.0245963773871965e-02
GS_349_12 0 NS_349 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 351/352
CS_351 NS_351 0 9.9999999999999998e-13
CS_352 NS_352 0 9.9999999999999998e-13
RS_351 NS_351 0 1.9398886873467703e+01
RS_352 NS_352 0 1.9398886873467703e+01
GL_351 0 NS_351 NS_352 0 5.0255945091433295e-02
GL_352 0 NS_352 NS_351 0 -5.0255945091433295e-02
GS_351_12 0 NS_351 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 353/354
CS_353 NS_353 0 9.9999999999999998e-13
CS_354 NS_354 0 9.9999999999999998e-13
RS_353 NS_353 0 4.6104523042200498e+01
RS_354 NS_354 0 4.6104523042200498e+01
GL_353 0 NS_353 NS_354 0 2.6612229878385272e-02
GL_354 0 NS_354 NS_353 0 -2.6612229878385272e-02
GS_353_12 0 NS_353 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 355/356
CS_355 NS_355 0 9.9999999999999998e-13
CS_356 NS_356 0 9.9999999999999998e-13
RS_355 NS_355 0 5.0459916965113045e+01
RS_356 NS_356 0 5.0459916965113038e+01
GL_355 0 NS_355 NS_356 0 3.3991465082001564e-02
GL_356 0 NS_356 NS_355 0 -3.3991465082001564e-02
GS_355_12 0 NS_355 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 357/358
CS_357 NS_357 0 9.9999999999999998e-13
CS_358 NS_358 0 9.9999999999999998e-13
RS_357 NS_357 0 1.4140189915393535e+03
RS_358 NS_358 0 1.4140189915393535e+03
GL_357 0 NS_357 NS_358 0 1.8736958636705965e-03
GL_358 0 NS_358 NS_357 0 -1.8736958636705965e-03
GS_357_12 0 NS_357 NA_12 0 7.3338024411935532e-01
*
* Complex pair n. 359/360
CS_359 NS_359 0 9.9999999999999998e-13
CS_360 NS_360 0 9.9999999999999998e-13
RS_359 NS_359 0 9.6884954140421924e+03
RS_360 NS_360 0 9.6884954140421905e+03
GL_359 0 NS_359 NS_360 0 7.9053621147275857e-05
GL_360 0 NS_360 NS_359 0 -7.9053621147275857e-05
GS_359_12 0 NS_359 NA_12 0 7.3338024411935532e-01
*
******************************


.ends
*******************
* End of subcircuit
*******************
