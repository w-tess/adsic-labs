**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [6 4 32] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_7_Module_via
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 -2.3476190152481161e-01
GC_1_2 b_1 NI_1 NS_2 0 5.7313802404226920e-02
GC_1_3 b_1 NI_1 NS_3 0 3.5070557596673506e-05
GC_1_4 b_1 NI_1 NS_4 0 -5.7550637103894193e-08
GC_1_5 b_1 NI_1 NS_5 0 8.4792708509077094e-02
GC_1_6 b_1 NI_1 NS_6 0 1.8302708641802974e-03
GC_1_7 b_1 NI_1 NS_7 0 1.1912200922952142e-04
GC_1_8 b_1 NI_1 NS_8 0 1.8099707981580474e-03
GC_1_9 b_1 NI_1 NS_9 0 6.3553819087257260e-03
GC_1_10 b_1 NI_1 NS_10 0 5.6406106277975213e-03
GC_1_11 b_1 NI_1 NS_11 0 -6.6967051856477696e-03
GC_1_12 b_1 NI_1 NS_12 0 3.2003725177471671e-03
GC_1_13 b_1 NI_1 NS_13 0 -1.1790878424069107e-05
GC_1_14 b_1 NI_1 NS_14 0 3.8503755691126717e-06
GC_1_15 b_1 NI_1 NS_15 0 3.0535255299386479e-06
GC_1_16 b_1 NI_1 NS_16 0 -3.8681003358483419e-06
GC_1_17 b_1 NI_1 NS_17 0 1.4466936754852926e-04
GC_1_18 b_1 NI_1 NS_18 0 -3.2847423884007327e-05
GC_1_19 b_1 NI_1 NS_19 0 3.5556387841469212e-06
GC_1_20 b_1 NI_1 NS_20 0 2.2733405913017598e-05
GC_1_21 b_1 NI_1 NS_21 0 2.9017389421552667e-04
GC_1_22 b_1 NI_1 NS_22 0 1.2279194976957467e-05
GC_1_23 b_1 NI_1 NS_23 0 2.1618327386417936e-06
GC_1_24 b_1 NI_1 NS_24 0 -6.7715212038482963e-07
GC_1_25 b_1 NI_1 NS_25 0 5.2748502844588091e-04
GC_1_26 b_1 NI_1 NS_26 0 -7.0275726374697904e-04
GC_1_27 b_1 NI_1 NS_27 0 -1.7106643364005989e-05
GC_1_28 b_1 NI_1 NS_28 0 -7.4930472481771201e-06
GC_1_29 b_1 NI_1 NS_29 0 -1.0676140772074840e-05
GC_1_30 b_1 NI_1 NS_30 0 3.0232130735855309e-05
GC_1_31 b_1 NI_1 NS_31 0 3.4290849583272460e-04
GC_1_32 b_1 NI_1 NS_32 0 3.1767472901836745e-05
GC_1_33 b_1 NI_1 NS_33 0 5.4902060238711157e-06
GC_1_34 b_1 NI_1 NS_34 0 -2.4650151058302983e-06
GC_1_35 b_1 NI_1 NS_35 0 3.2009959771444330e-02
GC_1_36 b_1 NI_1 NS_36 0 3.2719696476615920e-02
GC_1_37 b_1 NI_1 NS_37 0 1.6804908864368286e-04
GC_1_38 b_1 NI_1 NS_38 0 2.5135580356528736e-07
GC_1_39 b_1 NI_1 NS_39 0 -6.1874393326584481e-02
GC_1_40 b_1 NI_1 NS_40 0 -1.7409431503948192e-02
GC_1_41 b_1 NI_1 NS_41 0 -1.6877754454860845e-03
GC_1_42 b_1 NI_1 NS_42 0 5.1408019541974818e-03
GC_1_43 b_1 NI_1 NS_43 0 1.3108823115615131e-02
GC_1_44 b_1 NI_1 NS_44 0 1.6480821881009647e-02
GC_1_45 b_1 NI_1 NS_45 0 7.1536705640909302e-03
GC_1_46 b_1 NI_1 NS_46 0 -5.5301145380985716e-04
GC_1_47 b_1 NI_1 NS_47 0 -2.0884666125041100e-07
GC_1_48 b_1 NI_1 NS_48 0 -1.2705593496916481e-05
GC_1_49 b_1 NI_1 NS_49 0 3.5756476785548223e-06
GC_1_50 b_1 NI_1 NS_50 0 -1.8243789682008299e-05
GC_1_51 b_1 NI_1 NS_51 0 2.1814587672990690e-04
GC_1_52 b_1 NI_1 NS_52 0 1.6868740886348145e-04
GC_1_53 b_1 NI_1 NS_53 0 2.1960598062228721e-05
GC_1_54 b_1 NI_1 NS_54 0 -1.3836493289683241e-05
GC_1_55 b_1 NI_1 NS_55 0 3.2700138590341875e-04
GC_1_56 b_1 NI_1 NS_56 0 1.2486984015495982e-04
GC_1_57 b_1 NI_1 NS_57 0 -1.5125494660833857e-06
GC_1_58 b_1 NI_1 NS_58 0 -8.5171698370654821e-07
GC_1_59 b_1 NI_1 NS_59 0 2.9501617851636119e-04
GC_1_60 b_1 NI_1 NS_60 0 -6.1850003944988999e-04
GC_1_61 b_1 NI_1 NS_61 0 -6.1343331393865154e-06
GC_1_62 b_1 NI_1 NS_62 0 -2.2845404691796166e-05
GC_1_63 b_1 NI_1 NS_63 0 2.6437637254900810e-06
GC_1_64 b_1 NI_1 NS_64 0 -3.3486942178224434e-05
GC_1_65 b_1 NI_1 NS_65 0 4.3699590982081886e-04
GC_1_66 b_1 NI_1 NS_66 0 -3.1731305243606438e-05
GC_1_67 b_1 NI_1 NS_67 0 -1.1620538838658802e-05
GC_1_68 b_1 NI_1 NS_68 0 -1.8575138292907603e-05
GC_1_69 b_1 NI_1 NS_69 0 -3.1657118188169263e-02
GC_1_70 b_1 NI_1 NS_70 0 3.1159948802310278e-03
GC_1_71 b_1 NI_1 NS_71 0 -1.5426912768139085e-05
GC_1_72 b_1 NI_1 NS_72 0 -5.7358729582158904e-09
GC_1_73 b_1 NI_1 NS_73 0 1.0270010214037605e-02
GC_1_74 b_1 NI_1 NS_74 0 -9.5200833833707990e-03
GC_1_75 b_1 NI_1 NS_75 0 -1.9101991775227940e-03
GC_1_76 b_1 NI_1 NS_76 0 2.9132725826606887e-04
GC_1_77 b_1 NI_1 NS_77 0 5.1554691670436048e-03
GC_1_78 b_1 NI_1 NS_78 0 3.4628276666187996e-03
GC_1_79 b_1 NI_1 NS_79 0 1.8666620287616916e-03
GC_1_80 b_1 NI_1 NS_80 0 -1.9705655092230398e-04
GC_1_81 b_1 NI_1 NS_81 0 -1.0059794402394579e-05
GC_1_82 b_1 NI_1 NS_82 0 2.1296775407908357e-06
GC_1_83 b_1 NI_1 NS_83 0 2.2299472042933832e-06
GC_1_84 b_1 NI_1 NS_84 0 -3.8458737633432268e-06
GC_1_85 b_1 NI_1 NS_85 0 1.5685599919711008e-04
GC_1_86 b_1 NI_1 NS_86 0 -3.8577869910971789e-05
GC_1_87 b_1 NI_1 NS_87 0 3.7221189058105502e-06
GC_1_88 b_1 NI_1 NS_88 0 1.5529487530100197e-05
GC_1_89 b_1 NI_1 NS_89 0 1.9027272124624468e-04
GC_1_90 b_1 NI_1 NS_90 0 -6.9065617389403311e-06
GC_1_91 b_1 NI_1 NS_91 0 7.6357258399578332e-07
GC_1_92 b_1 NI_1 NS_92 0 2.2263199358143584e-06
GC_1_93 b_1 NI_1 NS_93 0 8.1868974820227276e-05
GC_1_94 b_1 NI_1 NS_94 0 -3.6498797477095741e-04
GC_1_95 b_1 NI_1 NS_95 0 1.1751038235879870e-05
GC_1_96 b_1 NI_1 NS_96 0 -1.7260291347903923e-05
GC_1_97 b_1 NI_1 NS_97 0 -3.1467610565500775e-06
GC_1_98 b_1 NI_1 NS_98 0 1.7248352465372574e-05
GC_1_99 b_1 NI_1 NS_99 0 4.4073178007147506e-04
GC_1_100 b_1 NI_1 NS_100 0 8.2753916500390119e-05
GC_1_101 b_1 NI_1 NS_101 0 3.0246262348264537e-06
GC_1_102 b_1 NI_1 NS_102 0 -1.7723129126214380e-06
GC_1_103 b_1 NI_1 NS_103 0 3.0722076756179034e-02
GC_1_104 b_1 NI_1 NS_104 0 -3.3971232756807067e-03
GC_1_105 b_1 NI_1 NS_105 0 -2.2139581244340832e-06
GC_1_106 b_1 NI_1 NS_106 0 9.6182806071163380e-09
GC_1_107 b_1 NI_1 NS_107 0 -1.5126270987009881e-02
GC_1_108 b_1 NI_1 NS_108 0 1.1482604009742884e-02
GC_1_109 b_1 NI_1 NS_109 0 2.1544010414953148e-04
GC_1_110 b_1 NI_1 NS_110 0 1.2701205364119576e-03
GC_1_111 b_1 NI_1 NS_111 0 4.1823048363005587e-03
GC_1_112 b_1 NI_1 NS_112 0 -9.1192589709208557e-03
GC_1_113 b_1 NI_1 NS_113 0 -8.5233548374701353e-03
GC_1_114 b_1 NI_1 NS_114 0 -2.2575176331694445e-03
GC_1_115 b_1 NI_1 NS_115 0 9.9919989641262950e-07
GC_1_116 b_1 NI_1 NS_116 0 -8.2328495336148385e-06
GC_1_117 b_1 NI_1 NS_117 0 5.0968714734522296e-06
GC_1_118 b_1 NI_1 NS_118 0 -1.8071168713222243e-05
GC_1_119 b_1 NI_1 NS_119 0 2.1316992291480814e-04
GC_1_120 b_1 NI_1 NS_120 0 1.6257790788322461e-04
GC_1_121 b_1 NI_1 NS_121 0 1.3372192844490680e-05
GC_1_122 b_1 NI_1 NS_122 0 -1.5186621284457262e-05
GC_1_123 b_1 NI_1 NS_123 0 2.2701577352584720e-04
GC_1_124 b_1 NI_1 NS_124 0 9.9626794763142367e-05
GC_1_125 b_1 NI_1 NS_125 0 6.3112230389332725e-06
GC_1_126 b_1 NI_1 NS_126 0 1.1906427351759709e-06
GC_1_127 b_1 NI_1 NS_127 0 -1.3911523292452308e-04
GC_1_128 b_1 NI_1 NS_128 0 -3.4321117031549934e-04
GC_1_129 b_1 NI_1 NS_129 0 -7.7109193063468698e-06
GC_1_130 b_1 NI_1 NS_130 0 1.5730406447191251e-06
GC_1_131 b_1 NI_1 NS_131 0 2.3059563822539316e-06
GC_1_132 b_1 NI_1 NS_132 0 -1.5363955718861674e-05
GC_1_133 b_1 NI_1 NS_133 0 2.7812191494932810e-04
GC_1_134 b_1 NI_1 NS_134 0 -2.0109752935072589e-04
GC_1_135 b_1 NI_1 NS_135 0 -8.1291670267429272e-06
GC_1_136 b_1 NI_1 NS_136 0 -1.7189984520096298e-05
GC_1_137 b_1 NI_1 NS_137 0 -1.1373952718728340e-02
GC_1_138 b_1 NI_1 NS_138 0 1.4503987994998783e-03
GC_1_139 b_1 NI_1 NS_139 0 -2.8391792384441965e-06
GC_1_140 b_1 NI_1 NS_140 0 -2.7604371030460235e-09
GC_1_141 b_1 NI_1 NS_141 0 2.7030250748053919e-03
GC_1_142 b_1 NI_1 NS_142 0 -1.9543051266785291e-03
GC_1_143 b_1 NI_1 NS_143 0 -5.1294702900277537e-04
GC_1_144 b_1 NI_1 NS_144 0 1.0720016452352519e-03
GC_1_145 b_1 NI_1 NS_145 0 2.1084998121009843e-03
GC_1_146 b_1 NI_1 NS_146 0 -1.3339213356450205e-03
GC_1_147 b_1 NI_1 NS_147 0 -1.7860731193748691e-04
GC_1_148 b_1 NI_1 NS_148 0 -1.8464750817505067e-04
GC_1_149 b_1 NI_1 NS_149 0 -1.0345534436395367e-07
GC_1_150 b_1 NI_1 NS_150 0 -3.5620347634570140e-06
GC_1_151 b_1 NI_1 NS_151 0 1.5640164038560664e-06
GC_1_152 b_1 NI_1 NS_152 0 -4.0672528324346685e-06
GC_1_153 b_1 NI_1 NS_153 0 1.6047617895642300e-04
GC_1_154 b_1 NI_1 NS_154 0 -3.8695788776782315e-05
GC_1_155 b_1 NI_1 NS_155 0 -2.2024897944514057e-07
GC_1_156 b_1 NI_1 NS_156 0 4.8750055925570045e-06
GC_1_157 b_1 NI_1 NS_157 0 6.5188407815969620e-05
GC_1_158 b_1 NI_1 NS_158 0 -1.3628769704935285e-05
GC_1_159 b_1 NI_1 NS_159 0 -8.3678823679172138e-08
GC_1_160 b_1 NI_1 NS_160 0 8.8498249358898194e-07
GC_1_161 b_1 NI_1 NS_161 0 -2.4621096722935175e-04
GC_1_162 b_1 NI_1 NS_162 0 -5.8824824351543568e-05
GC_1_163 b_1 NI_1 NS_163 0 3.4336697720496787e-05
GC_1_164 b_1 NI_1 NS_164 0 -2.2968762631857196e-05
GC_1_165 b_1 NI_1 NS_165 0 -3.9120140699970341e-06
GC_1_166 b_1 NI_1 NS_166 0 3.8121766916795109e-06
GC_1_167 b_1 NI_1 NS_167 0 5.5044278828542766e-04
GC_1_168 b_1 NI_1 NS_168 0 4.7189603956619069e-05
GC_1_169 b_1 NI_1 NS_169 0 1.7903955014165481e-06
GC_1_170 b_1 NI_1 NS_170 0 -5.0008925795479532e-07
GC_1_171 b_1 NI_1 NS_171 0 1.0923923846753357e-02
GC_1_172 b_1 NI_1 NS_172 0 -9.9093547233804636e-04
GC_1_173 b_1 NI_1 NS_173 0 -5.0420318761983594e-07
GC_1_174 b_1 NI_1 NS_174 0 4.0613332842324266e-09
GC_1_175 b_1 NI_1 NS_175 0 -4.6032555066704527e-03
GC_1_176 b_1 NI_1 NS_176 0 4.7075079694364093e-03
GC_1_177 b_1 NI_1 NS_177 0 1.0470823129737126e-04
GC_1_178 b_1 NI_1 NS_178 0 1.2216823608871741e-03
GC_1_179 b_1 NI_1 NS_179 0 1.2341744570448748e-03
GC_1_180 b_1 NI_1 NS_180 0 -4.5722213131294352e-03
GC_1_181 b_1 NI_1 NS_181 0 -3.8831213595553562e-03
GC_1_182 b_1 NI_1 NS_182 0 -3.5043686899488601e-04
GC_1_183 b_1 NI_1 NS_183 0 -1.9925457661667509e-06
GC_1_184 b_1 NI_1 NS_184 0 -1.8025931211575755e-07
GC_1_185 b_1 NI_1 NS_185 0 5.4110874899155244e-06
GC_1_186 b_1 NI_1 NS_186 0 -1.8433002172691014e-05
GC_1_187 b_1 NI_1 NS_187 0 2.1095218456431417e-04
GC_1_188 b_1 NI_1 NS_188 0 1.5828722460595708e-04
GC_1_189 b_1 NI_1 NS_189 0 6.9360686965348669e-06
GC_1_190 b_1 NI_1 NS_190 0 -2.5853831125879201e-06
GC_1_191 b_1 NI_1 NS_191 0 6.2305608493093160e-05
GC_1_192 b_1 NI_1 NS_192 0 3.3611621446890042e-05
GC_1_193 b_1 NI_1 NS_193 0 1.3262876435067759e-06
GC_1_194 b_1 NI_1 NS_194 0 -7.8071333391301999e-08
GC_1_195 b_1 NI_1 NS_195 0 -1.7782476325983455e-04
GC_1_196 b_1 NI_1 NS_196 0 -2.4741239587442770e-05
GC_1_197 b_1 NI_1 NS_197 0 6.7187772040314824e-07
GC_1_198 b_1 NI_1 NS_198 0 1.2257205215788823e-05
GC_1_199 b_1 NI_1 NS_199 0 1.1931166701003403e-06
GC_1_200 b_1 NI_1 NS_200 0 -1.1017135045293321e-05
GC_1_201 b_1 NI_1 NS_201 0 3.9572249699441339e-04
GC_1_202 b_1 NI_1 NS_202 0 -1.5734619797388028e-04
GC_1_203 b_1 NI_1 NS_203 0 -1.1966920564689842e-05
GC_1_204 b_1 NI_1 NS_204 0 -1.9429578593684316e-05
GC_1_205 b_1 NI_1 NS_205 0 -3.0412032029685475e-03
GC_1_206 b_1 NI_1 NS_206 0 5.6947557399680230e-04
GC_1_207 b_1 NI_1 NS_207 0 -9.6944960983608573e-07
GC_1_208 b_1 NI_1 NS_208 0 -1.1830912794069074e-09
GC_1_209 b_1 NI_1 NS_209 0 1.4261246104470212e-03
GC_1_210 b_1 NI_1 NS_210 0 -3.4967948768265461e-04
GC_1_211 b_1 NI_1 NS_211 0 -7.0604122291234919e-04
GC_1_212 b_1 NI_1 NS_212 0 2.7752912413732156e-04
GC_1_213 b_1 NI_1 NS_213 0 2.1133722932028791e-05
GC_1_214 b_1 NI_1 NS_214 0 1.3191327557761167e-04
GC_1_215 b_1 NI_1 NS_215 0 4.8294649307297898e-04
GC_1_216 b_1 NI_1 NS_216 0 1.3021460783595772e-04
GC_1_217 b_1 NI_1 NS_217 0 4.6795677933238472e-08
GC_1_218 b_1 NI_1 NS_218 0 1.5979265938679379e-06
GC_1_219 b_1 NI_1 NS_219 0 1.5105287843698764e-06
GC_1_220 b_1 NI_1 NS_220 0 -3.7040427436798161e-06
GC_1_221 b_1 NI_1 NS_221 0 1.5909935337923086e-04
GC_1_222 b_1 NI_1 NS_222 0 -4.2454103402633932e-05
GC_1_223 b_1 NI_1 NS_223 0 -1.2405611744357635e-06
GC_1_224 b_1 NI_1 NS_224 0 -7.6111416101028372e-06
GC_1_225 b_1 NI_1 NS_225 0 -8.6255185722256361e-05
GC_1_226 b_1 NI_1 NS_226 0 -8.2379059073955117e-06
GC_1_227 b_1 NI_1 NS_227 0 3.9895794428205411e-07
GC_1_228 b_1 NI_1 NS_228 0 1.4327494557923282e-06
GC_1_229 b_1 NI_1 NS_229 0 -5.5169339334113410e-04
GC_1_230 b_1 NI_1 NS_230 0 2.4925963257606525e-04
GC_1_231 b_1 NI_1 NS_231 0 3.1983861960409273e-05
GC_1_232 b_1 NI_1 NS_232 0 -8.8753280517954899e-06
GC_1_233 b_1 NI_1 NS_233 0 5.6251791802242378e-06
GC_1_234 b_1 NI_1 NS_234 0 -1.1560722795681317e-05
GC_1_235 b_1 NI_1 NS_235 0 6.1009966335509786e-04
GC_1_236 b_1 NI_1 NS_236 0 -1.7156159070872000e-05
GC_1_237 b_1 NI_1 NS_237 0 3.0105783900507777e-06
GC_1_238 b_1 NI_1 NS_238 0 8.8667496772094124e-07
GC_1_239 b_1 NI_1 NS_239 0 6.4456076140368343e-03
GC_1_240 b_1 NI_1 NS_240 0 -5.3498891388806366e-04
GC_1_241 b_1 NI_1 NS_241 0 -1.5274967685217476e-07
GC_1_242 b_1 NI_1 NS_242 0 1.9703665412226863e-09
GC_1_243 b_1 NI_1 NS_243 0 -1.8570169290050322e-03
GC_1_244 b_1 NI_1 NS_244 0 2.2024766094942399e-03
GC_1_245 b_1 NI_1 NS_245 0 -3.9584143002304307e-04
GC_1_246 b_1 NI_1 NS_246 0 8.9321588536718283e-04
GC_1_247 b_1 NI_1 NS_247 0 9.6371897394787050e-04
GC_1_248 b_1 NI_1 NS_248 0 -1.7581737681820657e-03
GC_1_249 b_1 NI_1 NS_249 0 -1.6761462196828003e-03
GC_1_250 b_1 NI_1 NS_250 0 -1.3762077856964940e-04
GC_1_251 b_1 NI_1 NS_251 0 2.9027670956539026e-07
GC_1_252 b_1 NI_1 NS_252 0 1.3250059375620820e-06
GC_1_253 b_1 NI_1 NS_253 0 4.8630162301243331e-06
GC_1_254 b_1 NI_1 NS_254 0 -1.7947927853710601e-05
GC_1_255 b_1 NI_1 NS_255 0 2.1644136384353126e-04
GC_1_256 b_1 NI_1 NS_256 0 1.5536782872127474e-04
GC_1_257 b_1 NI_1 NS_257 0 -8.1691623069295381e-06
GC_1_258 b_1 NI_1 NS_258 0 1.5866622651224244e-06
GC_1_259 b_1 NI_1 NS_259 0 -8.3115441776817974e-05
GC_1_260 b_1 NI_1 NS_260 0 -4.1380887793063904e-05
GC_1_261 b_1 NI_1 NS_261 0 2.2215011797082572e-06
GC_1_262 b_1 NI_1 NS_262 0 -8.9785794975108142e-08
GC_1_263 b_1 NI_1 NS_263 0 -3.1780949669871005e-04
GC_1_264 b_1 NI_1 NS_264 0 2.2472202088774356e-04
GC_1_265 b_1 NI_1 NS_265 0 1.6263470630039532e-06
GC_1_266 b_1 NI_1 NS_266 0 2.0683364638883891e-05
GC_1_267 b_1 NI_1 NS_267 0 -1.7045418288327103e-06
GC_1_268 b_1 NI_1 NS_268 0 1.2689147420373884e-05
GC_1_269 b_1 NI_1 NS_269 0 4.2602826978879439e-04
GC_1_270 b_1 NI_1 NS_270 0 -2.1085468106708349e-04
GC_1_271 b_1 NI_1 NS_271 0 -1.0779384947541552e-05
GC_1_272 b_1 NI_1 NS_272 0 -1.8806989572204151e-05
GC_1_273 b_1 NI_1 NS_273 0 4.2780760341808114e-03
GC_1_274 b_1 NI_1 NS_274 0 -2.4442290758634530e-05
GC_1_275 b_1 NI_1 NS_275 0 2.2728553725897993e-07
GC_1_276 b_1 NI_1 NS_276 0 -8.6800924971699220e-10
GC_1_277 b_1 NI_1 NS_277 0 1.6291288342388660e-03
GC_1_278 b_1 NI_1 NS_278 0 1.5105402678325479e-03
GC_1_279 b_1 NI_1 NS_279 0 9.5865243964358689e-04
GC_1_280 b_1 NI_1 NS_280 0 -8.7359934453526495e-05
GC_1_281 b_1 NI_1 NS_281 0 -5.6543789084542075e-03
GC_1_282 b_1 NI_1 NS_282 0 -9.5774020416230610e-04
GC_1_283 b_1 NI_1 NS_283 0 1.4993384049315146e-03
GC_1_284 b_1 NI_1 NS_284 0 2.3679275184751705e-03
GC_1_285 b_1 NI_1 NS_285 0 1.0637145990507123e-05
GC_1_286 b_1 NI_1 NS_286 0 -2.9607303019201653e-06
GC_1_287 b_1 NI_1 NS_287 0 1.2804731468468340e-06
GC_1_288 b_1 NI_1 NS_288 0 -3.5278308538594135e-06
GC_1_289 b_1 NI_1 NS_289 0 1.6382644626205151e-04
GC_1_290 b_1 NI_1 NS_290 0 -4.1962138597130696e-05
GC_1_291 b_1 NI_1 NS_291 0 -4.1065361891461702e-06
GC_1_292 b_1 NI_1 NS_292 0 -1.8042520909516444e-05
GC_1_293 b_1 NI_1 NS_293 0 -2.1791303611820348e-04
GC_1_294 b_1 NI_1 NS_294 0 -1.3664068540154773e-05
GC_1_295 b_1 NI_1 NS_295 0 6.1487022806387966e-08
GC_1_296 b_1 NI_1 NS_296 0 4.3404359870729357e-06
GC_1_297 b_1 NI_1 NS_297 0 -3.4339547683755694e-04
GC_1_298 b_1 NI_1 NS_298 0 4.2457526838999519e-04
GC_1_299 b_1 NI_1 NS_299 0 1.3347171761893207e-05
GC_1_300 b_1 NI_1 NS_300 0 8.9637008189670122e-06
GC_1_301 b_1 NI_1 NS_301 0 5.0120627958345473e-06
GC_1_302 b_1 NI_1 NS_302 0 -2.3884498525880083e-05
GC_1_303 b_1 NI_1 NS_303 0 5.8616816465808510e-04
GC_1_304 b_1 NI_1 NS_304 0 2.9526525728560757e-05
GC_1_305 b_1 NI_1 NS_305 0 2.6951042954639914e-06
GC_1_306 b_1 NI_1 NS_306 0 2.4424435517215271e-07
GC_1_307 b_1 NI_1 NS_307 0 4.7345918870848134e-03
GC_1_308 b_1 NI_1 NS_308 0 -3.4366385291377717e-04
GC_1_309 b_1 NI_1 NS_309 0 1.5106440629448694e-07
GC_1_310 b_1 NI_1 NS_310 0 9.4137862306373364e-10
GC_1_311 b_1 NI_1 NS_311 0 -4.3449911830012396e-04
GC_1_312 b_1 NI_1 NS_312 0 8.6125765249453565e-04
GC_1_313 b_1 NI_1 NS_313 0 6.2368399924161945e-04
GC_1_314 b_1 NI_1 NS_314 0 -2.1825008504636770e-04
GC_1_315 b_1 NI_1 NS_315 0 -3.2458427885253107e-03
GC_1_316 b_1 NI_1 NS_316 0 3.0259901352955803e-04
GC_1_317 b_1 NI_1 NS_317 0 1.1838453871631511e-03
GC_1_318 b_1 NI_1 NS_318 0 5.8640889715367824e-04
GC_1_319 b_1 NI_1 NS_319 0 -1.2006609199176982e-06
GC_1_320 b_1 NI_1 NS_320 0 9.7221989483725732e-06
GC_1_321 b_1 NI_1 NS_321 0 5.2673962464673876e-06
GC_1_322 b_1 NI_1 NS_322 0 -1.8464037416190329e-05
GC_1_323 b_1 NI_1 NS_323 0 2.1399819726734937e-04
GC_1_324 b_1 NI_1 NS_324 0 1.5993556827673710e-04
GC_1_325 b_1 NI_1 NS_325 0 -1.3115166340991371e-05
GC_1_326 b_1 NI_1 NS_326 0 1.3797167816642410e-05
GC_1_327 b_1 NI_1 NS_327 0 -2.5483635044377218e-04
GC_1_328 b_1 NI_1 NS_328 0 -1.0341574861566638e-04
GC_1_329 b_1 NI_1 NS_329 0 2.8834982645030720e-06
GC_1_330 b_1 NI_1 NS_330 0 2.4756078762494141e-07
GC_1_331 b_1 NI_1 NS_331 0 -1.1059814998726671e-04
GC_1_332 b_1 NI_1 NS_332 0 3.2429607600523776e-04
GC_1_333 b_1 NI_1 NS_333 0 5.9064427067465109e-06
GC_1_334 b_1 NI_1 NS_334 0 1.2326822722081881e-05
GC_1_335 b_1 NI_1 NS_335 0 -4.9392301249461981e-06
GC_1_336 b_1 NI_1 NS_336 0 1.7366727720232249e-05
GC_1_337 b_1 NI_1 NS_337 0 4.3369367808554303e-04
GC_1_338 b_1 NI_1 NS_338 0 -1.4839602266219847e-04
GC_1_339 b_1 NI_1 NS_339 0 -1.0122546035889219e-05
GC_1_340 b_1 NI_1 NS_340 0 -1.6813558864609795e-05
GC_1_341 b_1 NI_1 NS_341 0 6.5904807559503146e-03
GC_1_342 b_1 NI_1 NS_342 0 -2.5708472207197099e-04
GC_1_343 b_1 NI_1 NS_343 0 6.0979909172595430e-07
GC_1_344 b_1 NI_1 NS_344 0 -6.1616422512070754e-10
GC_1_345 b_1 NI_1 NS_345 0 1.5645500060145604e-03
GC_1_346 b_1 NI_1 NS_346 0 2.0017523425897099e-03
GC_1_347 b_1 NI_1 NS_347 0 1.8705666383419777e-03
GC_1_348 b_1 NI_1 NS_348 0 -6.5671343638962665e-04
GC_1_349 b_1 NI_1 NS_349 0 -7.8873481578922398e-03
GC_1_350 b_1 NI_1 NS_350 0 -7.2195387272748642e-04
GC_1_351 b_1 NI_1 NS_351 0 1.8083956569762919e-03
GC_1_352 b_1 NI_1 NS_352 0 2.8496888973924394e-03
GC_1_353 b_1 NI_1 NS_353 0 1.2293838459796900e-05
GC_1_354 b_1 NI_1 NS_354 0 -4.0951774069529110e-06
GC_1_355 b_1 NI_1 NS_355 0 1.0123922608883901e-06
GC_1_356 b_1 NI_1 NS_356 0 -3.0941621948816188e-06
GC_1_357 b_1 NI_1 NS_357 0 1.5883069648530752e-04
GC_1_358 b_1 NI_1 NS_358 0 -4.1862836720816466e-05
GC_1_359 b_1 NI_1 NS_359 0 -3.5225816775025924e-06
GC_1_360 b_1 NI_1 NS_360 0 -2.4785539958298296e-05
GC_1_361 b_1 NI_1 NS_361 0 -2.9916784754394174e-04
GC_1_362 b_1 NI_1 NS_362 0 -1.5012637009829682e-05
GC_1_363 b_1 NI_1 NS_363 0 -1.3306450229798607e-06
GC_1_364 b_1 NI_1 NS_364 0 2.2026980847962253e-06
GC_1_365 b_1 NI_1 NS_365 0 -1.7548031124937666e-04
GC_1_366 b_1 NI_1 NS_366 0 4.5531562528048936e-04
GC_1_367 b_1 NI_1 NS_367 0 -1.5540275044910584e-05
GC_1_368 b_1 NI_1 NS_368 0 2.7587091529911209e-05
GC_1_369 b_1 NI_1 NS_369 0 9.3391621522108936e-06
GC_1_370 b_1 NI_1 NS_370 0 -3.1663593970992628e-05
GC_1_371 b_1 NI_1 NS_371 0 6.5652996856274530e-04
GC_1_372 b_1 NI_1 NS_372 0 2.9008193251953811e-05
GC_1_373 b_1 NI_1 NS_373 0 3.5005990384637468e-06
GC_1_374 b_1 NI_1 NS_374 0 7.0858461139009653e-07
GC_1_375 b_1 NI_1 NS_375 0 7.0918358494062427e-03
GC_1_376 b_1 NI_1 NS_376 0 -4.6171480516182058e-04
GC_1_377 b_1 NI_1 NS_377 0 7.8397669280374594e-07
GC_1_378 b_1 NI_1 NS_378 0 2.7813146186906737e-10
GC_1_379 b_1 NI_1 NS_379 0 5.9929465320619692e-04
GC_1_380 b_1 NI_1 NS_380 0 1.5791845991903193e-03
GC_1_381 b_1 NI_1 NS_381 0 1.3769525366940155e-03
GC_1_382 b_1 NI_1 NS_382 0 -1.3596431318487190e-03
GC_1_383 b_1 NI_1 NS_383 0 -6.7299545117768013e-03
GC_1_384 b_1 NI_1 NS_384 0 8.7059752762137397e-04
GC_1_385 b_1 NI_1 NS_385 0 1.7678525617706871e-03
GC_1_386 b_1 NI_1 NS_386 0 2.0430349030950063e-03
GC_1_387 b_1 NI_1 NS_387 0 -2.0298660696732119e-06
GC_1_388 b_1 NI_1 NS_388 0 1.1883912239679369e-05
GC_1_389 b_1 NI_1 NS_389 0 4.7055762554206580e-06
GC_1_390 b_1 NI_1 NS_390 0 -1.7366819102459687e-05
GC_1_391 b_1 NI_1 NS_391 0 2.0850591022393902e-04
GC_1_392 b_1 NI_1 NS_392 0 1.5751372040710013e-04
GC_1_393 b_1 NI_1 NS_393 0 -2.2776421200741393e-05
GC_1_394 b_1 NI_1 NS_394 0 1.5281477255479038e-05
GC_1_395 b_1 NI_1 NS_395 0 -3.2850133508436578e-04
GC_1_396 b_1 NI_1 NS_396 0 -1.5665465959404450e-04
GC_1_397 b_1 NI_1 NS_397 0 3.0793703363037989e-07
GC_1_398 b_1 NI_1 NS_398 0 -2.2371641492830852e-07
GC_1_399 b_1 NI_1 NS_399 0 -5.0290360464067945e-06
GC_1_400 b_1 NI_1 NS_400 0 3.5547547929937526e-04
GC_1_401 b_1 NI_1 NS_401 0 5.4551206575307631e-06
GC_1_402 b_1 NI_1 NS_402 0 2.1525756243933596e-06
GC_1_403 b_1 NI_1 NS_403 0 -7.4406703190945325e-06
GC_1_404 b_1 NI_1 NS_404 0 2.9076697229700215e-05
GC_1_405 b_1 NI_1 NS_405 0 4.8737391569512046e-04
GC_1_406 b_1 NI_1 NS_406 0 -1.4037010527179100e-04
GC_1_407 b_1 NI_1 NS_407 0 -9.8137166636898801e-06
GC_1_408 b_1 NI_1 NS_408 0 -1.7335113658101149e-05
GD_1_1 b_1 NI_1 NA_1 0 1.0732684619642623e-01
GD_1_2 b_1 NI_1 NA_2 0 -3.4437675011807056e-02
GD_1_3 b_1 NI_1 NA_3 0 1.3894851320915055e-02
GD_1_4 b_1 NI_1 NA_4 0 -1.0656353922048056e-02
GD_1_5 b_1 NI_1 NA_5 0 6.2221544729821471e-03
GD_1_6 b_1 NI_1 NA_6 0 -3.9477678998526763e-03
GD_1_7 b_1 NI_1 NA_7 0 1.8204796529785162e-03
GD_1_8 b_1 NI_1 NA_8 0 -4.7377929509147178e-03
GD_1_9 b_1 NI_1 NA_9 0 -3.4471328115757011e-03
GD_1_10 b_1 NI_1 NA_10 0 -3.9608788045466499e-03
GD_1_11 b_1 NI_1 NA_11 0 -5.1252002380781812e-03
GD_1_12 b_1 NI_1 NA_12 0 -5.0035883883835421e-03
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 3.2009960082686952e-02
GC_2_2 b_2 NI_2 NS_2 0 3.2719696405743667e-02
GC_2_3 b_2 NI_2 NS_3 0 1.6804908934080331e-04
GC_2_4 b_2 NI_2 NS_4 0 2.5135580082319829e-07
GC_2_5 b_2 NI_2 NS_5 0 -6.1874393496143099e-02
GC_2_6 b_2 NI_2 NS_6 0 -1.7409431408426823e-02
GC_2_7 b_2 NI_2 NS_7 0 -1.6877754283437145e-03
GC_2_8 b_2 NI_2 NS_8 0 5.1408019653557185e-03
GC_2_9 b_2 NI_2 NS_9 0 1.3108823151100067e-02
GC_2_10 b_2 NI_2 NS_10 0 1.6480821761749524e-02
GC_2_11 b_2 NI_2 NS_11 0 7.1536704672391016e-03
GC_2_12 b_2 NI_2 NS_12 0 -5.5301149028248470e-04
GC_2_13 b_2 NI_2 NS_13 0 -2.0884666434877277e-07
GC_2_14 b_2 NI_2 NS_14 0 -1.2705593408129004e-05
GC_2_15 b_2 NI_2 NS_15 0 3.5756476675921844e-06
GC_2_16 b_2 NI_2 NS_16 0 -1.8243789593440759e-05
GC_2_17 b_2 NI_2 NS_17 0 2.1814587640441577e-04
GC_2_18 b_2 NI_2 NS_18 0 1.6868740842448799e-04
GC_2_19 b_2 NI_2 NS_19 0 2.1960598162960942e-05
GC_2_20 b_2 NI_2 NS_20 0 -1.3836493308320673e-05
GC_2_21 b_2 NI_2 NS_21 0 3.2700138542805129e-04
GC_2_22 b_2 NI_2 NS_22 0 1.2486984031317167e-04
GC_2_23 b_2 NI_2 NS_23 0 -1.5125494334404821e-06
GC_2_24 b_2 NI_2 NS_24 0 -8.5171701730460473e-07
GC_2_25 b_2 NI_2 NS_25 0 2.9501617777122417e-04
GC_2_26 b_2 NI_2 NS_26 0 -6.1850003991535218e-04
GC_2_27 b_2 NI_2 NS_27 0 -6.1343332312158721e-06
GC_2_28 b_2 NI_2 NS_28 0 -2.2845404588117331e-05
GC_2_29 b_2 NI_2 NS_29 0 2.6437637545091541e-06
GC_2_30 b_2 NI_2 NS_30 0 -3.3486942254259797e-05
GC_2_31 b_2 NI_2 NS_31 0 4.3699590896645844e-04
GC_2_32 b_2 NI_2 NS_32 0 -3.1731307089727079e-05
GC_2_33 b_2 NI_2 NS_33 0 -1.1620538747783134e-05
GC_2_34 b_2 NI_2 NS_34 0 -1.8575138250435423e-05
GC_2_35 b_2 NI_2 NS_35 0 1.8881342975304912e-03
GC_2_36 b_2 NI_2 NS_36 0 2.9906938804904040e-02
GC_2_37 b_2 NI_2 NS_37 0 5.8528431755688547e-05
GC_2_38 b_2 NI_2 NS_38 0 -7.0049119109049089e-08
GC_2_39 b_2 NI_2 NS_39 0 4.9715948785729928e-02
GC_2_40 b_2 NI_2 NS_40 0 3.7431481795238336e-02
GC_2_41 b_2 NI_2 NS_41 0 -4.4863900726984911e-03
GC_2_42 b_2 NI_2 NS_42 0 2.6701767278140523e-03
GC_2_43 b_2 NI_2 NS_43 0 -7.3877990156364318e-03
GC_2_44 b_2 NI_2 NS_44 0 1.4688684583857430e-02
GC_2_45 b_2 NI_2 NS_45 0 8.1520453610606984e-04
GC_2_46 b_2 NI_2 NS_46 0 4.9450887833921708e-03
GC_2_47 b_2 NI_2 NS_47 0 1.3711720568998400e-05
GC_2_48 b_2 NI_2 NS_48 0 2.6937194332246283e-06
GC_2_49 b_2 NI_2 NS_49 0 7.9200137337501960e-06
GC_2_50 b_2 NI_2 NS_50 0 -8.5773458562214236e-05
GC_2_51 b_2 NI_2 NS_51 0 2.8019481097243823e-06
GC_2_52 b_2 NI_2 NS_52 0 4.3086843792028044e-04
GC_2_53 b_2 NI_2 NS_53 0 -3.9300141262196391e-05
GC_2_54 b_2 NI_2 NS_54 0 -1.9929961342093711e-05
GC_2_55 b_2 NI_2 NS_55 0 3.1707989527429464e-04
GC_2_56 b_2 NI_2 NS_56 0 2.8008386774325489e-04
GC_2_57 b_2 NI_2 NS_57 0 -2.7542319599952974e-06
GC_2_58 b_2 NI_2 NS_58 0 1.6995234882018798e-06
GC_2_59 b_2 NI_2 NS_59 0 1.2881655766704996e-04
GC_2_60 b_2 NI_2 NS_60 0 -3.8235812228752317e-04
GC_2_61 b_2 NI_2 NS_61 0 -1.2660134551537130e-06
GC_2_62 b_2 NI_2 NS_62 0 -8.7522058561020470e-06
GC_2_63 b_2 NI_2 NS_63 0 -1.8791370529854795e-06
GC_2_64 b_2 NI_2 NS_64 0 2.0498222093756244e-05
GC_2_65 b_2 NI_2 NS_65 0 3.5642338818239641e-04
GC_2_66 b_2 NI_2 NS_66 0 -6.8440454802491161e-05
GC_2_67 b_2 NI_2 NS_67 0 -3.5827318573947375e-05
GC_2_68 b_2 NI_2 NS_68 0 4.5793604705509882e-05
GC_2_69 b_2 NI_2 NS_69 0 2.9370522612131481e-02
GC_2_70 b_2 NI_2 NS_70 0 -3.2161763880872939e-03
GC_2_71 b_2 NI_2 NS_71 0 -2.7622708734588186e-06
GC_2_72 b_2 NI_2 NS_72 0 9.7841448952529163e-09
GC_2_73 b_2 NI_2 NS_73 0 -1.4937047544501137e-02
GC_2_74 b_2 NI_2 NS_74 0 1.0982326699271865e-02
GC_2_75 b_2 NI_2 NS_75 0 9.3482999640182450e-05
GC_2_76 b_2 NI_2 NS_76 0 1.0424911114032837e-03
GC_2_77 b_2 NI_2 NS_77 0 3.9531745939806601e-03
GC_2_78 b_2 NI_2 NS_78 0 -8.3909700709851927e-03
GC_2_79 b_2 NI_2 NS_79 0 -7.8011654548330667e-03
GC_2_80 b_2 NI_2 NS_80 0 -2.4381530661474219e-03
GC_2_81 b_2 NI_2 NS_81 0 1.6886031692895535e-06
GC_2_82 b_2 NI_2 NS_82 0 -9.2850265136621189e-06
GC_2_83 b_2 NI_2 NS_83 0 5.4564606022707196e-06
GC_2_84 b_2 NI_2 NS_84 0 -1.7383572043712878e-05
GC_2_85 b_2 NI_2 NS_85 0 2.0973515188680951e-04
GC_2_86 b_2 NI_2 NS_86 0 1.5912617396931085e-04
GC_2_87 b_2 NI_2 NS_87 0 1.5865634078670285e-05
GC_2_88 b_2 NI_2 NS_88 0 -1.1907141102788260e-05
GC_2_89 b_2 NI_2 NS_89 0 2.1264910567180865e-04
GC_2_90 b_2 NI_2 NS_90 0 9.4137014311259002e-05
GC_2_91 b_2 NI_2 NS_91 0 4.4275833696888892e-06
GC_2_92 b_2 NI_2 NS_92 0 -3.4145382086495295e-07
GC_2_93 b_2 NI_2 NS_93 0 -1.3542607079450517e-04
GC_2_94 b_2 NI_2 NS_94 0 -3.3941687048874569e-04
GC_2_95 b_2 NI_2 NS_95 0 -8.4839353256329169e-06
GC_2_96 b_2 NI_2 NS_96 0 4.5246784357068218e-06
GC_2_97 b_2 NI_2 NS_97 0 -8.3032211100834007e-10
GC_2_98 b_2 NI_2 NS_98 0 -1.6739717813816514e-05
GC_2_99 b_2 NI_2 NS_99 0 2.8283216028301565e-04
GC_2_100 b_2 NI_2 NS_100 0 -1.8003605347199369e-04
GC_2_101 b_2 NI_2 NS_101 0 -6.3176620086581987e-06
GC_2_102 b_2 NI_2 NS_102 0 -1.6913493943998651e-05
GC_2_103 b_2 NI_2 NS_103 0 -1.5332093370748650e-02
GC_2_104 b_2 NI_2 NS_104 0 -1.2314667898533859e-03
GC_2_105 b_2 NI_2 NS_105 0 -1.6810069420903579e-05
GC_2_106 b_2 NI_2 NS_106 0 -4.9173208334374858e-09
GC_2_107 b_2 NI_2 NS_107 0 7.3474883609324368e-03
GC_2_108 b_2 NI_2 NS_108 0 -1.3076116995125443e-02
GC_2_109 b_2 NI_2 NS_109 0 -9.2764423413423287e-04
GC_2_110 b_2 NI_2 NS_110 0 1.5729459972767458e-03
GC_2_111 b_2 NI_2 NS_111 0 2.0262369004007243e-03
GC_2_112 b_2 NI_2 NS_112 0 3.0609941217618303e-03
GC_2_113 b_2 NI_2 NS_113 0 2.6098405314338947e-03
GC_2_114 b_2 NI_2 NS_114 0 2.2776607411206583e-03
GC_2_115 b_2 NI_2 NS_115 0 1.2288450709588903e-05
GC_2_116 b_2 NI_2 NS_116 0 3.2857666296868966e-06
GC_2_117 b_2 NI_2 NS_117 0 8.0201642780271958e-06
GC_2_118 b_2 NI_2 NS_118 0 -8.8850852064773425e-05
GC_2_119 b_2 NI_2 NS_119 0 9.8347725565516542e-06
GC_2_120 b_2 NI_2 NS_120 0 4.4338832889174730e-04
GC_2_121 b_2 NI_2 NS_121 0 -2.6828472407368918e-05
GC_2_122 b_2 NI_2 NS_122 0 -3.1731858434414485e-06
GC_2_123 b_2 NI_2 NS_123 0 2.3079223926651457e-04
GC_2_124 b_2 NI_2 NS_124 0 1.5691602379553767e-04
GC_2_125 b_2 NI_2 NS_125 0 5.7164347992835067e-07
GC_2_126 b_2 NI_2 NS_126 0 1.4167287151866778e-06
GC_2_127 b_2 NI_2 NS_127 0 -8.7603650681209930e-05
GC_2_128 b_2 NI_2 NS_128 0 -1.5897446898922475e-04
GC_2_129 b_2 NI_2 NS_129 0 -4.0092218938830947e-06
GC_2_130 b_2 NI_2 NS_130 0 -5.3004052263748386e-06
GC_2_131 b_2 NI_2 NS_131 0 -1.1048630116668595e-06
GC_2_132 b_2 NI_2 NS_132 0 1.3873149167480591e-05
GC_2_133 b_2 NI_2 NS_133 0 2.6118491015722945e-04
GC_2_134 b_2 NI_2 NS_134 0 -1.2534189742104639e-04
GC_2_135 b_2 NI_2 NS_135 0 -3.1410330573737742e-05
GC_2_136 b_2 NI_2 NS_136 0 4.5292397690485394e-05
GC_2_137 b_2 NI_2 NS_137 0 1.4777411218390995e-02
GC_2_138 b_2 NI_2 NS_138 0 -1.2746317991792614e-03
GC_2_139 b_2 NI_2 NS_139 0 4.1498022318734594e-07
GC_2_140 b_2 NI_2 NS_140 0 3.7348089151371698e-09
GC_2_141 b_2 NI_2 NS_141 0 -4.5503750921080353e-03
GC_2_142 b_2 NI_2 NS_142 0 5.9428470175790444e-03
GC_2_143 b_2 NI_2 NS_143 0 4.1983360686881723e-05
GC_2_144 b_2 NI_2 NS_144 0 9.2106433842221828e-04
GC_2_145 b_2 NI_2 NS_145 0 4.9507564676364638e-06
GC_2_146 b_2 NI_2 NS_146 0 -4.6539423743250817e-03
GC_2_147 b_2 NI_2 NS_147 0 -4.0485848193170734e-03
GC_2_148 b_2 NI_2 NS_148 0 4.6166240711193482e-04
GC_2_149 b_2 NI_2 NS_149 0 1.7712048187589303e-06
GC_2_150 b_2 NI_2 NS_150 0 2.7004233235620407e-06
GC_2_151 b_2 NI_2 NS_151 0 5.4235971553718636e-06
GC_2_152 b_2 NI_2 NS_152 0 -1.9024513216974821e-05
GC_2_153 b_2 NI_2 NS_153 0 2.1142228132154110e-04
GC_2_154 b_2 NI_2 NS_154 0 1.6341038446428653e-04
GC_2_155 b_2 NI_2 NS_155 0 4.5972252172079780e-06
GC_2_156 b_2 NI_2 NS_156 0 -1.3993519538466948e-06
GC_2_157 b_2 NI_2 NS_157 0 7.2473883541498870e-05
GC_2_158 b_2 NI_2 NS_158 0 2.0858671634232289e-05
GC_2_159 b_2 NI_2 NS_159 0 1.0538877426639567e-06
GC_2_160 b_2 NI_2 NS_160 0 -8.5106795204570240e-07
GC_2_161 b_2 NI_2 NS_161 0 -2.2653222866113315e-04
GC_2_162 b_2 NI_2 NS_162 0 -6.0344532015937344e-05
GC_2_163 b_2 NI_2 NS_163 0 -5.3089421499372127e-06
GC_2_164 b_2 NI_2 NS_164 0 1.7532060185611002e-05
GC_2_165 b_2 NI_2 NS_165 0 4.0652306457326519e-06
GC_2_166 b_2 NI_2 NS_166 0 -6.8897672162538619e-06
GC_2_167 b_2 NI_2 NS_167 0 3.8581776448301047e-04
GC_2_168 b_2 NI_2 NS_168 0 -1.6008857623391382e-04
GC_2_169 b_2 NI_2 NS_169 0 -6.4882529109477662e-06
GC_2_170 b_2 NI_2 NS_170 0 -1.6113659420129500e-05
GC_2_171 b_2 NI_2 NS_171 0 -4.1956145668695047e-03
GC_2_172 b_2 NI_2 NS_172 0 -1.1458353058879222e-03
GC_2_173 b_2 NI_2 NS_173 0 -2.4677847788672626e-06
GC_2_174 b_2 NI_2 NS_174 0 -3.8011455716095133e-09
GC_2_175 b_2 NI_2 NS_175 0 1.1173785669968638e-03
GC_2_176 b_2 NI_2 NS_176 0 -5.7754595526868426e-03
GC_2_177 b_2 NI_2 NS_177 0 -9.8345746222051552e-05
GC_2_178 b_2 NI_2 NS_178 0 7.8634017092951475e-04
GC_2_179 b_2 NI_2 NS_179 0 7.6123439616810663e-04
GC_2_180 b_2 NI_2 NS_180 0 4.6511991331836858e-04
GC_2_181 b_2 NI_2 NS_181 0 9.8823757173222330e-04
GC_2_182 b_2 NI_2 NS_182 0 6.1309237601857086e-04
GC_2_183 b_2 NI_2 NS_183 0 5.7881496986000574e-07
GC_2_184 b_2 NI_2 NS_184 0 -5.6832260877519755e-07
GC_2_185 b_2 NI_2 NS_185 0 6.7453557300145655e-06
GC_2_186 b_2 NI_2 NS_186 0 -8.8697761168778609e-05
GC_2_187 b_2 NI_2 NS_187 0 2.6191843879482410e-05
GC_2_188 b_2 NI_2 NS_188 0 4.4564360039789819e-04
GC_2_189 b_2 NI_2 NS_189 0 -1.1135891111836647e-05
GC_2_190 b_2 NI_2 NS_190 0 -9.6642851707935980e-06
GC_2_191 b_2 NI_2 NS_191 0 7.3630295514289808e-05
GC_2_192 b_2 NI_2 NS_192 0 7.8419787085046535e-05
GC_2_193 b_2 NI_2 NS_193 0 -6.7665874357261425e-07
GC_2_194 b_2 NI_2 NS_194 0 8.6731415930141588e-07
GC_2_195 b_2 NI_2 NS_195 0 -7.8883105646294159e-05
GC_2_196 b_2 NI_2 NS_196 0 1.4107884863944540e-05
GC_2_197 b_2 NI_2 NS_197 0 -5.5273122622701411e-06
GC_2_198 b_2 NI_2 NS_198 0 -8.0874434965310025e-06
GC_2_199 b_2 NI_2 NS_199 0 5.2661923028145237e-07
GC_2_200 b_2 NI_2 NS_200 0 7.7064753772509595e-06
GC_2_201 b_2 NI_2 NS_201 0 3.3034061777121703e-04
GC_2_202 b_2 NI_2 NS_202 0 -1.9723433255253614e-04
GC_2_203 b_2 NI_2 NS_203 0 -3.3640832561792243e-05
GC_2_204 b_2 NI_2 NS_204 0 5.3584372411330792e-05
GC_2_205 b_2 NI_2 NS_205 0 6.3021193745604357e-03
GC_2_206 b_2 NI_2 NS_206 0 -4.8523184538031586e-04
GC_2_207 b_2 NI_2 NS_207 0 -2.3563500297886466e-07
GC_2_208 b_2 NI_2 NS_208 0 2.0297677129969705e-09
GC_2_209 b_2 NI_2 NS_209 0 -1.7529292316191053e-03
GC_2_210 b_2 NI_2 NS_210 0 1.9670467517206710e-03
GC_2_211 b_2 NI_2 NS_211 0 -5.9233314182700111e-04
GC_2_212 b_2 NI_2 NS_212 0 8.6220036721166259e-04
GC_2_213 b_2 NI_2 NS_213 0 1.0952544920719118e-03
GC_2_214 b_2 NI_2 NS_214 0 -1.0969413964459994e-03
GC_2_215 b_2 NI_2 NS_215 0 -1.2933336472805599e-03
GC_2_216 b_2 NI_2 NS_216 0 -3.1772184772237057e-04
GC_2_217 b_2 NI_2 NS_217 0 -1.5279832657004751e-06
GC_2_218 b_2 NI_2 NS_218 0 3.3437123078645888e-07
GC_2_219 b_2 NI_2 NS_219 0 5.1384322693682593e-06
GC_2_220 b_2 NI_2 NS_220 0 -1.8057624125964127e-05
GC_2_221 b_2 NI_2 NS_221 0 2.1377371117873247e-04
GC_2_222 b_2 NI_2 NS_222 0 1.5569633035190006e-04
GC_2_223 b_2 NI_2 NS_223 0 -6.8565111845632433e-06
GC_2_224 b_2 NI_2 NS_224 0 5.3984649349903595e-06
GC_2_225 b_2 NI_2 NS_225 0 -9.2285333811078729e-05
GC_2_226 b_2 NI_2 NS_226 0 -5.0608525674318874e-05
GC_2_227 b_2 NI_2 NS_227 0 1.3333684336616394e-06
GC_2_228 b_2 NI_2 NS_228 0 -8.2508078747381681e-07
GC_2_229 b_2 NI_2 NS_229 0 -3.2746502079067342e-04
GC_2_230 b_2 NI_2 NS_230 0 2.0147154297703711e-04
GC_2_231 b_2 NI_2 NS_231 0 -4.8480663739177756e-06
GC_2_232 b_2 NI_2 NS_232 0 2.3607231756869185e-05
GC_2_233 b_2 NI_2 NS_233 0 -4.0408717697132722e-06
GC_2_234 b_2 NI_2 NS_234 0 1.4044851740334683e-05
GC_2_235 b_2 NI_2 NS_235 0 4.2754546650300353e-04
GC_2_236 b_2 NI_2 NS_236 0 -2.1230034488666641e-04
GC_2_237 b_2 NI_2 NS_237 0 -5.7389550081172496e-06
GC_2_238 b_2 NI_2 NS_238 0 -1.5729883474631778e-05
GC_2_239 b_2 NI_2 NS_239 0 -5.7896326627681870e-03
GC_2_240 b_2 NI_2 NS_240 0 -2.7497930466310836e-05
GC_2_241 b_2 NI_2 NS_241 0 -2.5204434100312248e-06
GC_2_242 b_2 NI_2 NS_242 0 -7.2602404183262800e-10
GC_2_243 b_2 NI_2 NS_243 0 1.6323979877156268e-03
GC_2_244 b_2 NI_2 NS_244 0 -4.3337486922215215e-03
GC_2_245 b_2 NI_2 NS_245 0 -2.9015460739158574e-04
GC_2_246 b_2 NI_2 NS_246 0 5.8974313625336525e-04
GC_2_247 b_2 NI_2 NS_247 0 7.3788847139375315e-04
GC_2_248 b_2 NI_2 NS_248 0 1.3739475276262122e-03
GC_2_249 b_2 NI_2 NS_249 0 1.7166815775903192e-03
GC_2_250 b_2 NI_2 NS_250 0 -5.7801686894013305e-05
GC_2_251 b_2 NI_2 NS_251 0 -3.0733731778110001e-07
GC_2_252 b_2 NI_2 NS_252 0 6.6872137443764009e-07
GC_2_253 b_2 NI_2 NS_253 0 7.8606292744132300e-06
GC_2_254 b_2 NI_2 NS_254 0 -8.7460138535050083e-05
GC_2_255 b_2 NI_2 NS_255 0 1.9144431467671045e-05
GC_2_256 b_2 NI_2 NS_256 0 4.3309099689978832e-04
GC_2_257 b_2 NI_2 NS_257 0 1.0851083323680588e-05
GC_2_258 b_2 NI_2 NS_258 0 1.3094907606405024e-05
GC_2_259 b_2 NI_2 NS_259 0 -9.0554755709245738e-05
GC_2_260 b_2 NI_2 NS_260 0 -1.0588300647751087e-04
GC_2_261 b_2 NI_2 NS_261 0 -2.7377707698362557e-07
GC_2_262 b_2 NI_2 NS_262 0 -1.4854770998596593e-07
GC_2_263 b_2 NI_2 NS_263 0 -1.2193567196466724e-04
GC_2_264 b_2 NI_2 NS_264 0 2.2194778804342639e-04
GC_2_265 b_2 NI_2 NS_265 0 -3.8811156898902025e-06
GC_2_266 b_2 NI_2 NS_266 0 -1.6252244749457199e-06
GC_2_267 b_2 NI_2 NS_267 0 1.1926466344612608e-07
GC_2_268 b_2 NI_2 NS_268 0 -7.9284292043698305e-06
GC_2_269 b_2 NI_2 NS_269 0 3.2983686805244570e-04
GC_2_270 b_2 NI_2 NS_270 0 -2.2758408605247842e-04
GC_2_271 b_2 NI_2 NS_271 0 -3.3402909283911169e-05
GC_2_272 b_2 NI_2 NS_272 0 5.3566444844200323e-05
GC_2_273 b_2 NI_2 NS_273 0 6.2643030333459559e-03
GC_2_274 b_2 NI_2 NS_274 0 -4.6635244069984425e-04
GC_2_275 b_2 NI_2 NS_275 0 5.2644397786840213e-07
GC_2_276 b_2 NI_2 NS_276 0 8.5732329735157252e-10
GC_2_277 b_2 NI_2 NS_277 0 -4.4023374906994539e-04
GC_2_278 b_2 NI_2 NS_278 0 1.4050092207633902e-03
GC_2_279 b_2 NI_2 NS_279 0 7.1670779615123383e-04
GC_2_280 b_2 NI_2 NS_280 0 -1.6614218074441017e-04
GC_2_281 b_2 NI_2 NS_281 0 -3.5734917940475406e-03
GC_2_282 b_2 NI_2 NS_282 0 -1.3823862435296671e-04
GC_2_283 b_2 NI_2 NS_283 0 8.7967988246101590e-04
GC_2_284 b_2 NI_2 NS_284 0 9.8463304596126643e-04
GC_2_285 b_2 NI_2 NS_285 0 -2.1142383888907148e-06
GC_2_286 b_2 NI_2 NS_286 0 1.1689092228117409e-05
GC_2_287 b_2 NI_2 NS_287 0 4.7477589114343418e-06
GC_2_288 b_2 NI_2 NS_288 0 -1.8050486241737617e-05
GC_2_289 b_2 NI_2 NS_289 0 2.1686576659029217e-04
GC_2_290 b_2 NI_2 NS_290 0 1.6156568867520705e-04
GC_2_291 b_2 NI_2 NS_291 0 -1.6486314380926278e-05
GC_2_292 b_2 NI_2 NS_292 0 1.5243506841843172e-05
GC_2_293 b_2 NI_2 NS_293 0 -2.4229882672371060e-04
GC_2_294 b_2 NI_2 NS_294 0 -1.2113166821211889e-04
GC_2_295 b_2 NI_2 NS_295 0 2.0521152931681823e-06
GC_2_296 b_2 NI_2 NS_296 0 -6.6686304478234738e-07
GC_2_297 b_2 NI_2 NS_297 0 -1.3208029536861731e-04
GC_2_298 b_2 NI_2 NS_298 0 3.1764827266894473e-04
GC_2_299 b_2 NI_2 NS_299 0 -6.6161059227002345e-07
GC_2_300 b_2 NI_2 NS_300 0 1.1199387954725186e-05
GC_2_301 b_2 NI_2 NS_301 0 -1.9951507771819995e-06
GC_2_302 b_2 NI_2 NS_302 0 2.3329564554613439e-05
GC_2_303 b_2 NI_2 NS_303 0 4.2464534274951282e-04
GC_2_304 b_2 NI_2 NS_304 0 -1.5506489125482621e-04
GC_2_305 b_2 NI_2 NS_305 0 -7.3055960645482667e-06
GC_2_306 b_2 NI_2 NS_306 0 -1.4769053423738551e-05
GC_2_307 b_2 NI_2 NS_307 0 -4.6173112964067125e-04
GC_2_308 b_2 NI_2 NS_308 0 -1.1208617505346468e-04
GC_2_309 b_2 NI_2 NS_309 0 -8.0019719883010031e-07
GC_2_310 b_2 NI_2 NS_310 0 -5.5567216346215009e-10
GC_2_311 b_2 NI_2 NS_311 0 1.5551337129657591e-03
GC_2_312 b_2 NI_2 NS_312 0 -1.5631976287212310e-03
GC_2_313 b_2 NI_2 NS_313 0 2.9645586213900298e-04
GC_2_314 b_2 NI_2 NS_314 0 -4.4836037394161159e-04
GC_2_315 b_2 NI_2 NS_315 0 -2.3601669476225975e-03
GC_2_316 b_2 NI_2 NS_316 0 1.9282172305931770e-03
GC_2_317 b_2 NI_2 NS_317 0 1.8153468983205185e-03
GC_2_318 b_2 NI_2 NS_318 0 3.8370445195764916e-04
GC_2_319 b_2 NI_2 NS_319 0 -1.2365186512479392e-05
GC_2_320 b_2 NI_2 NS_320 0 -2.8898136156571199e-06
GC_2_321 b_2 NI_2 NS_321 0 6.9308393482756040e-06
GC_2_322 b_2 NI_2 NS_322 0 -8.9428339921494894e-05
GC_2_323 b_2 NI_2 NS_323 0 1.7788896153279845e-05
GC_2_324 b_2 NI_2 NS_324 0 4.4732108414555590e-04
GC_2_325 b_2 NI_2 NS_325 0 2.6645754409418229e-05
GC_2_326 b_2 NI_2 NS_326 0 5.5947523404033525e-06
GC_2_327 b_2 NI_2 NS_327 0 -2.4952494090434510e-04
GC_2_328 b_2 NI_2 NS_328 0 -1.7932622787370721e-04
GC_2_329 b_2 NI_2 NS_329 0 -9.2902838594549157e-08
GC_2_330 b_2 NI_2 NS_330 0 2.8214125476651691e-06
GC_2_331 b_2 NI_2 NS_331 0 1.4313751587668671e-05
GC_2_332 b_2 NI_2 NS_332 0 2.3791382993152807e-04
GC_2_333 b_2 NI_2 NS_333 0 6.7360423483810046e-07
GC_2_334 b_2 NI_2 NS_334 0 2.4254125658450884e-06
GC_2_335 b_2 NI_2 NS_335 0 2.2085230457695050e-06
GC_2_336 b_2 NI_2 NS_336 0 -1.3837913852233681e-05
GC_2_337 b_2 NI_2 NS_337 0 3.1315540108957954e-04
GC_2_338 b_2 NI_2 NS_338 0 -2.0751176472124077e-04
GC_2_339 b_2 NI_2 NS_339 0 -3.0450876876356135e-05
GC_2_340 b_2 NI_2 NS_340 0 4.6772907033801304e-05
GC_2_341 b_2 NI_2 NS_341 0 7.0745965332746326e-03
GC_2_342 b_2 NI_2 NS_342 0 -4.6533964544764384e-04
GC_2_343 b_2 NI_2 NS_343 0 7.9558583950628667e-07
GC_2_344 b_2 NI_2 NS_344 0 2.7021860213735746e-10
GC_2_345 b_2 NI_2 NS_345 0 5.8203079945171174e-04
GC_2_346 b_2 NI_2 NS_346 0 1.6089572296772159e-03
GC_2_347 b_2 NI_2 NS_347 0 1.4710529782290410e-03
GC_2_348 b_2 NI_2 NS_348 0 -1.3561538919308696e-03
GC_2_349 b_2 NI_2 NS_349 0 -6.8784146895513381e-03
GC_2_350 b_2 NI_2 NS_350 0 6.8762290065519857e-04
GC_2_351 b_2 NI_2 NS_351 0 1.7513892184711820e-03
GC_2_352 b_2 NI_2 NS_352 0 2.1300702587493414e-03
GC_2_353 b_2 NI_2 NS_353 0 -1.2009240721659044e-06
GC_2_354 b_2 NI_2 NS_354 0 1.2906686287505498e-05
GC_2_355 b_2 NI_2 NS_355 0 3.9210510142348941e-06
GC_2_356 b_2 NI_2 NS_356 0 -1.6465798758076340e-05
GC_2_357 b_2 NI_2 NS_357 0 2.1124397459282572e-04
GC_2_358 b_2 NI_2 NS_358 0 1.5297126786804606e-04
GC_2_359 b_2 NI_2 NS_359 0 -2.4085319515609582e-05
GC_2_360 b_2 NI_2 NS_360 0 1.7724140247805053e-05
GC_2_361 b_2 NI_2 NS_361 0 -3.2648903707968992e-04
GC_2_362 b_2 NI_2 NS_362 0 -1.6305722216264736e-04
GC_2_363 b_2 NI_2 NS_363 0 1.3020936135731586e-07
GC_2_364 b_2 NI_2 NS_364 0 -3.6100324271855756e-07
GC_2_365 b_2 NI_2 NS_365 0 5.9197033570109594e-06
GC_2_366 b_2 NI_2 NS_366 0 3.7180671606473027e-04
GC_2_367 b_2 NI_2 NS_367 0 2.0490347592832806e-06
GC_2_368 b_2 NI_2 NS_368 0 -2.2602787331038175e-06
GC_2_369 b_2 NI_2 NS_369 0 -7.6497684958098090e-06
GC_2_370 b_2 NI_2 NS_370 0 3.1776633370321741e-05
GC_2_371 b_2 NI_2 NS_371 0 4.8282715419701119e-04
GC_2_372 b_2 NI_2 NS_372 0 -1.4040043237279791e-04
GC_2_373 b_2 NI_2 NS_373 0 -9.6615558250150400e-06
GC_2_374 b_2 NI_2 NS_374 0 -1.6431033988288609e-05
GC_2_375 b_2 NI_2 NS_375 0 2.4229917486743068e-03
GC_2_376 b_2 NI_2 NS_376 0 -9.8386083651892274e-05
GC_2_377 b_2 NI_2 NS_377 0 -4.3918588400225597e-07
GC_2_378 b_2 NI_2 NS_378 0 -2.3795368037009932e-10
GC_2_379 b_2 NI_2 NS_379 0 1.9634686358312825e-03
GC_2_380 b_2 NI_2 NS_380 0 -3.3510140910321726e-04
GC_2_381 b_2 NI_2 NS_381 0 5.4668581571556659e-04
GC_2_382 b_2 NI_2 NS_382 0 -1.2699744739749373e-03
GC_2_383 b_2 NI_2 NS_383 0 -4.6180370717010350e-03
GC_2_384 b_2 NI_2 NS_384 0 2.4918473347623304e-03
GC_2_385 b_2 NI_2 NS_385 0 2.2235353422522448e-03
GC_2_386 b_2 NI_2 NS_386 0 1.4004576540005550e-03
GC_2_387 b_2 NI_2 NS_387 0 -1.4840253418448835e-05
GC_2_388 b_2 NI_2 NS_388 0 -5.1143436791844770e-06
GC_2_389 b_2 NI_2 NS_389 0 7.9411387917114686e-06
GC_2_390 b_2 NI_2 NS_390 0 -8.5623185787044877e-05
GC_2_391 b_2 NI_2 NS_391 0 5.9387476085278704e-06
GC_2_392 b_2 NI_2 NS_392 0 4.2775703462745755e-04
GC_2_393 b_2 NI_2 NS_393 0 3.8912322371223130e-05
GC_2_394 b_2 NI_2 NS_394 0 2.2642834863453080e-05
GC_2_395 b_2 NI_2 NS_395 0 -3.2645316557399200e-04
GC_2_396 b_2 NI_2 NS_396 0 -3.0819343960575599e-04
GC_2_397 b_2 NI_2 NS_397 0 1.8761244718455248e-08
GC_2_398 b_2 NI_2 NS_398 0 1.7867164325333027e-07
GC_2_399 b_2 NI_2 NS_399 0 7.5346705127689385e-05
GC_2_400 b_2 NI_2 NS_400 0 2.4783108591084545e-04
GC_2_401 b_2 NI_2 NS_401 0 4.4739637087097636e-06
GC_2_402 b_2 NI_2 NS_402 0 1.0116692952580731e-05
GC_2_403 b_2 NI_2 NS_403 0 1.3524351932588264e-06
GC_2_404 b_2 NI_2 NS_404 0 -2.3185504240116467e-05
GC_2_405 b_2 NI_2 NS_405 0 3.3336081576961499e-04
GC_2_406 b_2 NI_2 NS_406 0 -2.1080812504551294e-04
GC_2_407 b_2 NI_2 NS_407 0 -3.2992078930877376e-05
GC_2_408 b_2 NI_2 NS_408 0 4.6785746683792454e-05
GD_2_1 b_2 NI_2 NA_1 0 -3.4437674971680821e-02
GD_2_2 b_2 NI_2 NA_2 0 -2.5209745917522192e-01
GD_2_3 b_2 NI_2 NA_3 0 -9.6256403331112760e-03
GD_2_4 b_2 NI_2 NA_4 0 7.0252725790054217e-03
GD_2_5 b_2 NI_2 NA_5 0 -6.6284202906489124e-03
GD_2_6 b_2 NI_2 NA_6 0 2.9032615388974170e-03
GD_2_7 b_2 NI_2 NA_7 0 -5.3303552120016326e-03
GD_2_8 b_2 NI_2 NA_8 0 1.6709457763681255e-03
GD_2_9 b_2 NI_2 NA_9 0 -5.1900717912031543e-03
GD_2_10 b_2 NI_2 NA_10 0 -1.5923225299925502e-03
GD_2_11 b_2 NI_2 NA_11 0 -4.8175188613905490e-03
GD_2_12 b_2 NI_2 NA_12 0 -3.5936774311335186e-03
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 -3.1657117757508395e-02
GC_3_2 b_3 NI_3 NS_2 0 3.1159948135554712e-03
GC_3_3 b_3 NI_3 NS_3 0 -1.5426912488858834e-05
GC_3_4 b_3 NI_3 NS_4 0 -5.7358684544272579e-09
GC_3_5 b_3 NI_3 NS_5 0 1.0270010073742059e-02
GC_3_6 b_3 NI_3 NS_6 0 -9.5200833260637510e-03
GC_3_7 b_3 NI_3 NS_7 0 -1.9101992232935891e-03
GC_3_8 b_3 NI_3 NS_8 0 2.9132725522751406e-04
GC_3_9 b_3 NI_3 NS_9 0 5.1554692831192019e-03
GC_3_10 b_3 NI_3 NS_10 0 3.4628277995554335e-03
GC_3_11 b_3 NI_3 NS_11 0 1.8666619998889561e-03
GC_3_12 b_3 NI_3 NS_12 0 -1.9705667738551281e-04
GC_3_13 b_3 NI_3 NS_13 0 -1.0059794431861403e-05
GC_3_14 b_3 NI_3 NS_14 0 2.1296774084557837e-06
GC_3_15 b_3 NI_3 NS_15 0 2.2299472636128771e-06
GC_3_16 b_3 NI_3 NS_16 0 -3.8458737448121965e-06
GC_3_17 b_3 NI_3 NS_17 0 1.5685599857109196e-04
GC_3_18 b_3 NI_3 NS_18 0 -3.8577870066370100e-05
GC_3_19 b_3 NI_3 NS_19 0 3.7221189803450725e-06
GC_3_20 b_3 NI_3 NS_20 0 1.5529487456155478e-05
GC_3_21 b_3 NI_3 NS_21 0 1.9027272068303878e-04
GC_3_22 b_3 NI_3 NS_22 0 -6.9065612294176880e-06
GC_3_23 b_3 NI_3 NS_23 0 7.6357266655795430e-07
GC_3_24 b_3 NI_3 NS_24 0 2.2263199888623048e-06
GC_3_25 b_3 NI_3 NS_25 0 8.1868982386856199e-05
GC_3_26 b_3 NI_3 NS_26 0 -3.6498798093902065e-04
GC_3_27 b_3 NI_3 NS_27 0 1.1751037517230032e-05
GC_3_28 b_3 NI_3 NS_28 0 -1.7260292613885041e-05
GC_3_29 b_3 NI_3 NS_29 0 -3.1467618332847539e-06
GC_3_30 b_3 NI_3 NS_30 0 1.7248353022619263e-05
GC_3_31 b_3 NI_3 NS_31 0 4.4073178307715865e-04
GC_3_32 b_3 NI_3 NS_32 0 8.2753910937013306e-05
GC_3_33 b_3 NI_3 NS_33 0 3.0246263327949095e-06
GC_3_34 b_3 NI_3 NS_34 0 -1.7723127948143982e-06
GC_3_35 b_3 NI_3 NS_35 0 2.9370522203007125e-02
GC_3_36 b_3 NI_3 NS_36 0 -3.2161763072070795e-03
GC_3_37 b_3 NI_3 NS_37 0 -2.7622716728261531e-06
GC_3_38 b_3 NI_3 NS_38 0 9.7841499432227165e-09
GC_3_39 b_3 NI_3 NS_39 0 -1.4937047353908750e-02
GC_3_40 b_3 NI_3 NS_40 0 1.0982326490676089e-02
GC_3_41 b_3 NI_3 NS_41 0 9.3482938207771737e-05
GC_3_42 b_3 NI_3 NS_42 0 1.0424910912318851e-03
GC_3_43 b_3 NI_3 NS_43 0 3.9531746181320172e-03
GC_3_44 b_3 NI_3 NS_44 0 -8.3909697451751263e-03
GC_3_45 b_3 NI_3 NS_45 0 -7.8011652539187858e-03
GC_3_46 b_3 NI_3 NS_46 0 -2.4381531061268354e-03
GC_3_47 b_3 NI_3 NS_47 0 1.6886031528493663e-06
GC_3_48 b_3 NI_3 NS_48 0 -9.2850266963327123e-06
GC_3_49 b_3 NI_3 NS_49 0 5.4564605108785768e-06
GC_3_50 b_3 NI_3 NS_50 0 -1.7383572019839969e-05
GC_3_51 b_3 NI_3 NS_51 0 2.0973515263258995e-04
GC_3_52 b_3 NI_3 NS_52 0 1.5912617355570282e-04
GC_3_53 b_3 NI_3 NS_53 0 1.5865633971151659e-05
GC_3_54 b_3 NI_3 NS_54 0 -1.1907141014102599e-05
GC_3_55 b_3 NI_3 NS_55 0 2.1264910626884892e-04
GC_3_56 b_3 NI_3 NS_56 0 9.4137013561850072e-05
GC_3_57 b_3 NI_3 NS_57 0 4.4275834541720325e-06
GC_3_58 b_3 NI_3 NS_58 0 -3.4145374084170214e-07
GC_3_59 b_3 NI_3 NS_59 0 -1.3542606351372232e-04
GC_3_60 b_3 NI_3 NS_60 0 -3.3941687203123248e-04
GC_3_61 b_3 NI_3 NS_61 0 -8.4839355767365829e-06
GC_3_62 b_3 NI_3 NS_62 0 4.5246781818230666e-06
GC_3_63 b_3 NI_3 NS_63 0 -8.3044336409237884e-10
GC_3_64 b_3 NI_3 NS_64 0 -1.6739718101966955e-05
GC_3_65 b_3 NI_3 NS_65 0 2.8283216418212217e-04
GC_3_66 b_3 NI_3 NS_66 0 -1.8003605427310138e-04
GC_3_67 b_3 NI_3 NS_67 0 -6.3176618693979684e-06
GC_3_68 b_3 NI_3 NS_68 0 -1.6913493780313772e-05
GC_3_69 b_3 NI_3 NS_69 0 -2.2863723288039062e-01
GC_3_70 b_3 NI_3 NS_70 0 5.7019950544015652e-02
GC_3_71 b_3 NI_3 NS_71 0 3.4993239880630193e-05
GC_3_72 b_3 NI_3 NS_72 0 -5.4777939538711366e-08
GC_3_73 b_3 NI_3 NS_73 0 8.5039250860860768e-02
GC_3_74 b_3 NI_3 NS_74 0 2.3147362872968230e-03
GC_3_75 b_3 NI_3 NS_75 0 9.2182115844725431e-04
GC_3_76 b_3 NI_3 NS_76 0 1.8190613745658910e-03
GC_3_77 b_3 NI_3 NS_77 0 2.5182122690364972e-03
GC_3_78 b_3 NI_3 NS_78 0 7.2892234500414408e-03
GC_3_79 b_3 NI_3 NS_79 0 -3.7744417432746028e-03
GC_3_80 b_3 NI_3 NS_80 0 4.0982639544739092e-03
GC_3_81 b_3 NI_3 NS_81 0 -8.0029252937999178e-06
GC_3_82 b_3 NI_3 NS_82 0 3.6778392007231163e-06
GC_3_83 b_3 NI_3 NS_83 0 3.5302330643724880e-06
GC_3_84 b_3 NI_3 NS_84 0 -3.6287407451989922e-06
GC_3_85 b_3 NI_3 NS_85 0 1.4685371368891703e-04
GC_3_86 b_3 NI_3 NS_86 0 -4.6461707087721289e-05
GC_3_87 b_3 NI_3 NS_87 0 4.3219352698077899e-06
GC_3_88 b_3 NI_3 NS_88 0 7.4079997894560663e-06
GC_3_89 b_3 NI_3 NS_89 0 1.2388336159877754e-04
GC_3_90 b_3 NI_3 NS_90 0 9.6434516584336138e-06
GC_3_91 b_3 NI_3 NS_91 0 8.5798816608085647e-06
GC_3_92 b_3 NI_3 NS_92 0 9.0206517659612411e-06
GC_3_93 b_3 NI_3 NS_93 0 1.8130929021689993e-04
GC_3_94 b_3 NI_3 NS_94 0 -2.6159807050808807e-04
GC_3_95 b_3 NI_3 NS_95 0 -1.5784081491820274e-05
GC_3_96 b_3 NI_3 NS_96 0 1.3269459896287784e-06
GC_3_97 b_3 NI_3 NS_97 0 -4.0285556160230622e-07
GC_3_98 b_3 NI_3 NS_98 0 1.3306032025631258e-05
GC_3_99 b_3 NI_3 NS_99 0 3.7617602086522810e-04
GC_3_100 b_3 NI_3 NS_100 0 4.1011914338179406e-05
GC_3_101 b_3 NI_3 NS_101 0 4.2676244613633493e-06
GC_3_102 b_3 NI_3 NS_102 0 -1.2354960392477773e-06
GC_3_103 b_3 NI_3 NS_103 0 2.4153574019465759e-02
GC_3_104 b_3 NI_3 NS_104 0 3.4113441834442655e-02
GC_3_105 b_3 NI_3 NS_105 0 1.5538821673079565e-04
GC_3_106 b_3 NI_3 NS_106 0 2.7164887541789786e-07
GC_3_107 b_3 NI_3 NS_107 0 -5.7083046540564467e-02
GC_3_108 b_3 NI_3 NS_108 0 -2.0359477079490741e-02
GC_3_109 b_3 NI_3 NS_109 0 -8.3340879484709938e-04
GC_3_110 b_3 NI_3 NS_110 0 4.5815200088597744e-03
GC_3_111 b_3 NI_3 NS_111 0 9.5948955766218518e-03
GC_3_112 b_3 NI_3 NS_112 0 1.8374942527255481e-02
GC_3_113 b_3 NI_3 NS_113 0 1.0676602707385022e-02
GC_3_114 b_3 NI_3 NS_114 0 1.5782093350953665e-03
GC_3_115 b_3 NI_3 NS_115 0 -3.5966754946020723e-07
GC_3_116 b_3 NI_3 NS_116 0 -8.1905976674332100e-06
GC_3_117 b_3 NI_3 NS_117 0 3.5730132929068854e-06
GC_3_118 b_3 NI_3 NS_118 0 -1.8337433254482916e-05
GC_3_119 b_3 NI_3 NS_119 0 2.3904684266906441e-04
GC_3_120 b_3 NI_3 NS_120 0 1.6136187959046939e-04
GC_3_121 b_3 NI_3 NS_121 0 7.5552583145700639e-06
GC_3_122 b_3 NI_3 NS_122 0 -1.0381676665669700e-05
GC_3_123 b_3 NI_3 NS_123 0 1.7938391659878496e-04
GC_3_124 b_3 NI_3 NS_124 0 4.0757853550050168e-05
GC_3_125 b_3 NI_3 NS_125 0 9.8936344564279669e-06
GC_3_126 b_3 NI_3 NS_126 0 -1.1970241580643022e-06
GC_3_127 b_3 NI_3 NS_127 0 1.3664941069233349e-04
GC_3_128 b_3 NI_3 NS_128 0 -2.5915661808407787e-04
GC_3_129 b_3 NI_3 NS_129 0 -3.6704441983276794e-06
GC_3_130 b_3 NI_3 NS_130 0 -1.1067836993169835e-05
GC_3_131 b_3 NI_3 NS_131 0 -6.4559234562571338e-07
GC_3_132 b_3 NI_3 NS_132 0 -1.3010790722563894e-05
GC_3_133 b_3 NI_3 NS_133 0 3.9174723114269511e-04
GC_3_134 b_3 NI_3 NS_134 0 -3.3277527051566277e-05
GC_3_135 b_3 NI_3 NS_135 0 -8.9518129753282191e-06
GC_3_136 b_3 NI_3 NS_136 0 -1.6433883711657975e-05
GC_3_137 b_3 NI_3 NS_137 0 -1.7988308561269293e-02
GC_3_138 b_3 NI_3 NS_138 0 2.1699347258428933e-03
GC_3_139 b_3 NI_3 NS_139 0 -6.6258503152992235e-06
GC_3_140 b_3 NI_3 NS_140 0 -4.2996878687810789e-09
GC_3_141 b_3 NI_3 NS_141 0 5.4814728198173167e-03
GC_3_142 b_3 NI_3 NS_142 0 -4.4066954945721909e-03
GC_3_143 b_3 NI_3 NS_143 0 7.6074209005561012e-04
GC_3_144 b_3 NI_3 NS_144 0 4.5990183160508484e-04
GC_3_145 b_3 NI_3 NS_145 0 2.5334403294301590e-04
GC_3_146 b_3 NI_3 NS_146 0 -3.9557310379306282e-04
GC_3_147 b_3 NI_3 NS_147 0 1.2502222137282448e-03
GC_3_148 b_3 NI_3 NS_148 0 6.0862049130588230e-04
GC_3_149 b_3 NI_3 NS_149 0 4.0974455766254507e-07
GC_3_150 b_3 NI_3 NS_150 0 -2.8059484855499151e-06
GC_3_151 b_3 NI_3 NS_151 0 1.6384731380644622e-06
GC_3_152 b_3 NI_3 NS_152 0 -3.9550075009900925e-06
GC_3_153 b_3 NI_3 NS_153 0 1.6311331941021529e-04
GC_3_154 b_3 NI_3 NS_154 0 -4.4407222773175412e-05
GC_3_155 b_3 NI_3 NS_155 0 5.5300333223925817e-07
GC_3_156 b_3 NI_3 NS_156 0 3.3485650924491363e-06
GC_3_157 b_3 NI_3 NS_157 0 3.0871233032454359e-05
GC_3_158 b_3 NI_3 NS_158 0 -1.0358839781530930e-05
GC_3_159 b_3 NI_3 NS_159 0 2.3495751483790722e-06
GC_3_160 b_3 NI_3 NS_160 0 3.7407058430685886e-06
GC_3_161 b_3 NI_3 NS_161 0 4.3100676859597376e-04
GC_3_162 b_3 NI_3 NS_162 0 -9.3737008995038805e-05
GC_3_163 b_3 NI_3 NS_163 0 -3.2130285924590013e-05
GC_3_164 b_3 NI_3 NS_164 0 7.9641338794722720e-06
GC_3_165 b_3 NI_3 NS_165 0 -2.0462564694764825e-06
GC_3_166 b_3 NI_3 NS_166 0 2.5258388673542843e-06
GC_3_167 b_3 NI_3 NS_167 0 5.5498322400417881e-04
GC_3_168 b_3 NI_3 NS_168 0 6.9387169684034650e-05
GC_3_169 b_3 NI_3 NS_169 0 1.0955904194669451e-06
GC_3_170 b_3 NI_3 NS_170 0 -1.9584958873595123e-07
GC_3_171 b_3 NI_3 NS_171 0 2.4281996779761821e-02
GC_3_172 b_3 NI_3 NS_172 0 -1.9476110494428328e-03
GC_3_173 b_3 NI_3 NS_173 0 -1.6180031917497762e-06
GC_3_174 b_3 NI_3 NS_174 0 7.3122406457547198e-09
GC_3_175 b_3 NI_3 NS_175 0 -6.7212766715831996e-03
GC_3_176 b_3 NI_3 NS_176 0 9.7809334996590610e-03
GC_3_177 b_3 NI_3 NS_177 0 1.5286347352414385e-03
GC_3_178 b_3 NI_3 NS_178 0 -8.3858689792331036e-04
GC_3_179 b_3 NI_3 NS_179 0 -4.9878050104326709e-03
GC_3_180 b_3 NI_3 NS_180 0 -5.9445639401112917e-03
GC_3_181 b_3 NI_3 NS_181 0 -4.8684732795332029e-03
GC_3_182 b_3 NI_3 NS_182 0 2.0734958115279532e-03
GC_3_183 b_3 NI_3 NS_183 0 -3.6686143785943824e-07
GC_3_184 b_3 NI_3 NS_184 0 -4.4756343168594027e-07
GC_3_185 b_3 NI_3 NS_185 0 5.3414430461050523e-06
GC_3_186 b_3 NI_3 NS_186 0 -1.8401455758533885e-05
GC_3_187 b_3 NI_3 NS_187 0 2.2054589661227794e-04
GC_3_188 b_3 NI_3 NS_188 0 1.5572914576443547e-04
GC_3_189 b_3 NI_3 NS_189 0 5.3297366771012797e-06
GC_3_190 b_3 NI_3 NS_190 0 -1.3838197230834843e-06
GC_3_191 b_3 NI_3 NS_191 0 2.8854638660833788e-05
GC_3_192 b_3 NI_3 NS_192 0 2.0729405322491073e-05
GC_3_193 b_3 NI_3 NS_193 0 5.0055942122935737e-06
GC_3_194 b_3 NI_3 NS_194 0 -3.6969473328624445e-07
GC_3_195 b_3 NI_3 NS_195 0 2.0210339141725402e-04
GC_3_196 b_3 NI_3 NS_196 0 -1.4138930233527670e-04
GC_3_197 b_3 NI_3 NS_197 0 -1.3115632901183859e-06
GC_3_198 b_3 NI_3 NS_198 0 -1.7211248053411336e-05
GC_3_199 b_3 NI_3 NS_199 0 -1.8374434733432277e-06
GC_3_200 b_3 NI_3 NS_200 0 -7.5555487547511848e-06
GC_3_201 b_3 NI_3 NS_201 0 3.7706640009316157e-04
GC_3_202 b_3 NI_3 NS_202 0 -1.3393097500776047e-04
GC_3_203 b_3 NI_3 NS_203 0 -9.7619360895116050e-06
GC_3_204 b_3 NI_3 NS_204 0 -1.7941821729682132e-05
GC_3_205 b_3 NI_3 NS_205 0 -1.2182969228988807e-02
GC_3_206 b_3 NI_3 NS_206 0 1.5127463562491957e-03
GC_3_207 b_3 NI_3 NS_207 0 -3.3241719780191096e-06
GC_3_208 b_3 NI_3 NS_208 0 -2.1976785160500734e-09
GC_3_209 b_3 NI_3 NS_209 0 2.9892912092979668e-03
GC_3_210 b_3 NI_3 NS_210 0 -2.4636885890959568e-03
GC_3_211 b_3 NI_3 NS_211 0 4.8879451525962302e-04
GC_3_212 b_3 NI_3 NS_212 0 -9.6542737656613741e-05
GC_3_213 b_3 NI_3 NS_213 0 -1.0400653824845292e-03
GC_3_214 b_3 NI_3 NS_214 0 -4.3708540384419564e-04
GC_3_215 b_3 NI_3 NS_215 0 1.1709985883047122e-03
GC_3_216 b_3 NI_3 NS_216 0 1.7045220385948940e-04
GC_3_217 b_3 NI_3 NS_217 0 2.9974081723653814e-07
GC_3_218 b_3 NI_3 NS_218 0 1.3651905644299013e-06
GC_3_219 b_3 NI_3 NS_219 0 1.6036026259832133e-06
GC_3_220 b_3 NI_3 NS_220 0 -3.7533198859083816e-06
GC_3_221 b_3 NI_3 NS_221 0 1.6137306375868356e-04
GC_3_222 b_3 NI_3 NS_222 0 -4.7713925459401349e-05
GC_3_223 b_3 NI_3 NS_223 0 -9.3179770150438731e-07
GC_3_224 b_3 NI_3 NS_224 0 -5.3192010391803357e-06
GC_3_225 b_3 NI_3 NS_225 0 -5.6222236101709694e-05
GC_3_226 b_3 NI_3 NS_226 0 -5.3174169549608365e-06
GC_3_227 b_3 NI_3 NS_227 0 2.7875372590343291e-06
GC_3_228 b_3 NI_3 NS_228 0 3.7719154432180725e-06
GC_3_229 b_3 NI_3 NS_229 0 2.2642360114855008e-04
GC_3_230 b_3 NI_3 NS_230 0 1.1810400039119380e-04
GC_3_231 b_3 NI_3 NS_231 0 -3.0719019068305686e-05
GC_3_232 b_3 NI_3 NS_232 0 1.3608512373027467e-05
GC_3_233 b_3 NI_3 NS_233 0 2.4674888059328027e-06
GC_3_234 b_3 NI_3 NS_234 0 -7.8408044786287796e-06
GC_3_235 b_3 NI_3 NS_235 0 5.9446189885350650e-04
GC_3_236 b_3 NI_3 NS_236 0 1.8328745161828219e-05
GC_3_237 b_3 NI_3 NS_237 0 1.8685430332392772e-06
GC_3_238 b_3 NI_3 NS_238 0 8.0899737166776477e-07
GC_3_239 b_3 NI_3 NS_239 0 1.9539864611530722e-02
GC_3_240 b_3 NI_3 NS_240 0 -1.4587579686731692e-03
GC_3_241 b_3 NI_3 NS_241 0 5.0631612550396456e-07
GC_3_242 b_3 NI_3 NS_242 0 3.5449491039195167e-09
GC_3_243 b_3 NI_3 NS_243 0 -2.8896458549953542e-03
GC_3_244 b_3 NI_3 NS_244 0 6.9183056891905593e-03
GC_3_245 b_3 NI_3 NS_245 0 6.4936763796171414e-04
GC_3_246 b_3 NI_3 NS_246 0 -1.0592189914524436e-03
GC_3_247 b_3 NI_3 NS_247 0 -5.9460610307966429e-03
GC_3_248 b_3 NI_3 NS_248 0 -2.6288933310616297e-03
GC_3_249 b_3 NI_3 NS_249 0 -2.2281767970423385e-03
GC_3_250 b_3 NI_3 NS_250 0 2.7254518507661449e-03
GC_3_251 b_3 NI_3 NS_251 0 1.4086371643842369e-06
GC_3_252 b_3 NI_3 NS_252 0 4.8155759468492565e-07
GC_3_253 b_3 NI_3 NS_253 0 4.8716948424988668e-06
GC_3_254 b_3 NI_3 NS_254 0 -1.8248516158585497e-05
GC_3_255 b_3 NI_3 NS_255 0 2.2516092969099001e-04
GC_3_256 b_3 NI_3 NS_256 0 1.5520201555126141e-04
GC_3_257 b_3 NI_3 NS_257 0 -6.1722617554448537e-06
GC_3_258 b_3 NI_3 NS_258 0 6.6588212551494035e-07
GC_3_259 b_3 NI_3 NS_259 0 -4.6945677380748490e-05
GC_3_260 b_3 NI_3 NS_260 0 -2.4503295198768362e-05
GC_3_261 b_3 NI_3 NS_261 0 5.3163392679009403e-06
GC_3_262 b_3 NI_3 NS_262 0 -9.3506091399803344e-07
GC_3_263 b_3 NI_3 NS_263 0 1.3689602798587464e-04
GC_3_264 b_3 NI_3 NS_264 0 5.5135393206939088e-05
GC_3_265 b_3 NI_3 NS_265 0 -3.6746161124000197e-07
GC_3_266 b_3 NI_3 NS_266 0 -1.3497485687007430e-05
GC_3_267 b_3 NI_3 NS_267 0 -1.3785368525450560e-06
GC_3_268 b_3 NI_3 NS_268 0 6.6746579790493244e-06
GC_3_269 b_3 NI_3 NS_269 0 4.0169371322016083e-04
GC_3_270 b_3 NI_3 NS_270 0 -1.4649294247969137e-04
GC_3_271 b_3 NI_3 NS_271 0 -9.3748914465049285e-06
GC_3_272 b_3 NI_3 NS_272 0 -1.7858700642782657e-05
GC_3_273 b_3 NI_3 NS_273 0 1.0790889971644901e-03
GC_3_274 b_3 NI_3 NS_274 0 3.6986605813070245e-04
GC_3_275 b_3 NI_3 NS_275 0 -7.4221768883144274e-07
GC_3_276 b_3 NI_3 NS_276 0 -1.1520770632236326e-09
GC_3_277 b_3 NI_3 NS_277 0 2.5188278993296953e-03
GC_3_278 b_3 NI_3 NS_278 0 8.3574185049936341e-04
GC_3_279 b_3 NI_3 NS_279 0 9.4959848342309665e-04
GC_3_280 b_3 NI_3 NS_280 0 -6.6482076006255596e-04
GC_3_281 b_3 NI_3 NS_281 0 -7.3156004179463783e-03
GC_3_282 b_3 NI_3 NS_282 0 -8.6890688802976508e-04
GC_3_283 b_3 NI_3 NS_283 0 2.4824479535484364e-03
GC_3_284 b_3 NI_3 NS_284 0 2.9941122875905184e-03
GC_3_285 b_3 NI_3 NS_285 0 9.5599116680565133e-06
GC_3_286 b_3 NI_3 NS_286 0 -2.8930231677559654e-06
GC_3_287 b_3 NI_3 NS_287 0 1.5618302927671878e-06
GC_3_288 b_3 NI_3 NS_288 0 -3.3663602023493332e-06
GC_3_289 b_3 NI_3 NS_289 0 1.6490364942202198e-04
GC_3_290 b_3 NI_3 NS_290 0 -4.8937687389983200e-05
GC_3_291 b_3 NI_3 NS_291 0 -1.9579644001512383e-06
GC_3_292 b_3 NI_3 NS_292 0 -1.1770668325909755e-05
GC_3_293 b_3 NI_3 NS_293 0 -1.7597065964091647e-04
GC_3_294 b_3 NI_3 NS_294 0 -2.7651154178221741e-06
GC_3_295 b_3 NI_3 NS_295 0 5.2963551405886423e-06
GC_3_296 b_3 NI_3 NS_296 0 1.0703069222050695e-05
GC_3_297 b_3 NI_3 NS_297 0 -4.0449058480004183e-05
GC_3_298 b_3 NI_3 NS_298 0 3.3603200152406310e-04
GC_3_299 b_3 NI_3 NS_299 0 -4.8728454200754302e-06
GC_3_300 b_3 NI_3 NS_300 0 6.8159908381299031e-06
GC_3_301 b_3 NI_3 NS_301 0 3.1009172998685184e-06
GC_3_302 b_3 NI_3 NS_302 0 -1.5270704235887292e-05
GC_3_303 b_3 NI_3 NS_303 0 5.1361892175329096e-04
GC_3_304 b_3 NI_3 NS_304 0 9.9783709623546925e-05
GC_3_305 b_3 NI_3 NS_305 0 2.0115067301695144e-06
GC_3_306 b_3 NI_3 NS_306 0 -1.2198646383060137e-06
GC_3_307 b_3 NI_3 NS_307 0 1.2357086339855581e-02
GC_3_308 b_3 NI_3 NS_308 0 -8.3524087854587928e-04
GC_3_309 b_3 NI_3 NS_309 0 7.9833571176064151e-07
GC_3_310 b_3 NI_3 NS_310 0 1.3506172179123577e-09
GC_3_311 b_3 NI_3 NS_311 0 -3.3438270750758424e-04
GC_3_312 b_3 NI_3 NS_312 0 3.1464948150181672e-03
GC_3_313 b_3 NI_3 NS_313 0 5.4102972439530887e-04
GC_3_314 b_3 NI_3 NS_314 0 -8.2844812342152080e-04
GC_3_315 b_3 NI_3 NS_315 0 -6.5662373248325497e-03
GC_3_316 b_3 NI_3 NS_316 0 1.8740076985933069e-04
GC_3_317 b_3 NI_3 NS_317 0 1.2913378079246118e-03
GC_3_318 b_3 NI_3 NS_318 0 2.4130251996781174e-03
GC_3_319 b_3 NI_3 NS_319 0 -5.9103006914250901e-07
GC_3_320 b_3 NI_3 NS_320 0 8.0114927769721748e-06
GC_3_321 b_3 NI_3 NS_321 0 4.9765819192984352e-06
GC_3_322 b_3 NI_3 NS_322 0 -1.8625746490943209e-05
GC_3_323 b_3 NI_3 NS_323 0 2.2553292365912918e-04
GC_3_324 b_3 NI_3 NS_324 0 1.5925064755759356e-04
GC_3_325 b_3 NI_3 NS_325 0 -6.9114931478369402e-06
GC_3_326 b_3 NI_3 NS_326 0 1.1731554776897529e-05
GC_3_327 b_3 NI_3 NS_327 0 -2.0665041067015739e-04
GC_3_328 b_3 NI_3 NS_328 0 -7.2190629439801752e-05
GC_3_329 b_3 NI_3 NS_329 0 1.0482418841015882e-05
GC_3_330 b_3 NI_3 NS_330 0 -4.2889886801568430e-07
GC_3_331 b_3 NI_3 NS_331 0 6.1794823611424448e-05
GC_3_332 b_3 NI_3 NS_332 0 2.3789647674355311e-04
GC_3_333 b_3 NI_3 NS_333 0 2.0787884987935656e-06
GC_3_334 b_3 NI_3 NS_334 0 -3.3484113371032600e-06
GC_3_335 b_3 NI_3 NS_335 0 -1.5157136751309260e-06
GC_3_336 b_3 NI_3 NS_336 0 1.0569425662517569e-05
GC_3_337 b_3 NI_3 NS_337 0 3.6571859357000978e-04
GC_3_338 b_3 NI_3 NS_338 0 -9.1099376693094526e-05
GC_3_339 b_3 NI_3 NS_339 0 -8.1607272119721009e-06
GC_3_340 b_3 NI_3 NS_340 0 -1.6472603763361956e-05
GC_3_341 b_3 NI_3 NS_341 0 4.7652784139005089e-03
GC_3_342 b_3 NI_3 NS_342 0 -3.6921304758992362e-05
GC_3_343 b_3 NI_3 NS_343 0 2.5169146273236444e-07
GC_3_344 b_3 NI_3 NS_344 0 -8.9150570836021315e-10
GC_3_345 b_3 NI_3 NS_345 0 1.7124153833516860e-03
GC_3_346 b_3 NI_3 NS_346 0 1.5475794148264066e-03
GC_3_347 b_3 NI_3 NS_347 0 7.4430431749143776e-04
GC_3_348 b_3 NI_3 NS_348 0 -1.6023125801478393e-04
GC_3_349 b_3 NI_3 NS_349 0 -5.5314485356319403e-03
GC_3_350 b_3 NI_3 NS_350 0 -4.4655700561169355e-04
GC_3_351 b_3 NI_3 NS_351 0 1.6138143949288701e-03
GC_3_352 b_3 NI_3 NS_352 0 2.2938437783428080e-03
GC_3_353 b_3 NI_3 NS_353 0 1.0323274411054598e-05
GC_3_354 b_3 NI_3 NS_354 0 -3.6656006988749180e-06
GC_3_355 b_3 NI_3 NS_355 0 1.0985201637522789e-06
GC_3_356 b_3 NI_3 NS_356 0 -3.3395124637520399e-06
GC_3_357 b_3 NI_3 NS_357 0 1.6102096917897354e-04
GC_3_358 b_3 NI_3 NS_358 0 -4.5218442414686130e-05
GC_3_359 b_3 NI_3 NS_359 0 -3.1585124585837798e-06
GC_3_360 b_3 NI_3 NS_360 0 -1.6482095724367912e-05
GC_3_361 b_3 NI_3 NS_361 0 -2.0490222698067649e-04
GC_3_362 b_3 NI_3 NS_362 0 -4.3169615799872669e-06
GC_3_363 b_3 NI_3 NS_363 0 4.0857935313704337e-07
GC_3_364 b_3 NI_3 NS_364 0 4.2656657860943983e-06
GC_3_365 b_3 NI_3 NS_365 0 -3.9050387612390845e-04
GC_3_366 b_3 NI_3 NS_366 0 4.0661314238173076e-04
GC_3_367 b_3 NI_3 NS_367 0 1.9145330452590791e-05
GC_3_368 b_3 NI_3 NS_368 0 -1.9537005297112207e-06
GC_3_369 b_3 NI_3 NS_369 0 4.3210307197001049e-06
GC_3_370 b_3 NI_3 NS_370 0 -2.1205015463838483e-05
GC_3_371 b_3 NI_3 NS_371 0 5.8047115354177938e-04
GC_3_372 b_3 NI_3 NS_372 0 2.7934939342932926e-05
GC_3_373 b_3 NI_3 NS_373 0 2.9211804608507179e-06
GC_3_374 b_3 NI_3 NS_374 0 2.0872343116634177e-07
GC_3_375 b_3 NI_3 NS_375 0 5.6565050872628524e-03
GC_3_376 b_3 NI_3 NS_376 0 -4.4119086380877814e-04
GC_3_377 b_3 NI_3 NS_377 0 4.6096104420739040e-07
GC_3_378 b_3 NI_3 NS_378 0 8.8254120824108671e-10
GC_3_379 b_3 NI_3 NS_379 0 -5.8577980348730634e-04
GC_3_380 b_3 NI_3 NS_380 0 1.2278727387525327e-03
GC_3_381 b_3 NI_3 NS_381 0 5.9221018412023503e-04
GC_3_382 b_3 NI_3 NS_382 0 -6.7901829734173417e-05
GC_3_383 b_3 NI_3 NS_383 0 -2.9555030611322099e-03
GC_3_384 b_3 NI_3 NS_384 0 -1.1020709617604483e-04
GC_3_385 b_3 NI_3 NS_385 0 7.6426817047968746e-04
GC_3_386 b_3 NI_3 NS_386 0 6.6649062419178804e-04
GC_3_387 b_3 NI_3 NS_387 0 -2.4629474417613138e-06
GC_3_388 b_3 NI_3 NS_388 0 1.0671816676241007e-05
GC_3_389 b_3 NI_3 NS_389 0 4.8800843891745524e-06
GC_3_390 b_3 NI_3 NS_390 0 -1.7866073673697156e-05
GC_3_391 b_3 NI_3 NS_391 0 2.1554385295855587e-04
GC_3_392 b_3 NI_3 NS_392 0 1.5960848110434356e-04
GC_3_393 b_3 NI_3 NS_393 0 -1.4650885555473925e-05
GC_3_394 b_3 NI_3 NS_394 0 1.1245295470411828e-05
GC_3_395 b_3 NI_3 NS_395 0 -2.3255592881209512e-04
GC_3_396 b_3 NI_3 NS_396 0 -9.8410687662910327e-05
GC_3_397 b_3 NI_3 NS_397 0 2.5120256159146356e-06
GC_3_398 b_3 NI_3 NS_398 0 -5.6360441608942203e-07
GC_3_399 b_3 NI_3 NS_399 0 -1.5371761147628575e-04
GC_3_400 b_3 NI_3 NS_400 0 3.2102334139093460e-04
GC_3_401 b_3 NI_3 NS_401 0 -4.5645802659496884e-07
GC_3_402 b_3 NI_3 NS_402 0 1.2225113317029522e-05
GC_3_403 b_3 NI_3 NS_403 0 -1.5482971368152968e-06
GC_3_404 b_3 NI_3 NS_404 0 1.9004480054758484e-05
GC_3_405 b_3 NI_3 NS_405 0 4.2222587711979452e-04
GC_3_406 b_3 NI_3 NS_406 0 -1.5487113775876273e-04
GC_3_407 b_3 NI_3 NS_407 0 -7.6611110517437370e-06
GC_3_408 b_3 NI_3 NS_408 0 -1.6383416882241434e-05
GD_3_1 b_3 NI_3 NA_1 0 1.3894850786047967e-02
GD_3_2 b_3 NI_3 NA_2 0 -9.6256405664372595e-03
GD_3_3 b_3 NI_3 NA_3 0 9.9246764772710230e-02
GD_3_4 b_3 NI_3 NA_4 0 -3.4400077369887663e-02
GD_3_5 b_3 NI_3 NA_5 0 6.4410711556076566e-03
GD_3_6 b_3 NI_3 NA_6 0 -8.8109994477151860e-03
GD_3_7 b_3 NI_3 NA_7 0 7.7119977934510722e-03
GD_3_8 b_3 NI_3 NA_8 0 -9.8543399336702663e-03
GD_3_9 b_3 NI_3 NA_9 0 6.5939179130067164e-04
GD_3_10 b_3 NI_3 NA_10 0 -8.9344800400741400e-03
GD_3_11 b_3 NI_3 NA_11 0 -4.2636923307316213e-03
GD_3_12 b_3 NI_3 NA_12 0 -4.7388103356727366e-03
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 3.0722075314258811e-02
GC_4_2 b_4 NI_4 NS_2 0 -3.3971231356417857e-03
GC_4_3 b_4 NI_4 NS_3 0 -2.2139591079784076e-06
GC_4_4 b_4 NI_4 NS_4 0 9.6182855343929478e-09
GC_4_5 b_4 NI_4 NS_5 0 -1.5126270898170117e-02
GC_4_6 b_4 NI_4 NS_6 0 1.1482603565857782e-02
GC_4_7 b_4 NI_4 NS_7 0 2.1544009783246173e-04
GC_4_8 b_4 NI_4 NS_8 0 1.2701205829975819e-03
GC_4_9 b_4 NI_4 NS_9 0 4.1823050889618872e-03
GC_4_10 b_4 NI_4 NS_10 0 -9.1192588514681077e-03
GC_4_11 b_4 NI_4 NS_11 0 -8.5233546600576165e-03
GC_4_12 b_4 NI_4 NS_12 0 -2.2575178158350862e-03
GC_4_13 b_4 NI_4 NS_13 0 9.9919983573866380e-07
GC_4_14 b_4 NI_4 NS_14 0 -8.2328494910719091e-06
GC_4_15 b_4 NI_4 NS_15 0 5.0968714436143836e-06
GC_4_16 b_4 NI_4 NS_16 0 -1.8071168649416196e-05
GC_4_17 b_4 NI_4 NS_17 0 2.1316992321544564e-04
GC_4_18 b_4 NI_4 NS_18 0 1.6257790722779477e-04
GC_4_19 b_4 NI_4 NS_19 0 1.3372192913994090e-05
GC_4_20 b_4 NI_4 NS_20 0 -1.5186621201287107e-05
GC_4_21 b_4 NI_4 NS_21 0 2.2701577283860342e-04
GC_4_22 b_4 NI_4 NS_22 0 9.9626794059669592e-05
GC_4_23 b_4 NI_4 NS_23 0 6.3112230088680769e-06
GC_4_24 b_4 NI_4 NS_24 0 1.1906427234529697e-06
GC_4_25 b_4 NI_4 NS_25 0 -1.3911523222983073e-04
GC_4_26 b_4 NI_4 NS_26 0 -3.4321116909448169e-04
GC_4_27 b_4 NI_4 NS_27 0 -7.7109189771243045e-06
GC_4_28 b_4 NI_4 NS_28 0 1.5730404857834399e-06
GC_4_29 b_4 NI_4 NS_29 0 2.3059562705161628e-06
GC_4_30 b_4 NI_4 NS_30 0 -1.5363955755154881e-05
GC_4_31 b_4 NI_4 NS_31 0 2.7812192018730850e-04
GC_4_32 b_4 NI_4 NS_32 0 -2.0109752586805075e-04
GC_4_33 b_4 NI_4 NS_33 0 -8.1291674464243236e-06
GC_4_34 b_4 NI_4 NS_34 0 -1.7189984830515123e-05
GC_4_35 b_4 NI_4 NS_35 0 -1.5332094972989216e-02
GC_4_36 b_4 NI_4 NS_36 0 -1.2314666001420498e-03
GC_4_37 b_4 NI_4 NS_37 0 -1.6810071032280359e-05
GC_4_38 b_4 NI_4 NS_38 0 -4.9173158125438772e-09
GC_4_39 b_4 NI_4 NS_39 0 7.3474885538126287e-03
GC_4_40 b_4 NI_4 NS_40 0 -1.3076117482014666e-02
GC_4_41 b_4 NI_4 NS_41 0 -9.2764425207295901e-04
GC_4_42 b_4 NI_4 NS_42 0 1.5729460149960814e-03
GC_4_43 b_4 NI_4 NS_43 0 2.0262370733075863e-03
GC_4_44 b_4 NI_4 NS_44 0 3.0609943770552608e-03
GC_4_45 b_4 NI_4 NS_45 0 2.6098408042121660e-03
GC_4_46 b_4 NI_4 NS_46 0 2.2776605650013924e-03
GC_4_47 b_4 NI_4 NS_47 0 1.2288450781081831e-05
GC_4_48 b_4 NI_4 NS_48 0 3.2857665885427930e-06
GC_4_49 b_4 NI_4 NS_49 0 8.0201642338417577e-06
GC_4_50 b_4 NI_4 NS_50 0 -8.8850851891836619e-05
GC_4_51 b_4 NI_4 NS_51 0 9.8347727389363232e-06
GC_4_52 b_4 NI_4 NS_52 0 4.4338832798377769e-04
GC_4_53 b_4 NI_4 NS_53 0 -2.6828472173913132e-05
GC_4_54 b_4 NI_4 NS_54 0 -3.1731855702128792e-06
GC_4_55 b_4 NI_4 NS_55 0 2.3079223782653330e-04
GC_4_56 b_4 NI_4 NS_56 0 1.5691602282530721e-04
GC_4_57 b_4 NI_4 NS_57 0 5.7164335899168617e-07
GC_4_58 b_4 NI_4 NS_58 0 1.4167287445199114e-06
GC_4_59 b_4 NI_4 NS_59 0 -8.7603645830909444e-05
GC_4_60 b_4 NI_4 NS_60 0 -1.5897446547853469e-04
GC_4_61 b_4 NI_4 NS_61 0 -4.0092215732092280e-06
GC_4_62 b_4 NI_4 NS_62 0 -5.3004053224828297e-06
GC_4_63 b_4 NI_4 NS_63 0 -1.1048628316109898e-06
GC_4_64 b_4 NI_4 NS_64 0 1.3873148943323914e-05
GC_4_65 b_4 NI_4 NS_65 0 2.6118491986014896e-04
GC_4_66 b_4 NI_4 NS_66 0 -1.2534189331504797e-04
GC_4_67 b_4 NI_4 NS_67 0 -3.1410331220844892e-05
GC_4_68 b_4 NI_4 NS_68 0 4.5292397812703771e-05
GC_4_69 b_4 NI_4 NS_69 0 2.4153570683015310e-02
GC_4_70 b_4 NI_4 NS_70 0 3.4113442222253418e-02
GC_4_71 b_4 NI_4 NS_71 0 1.5538821398222458e-04
GC_4_72 b_4 NI_4 NS_72 0 2.7164888932076182e-07
GC_4_73 b_4 NI_4 NS_73 0 -5.7083046136506346e-02
GC_4_74 b_4 NI_4 NS_74 0 -2.0359478078410567e-02
GC_4_75 b_4 NI_4 NS_75 0 -8.3340887224729403e-04
GC_4_76 b_4 NI_4 NS_76 0 4.5815201503527523e-03
GC_4_77 b_4 NI_4 NS_77 0 9.5948962966375863e-03
GC_4_78 b_4 NI_4 NS_78 0 1.8374942867699647e-02
GC_4_79 b_4 NI_4 NS_79 0 1.0676603059133219e-02
GC_4_80 b_4 NI_4 NS_80 0 1.5782089851961341e-03
GC_4_81 b_4 NI_4 NS_81 0 -3.5966773994184732e-07
GC_4_82 b_4 NI_4 NS_82 0 -8.1905976306940690e-06
GC_4_83 b_4 NI_4 NS_83 0 3.5730130882450906e-06
GC_4_84 b_4 NI_4 NS_84 0 -1.8337433341917401e-05
GC_4_85 b_4 NI_4 NS_85 0 2.3904684469989749e-04
GC_4_86 b_4 NI_4 NS_86 0 1.6136187931353949e-04
GC_4_87 b_4 NI_4 NS_87 0 7.5552581336031560e-06
GC_4_88 b_4 NI_4 NS_88 0 -1.0381676439990689e-05
GC_4_89 b_4 NI_4 NS_89 0 1.7938391775592700e-04
GC_4_90 b_4 NI_4 NS_90 0 4.0757851960815511e-05
GC_4_91 b_4 NI_4 NS_91 0 9.8936354394581660e-06
GC_4_92 b_4 NI_4 NS_92 0 -1.1970237673332249e-06
GC_4_93 b_4 NI_4 NS_93 0 1.3664941078384802e-04
GC_4_94 b_4 NI_4 NS_94 0 -2.5915662712819353e-04
GC_4_95 b_4 NI_4 NS_95 0 -3.6704448095459626e-06
GC_4_96 b_4 NI_4 NS_96 0 -1.1067836862657189e-05
GC_4_97 b_4 NI_4 NS_97 0 -6.4559252368353430e-07
GC_4_98 b_4 NI_4 NS_98 0 -1.3010790557374381e-05
GC_4_99 b_4 NI_4 NS_99 0 3.9174723386299371e-04
GC_4_100 b_4 NI_4 NS_100 0 -3.3277525731109437e-05
GC_4_101 b_4 NI_4 NS_101 0 -8.9518126536054359e-06
GC_4_102 b_4 NI_4 NS_102 0 -1.6433884589119209e-05
GC_4_103 b_4 NI_4 NS_103 0 9.3446004842317448e-03
GC_4_104 b_4 NI_4 NS_104 0 2.9665631886965995e-02
GC_4_105 b_4 NI_4 NS_105 0 5.7490952198826847e-05
GC_4_106 b_4 NI_4 NS_106 0 -6.6547552553303955e-08
GC_4_107 b_4 NI_4 NS_107 0 5.0186709636858930e-02
GC_4_108 b_4 NI_4 NS_108 0 3.9347797321146169e-02
GC_4_109 b_4 NI_4 NS_109 0 -3.6821452735486828e-03
GC_4_110 b_4 NI_4 NS_110 0 1.3145965825615221e-03
GC_4_111 b_4 NI_4 NS_111 0 -1.3505258112321127e-02
GC_4_112 b_4 NI_4 NS_112 0 1.5006209127992359e-02
GC_4_113 b_4 NI_4 NS_113 0 3.2684233515942710e-03
GC_4_114 b_4 NI_4 NS_114 0 7.8704509438946250e-03
GC_4_115 b_4 NI_4 NS_115 0 1.0012240604945117e-05
GC_4_116 b_4 NI_4 NS_116 0 5.8994647933695288e-07
GC_4_117 b_4 NI_4 NS_117 0 7.9765583160825848e-06
GC_4_118 b_4 NI_4 NS_118 0 -9.0403643125097876e-05
GC_4_119 b_4 NI_4 NS_119 0 1.6566064245599580e-05
GC_4_120 b_4 NI_4 NS_120 0 4.4118146628215402e-04
GC_4_121 b_4 NI_4 NS_121 0 -2.1167015567885498e-05
GC_4_122 b_4 NI_4 NS_122 0 5.4692059816498306e-06
GC_4_123 b_4 NI_4 NS_123 0 1.6721684513831543e-04
GC_4_124 b_4 NI_4 NS_124 0 7.8173631154193727e-05
GC_4_125 b_4 NI_4 NS_125 0 9.1810370648538592e-07
GC_4_126 b_4 NI_4 NS_126 0 2.8804847605870218e-06
GC_4_127 b_4 NI_4 NS_127 0 4.4439816797169911e-05
GC_4_128 b_4 NI_4 NS_128 0 -6.9838537494206130e-05
GC_4_129 b_4 NI_4 NS_129 0 1.9641536386796837e-06
GC_4_130 b_4 NI_4 NS_130 0 -2.3220455865847856e-06
GC_4_131 b_4 NI_4 NS_131 0 6.3170858774116690e-07
GC_4_132 b_4 NI_4 NS_132 0 6.7684363464841858e-06
GC_4_133 b_4 NI_4 NS_133 0 2.2992173133953327e-04
GC_4_134 b_4 NI_4 NS_134 0 -8.9978192247207928e-06
GC_4_135 b_4 NI_4 NS_135 0 -2.9623190339152481e-05
GC_4_136 b_4 NI_4 NS_136 0 4.3417829086474463e-05
GC_4_137 b_4 NI_4 NS_137 0 2.6808497473440867e-02
GC_4_138 b_4 NI_4 NS_138 0 -2.1456648481799211e-03
GC_4_139 b_4 NI_4 NS_139 0 -6.3608693190554912e-07
GC_4_140 b_4 NI_4 NS_140 0 6.9687230279565288e-09
GC_4_141 b_4 NI_4 NS_141 0 -6.7116968242341216e-03
GC_4_142 b_4 NI_4 NS_142 0 1.0915637441821051e-02
GC_4_143 b_4 NI_4 NS_143 0 1.6915671138101299e-03
GC_4_144 b_4 NI_4 NS_144 0 -8.8619624655507205e-04
GC_4_145 b_4 NI_4 NS_145 0 -5.7603044632328097e-03
GC_4_146 b_4 NI_4 NS_146 0 -6.9751314679929316e-03
GC_4_147 b_4 NI_4 NS_147 0 -5.5148046725129428e-03
GC_4_148 b_4 NI_4 NS_148 0 2.8907334094179821e-03
GC_4_149 b_4 NI_4 NS_149 0 2.8006732670861147e-06
GC_4_150 b_4 NI_4 NS_150 0 2.0496894214756603e-06
GC_4_151 b_4 NI_4 NS_151 0 5.4520604666497423e-06
GC_4_152 b_4 NI_4 NS_152 0 -1.9600872673666493e-05
GC_4_153 b_4 NI_4 NS_153 0 2.2080904573660827e-04
GC_4_154 b_4 NI_4 NS_154 0 1.6300103678714388e-04
GC_4_155 b_4 NI_4 NS_155 0 3.5514153140145637e-06
GC_4_156 b_4 NI_4 NS_156 0 -1.2902531217373433e-06
GC_4_157 b_4 NI_4 NS_157 0 3.8000857785363270e-05
GC_4_158 b_4 NI_4 NS_158 0 1.2464320268830883e-05
GC_4_159 b_4 NI_4 NS_159 0 5.3911804473666713e-06
GC_4_160 b_4 NI_4 NS_160 0 -1.4941783248950510e-06
GC_4_161 b_4 NI_4 NS_161 0 1.6202642563709619e-04
GC_4_162 b_4 NI_4 NS_162 0 -1.4467765933192368e-04
GC_4_163 b_4 NI_4 NS_163 0 -1.2277198879988602e-06
GC_4_164 b_4 NI_4 NS_164 0 -1.3506144795545922e-05
GC_4_165 b_4 NI_4 NS_165 0 8.3621397045922272e-07
GC_4_166 b_4 NI_4 NS_166 0 -4.4549031192458965e-06
GC_4_167 b_4 NI_4 NS_167 0 3.5383690603749297e-04
GC_4_168 b_4 NI_4 NS_168 0 -1.4762921911747257e-04
GC_4_169 b_4 NI_4 NS_169 0 -6.3673926484705783e-06
GC_4_170 b_4 NI_4 NS_170 0 -1.5336816576623976e-05
GC_4_171 b_4 NI_4 NS_171 0 -2.0337159877228160e-03
GC_4_172 b_4 NI_4 NS_172 0 -2.1357296269959567e-03
GC_4_173 b_4 NI_4 NS_173 0 -5.6524226802080097e-06
GC_4_174 b_4 NI_4 NS_174 0 -6.5335630409099225e-09
GC_4_175 b_4 NI_4 NS_175 0 1.9288705912478955e-03
GC_4_176 b_4 NI_4 NS_176 0 -8.0450980161637375e-03
GC_4_177 b_4 NI_4 NS_177 0 -6.0985647077895155e-06
GC_4_178 b_4 NI_4 NS_178 0 -2.5130574391787528e-04
GC_4_179 b_4 NI_4 NS_179 0 -2.1480707438443270e-03
GC_4_180 b_4 NI_4 NS_180 0 2.4950810917601903e-03
GC_4_181 b_4 NI_4 NS_181 0 2.8951289687664996e-03
GC_4_182 b_4 NI_4 NS_182 0 2.3490674048024232e-03
GC_4_183 b_4 NI_4 NS_183 0 9.3826852592950023e-07
GC_4_184 b_4 NI_4 NS_184 0 -9.5971190058673725e-07
GC_4_185 b_4 NI_4 NS_185 0 6.2429055711135058e-06
GC_4_186 b_4 NI_4 NS_186 0 -9.1563845703912340e-05
GC_4_187 b_4 NI_4 NS_187 0 3.7472477375467752e-05
GC_4_188 b_4 NI_4 NS_188 0 4.5629215258785008e-04
GC_4_189 b_4 NI_4 NS_189 0 -4.5912167548148616e-06
GC_4_190 b_4 NI_4 NS_190 0 -3.5072177189504715e-06
GC_4_191 b_4 NI_4 NS_191 0 4.0980305640960475e-05
GC_4_192 b_4 NI_4 NS_192 0 3.6946404847684248e-05
GC_4_193 b_4 NI_4 NS_193 0 3.8394640150732262e-07
GC_4_194 b_4 NI_4 NS_194 0 8.4893468795211096e-07
GC_4_195 b_4 NI_4 NS_195 0 1.1790753469106534e-04
GC_4_196 b_4 NI_4 NS_196 0 -1.3574155106168458e-04
GC_4_197 b_4 NI_4 NS_197 0 2.1281863282821384e-06
GC_4_198 b_4 NI_4 NS_198 0 -6.5417413855339555e-07
GC_4_199 b_4 NI_4 NS_199 0 -2.0264628258535310e-09
GC_4_200 b_4 NI_4 NS_200 0 3.9772447665736274e-06
GC_4_201 b_4 NI_4 NS_201 0 3.1314220767489549e-04
GC_4_202 b_4 NI_4 NS_202 0 -1.5974369642820835e-04
GC_4_203 b_4 NI_4 NS_203 0 -3.1294895718493689e-05
GC_4_204 b_4 NI_4 NS_204 0 5.2890711046416594e-05
GC_4_205 b_4 NI_4 NS_205 0 1.6300901698479069e-02
GC_4_206 b_4 NI_4 NS_206 0 -1.1352095043679351e-03
GC_4_207 b_4 NI_4 NS_207 0 -3.5750744015186862e-07
GC_4_208 b_4 NI_4 NS_208 0 3.7690177036544024e-09
GC_4_209 b_4 NI_4 NS_209 0 -2.7066876250150264e-03
GC_4_210 b_4 NI_4 NS_210 0 5.8402545191149208e-03
GC_4_211 b_4 NI_4 NS_211 0 5.1197852693886739e-04
GC_4_212 b_4 NI_4 NS_212 0 -8.9615443566083957e-04
GC_4_213 b_4 NI_4 NS_213 0 -5.1273459350995474e-03
GC_4_214 b_4 NI_4 NS_214 0 -2.0836614677236282e-03
GC_4_215 b_4 NI_4 NS_215 0 -1.6635040437122507e-03
GC_4_216 b_4 NI_4 NS_216 0 2.1256904024087161e-03
GC_4_217 b_4 NI_4 NS_217 0 -6.3217970092459471e-08
GC_4_218 b_4 NI_4 NS_218 0 -2.7912612243588702e-07
GC_4_219 b_4 NI_4 NS_219 0 5.4974348847932768e-06
GC_4_220 b_4 NI_4 NS_220 0 -1.8741474226699548e-05
GC_4_221 b_4 NI_4 NS_221 0 2.2025717424868207e-04
GC_4_222 b_4 NI_4 NS_222 0 1.5559196222018659e-04
GC_4_223 b_4 NI_4 NS_223 0 -3.2405083782121384e-06
GC_4_224 b_4 NI_4 NS_224 0 4.3866653677401926e-06
GC_4_225 b_4 NI_4 NS_225 0 -6.3858212993140768e-05
GC_4_226 b_4 NI_4 NS_226 0 -3.3516334861556001e-05
GC_4_227 b_4 NI_4 NS_227 0 4.1296704746278868e-06
GC_4_228 b_4 NI_4 NS_228 0 -1.8922745394879481e-06
GC_4_229 b_4 NI_4 NS_229 0 1.3105259088879315e-04
GC_4_230 b_4 NI_4 NS_230 0 5.3620918867566533e-05
GC_4_231 b_4 NI_4 NS_231 0 1.9051504390154989e-06
GC_4_232 b_4 NI_4 NS_232 0 -9.5269217969803975e-06
GC_4_233 b_4 NI_4 NS_233 0 -3.6347726391009882e-06
GC_4_234 b_4 NI_4 NS_234 0 6.5922656811783232e-06
GC_4_235 b_4 NI_4 NS_235 0 4.0826134301463990e-04
GC_4_236 b_4 NI_4 NS_236 0 -1.4713924758261176e-04
GC_4_237 b_4 NI_4 NS_237 0 -6.8246003823444254e-06
GC_4_238 b_4 NI_4 NS_238 0 -1.5527401917561609e-05
GC_4_239 b_4 NI_4 NS_239 0 -4.9127780124649844e-03
GC_4_240 b_4 NI_4 NS_240 0 -7.5207588437598417e-04
GC_4_241 b_4 NI_4 NS_241 0 -4.5512763403432280e-06
GC_4_242 b_4 NI_4 NS_242 0 -2.4409720358369519e-09
GC_4_243 b_4 NI_4 NS_243 0 2.3205563059181355e-03
GC_4_244 b_4 NI_4 NS_244 0 -6.8635248834428087e-03
GC_4_245 b_4 NI_4 NS_245 0 -3.5597553905903040e-04
GC_4_246 b_4 NI_4 NS_246 0 -2.1653021691759897e-04
GC_4_247 b_4 NI_4 NS_247 0 -1.6737844657150008e-03
GC_4_248 b_4 NI_4 NS_248 0 3.5898851008677847e-03
GC_4_249 b_4 NI_4 NS_249 0 3.7506862133868659e-03
GC_4_250 b_4 NI_4 NS_250 0 1.1601539027974908e-03
GC_4_251 b_4 NI_4 NS_251 0 7.4442179929927244e-08
GC_4_252 b_4 NI_4 NS_252 0 -8.8681900622742508e-08
GC_4_253 b_4 NI_4 NS_253 0 7.4438665524512193e-06
GC_4_254 b_4 NI_4 NS_254 0 -9.0632568593423737e-05
GC_4_255 b_4 NI_4 NS_255 0 2.8998835932722720e-05
GC_4_256 b_4 NI_4 NS_256 0 4.4602407587315238e-04
GC_4_257 b_4 NI_4 NS_257 0 5.6027059987555488e-06
GC_4_258 b_4 NI_4 NS_258 0 6.3752437621534524e-06
GC_4_259 b_4 NI_4 NS_259 0 -6.1282032126884527e-05
GC_4_260 b_4 NI_4 NS_260 0 -6.4161656854356197e-05
GC_4_261 b_4 NI_4 NS_261 0 -1.4468290414238615e-07
GC_4_262 b_4 NI_4 NS_262 0 -1.0445763274802080e-07
GC_4_263 b_4 NI_4 NS_263 0 1.1598003208037533e-04
GC_4_264 b_4 NI_4 NS_264 0 1.2163958285722479e-05
GC_4_265 b_4 NI_4 NS_265 0 4.8641710296447062e-06
GC_4_266 b_4 NI_4 NS_266 0 2.4934865247656159e-06
GC_4_267 b_4 NI_4 NS_267 0 4.2042019119564085e-07
GC_4_268 b_4 NI_4 NS_268 0 -5.8406543585383924e-06
GC_4_269 b_4 NI_4 NS_269 0 3.2454858434682188e-04
GC_4_270 b_4 NI_4 NS_270 0 -1.7111048163854557e-04
GC_4_271 b_4 NI_4 NS_271 0 -3.1502439793373693e-05
GC_4_272 b_4 NI_4 NS_272 0 5.2850961567763236e-05
GC_4_273 b_4 NI_4 NS_273 0 1.2731600965525726e-02
GC_4_274 b_4 NI_4 NS_274 0 -8.4088907648825284e-04
GC_4_275 b_4 NI_4 NS_275 0 8.3150589298122233e-07
GC_4_276 b_4 NI_4 NS_276 0 1.3529900424570534e-09
GC_4_277 b_4 NI_4 NS_277 0 -2.5330497958644119e-04
GC_4_278 b_4 NI_4 NS_278 0 3.2320864122986127e-03
GC_4_279 b_4 NI_4 NS_279 0 5.3010342644777377e-04
GC_4_280 b_4 NI_4 NS_280 0 -8.1327874031860792e-04
GC_4_281 b_4 NI_4 NS_281 0 -6.6985396016705908e-03
GC_4_282 b_4 NI_4 NS_282 0 2.1814962809837369e-04
GC_4_283 b_4 NI_4 NS_283 0 1.3645734794134336e-03
GC_4_284 b_4 NI_4 NS_284 0 2.5519260213338305e-03
GC_4_285 b_4 NI_4 NS_285 0 -7.8161741520911531e-07
GC_4_286 b_4 NI_4 NS_286 0 8.8972168612939045e-06
GC_4_287 b_4 NI_4 NS_287 0 4.9389978753472544e-06
GC_4_288 b_4 NI_4 NS_288 0 -1.8813917016470911e-05
GC_4_289 b_4 NI_4 NS_289 0 2.2493266496317825e-04
GC_4_290 b_4 NI_4 NS_290 0 1.6206128524120307e-04
GC_4_291 b_4 NI_4 NS_291 0 -6.6593406332838952e-06
GC_4_292 b_4 NI_4 NS_292 0 1.5108013507311004e-05
GC_4_293 b_4 NI_4 NS_293 0 -2.1050272587573379e-04
GC_4_294 b_4 NI_4 NS_294 0 -8.7765546508914536e-05
GC_4_295 b_4 NI_4 NS_295 0 1.0354574180534669e-05
GC_4_296 b_4 NI_4 NS_296 0 -8.1155600816056830e-07
GC_4_297 b_4 NI_4 NS_297 0 3.1102225728082074e-05
GC_4_298 b_4 NI_4 NS_298 0 2.2468720029111130e-04
GC_4_299 b_4 NI_4 NS_299 0 5.2817782934064775e-06
GC_4_300 b_4 NI_4 NS_300 0 2.5308917563681829e-07
GC_4_301 b_4 NI_4 NS_301 0 -1.1577824595747076e-06
GC_4_302 b_4 NI_4 NS_302 0 1.2849329769655656e-05
GC_4_303 b_4 NI_4 NS_303 0 3.6363087111687106e-04
GC_4_304 b_4 NI_4 NS_304 0 -9.4572866249596104e-05
GC_4_305 b_4 NI_4 NS_305 0 -7.6350519149002866e-06
GC_4_306 b_4 NI_4 NS_306 0 -1.5070718321688663e-05
GC_4_307 b_4 NI_4 NS_307 0 1.2332901948537717e-03
GC_4_308 b_4 NI_4 NS_308 0 -4.6498878836827729e-04
GC_4_309 b_4 NI_4 NS_309 0 -9.8632422644383170e-07
GC_4_310 b_4 NI_4 NS_310 0 -1.1652952841677422e-09
GC_4_311 b_4 NI_4 NS_311 0 2.0799342473908460e-03
GC_4_312 b_4 NI_4 NS_312 0 -2.1873216795998108e-03
GC_4_313 b_4 NI_4 NS_313 0 1.8471843078082838e-04
GC_4_314 b_4 NI_4 NS_314 0 -5.2135530022929090e-04
GC_4_315 b_4 NI_4 NS_315 0 -3.6465030621109966e-03
GC_4_316 b_4 NI_4 NS_316 0 2.3603705526559059e-03
GC_4_317 b_4 NI_4 NS_317 0 2.5594550993733745e-03
GC_4_318 b_4 NI_4 NS_318 0 1.3026060306810044e-03
GC_4_319 b_4 NI_4 NS_319 0 -9.6684348727147746e-06
GC_4_320 b_4 NI_4 NS_320 0 -1.9351402080353429e-06
GC_4_321 b_4 NI_4 NS_321 0 6.1010352659656218e-06
GC_4_322 b_4 NI_4 NS_322 0 -9.2664054121075154e-05
GC_4_323 b_4 NI_4 NS_323 0 3.0550624566591442e-05
GC_4_324 b_4 NI_4 NS_324 0 4.6219133466714868e-04
GC_4_325 b_4 NI_4 NS_325 0 2.4328099985845061e-05
GC_4_326 b_4 NI_4 NS_326 0 -3.1911981446737983e-06
GC_4_327 b_4 NI_4 NS_327 0 -2.1045952477054332e-04
GC_4_328 b_4 NI_4 NS_328 0 -1.0665595937500303e-04
GC_4_329 b_4 NI_4 NS_329 0 1.1242571263879393e-06
GC_4_330 b_4 NI_4 NS_330 0 6.6237957867612045e-06
GC_4_331 b_4 NI_4 NS_331 0 8.9366512850646442e-05
GC_4_332 b_4 NI_4 NS_332 0 1.4423243467850621e-04
GC_4_333 b_4 NI_4 NS_333 0 5.0242071767232703e-06
GC_4_334 b_4 NI_4 NS_334 0 2.3546879792860631e-06
GC_4_335 b_4 NI_4 NS_335 0 2.3010161282788980e-06
GC_4_336 b_4 NI_4 NS_336 0 -8.3740560135141393e-06
GC_4_337 b_4 NI_4 NS_337 0 2.6520154112004988e-04
GC_4_338 b_4 NI_4 NS_338 0 -1.5544770550869784e-04
GC_4_339 b_4 NI_4 NS_339 0 -2.8175362138204187e-05
GC_4_340 b_4 NI_4 NS_340 0 4.5776748979313733e-05
GC_4_341 b_4 NI_4 NS_341 0 3.9364504897553597e-03
GC_4_342 b_4 NI_4 NS_342 0 -2.9699639280753590e-04
GC_4_343 b_4 NI_4 NS_343 0 2.1277225867071449e-08
GC_4_344 b_4 NI_4 NS_344 0 1.0072970849020779e-09
GC_4_345 b_4 NI_4 NS_345 0 -6.0188217953505564e-04
GC_4_346 b_4 NI_4 NS_346 0 6.3457773918126740e-04
GC_4_347 b_4 NI_4 NS_347 0 5.9730468935422323e-04
GC_4_348 b_4 NI_4 NS_348 0 -1.8891344487168513e-05
GC_4_349 b_4 NI_4 NS_349 0 -2.6175278715475396e-03
GC_4_350 b_4 NI_4 NS_350 0 1.4294134387329320e-04
GC_4_351 b_4 NI_4 NS_351 0 1.0967118979345761e-03
GC_4_352 b_4 NI_4 NS_352 0 3.2349808974249932e-04
GC_4_353 b_4 NI_4 NS_353 0 -1.1429479384830232e-06
GC_4_354 b_4 NI_4 NS_354 0 1.0601000856992310e-05
GC_4_355 b_4 NI_4 NS_355 0 4.6084310233578903e-06
GC_4_356 b_4 NI_4 NS_356 0 -1.7489066471839153e-05
GC_4_357 b_4 NI_4 NS_357 0 2.1443604779410738e-04
GC_4_358 b_4 NI_4 NS_358 0 1.5572073072420790e-04
GC_4_359 b_4 NI_4 NS_359 0 -1.2547826690749066e-05
GC_4_360 b_4 NI_4 NS_360 0 1.6348273104798786e-05
GC_4_361 b_4 NI_4 NS_361 0 -2.4668938100828593e-04
GC_4_362 b_4 NI_4 NS_362 0 -1.0716621007874144e-04
GC_4_363 b_4 NI_4 NS_363 0 2.8564357313177077e-06
GC_4_364 b_4 NI_4 NS_364 0 -1.6180569437449356e-07
GC_4_365 b_4 NI_4 NS_365 0 -1.5020941678503349e-04
GC_4_366 b_4 NI_4 NS_366 0 3.2792648321525446e-04
GC_4_367 b_4 NI_4 NS_367 0 3.9939776526727949e-06
GC_4_368 b_4 NI_4 NS_368 0 1.2466440144670406e-05
GC_4_369 b_4 NI_4 NS_369 0 -4.2364884298846940e-06
GC_4_370 b_4 NI_4 NS_370 0 1.8937067716223001e-05
GC_4_371 b_4 NI_4 NS_371 0 4.2604239131957989e-04
GC_4_372 b_4 NI_4 NS_372 0 -1.5478303033432590e-04
GC_4_373 b_4 NI_4 NS_373 0 -9.7361841053690331e-06
GC_4_374 b_4 NI_4 NS_374 0 -1.6103565246464250e-05
GC_4_375 b_4 NI_4 NS_375 0 -7.1107908576954911e-04
GC_4_376 b_4 NI_4 NS_376 0 -1.0886719942082317e-04
GC_4_377 b_4 NI_4 NS_377 0 -8.1091852163688544e-07
GC_4_378 b_4 NI_4 NS_378 0 -5.8885706415570743e-10
GC_4_379 b_4 NI_4 NS_379 0 1.5100179670380518e-03
GC_4_380 b_4 NI_4 NS_380 0 -1.5895082833280768e-03
GC_4_381 b_4 NI_4 NS_381 0 3.5732118147432088e-04
GC_4_382 b_4 NI_4 NS_382 0 -4.0707420617954322e-04
GC_4_383 b_4 NI_4 NS_383 0 -2.3298827804190195e-03
GC_4_384 b_4 NI_4 NS_384 0 1.6988274719662761e-03
GC_4_385 b_4 NI_4 NS_385 0 1.7485513539714889e-03
GC_4_386 b_4 NI_4 NS_386 0 3.8653366267782374e-04
GC_4_387 b_4 NI_4 NS_387 0 -1.2185526935187940e-05
GC_4_388 b_4 NI_4 NS_388 0 -3.3252704024345802e-06
GC_4_389 b_4 NI_4 NS_389 0 7.3132802124413556e-06
GC_4_390 b_4 NI_4 NS_390 0 -8.9166320989853045e-05
GC_4_391 b_4 NI_4 NS_391 0 1.5646764153868870e-05
GC_4_392 b_4 NI_4 NS_392 0 4.4586684777388121e-04
GC_4_393 b_4 NI_4 NS_393 0 2.7022163034303749e-05
GC_4_394 b_4 NI_4 NS_394 0 4.4550583367789963e-06
GC_4_395 b_4 NI_4 NS_395 0 -2.4050569214358660e-04
GC_4_396 b_4 NI_4 NS_396 0 -1.7353534069734799e-04
GC_4_397 b_4 NI_4 NS_397 0 -1.3726795388434419e-07
GC_4_398 b_4 NI_4 NS_398 0 2.5285104845514264e-06
GC_4_399 b_4 NI_4 NS_399 0 3.6206584370512745e-06
GC_4_400 b_4 NI_4 NS_400 0 2.5996817897094913e-04
GC_4_401 b_4 NI_4 NS_401 0 3.1493547510026027e-06
GC_4_402 b_4 NI_4 NS_402 0 1.6102215091438779e-06
GC_4_403 b_4 NI_4 NS_403 0 1.7946355724706274e-06
GC_4_404 b_4 NI_4 NS_404 0 -1.3999347419251448e-05
GC_4_405 b_4 NI_4 NS_405 0 3.1093346184722355e-04
GC_4_406 b_4 NI_4 NS_406 0 -2.0352141778749483e-04
GC_4_407 b_4 NI_4 NS_407 0 -3.1096403855123119e-05
GC_4_408 b_4 NI_4 NS_408 0 4.6536348612960300e-05
GD_4_1 b_4 NI_4 NA_1 0 -1.0656352760186732e-02
GD_4_2 b_4 NI_4 NA_2 0 7.0252737429824137e-03
GD_4_3 b_4 NI_4 NA_3 0 -3.4400075371363095e-02
GD_4_4 b_4 NI_4 NA_4 0 -2.5812945306205354e-01
GD_4_5 b_4 NI_4 NA_5 0 -9.9818559582661327e-03
GD_4_6 b_4 NI_4 NA_6 0 2.3321051237280331e-03
GD_4_7 b_4 NI_4 NA_7 0 -7.9128318515889334e-03
GD_4_8 b_4 NI_4 NA_8 0 1.3409619415898296e-03
GD_4_9 b_4 NI_4 NA_9 0 -9.4804141917115854e-03
GD_4_10 b_4 NI_4 NA_10 0 -3.4066751219005735e-03
GD_4_11 b_4 NI_4 NA_11 0 -3.4892373072068815e-03
GD_4_12 b_4 NI_4 NA_12 0 -1.1462971442531176e-03
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 -1.1373952619694714e-02
GC_5_2 b_5 NI_5 NS_2 0 1.4503987860879806e-03
GC_5_3 b_5 NI_5 NS_3 0 -2.8391791813589468e-06
GC_5_4 b_5 NI_5 NS_4 0 -2.7604360920578030e-09
GC_5_5 b_5 NI_5 NS_5 0 2.7030250396707367e-03
GC_5_6 b_5 NI_5 NS_6 0 -1.9543050946232263e-03
GC_5_7 b_5 NI_5 NS_7 0 -5.1294703302199511e-04
GC_5_8 b_5 NI_5 NS_8 0 1.0720016403890106e-03
GC_5_9 b_5 NI_5 NS_9 0 2.1084998194546589e-03
GC_5_10 b_5 NI_5 NS_10 0 -1.3339213174668877e-03
GC_5_11 b_5 NI_5 NS_11 0 -1.7860732625268812e-04
GC_5_12 b_5 NI_5 NS_12 0 -1.8464754032266614e-04
GC_5_13 b_5 NI_5 NS_13 0 -1.0345536492732153e-07
GC_5_14 b_5 NI_5 NS_14 0 -3.5620347771351430e-06
GC_5_15 b_5 NI_5 NS_15 0 1.5640164329728117e-06
GC_5_16 b_5 NI_5 NS_16 0 -4.0672527979803430e-06
GC_5_17 b_5 NI_5 NS_17 0 1.6047617862265380e-04
GC_5_18 b_5 NI_5 NS_18 0 -3.8695788762466835e-05
GC_5_19 b_5 NI_5 NS_19 0 -2.2024897561656422e-07
GC_5_20 b_5 NI_5 NS_20 0 4.8750054952681131e-06
GC_5_21 b_5 NI_5 NS_21 0 6.5188407652049188e-05
GC_5_22 b_5 NI_5 NS_22 0 -1.3628769100637634e-05
GC_5_23 b_5 NI_5 NS_23 0 -8.3678806601487759e-08
GC_5_24 b_5 NI_5 NS_24 0 8.8498255285311604e-07
GC_5_25 b_5 NI_5 NS_25 0 -2.4621096584338700e-04
GC_5_26 b_5 NI_5 NS_26 0 -5.8824823850674148e-05
GC_5_27 b_5 NI_5 NS_27 0 3.4336697802084451e-05
GC_5_28 b_5 NI_5 NS_28 0 -2.2968762756585050e-05
GC_5_29 b_5 NI_5 NS_29 0 -3.9120140790120396e-06
GC_5_30 b_5 NI_5 NS_30 0 3.8121766244058309e-06
GC_5_31 b_5 NI_5 NS_31 0 5.5044279082521852e-04
GC_5_32 b_5 NI_5 NS_32 0 4.7189603436459911e-05
GC_5_33 b_5 NI_5 NS_33 0 1.7903954363179023e-06
GC_5_34 b_5 NI_5 NS_34 0 -5.0008919519655333e-07
GC_5_35 b_5 NI_5 NS_35 0 1.4777411354322388e-02
GC_5_36 b_5 NI_5 NS_36 0 -1.2746318048243099e-03
GC_5_37 b_5 NI_5 NS_37 0 4.1498024572012541e-07
GC_5_38 b_5 NI_5 NS_38 0 3.7348098693534627e-09
GC_5_39 b_5 NI_5 NS_39 0 -4.5503750621285191e-03
GC_5_40 b_5 NI_5 NS_40 0 5.9428470451035140e-03
GC_5_41 b_5 NI_5 NS_41 0 4.1983357405772744e-05
GC_5_42 b_5 NI_5 NS_42 0 9.2106432408606536e-04
GC_5_43 b_5 NI_5 NS_43 0 4.9506859739150697e-06
GC_5_44 b_5 NI_5 NS_44 0 -4.6539423543612594e-03
GC_5_45 b_5 NI_5 NS_45 0 -4.0485847962685910e-03
GC_5_46 b_5 NI_5 NS_46 0 4.6166245362405119e-04
GC_5_47 b_5 NI_5 NS_47 0 1.7712047634356537e-06
GC_5_48 b_5 NI_5 NS_48 0 2.7004233313911611e-06
GC_5_49 b_5 NI_5 NS_49 0 5.4235971487935482e-06
GC_5_50 b_5 NI_5 NS_50 0 -1.9024513177904450e-05
GC_5_51 b_5 NI_5 NS_51 0 2.1142228134967780e-04
GC_5_52 b_5 NI_5 NS_52 0 1.6341038427156000e-04
GC_5_53 b_5 NI_5 NS_53 0 4.5972252272316287e-06
GC_5_54 b_5 NI_5 NS_54 0 -1.3993518992380129e-06
GC_5_55 b_5 NI_5 NS_55 0 7.2473883566981918e-05
GC_5_56 b_5 NI_5 NS_56 0 2.0858671218377780e-05
GC_5_57 b_5 NI_5 NS_57 0 1.0538877427752441e-06
GC_5_58 b_5 NI_5 NS_58 0 -8.5106804651037030e-07
GC_5_59 b_5 NI_5 NS_59 0 -2.2653222963131968e-04
GC_5_60 b_5 NI_5 NS_60 0 -6.0344530525570222e-05
GC_5_61 b_5 NI_5 NS_61 0 -5.3089419813505825e-06
GC_5_62 b_5 NI_5 NS_62 0 1.7532060213009581e-05
GC_5_63 b_5 NI_5 NS_63 0 4.0652307074509453e-06
GC_5_64 b_5 NI_5 NS_64 0 -6.8897672412253774e-06
GC_5_65 b_5 NI_5 NS_65 0 3.8581776411589181e-04
GC_5_66 b_5 NI_5 NS_66 0 -1.6008857467453993e-04
GC_5_67 b_5 NI_5 NS_67 0 -6.4882529691555036e-06
GC_5_68 b_5 NI_5 NS_68 0 -1.6113659446939912e-05
GC_5_69 b_5 NI_5 NS_69 0 -1.7988308673438966e-02
GC_5_70 b_5 NI_5 NS_70 0 2.1699347544023519e-03
GC_5_71 b_5 NI_5 NS_71 0 -6.6258507206228381e-06
GC_5_72 b_5 NI_5 NS_72 0 -4.2996776411726075e-09
GC_5_73 b_5 NI_5 NS_73 0 5.4814729014706310e-03
GC_5_74 b_5 NI_5 NS_74 0 -4.4066955241552595e-03
GC_5_75 b_5 NI_5 NS_75 0 7.6074209655494754e-04
GC_5_76 b_5 NI_5 NS_76 0 4.5990183029293865e-04
GC_5_77 b_5 NI_5 NS_77 0 2.5334398299169217e-04
GC_5_78 b_5 NI_5 NS_78 0 -3.9557311193641676e-04
GC_5_79 b_5 NI_5 NS_79 0 1.2502222479137627e-03
GC_5_80 b_5 NI_5 NS_80 0 6.0862055835711286e-04
GC_5_81 b_5 NI_5 NS_81 0 4.0974456409234411e-07
GC_5_82 b_5 NI_5 NS_82 0 -2.8059484954441285e-06
GC_5_83 b_5 NI_5 NS_83 0 1.6384731788397448e-06
GC_5_84 b_5 NI_5 NS_84 0 -3.9550077718094795e-06
GC_5_85 b_5 NI_5 NS_85 0 1.6311331976470318e-04
GC_5_86 b_5 NI_5 NS_86 0 -4.4407222115376598e-05
GC_5_87 b_5 NI_5 NS_87 0 5.5300344106366811e-07
GC_5_88 b_5 NI_5 NS_88 0 3.3485652216131887e-06
GC_5_89 b_5 NI_5 NS_89 0 3.0871232771302006e-05
GC_5_90 b_5 NI_5 NS_90 0 -1.0358840517402062e-05
GC_5_91 b_5 NI_5 NS_91 0 2.3495749736117798e-06
GC_5_92 b_5 NI_5 NS_92 0 3.7407058717524671e-06
GC_5_93 b_5 NI_5 NS_93 0 4.3100676805607143e-04
GC_5_94 b_5 NI_5 NS_94 0 -9.3737009177919371e-05
GC_5_95 b_5 NI_5 NS_95 0 -3.2130286112603091e-05
GC_5_96 b_5 NI_5 NS_96 0 7.9641339521191827e-06
GC_5_97 b_5 NI_5 NS_97 0 -2.0462564882336603e-06
GC_5_98 b_5 NI_5 NS_98 0 2.5258388370541891e-06
GC_5_99 b_5 NI_5 NS_99 0 5.5498321909279913e-04
GC_5_100 b_5 NI_5 NS_100 0 6.9387170117743505e-05
GC_5_101 b_5 NI_5 NS_101 0 1.0955906515088025e-06
GC_5_102 b_5 NI_5 NS_102 0 -1.9584963333322497e-07
GC_5_103 b_5 NI_5 NS_103 0 2.6808497437250233e-02
GC_5_104 b_5 NI_5 NS_104 0 -2.1456648171618072e-03
GC_5_105 b_5 NI_5 NS_105 0 -6.3608727842348021e-07
GC_5_106 b_5 NI_5 NS_106 0 6.9687320369572759e-09
GC_5_107 b_5 NI_5 NS_107 0 -6.7116967109261197e-03
GC_5_108 b_5 NI_5 NS_108 0 1.0915637379326526e-02
GC_5_109 b_5 NI_5 NS_109 0 1.6915670809531716e-03
GC_5_110 b_5 NI_5 NS_110 0 -8.8619627630288249e-04
GC_5_111 b_5 NI_5 NS_111 0 -5.7603045209865819e-03
GC_5_112 b_5 NI_5 NS_112 0 -6.9751312649594856e-03
GC_5_113 b_5 NI_5 NS_113 0 -5.5148045590032394e-03
GC_5_114 b_5 NI_5 NS_114 0 2.8907334144874391e-03
GC_5_115 b_5 NI_5 NS_115 0 2.8006733216958598e-06
GC_5_116 b_5 NI_5 NS_116 0 2.0496892586117020e-06
GC_5_117 b_5 NI_5 NS_117 0 5.4520603960198085e-06
GC_5_118 b_5 NI_5 NS_118 0 -1.9600872674085693e-05
GC_5_119 b_5 NI_5 NS_119 0 2.2080904619310130e-04
GC_5_120 b_5 NI_5 NS_120 0 1.6300103669516323e-04
GC_5_121 b_5 NI_5 NS_121 0 3.5514152941854750e-06
GC_5_122 b_5 NI_5 NS_122 0 -1.2902531142983300e-06
GC_5_123 b_5 NI_5 NS_123 0 3.8000857968413866e-05
GC_5_124 b_5 NI_5 NS_124 0 1.2464320063848873e-05
GC_5_125 b_5 NI_5 NS_125 0 5.3911805846887886e-06
GC_5_126 b_5 NI_5 NS_126 0 -1.4941785052773674e-06
GC_5_127 b_5 NI_5 NS_127 0 1.6202643153821820e-04
GC_5_128 b_5 NI_5 NS_128 0 -1.4467765954629305e-04
GC_5_129 b_5 NI_5 NS_129 0 -1.2277201464194151e-06
GC_5_130 b_5 NI_5 NS_130 0 -1.3506145219188456e-05
GC_5_131 b_5 NI_5 NS_131 0 8.3621380110255263e-07
GC_5_132 b_5 NI_5 NS_132 0 -4.4549030688257352e-06
GC_5_133 b_5 NI_5 NS_133 0 3.5383690968988262e-04
GC_5_134 b_5 NI_5 NS_134 0 -1.4762921956976889e-04
GC_5_135 b_5 NI_5 NS_135 0 -6.3673927274417359e-06
GC_5_136 b_5 NI_5 NS_136 0 -1.5336816355691997e-05
GC_5_137 b_5 NI_5 NS_137 0 -2.2384059328012385e-01
GC_5_138 b_5 NI_5 NS_138 0 5.6277263399484238e-02
GC_5_139 b_5 NI_5 NS_139 0 4.0204584830929842e-05
GC_5_140 b_5 NI_5 NS_140 0 -5.8184993061757280e-08
GC_5_141 b_5 NI_5 NS_141 0 8.5015052539382213e-02
GC_5_142 b_5 NI_5 NS_142 0 4.4855378050876107e-03
GC_5_143 b_5 NI_5 NS_143 0 3.0089237294974001e-03
GC_5_144 b_5 NI_5 NS_144 0 1.3392399576763209e-03
GC_5_145 b_5 NI_5 NS_145 0 -2.3436100439199132e-03
GC_5_146 b_5 NI_5 NS_146 0 3.6745356432494932e-03
GC_5_147 b_5 NI_5 NS_147 0 -5.4829205665705800e-03
GC_5_148 b_5 NI_5 NS_148 0 6.3910231487295998e-03
GC_5_149 b_5 NI_5 NS_149 0 7.8192220425951645e-07
GC_5_150 b_5 NI_5 NS_150 0 2.3061017404127788e-06
GC_5_151 b_5 NI_5 NS_151 0 2.8116857336863939e-06
GC_5_152 b_5 NI_5 NS_152 0 -4.2808307599375046e-06
GC_5_153 b_5 NI_5 NS_153 0 1.5005058667003020e-04
GC_5_154 b_5 NI_5 NS_154 0 -4.2248917052305634e-05
GC_5_155 b_5 NI_5 NS_155 0 -9.7333666799337312e-08
GC_5_156 b_5 NI_5 NS_156 0 -3.9689634615520968e-07
GC_5_157 b_5 NI_5 NS_157 0 1.7112258288386232e-05
GC_5_158 b_5 NI_5 NS_158 0 6.9802227295704753e-06
GC_5_159 b_5 NI_5 NS_159 0 2.8379236976055318e-06
GC_5_160 b_5 NI_5 NS_160 0 1.3406329953724726e-06
GC_5_161 b_5 NI_5 NS_161 0 8.9102787161316800e-04
GC_5_162 b_5 NI_5 NS_162 0 -1.4073766285681161e-04
GC_5_163 b_5 NI_5 NS_163 0 -8.4753224536744293e-05
GC_5_164 b_5 NI_5 NS_164 0 3.1307231977608797e-05
GC_5_165 b_5 NI_5 NS_165 0 -2.7558506331272744e-06
GC_5_166 b_5 NI_5 NS_166 0 1.4931960608358469e-06
GC_5_167 b_5 NI_5 NS_167 0 5.8917173521732223e-04
GC_5_168 b_5 NI_5 NS_168 0 -1.5435494019324560e-05
GC_5_169 b_5 NI_5 NS_169 0 1.5103402500662558e-06
GC_5_170 b_5 NI_5 NS_170 0 1.0664430709024560e-06
GC_5_171 b_5 NI_5 NS_171 0 3.7890982846856158e-02
GC_5_172 b_5 NI_5 NS_172 0 3.2803455045768488e-02
GC_5_173 b_5 NI_5 NS_173 0 1.6630724839388164e-04
GC_5_174 b_5 NI_5 NS_174 0 2.5381250441336865e-07
GC_5_175 b_5 NI_5 NS_175 0 -5.7809488157756196e-02
GC_5_176 b_5 NI_5 NS_176 0 -1.5960464929923812e-02
GC_5_177 b_5 NI_5 NS_177 0 4.5741914908167618e-04
GC_5_178 b_5 NI_5 NS_178 0 2.6796339350366682e-03
GC_5_179 b_5 NI_5 NS_179 0 2.2482608369490953e-03
GC_5_180 b_5 NI_5 NS_180 0 1.8396447667934877e-02
GC_5_181 b_5 NI_5 NS_181 0 1.0464378986743668e-02
GC_5_182 b_5 NI_5 NS_182 0 3.8575376010025336e-03
GC_5_183 b_5 NI_5 NS_183 0 -5.2976107630249679e-07
GC_5_184 b_5 NI_5 NS_184 0 -6.7783871423220639e-07
GC_5_185 b_5 NI_5 NS_185 0 3.7271214696358449e-06
GC_5_186 b_5 NI_5 NS_186 0 -2.0018565207425974e-05
GC_5_187 b_5 NI_5 NS_187 0 2.3831405386803440e-04
GC_5_188 b_5 NI_5 NS_188 0 1.5923921145376797e-04
GC_5_189 b_5 NI_5 NS_189 0 4.6997270937389599e-08
GC_5_190 b_5 NI_5 NS_190 0 1.6571687364669641e-06
GC_5_191 b_5 NI_5 NS_191 0 3.0930437217421695e-05
GC_5_192 b_5 NI_5 NS_192 0 -1.7009662788574149e-05
GC_5_193 b_5 NI_5 NS_193 0 -1.3790251855134380e-06
GC_5_194 b_5 NI_5 NS_194 0 -1.9145348732909942e-06
GC_5_195 b_5 NI_5 NS_195 0 6.4905409392518310e-04
GC_5_196 b_5 NI_5 NS_196 0 -2.7202673886637192e-04
GC_5_197 b_5 NI_5 NS_197 0 -1.9557006815273407e-06
GC_5_198 b_5 NI_5 NS_198 0 -4.5839125377968796e-05
GC_5_199 b_5 NI_5 NS_199 0 -3.6227104727325928e-06
GC_5_200 b_5 NI_5 NS_200 0 -7.9447624327175570e-06
GC_5_201 b_5 NI_5 NS_201 0 5.9098869013214878e-04
GC_5_202 b_5 NI_5 NS_202 0 -6.5483927468155698e-05
GC_5_203 b_5 NI_5 NS_203 0 -1.1190985011362545e-05
GC_5_204 b_5 NI_5 NS_204 0 -1.6212926580233100e-05
GC_5_205 b_5 NI_5 NS_205 0 -2.4578684303094355e-02
GC_5_206 b_5 NI_5 NS_206 0 2.3109325422858585e-03
GC_5_207 b_5 NI_5 NS_207 0 -1.1969289320169429e-05
GC_5_208 b_5 NI_5 NS_208 0 -6.5212476367936964e-09
GC_5_209 b_5 NI_5 NS_209 0 9.9904325783141054e-03
GC_5_210 b_5 NI_5 NS_210 0 -7.1631520607390465e-03
GC_5_211 b_5 NI_5 NS_211 0 8.9129181490204808e-04
GC_5_212 b_5 NI_5 NS_212 0 -5.5497974867383185e-04
GC_5_213 b_5 NI_5 NS_213 0 -2.1589312700067242e-03
GC_5_214 b_5 NI_5 NS_214 0 8.3730781085390781e-04
GC_5_215 b_5 NI_5 NS_215 0 1.8697579300424141e-03
GC_5_216 b_5 NI_5 NS_216 0 2.1874797141119202e-03
GC_5_217 b_5 NI_5 NS_217 0 -9.6504215332428431e-08
GC_5_218 b_5 NI_5 NS_218 0 -3.2649106384260148e-07
GC_5_219 b_5 NI_5 NS_219 0 1.7081423737579245e-06
GC_5_220 b_5 NI_5 NS_220 0 -4.4546909613499894e-06
GC_5_221 b_5 NI_5 NS_221 0 1.5966999094929078e-04
GC_5_222 b_5 NI_5 NS_222 0 -4.2446823739653704e-05
GC_5_223 b_5 NI_5 NS_223 0 -7.7544182211576278e-08
GC_5_224 b_5 NI_5 NS_224 0 -1.4563104477215315e-06
GC_5_225 b_5 NI_5 NS_225 0 -2.0936780368262740e-05
GC_5_226 b_5 NI_5 NS_226 0 1.4234189436556967e-06
GC_5_227 b_5 NI_5 NS_227 0 9.3960759087522684e-07
GC_5_228 b_5 NI_5 NS_228 0 1.2655888809931691e-06
GC_5_229 b_5 NI_5 NS_229 0 8.2956417969895133e-04
GC_5_230 b_5 NI_5 NS_230 0 -1.9269097226843602e-05
GC_5_231 b_5 NI_5 NS_231 0 -8.0481899687617447e-05
GC_5_232 b_5 NI_5 NS_232 0 2.7088140932301320e-05
GC_5_233 b_5 NI_5 NS_233 0 1.0654380776271832e-06
GC_5_234 b_5 NI_5 NS_234 0 -3.4209768754471542e-06
GC_5_235 b_5 NI_5 NS_235 0 6.7614907788987784e-04
GC_5_236 b_5 NI_5 NS_236 0 1.7111326589894725e-05
GC_5_237 b_5 NI_5 NS_237 0 3.6397607898549644e-07
GC_5_238 b_5 NI_5 NS_238 0 1.4601820025814580e-06
GC_5_239 b_5 NI_5 NS_239 0 3.8454741459380659e-02
GC_5_240 b_5 NI_5 NS_240 0 -3.7520079819583448e-03
GC_5_241 b_5 NI_5 NS_241 0 -5.5177184432755324e-07
GC_5_242 b_5 NI_5 NS_242 0 7.7763443073349200e-09
GC_5_243 b_5 NI_5 NS_243 0 -1.2629000868299215e-02
GC_5_244 b_5 NI_5 NS_244 0 1.3572289280951515e-02
GC_5_245 b_5 NI_5 NS_245 0 2.0569629636937800e-03
GC_5_246 b_5 NI_5 NS_246 0 -1.6516363777757603e-03
GC_5_247 b_5 NI_5 NS_247 0 -6.5723456049894746e-03
GC_5_248 b_5 NI_5 NS_248 0 -6.8978475179837379e-03
GC_5_249 b_5 NI_5 NS_249 0 -5.7915729333336179e-03
GC_5_250 b_5 NI_5 NS_250 0 1.3642169118043941e-03
GC_5_251 b_5 NI_5 NS_251 0 1.0765546382808655e-06
GC_5_252 b_5 NI_5 NS_252 0 5.5287467480634102e-07
GC_5_253 b_5 NI_5 NS_253 0 5.2734393812488259e-06
GC_5_254 b_5 NI_5 NS_254 0 -1.9056269327845706e-05
GC_5_255 b_5 NI_5 NS_255 0 2.2164006507818370e-04
GC_5_256 b_5 NI_5 NS_256 0 1.5206293026416630e-04
GC_5_257 b_5 NI_5 NS_257 0 -9.7582809898567478e-07
GC_5_258 b_5 NI_5 NS_258 0 -1.0091767250470007e-07
GC_5_259 b_5 NI_5 NS_259 0 -2.8383041938911456e-05
GC_5_260 b_5 NI_5 NS_260 0 -4.3744723028936984e-06
GC_5_261 b_5 NI_5 NS_261 0 2.4953799498321454e-06
GC_5_262 b_5 NI_5 NS_262 0 -3.1052403866579314e-07
GC_5_263 b_5 NI_5 NS_263 0 4.5430660614313592e-04
GC_5_264 b_5 NI_5 NS_264 0 -1.5640574983967633e-04
GC_5_265 b_5 NI_5 NS_265 0 -4.9385753981605250e-06
GC_5_266 b_5 NI_5 NS_266 0 -3.9842778640184558e-05
GC_5_267 b_5 NI_5 NS_267 0 -5.4037811396775799e-06
GC_5_268 b_5 NI_5 NS_268 0 1.8079694989551823e-06
GC_5_269 b_5 NI_5 NS_269 0 4.7145020162774824e-04
GC_5_270 b_5 NI_5 NS_270 0 -2.1130533638697536e-04
GC_5_271 b_5 NI_5 NS_271 0 -8.1755647788538270e-06
GC_5_272 b_5 NI_5 NS_272 0 -1.5839886173805105e-05
GC_5_273 b_5 NI_5 NS_273 0 -1.1524578436301086e-02
GC_5_274 b_5 NI_5 NS_274 0 1.5028382553084318e-03
GC_5_275 b_5 NI_5 NS_275 0 -3.3155460366826683e-06
GC_5_276 b_5 NI_5 NS_276 0 -2.1612924803635223e-09
GC_5_277 b_5 NI_5 NS_277 0 3.1885440194595605e-03
GC_5_278 b_5 NI_5 NS_278 0 -2.5019623507636884e-03
GC_5_279 b_5 NI_5 NS_279 0 2.4757069407907982e-04
GC_5_280 b_5 NI_5 NS_280 0 -2.7440477878107691e-04
GC_5_281 b_5 NI_5 NS_281 0 -9.9884794514421590e-04
GC_5_282 b_5 NI_5 NS_282 0 4.3453767329538226e-04
GC_5_283 b_5 NI_5 NS_283 0 1.4320859461342806e-03
GC_5_284 b_5 NI_5 NS_284 0 1.3282558218311903e-04
GC_5_285 b_5 NI_5 NS_285 0 -6.3884599466989454e-07
GC_5_286 b_5 NI_5 NS_286 0 3.0385879194264209e-06
GC_5_287 b_5 NI_5 NS_287 0 1.6337265808079873e-06
GC_5_288 b_5 NI_5 NS_288 0 -3.8354230114479621e-06
GC_5_289 b_5 NI_5 NS_289 0 1.6248306428631271e-04
GC_5_290 b_5 NI_5 NS_290 0 -4.7229210296690663e-05
GC_5_291 b_5 NI_5 NS_291 0 2.1173813099672803e-07
GC_5_292 b_5 NI_5 NS_292 0 -3.8697217804209968e-06
GC_5_293 b_5 NI_5 NS_293 0 -4.6869147246608937e-05
GC_5_294 b_5 NI_5 NS_294 0 3.4179080167437307e-06
GC_5_295 b_5 NI_5 NS_295 0 3.1486075162853268e-06
GC_5_296 b_5 NI_5 NS_296 0 4.7800364769519877e-06
GC_5_297 b_5 NI_5 NS_297 0 1.5357999797457379e-04
GC_5_298 b_5 NI_5 NS_298 0 9.4630137610421722e-05
GC_5_299 b_5 NI_5 NS_299 0 -2.5099752206444198e-05
GC_5_300 b_5 NI_5 NS_300 0 2.4893981736563356e-06
GC_5_301 b_5 NI_5 NS_301 0 2.2973686987618735e-06
GC_5_302 b_5 NI_5 NS_302 0 -5.4819246634115955e-06
GC_5_303 b_5 NI_5 NS_303 0 5.8775318514592051e-04
GC_5_304 b_5 NI_5 NS_304 0 -6.3349345795156892e-06
GC_5_305 b_5 NI_5 NS_305 0 1.6267956875039875e-06
GC_5_306 b_5 NI_5 NS_306 0 6.1434601437724829e-07
GC_5_307 b_5 NI_5 NS_307 0 1.5887108495273097e-02
GC_5_308 b_5 NI_5 NS_308 0 -1.1065483144161619e-03
GC_5_309 b_5 NI_5 NS_309 0 -6.9482752504075076e-07
GC_5_310 b_5 NI_5 NS_310 0 4.0370184123455574e-09
GC_5_311 b_5 NI_5 NS_311 0 -2.6793994950468410e-03
GC_5_312 b_5 NI_5 NS_312 0 5.7506103592184169e-03
GC_5_313 b_5 NI_5 NS_313 0 5.0127014080544700e-04
GC_5_314 b_5 NI_5 NS_314 0 -8.0585932464183807e-04
GC_5_315 b_5 NI_5 NS_315 0 -4.6410356713936975e-03
GC_5_316 b_5 NI_5 NS_316 0 -2.3166589507709000e-03
GC_5_317 b_5 NI_5 NS_317 0 -1.9437663321229710e-03
GC_5_318 b_5 NI_5 NS_318 0 2.0985168273425564e-03
GC_5_319 b_5 NI_5 NS_319 0 -1.3675635560827221e-06
GC_5_320 b_5 NI_5 NS_320 0 -9.4761363607222349e-07
GC_5_321 b_5 NI_5 NS_321 0 5.5591359724620619e-06
GC_5_322 b_5 NI_5 NS_322 0 -1.9042841612049693e-05
GC_5_323 b_5 NI_5 NS_323 0 2.2142554820817211e-04
GC_5_324 b_5 NI_5 NS_324 0 1.5402699205785132e-04
GC_5_325 b_5 NI_5 NS_325 0 -2.8123794987267385e-06
GC_5_326 b_5 NI_5 NS_326 0 1.1745248333082181e-06
GC_5_327 b_5 NI_5 NS_327 0 -5.0332746997837845e-05
GC_5_328 b_5 NI_5 NS_328 0 -1.4751892287749061e-05
GC_5_329 b_5 NI_5 NS_329 0 5.0029522462363425e-06
GC_5_330 b_5 NI_5 NS_330 0 -1.8290710720017121e-06
GC_5_331 b_5 NI_5 NS_331 0 1.1691826840955915e-04
GC_5_332 b_5 NI_5 NS_332 0 8.9643912944516611e-05
GC_5_333 b_5 NI_5 NS_333 0 -3.8140015006581376e-06
GC_5_334 b_5 NI_5 NS_334 0 -1.4295580930038154e-05
GC_5_335 b_5 NI_5 NS_335 0 -3.4180294893414710e-06
GC_5_336 b_5 NI_5 NS_336 0 4.3446193378284745e-06
GC_5_337 b_5 NI_5 NS_337 0 3.8469774604502337e-04
GC_5_338 b_5 NI_5 NS_338 0 -1.6609326384337374e-04
GC_5_339 b_5 NI_5 NS_339 0 -6.4782700022094963e-06
GC_5_340 b_5 NI_5 NS_340 0 -1.5188851888670150e-05
GC_5_341 b_5 NI_5 NS_341 0 -2.8622177022428401e-03
GC_5_342 b_5 NI_5 NS_342 0 5.8851327952333832e-04
GC_5_343 b_5 NI_5 NS_343 0 -1.0298864966763025e-06
GC_5_344 b_5 NI_5 NS_344 0 -1.2006998388796959e-09
GC_5_345 b_5 NI_5 NS_345 0 1.5323556776897485e-03
GC_5_346 b_5 NI_5 NS_346 0 -4.5397319873391418e-04
GC_5_347 b_5 NI_5 NS_347 0 -1.0401356492838801e-03
GC_5_348 b_5 NI_5 NS_348 0 5.4147232368960596e-05
GC_5_349 b_5 NI_5 NS_349 0 3.3884830478356611e-04
GC_5_350 b_5 NI_5 NS_350 0 1.1008726921009724e-03
GC_5_351 b_5 NI_5 NS_351 0 6.7206615338891965e-04
GC_5_352 b_5 NI_5 NS_352 0 -1.1552819054169662e-04
GC_5_353 b_5 NI_5 NS_353 0 -9.2189530336984108e-07
GC_5_354 b_5 NI_5 NS_354 0 3.4633228020464295e-06
GC_5_355 b_5 NI_5 NS_355 0 1.4049616997112588e-06
GC_5_356 b_5 NI_5 NS_356 0 -3.6180738115984488e-06
GC_5_357 b_5 NI_5 NS_357 0 1.5695188827668228e-04
GC_5_358 b_5 NI_5 NS_358 0 -4.4913653698191418e-05
GC_5_359 b_5 NI_5 NS_359 0 3.7329392491571135e-07
GC_5_360 b_5 NI_5 NS_360 0 -4.8331641295905602e-06
GC_5_361 b_5 NI_5 NS_361 0 -6.8575196568477288e-05
GC_5_362 b_5 NI_5 NS_362 0 7.6708108420227848e-06
GC_5_363 b_5 NI_5 NS_363 0 6.6535546912673386e-07
GC_5_364 b_5 NI_5 NS_364 0 1.7916865187024615e-06
GC_5_365 b_5 NI_5 NS_365 0 -6.1779644540159689e-04
GC_5_366 b_5 NI_5 NS_366 0 2.1697438728228113e-04
GC_5_367 b_5 NI_5 NS_367 0 4.0716317259721804e-05
GC_5_368 b_5 NI_5 NS_368 0 -2.3436322750626952e-05
GC_5_369 b_5 NI_5 NS_369 0 4.5511178592163331e-06
GC_5_370 b_5 NI_5 NS_370 0 -6.9727967488132211e-06
GC_5_371 b_5 NI_5 NS_371 0 5.9902873648373320e-04
GC_5_372 b_5 NI_5 NS_372 0 -4.6277938217044891e-05
GC_5_373 b_5 NI_5 NS_373 0 2.9055001949352739e-06
GC_5_374 b_5 NI_5 NS_374 0 6.8394115093016755e-07
GC_5_375 b_5 NI_5 NS_375 0 5.4021798308820246e-03
GC_5_376 b_5 NI_5 NS_376 0 -4.3346914070500680e-04
GC_5_377 b_5 NI_5 NS_377 0 -4.7317694739413073e-07
GC_5_378 b_5 NI_5 NS_378 0 2.1521514942869591e-09
GC_5_379 b_5 NI_5 NS_379 0 -1.9034790315051490e-03
GC_5_380 b_5 NI_5 NS_380 0 1.7235803106456359e-03
GC_5_381 b_5 NI_5 NS_381 0 -7.6963993710624831e-04
GC_5_382 b_5 NI_5 NS_382 0 9.4719002733915675e-04
GC_5_383 b_5 NI_5 NS_383 0 1.9703931574612771e-03
GC_5_384 b_5 NI_5 NS_384 0 -1.0335447002475752e-03
GC_5_385 b_5 NI_5 NS_385 0 -1.4931646151946950e-03
GC_5_386 b_5 NI_5 NS_386 0 -7.1922081734784524e-04
GC_5_387 b_5 NI_5 NS_387 0 -3.1306282871690516e-06
GC_5_388 b_5 NI_5 NS_388 0 -9.4461711789186468e-07
GC_5_389 b_5 NI_5 NS_389 0 5.4250480414665168e-06
GC_5_390 b_5 NI_5 NS_390 0 -1.8420695723537245e-05
GC_5_391 b_5 NI_5 NS_391 0 2.1202949979123685e-04
GC_5_392 b_5 NI_5 NS_392 0 1.5543281426769870e-04
GC_5_393 b_5 NI_5 NS_393 0 -4.1713392620949157e-06
GC_5_394 b_5 NI_5 NS_394 0 1.2719174555189891e-06
GC_5_395 b_5 NI_5 NS_395 0 -7.8345097337881363e-05
GC_5_396 b_5 NI_5 NS_396 0 -2.1931711040258326e-05
GC_5_397 b_5 NI_5 NS_397 0 1.6913553438384495e-06
GC_5_398 b_5 NI_5 NS_398 0 -7.6928513183719990e-07
GC_5_399 b_5 NI_5 NS_399 0 -3.4506704688041530e-04
GC_5_400 b_5 NI_5 NS_400 0 2.2281252126397168e-04
GC_5_401 b_5 NI_5 NS_401 0 -8.3649286992617884e-06
GC_5_402 b_5 NI_5 NS_402 0 2.0621716281937393e-05
GC_5_403 b_5 NI_5 NS_403 0 -3.2667044291044090e-06
GC_5_404 b_5 NI_5 NS_404 0 9.6005338366192016e-06
GC_5_405 b_5 NI_5 NS_405 0 4.1271430860975446e-04
GC_5_406 b_5 NI_5 NS_406 0 -2.3123693608877356e-04
GC_5_407 b_5 NI_5 NS_407 0 -5.5405075231165416e-06
GC_5_408 b_5 NI_5 NS_408 0 -1.5541170802666494e-05
GD_5_1 b_5 NI_5 NA_1 0 6.2221544138608455e-03
GD_5_2 b_5 NI_5 NA_2 0 -6.6284204565197572e-03
GD_5_3 b_5 NI_5 NA_3 0 6.4410711691190422e-03
GD_5_4 b_5 NI_5 NA_4 0 -9.9818562545322346e-03
GD_5_5 b_5 NI_5 NA_5 0 9.9837283571118610e-02
GD_5_6 b_5 NI_5 NA_6 0 -4.0969397149139442e-02
GD_5_7 b_5 NI_5 NA_7 0 1.1444632400471874e-02
GD_5_8 b_5 NI_5 NA_8 0 -1.4684082980540513e-02
GD_5_9 b_5 NI_5 NA_9 0 6.3443274442737457e-03
GD_5_10 b_5 NI_5 NA_10 0 -7.8366526450173654e-03
GD_5_11 b_5 NI_5 NA_11 0 1.2182002000193340e-03
GD_5_12 b_5 NI_5 NA_12 0 -4.6948877768767851e-03
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 1.0923923999200523e-02
GC_6_2 b_6 NI_6 NS_2 0 -9.9093547729459238e-04
GC_6_3 b_6 NI_6 NS_3 0 -5.0420317851012217e-07
GC_6_4 b_6 NI_6 NS_4 0 4.0613342278015129e-09
GC_6_5 b_6 NI_6 NS_5 0 -4.6032554652413946e-03
GC_6_6 b_6 NI_6 NS_6 0 4.7075079992328567e-03
GC_6_7 b_6 NI_6 NS_7 0 1.0470823039937682e-04
GC_6_8 b_6 NI_6 NS_8 0 1.2216823406147096e-03
GC_6_9 b_6 NI_6 NS_9 0 1.2341743622257745e-03
GC_6_10 b_6 NI_6 NS_10 0 -4.5722212799371243e-03
GC_6_11 b_6 NI_6 NS_11 0 -3.8831213288262239e-03
GC_6_12 b_6 NI_6 NS_12 0 -3.5043681490104712e-04
GC_6_13 b_6 NI_6 NS_13 0 -1.9925457460619525e-06
GC_6_14 b_6 NI_6 NS_14 0 -1.8025931504124768e-07
GC_6_15 b_6 NI_6 NS_15 0 5.4110874523071684e-06
GC_6_16 b_6 NI_6 NS_16 0 -1.8433002166919731e-05
GC_6_17 b_6 NI_6 NS_17 0 2.1095218482681340e-04
GC_6_18 b_6 NI_6 NS_18 0 1.5828722451434183e-04
GC_6_19 b_6 NI_6 NS_19 0 6.9360686670825428e-06
GC_6_20 b_6 NI_6 NS_20 0 -2.5853830712530519e-06
GC_6_21 b_6 NI_6 NS_21 0 6.2305608764986128e-05
GC_6_22 b_6 NI_6 NS_22 0 3.3611621124637868e-05
GC_6_23 b_6 NI_6 NS_23 0 1.3262876527726787e-06
GC_6_24 b_6 NI_6 NS_24 0 -7.8071328523980362e-08
GC_6_25 b_6 NI_6 NS_25 0 -1.7782476254548846e-04
GC_6_26 b_6 NI_6 NS_26 0 -2.4741237688533795e-05
GC_6_27 b_6 NI_6 NS_27 0 6.7187784184768681e-07
GC_6_28 b_6 NI_6 NS_28 0 1.2257205124332133e-05
GC_6_29 b_6 NI_6 NS_29 0 1.1931166884851907e-06
GC_6_30 b_6 NI_6 NS_30 0 -1.1017135117500821e-05
GC_6_31 b_6 NI_6 NS_31 0 3.9572249705983116e-04
GC_6_32 b_6 NI_6 NS_32 0 -1.5734619680536575e-04
GC_6_33 b_6 NI_6 NS_33 0 -1.1966920583434141e-05
GC_6_34 b_6 NI_6 NS_34 0 -1.9429578601501549e-05
GC_6_35 b_6 NI_6 NS_35 0 -4.1956147206903931e-03
GC_6_36 b_6 NI_6 NS_36 0 -1.1458352979102232e-03
GC_6_37 b_6 NI_6 NS_37 0 -2.4677847871682554e-06
GC_6_38 b_6 NI_6 NS_38 0 -3.8011446924284786e-09
GC_6_39 b_6 NI_6 NS_39 0 1.1173785434543131e-03
GC_6_40 b_6 NI_6 NS_40 0 -5.7754595921816164e-03
GC_6_41 b_6 NI_6 NS_41 0 -9.8345746687153373e-05
GC_6_42 b_6 NI_6 NS_42 0 7.8634018435441569e-04
GC_6_43 b_6 NI_6 NS_43 0 7.6123446135840109e-04
GC_6_44 b_6 NI_6 NS_44 0 4.6511990170919549e-04
GC_6_45 b_6 NI_6 NS_45 0 9.8823756561435992e-04
GC_6_46 b_6 NI_6 NS_46 0 6.1309233273465448e-04
GC_6_47 b_6 NI_6 NS_47 0 5.7881491882086522e-07
GC_6_48 b_6 NI_6 NS_48 0 -5.6832259446768229e-07
GC_6_49 b_6 NI_6 NS_49 0 6.7453557261610823e-06
GC_6_50 b_6 NI_6 NS_50 0 -8.8697761183805218e-05
GC_6_51 b_6 NI_6 NS_51 0 2.6191843823482805e-05
GC_6_52 b_6 NI_6 NS_52 0 4.4564360043875873e-04
GC_6_53 b_6 NI_6 NS_53 0 -1.1135891116589272e-05
GC_6_54 b_6 NI_6 NS_54 0 -9.6642852249766253e-06
GC_6_55 b_6 NI_6 NS_55 0 7.3630295379228805e-05
GC_6_56 b_6 NI_6 NS_56 0 7.8419787395061922e-05
GC_6_57 b_6 NI_6 NS_57 0 -6.7665876868779250e-07
GC_6_58 b_6 NI_6 NS_58 0 8.6731426069638316e-07
GC_6_59 b_6 NI_6 NS_59 0 -7.8883106395334339e-05
GC_6_60 b_6 NI_6 NS_60 0 1.4107884604987459e-05
GC_6_61 b_6 NI_6 NS_61 0 -5.5273121970138673e-06
GC_6_62 b_6 NI_6 NS_62 0 -8.0874434454234858e-06
GC_6_63 b_6 NI_6 NS_63 0 5.2661925289544451e-07
GC_6_64 b_6 NI_6 NS_64 0 7.7064753635570151e-06
GC_6_65 b_6 NI_6 NS_65 0 3.3034061841789891e-04
GC_6_66 b_6 NI_6 NS_66 0 -1.9723433247512039e-04
GC_6_67 b_6 NI_6 NS_67 0 -3.3640832604614048e-05
GC_6_68 b_6 NI_6 NS_68 0 5.3584372385966512e-05
GC_6_69 b_6 NI_6 NS_69 0 2.4281995731971640e-02
GC_6_70 b_6 NI_6 NS_70 0 -1.9476109567026379e-03
GC_6_71 b_6 NI_6 NS_71 0 -1.6180037787239025e-06
GC_6_72 b_6 NI_6 NS_72 0 7.3122494528776733e-09
GC_6_73 b_6 NI_6 NS_73 0 -6.7212766616745519e-03
GC_6_74 b_6 NI_6 NS_74 0 9.7809332401103816e-03
GC_6_75 b_6 NI_6 NS_75 0 1.5286347237941427e-03
GC_6_76 b_6 NI_6 NS_76 0 -8.3858681094445525e-04
GC_6_77 b_6 NI_6 NS_77 0 -4.9878046212613551e-03
GC_6_78 b_6 NI_6 NS_78 0 -5.9445640437262009e-03
GC_6_79 b_6 NI_6 NS_79 0 -4.8684733271041189e-03
GC_6_80 b_6 NI_6 NS_80 0 2.0734956931810285e-03
GC_6_81 b_6 NI_6 NS_81 0 -3.6686164774559454e-07
GC_6_82 b_6 NI_6 NS_82 0 -4.4756344326086615e-07
GC_6_83 b_6 NI_6 NS_83 0 5.3414429963074288e-06
GC_6_84 b_6 NI_6 NS_84 0 -1.8401455752188656e-05
GC_6_85 b_6 NI_6 NS_85 0 2.2054589696656639e-04
GC_6_86 b_6 NI_6 NS_86 0 1.5572914558961958e-04
GC_6_87 b_6 NI_6 NS_87 0 5.3297367012818502e-06
GC_6_88 b_6 NI_6 NS_88 0 -1.3838197013233019e-06
GC_6_89 b_6 NI_6 NS_89 0 2.8854638494654296e-05
GC_6_90 b_6 NI_6 NS_90 0 2.0729404933249622e-05
GC_6_91 b_6 NI_6 NS_91 0 5.0055940648486131e-06
GC_6_92 b_6 NI_6 NS_92 0 -3.6969528210215309e-07
GC_6_93 b_6 NI_6 NS_93 0 2.0210338363365026e-04
GC_6_94 b_6 NI_6 NS_94 0 -1.4138931789322350e-04
GC_6_95 b_6 NI_6 NS_95 0 -1.3115660866775028e-06
GC_6_96 b_6 NI_6 NS_96 0 -1.7211246834623777e-05
GC_6_97 b_6 NI_6 NS_97 0 -1.8374427792876613e-06
GC_6_98 b_6 NI_6 NS_98 0 -7.5555470224109131e-06
GC_6_99 b_6 NI_6 NS_99 0 3.7706639114235896e-04
GC_6_100 b_6 NI_6 NS_100 0 -1.3393097819466677e-04
GC_6_101 b_6 NI_6 NS_101 0 -9.7619359091794153e-06
GC_6_102 b_6 NI_6 NS_102 0 -1.7941821805486109e-05
GC_6_103 b_6 NI_6 NS_103 0 -2.0337120872231805e-03
GC_6_104 b_6 NI_6 NS_104 0 -2.1357301493801248e-03
GC_6_105 b_6 NI_6 NS_105 0 -5.6524192893720688e-06
GC_6_106 b_6 NI_6 NS_106 0 -6.5335535059067759e-09
GC_6_107 b_6 NI_6 NS_107 0 1.9288693860963785e-03
GC_6_108 b_6 NI_6 NS_108 0 -8.0450963967488142e-03
GC_6_109 b_6 NI_6 NS_109 0 -6.0988630557311424e-06
GC_6_110 b_6 NI_6 NS_110 0 -2.5130543323013970e-04
GC_6_111 b_6 NI_6 NS_111 0 -2.1480684973417419e-03
GC_6_112 b_6 NI_6 NS_112 0 2.4950805362850600e-03
GC_6_113 b_6 NI_6 NS_113 0 2.8951266075030184e-03
GC_6_114 b_6 NI_6 NS_114 0 2.3490665266702321e-03
GC_6_115 b_6 NI_6 NS_115 0 9.3826718635613887e-07
GC_6_116 b_6 NI_6 NS_116 0 -9.5971248024891572e-07
GC_6_117 b_6 NI_6 NS_117 0 6.2429052195427757e-06
GC_6_118 b_6 NI_6 NS_118 0 -9.1563846617065425e-05
GC_6_119 b_6 NI_6 NS_119 0 3.7472479092471678e-05
GC_6_120 b_6 NI_6 NS_120 0 4.5629216132262162e-04
GC_6_121 b_6 NI_6 NS_121 0 -4.5912183762172037e-06
GC_6_122 b_6 NI_6 NS_122 0 -3.5072184112487118e-06
GC_6_123 b_6 NI_6 NS_123 0 4.0980320621541588e-05
GC_6_124 b_6 NI_6 NS_124 0 3.6946414180773501e-05
GC_6_125 b_6 NI_6 NS_125 0 3.8394977797820011e-07
GC_6_126 b_6 NI_6 NS_126 0 8.4893024398459740e-07
GC_6_127 b_6 NI_6 NS_127 0 1.1790757977172788e-04
GC_6_128 b_6 NI_6 NS_128 0 -1.3574162367860926e-04
GC_6_129 b_6 NI_6 NS_129 0 2.1281851390541692e-06
GC_6_130 b_6 NI_6 NS_130 0 -6.5417577614200997e-07
GC_6_131 b_6 NI_6 NS_131 0 -2.0272263469956200e-09
GC_6_132 b_6 NI_6 NS_132 0 3.9772400478796834e-06
GC_6_133 b_6 NI_6 NS_133 0 3.1314226985137083e-04
GC_6_134 b_6 NI_6 NS_134 0 -1.5974390064248727e-04
GC_6_135 b_6 NI_6 NS_135 0 -3.1294897893067158e-05
GC_6_136 b_6 NI_6 NS_136 0 5.2890716848196115e-05
GC_6_137 b_6 NI_6 NS_137 0 3.7890983142164394e-02
GC_6_138 b_6 NI_6 NS_138 0 3.2803454991012913e-02
GC_6_139 b_6 NI_6 NS_139 0 1.6630724895000656e-04
GC_6_140 b_6 NI_6 NS_140 0 2.5381250084940330e-07
GC_6_141 b_6 NI_6 NS_141 0 -5.7809488267683957e-02
GC_6_142 b_6 NI_6 NS_142 0 -1.5960464828535952e-02
GC_6_143 b_6 NI_6 NS_143 0 4.5741916343203243e-04
GC_6_144 b_6 NI_6 NS_144 0 2.6796339392119901e-03
GC_6_145 b_6 NI_6 NS_145 0 2.2482608469633642e-03
GC_6_146 b_6 NI_6 NS_146 0 1.8396447566630229e-02
GC_6_147 b_6 NI_6 NS_147 0 1.0464378893282571e-02
GC_6_148 b_6 NI_6 NS_148 0 3.8575375940500941e-03
GC_6_149 b_6 NI_6 NS_149 0 -5.2976110752078576e-07
GC_6_150 b_6 NI_6 NS_150 0 -6.7783871844381365e-07
GC_6_151 b_6 NI_6 NS_151 0 3.7271214732683584e-06
GC_6_152 b_6 NI_6 NS_152 0 -2.0018565237964348e-05
GC_6_153 b_6 NI_6 NS_153 0 2.3831405368443694e-04
GC_6_154 b_6 NI_6 NS_154 0 1.5923921171147334e-04
GC_6_155 b_6 NI_6 NS_155 0 4.6997287336625415e-08
GC_6_156 b_6 NI_6 NS_156 0 1.6571686388408921e-06
GC_6_157 b_6 NI_6 NS_157 0 3.0930437117627437e-05
GC_6_158 b_6 NI_6 NS_158 0 -1.7009662204909498e-05
GC_6_159 b_6 NI_6 NS_159 0 -1.3790251521391542e-06
GC_6_160 b_6 NI_6 NS_160 0 -1.9145348058470617e-06
GC_6_161 b_6 NI_6 NS_161 0 6.4905409281740256e-04
GC_6_162 b_6 NI_6 NS_162 0 -2.7202673972104540e-04
GC_6_163 b_6 NI_6 NS_163 0 -1.9557007163513224e-06
GC_6_164 b_6 NI_6 NS_164 0 -4.5839125360628771e-05
GC_6_165 b_6 NI_6 NS_165 0 -3.6227105078499562e-06
GC_6_166 b_6 NI_6 NS_166 0 -7.9447624182447319e-06
GC_6_167 b_6 NI_6 NS_167 0 5.9098868931040821e-04
GC_6_168 b_6 NI_6 NS_168 0 -6.5483929130906920e-05
GC_6_169 b_6 NI_6 NS_169 0 -1.1190985033039956e-05
GC_6_170 b_6 NI_6 NS_170 0 -1.6212926617639376e-05
GC_6_171 b_6 NI_6 NS_171 0 1.3342016745102922e-02
GC_6_172 b_6 NI_6 NS_172 0 2.9250107218226112e-02
GC_6_173 b_6 NI_6 NS_173 0 6.2362648101517329e-05
GC_6_174 b_6 NI_6 NS_174 0 -6.9779639272115893e-08
GC_6_175 b_6 NI_6 NS_175 0 4.9139309349969379e-02
GC_6_176 b_6 NI_6 NS_176 0 4.1144000328233871e-02
GC_6_177 b_6 NI_6 NS_177 0 -3.5639203442905526e-03
GC_6_178 b_6 NI_6 NS_178 0 6.5882491845943580e-04
GC_6_179 b_6 NI_6 NS_179 0 -1.3894351670626024e-02
GC_6_180 b_6 NI_6 NS_180 0 1.6466706129650555e-02
GC_6_181 b_6 NI_6 NS_181 0 2.3133697667007064e-03
GC_6_182 b_6 NI_6 NS_182 0 6.6127394436194713e-03
GC_6_183 b_6 NI_6 NS_183 0 -9.5322334738644303e-07
GC_6_184 b_6 NI_6 NS_184 0 -2.5087324070172779e-06
GC_6_185 b_6 NI_6 NS_185 0 5.9720568557909761e-06
GC_6_186 b_6 NI_6 NS_186 0 -8.8927496810643010e-05
GC_6_187 b_6 NI_6 NS_187 0 4.4653144294022607e-05
GC_6_188 b_6 NI_6 NS_188 0 4.3638996098726874e-04
GC_6_189 b_6 NI_6 NS_189 0 -3.9629750866832105e-06
GC_6_190 b_6 NI_6 NS_190 0 -2.1080761521499474e-06
GC_6_191 b_6 NI_6 NS_191 0 1.6341752204190348e-05
GC_6_192 b_6 NI_6 NS_192 0 9.2371422399514235e-06
GC_6_193 b_6 NI_6 NS_193 0 -2.2192046681105241e-06
GC_6_194 b_6 NI_6 NS_194 0 1.3463621815330098e-08
GC_6_195 b_6 NI_6 NS_195 0 3.6546790781384186e-04
GC_6_196 b_6 NI_6 NS_196 0 -2.6173302506112857e-04
GC_6_197 b_6 NI_6 NS_197 0 1.0136519343792824e-05
GC_6_198 b_6 NI_6 NS_198 0 -4.4059327847435776e-07
GC_6_199 b_6 NI_6 NS_199 0 -5.4605915553575047e-07
GC_6_200 b_6 NI_6 NS_200 0 -1.1637641062224544e-06
GC_6_201 b_6 NI_6 NS_201 0 4.2656946480985506e-04
GC_6_202 b_6 NI_6 NS_202 0 -1.5087383097995991e-04
GC_6_203 b_6 NI_6 NS_203 0 -3.4667029340881692e-05
GC_6_204 b_6 NI_6 NS_204 0 6.1949345516929791e-05
GC_6_205 b_6 NI_6 NS_205 0 3.9398689366914041e-02
GC_6_206 b_6 NI_6 NS_206 0 -3.8027456410936679e-03
GC_6_207 b_6 NI_6 NS_207 0 -2.2108134114487555e-07
GC_6_208 b_6 NI_6 NS_208 0 7.6575934685440494e-09
GC_6_209 b_6 NI_6 NS_209 0 -1.2692397720930552e-02
GC_6_210 b_6 NI_6 NS_210 0 1.3989841253027253e-02
GC_6_211 b_6 NI_6 NS_211 0 2.0040860630008120e-03
GC_6_212 b_6 NI_6 NS_212 0 -1.7541344749119143e-03
GC_6_213 b_6 NI_6 NS_213 0 -6.8895796563513386e-03
GC_6_214 b_6 NI_6 NS_214 0 -6.9691632879346748e-03
GC_6_215 b_6 NI_6 NS_215 0 -5.8144425891092019e-03
GC_6_216 b_6 NI_6 NS_216 0 1.5417696669837346e-03
GC_6_217 b_6 NI_6 NS_217 0 1.0895417091455786e-06
GC_6_218 b_6 NI_6 NS_218 0 5.5556073563999872e-07
GC_6_219 b_6 NI_6 NS_219 0 4.8279231782139232e-06
GC_6_220 b_6 NI_6 NS_220 0 -1.8629319524865497e-05
GC_6_221 b_6 NI_6 NS_221 0 2.2422802931395248e-04
GC_6_222 b_6 NI_6 NS_222 0 1.4853378576340834e-04
GC_6_223 b_6 NI_6 NS_223 0 -1.8957991538499251e-06
GC_6_224 b_6 NI_6 NS_224 0 9.9824057958898643e-07
GC_6_225 b_6 NI_6 NS_225 0 -2.5684842002493103e-05
GC_6_226 b_6 NI_6 NS_226 0 -9.5445547036636145e-06
GC_6_227 b_6 NI_6 NS_227 0 2.5020812418024360e-06
GC_6_228 b_6 NI_6 NS_228 0 -3.5815133009204460e-07
GC_6_229 b_6 NI_6 NS_229 0 4.2655454678124788e-04
GC_6_230 b_6 NI_6 NS_230 0 -1.7189299558522105e-04
GC_6_231 b_6 NI_6 NS_231 0 -1.9651571489894842e-06
GC_6_232 b_6 NI_6 NS_232 0 -3.6011901352146402e-05
GC_6_233 b_6 NI_6 NS_233 0 -4.9733150174181302e-06
GC_6_234 b_6 NI_6 NS_234 0 3.4938481161674228e-06
GC_6_235 b_6 NI_6 NS_235 0 4.6661137455839609e-04
GC_6_236 b_6 NI_6 NS_236 0 -2.0891821401787004e-04
GC_6_237 b_6 NI_6 NS_237 0 -8.4037805194710131e-06
GC_6_238 b_6 NI_6 NS_238 0 -1.6195804985290001e-05
GC_6_239 b_6 NI_6 NS_239 0 -3.6774142583276882e-03
GC_6_240 b_6 NI_6 NS_240 0 -2.0338603084609956e-03
GC_6_241 b_6 NI_6 NS_241 0 -1.2217708599690424e-05
GC_6_242 b_6 NI_6 NS_242 0 -6.2794739644959556e-09
GC_6_243 b_6 NI_6 NS_243 0 6.9045378966442117e-03
GC_6_244 b_6 NI_6 NS_244 0 -9.3401851895370570e-03
GC_6_245 b_6 NI_6 NS_245 0 -3.6092172102635711e-04
GC_6_246 b_6 NI_6 NS_246 0 -2.9917285492014217e-04
GC_6_247 b_6 NI_6 NS_247 0 -3.6364345147392612e-03
GC_6_248 b_6 NI_6 NS_248 0 4.8358167457894672e-03
GC_6_249 b_6 NI_6 NS_249 0 3.2294594245785065e-03
GC_6_250 b_6 NI_6 NS_250 0 3.8338757600223658e-03
GC_6_251 b_6 NI_6 NS_251 0 1.9283571160520147e-07
GC_6_252 b_6 NI_6 NS_252 0 -4.0058206004823367e-07
GC_6_253 b_6 NI_6 NS_253 0 6.5086391977379008e-06
GC_6_254 b_6 NI_6 NS_254 0 -8.9957219622989465e-05
GC_6_255 b_6 NI_6 NS_255 0 4.3652196873770543e-05
GC_6_256 b_6 NI_6 NS_256 0 4.4486709223855766e-04
GC_6_257 b_6 NI_6 NS_257 0 3.6744129782696514e-06
GC_6_258 b_6 NI_6 NS_258 0 4.8664915917705327e-06
GC_6_259 b_6 NI_6 NS_259 0 -1.9158460226521493e-05
GC_6_260 b_6 NI_6 NS_260 0 -3.5878298239642588e-05
GC_6_261 b_6 NI_6 NS_261 0 -1.0708892837522199e-07
GC_6_262 b_6 NI_6 NS_262 0 -1.0085261869873894e-06
GC_6_263 b_6 NI_6 NS_263 0 2.5235126750942384e-04
GC_6_264 b_6 NI_6 NS_264 0 -2.0036362318822629e-04
GC_6_265 b_6 NI_6 NS_265 0 1.0238278233107007e-05
GC_6_266 b_6 NI_6 NS_266 0 4.6973424225915092e-06
GC_6_267 b_6 NI_6 NS_267 0 -1.4850965915180337e-06
GC_6_268 b_6 NI_6 NS_268 0 -4.2845934282747884e-06
GC_6_269 b_6 NI_6 NS_269 0 3.6102274771749877e-04
GC_6_270 b_6 NI_6 NS_270 0 -2.1690426323265464e-04
GC_6_271 b_6 NI_6 NS_271 0 -3.3168601378930410e-05
GC_6_272 b_6 NI_6 NS_272 0 6.2037108450309635e-05
GC_6_273 b_6 NI_6 NS_273 0 1.9252399373864328e-02
GC_6_274 b_6 NI_6 NS_274 0 -1.4019191745883520e-03
GC_6_275 b_6 NI_6 NS_275 0 2.9704686852451721e-07
GC_6_276 b_6 NI_6 NS_276 0 3.6651218875960764e-09
GC_6_277 b_6 NI_6 NS_277 0 -2.9344176703762471e-03
GC_6_278 b_6 NI_6 NS_278 0 6.9317189153136781e-03
GC_6_279 b_6 NI_6 NS_279 0 4.8453207872418828e-04
GC_6_280 b_6 NI_6 NS_280 0 -9.3438377383054001e-04
GC_6_281 b_6 NI_6 NS_281 0 -5.3627140964110894e-03
GC_6_282 b_6 NI_6 NS_282 0 -2.7018997709248975e-03
GC_6_283 b_6 NI_6 NS_283 0 -2.3571635780482414e-03
GC_6_284 b_6 NI_6 NS_284 0 2.6137202303906301e-03
GC_6_285 b_6 NI_6 NS_285 0 1.7829410513719259e-06
GC_6_286 b_6 NI_6 NS_286 0 1.3392131824125870e-06
GC_6_287 b_6 NI_6 NS_287 0 4.6156931914641437e-06
GC_6_288 b_6 NI_6 NS_288 0 -1.8386300393511748e-05
GC_6_289 b_6 NI_6 NS_289 0 2.2705407240919292e-04
GC_6_290 b_6 NI_6 NS_290 0 1.5334470533336504e-04
GC_6_291 b_6 NI_6 NS_291 0 -5.8952980872644831e-06
GC_6_292 b_6 NI_6 NS_292 0 1.9408004739950469e-06
GC_6_293 b_6 NI_6 NS_293 0 -3.7069794333158799e-05
GC_6_294 b_6 NI_6 NS_294 0 -2.4795825079858923e-05
GC_6_295 b_6 NI_6 NS_295 0 5.8375808336809502e-06
GC_6_296 b_6 NI_6 NS_296 0 -7.1649665643399934e-07
GC_6_297 b_6 NI_6 NS_297 0 5.2722614979527746e-05
GC_6_298 b_6 NI_6 NS_298 0 4.5308802344149217e-05
GC_6_299 b_6 NI_6 NS_299 0 3.5772893687455974e-06
GC_6_300 b_6 NI_6 NS_300 0 -7.1102903068567651e-06
GC_6_301 b_6 NI_6 NS_301 0 -3.9538089680439776e-07
GC_6_302 b_6 NI_6 NS_302 0 8.3386400260782330e-06
GC_6_303 b_6 NI_6 NS_303 0 3.8217129698771480e-04
GC_6_304 b_6 NI_6 NS_304 0 -1.6632278197421303e-04
GC_6_305 b_6 NI_6 NS_305 0 -8.8253403780796183e-06
GC_6_306 b_6 NI_6 NS_306 0 -1.6230668438016593e-05
GC_6_307 b_6 NI_6 NS_307 0 -4.9892365757837993e-03
GC_6_308 b_6 NI_6 NS_308 0 -7.7323317557513105e-04
GC_6_309 b_6 NI_6 NS_309 0 -4.5212466265816156e-06
GC_6_310 b_6 NI_6 NS_310 0 -2.5022878588523312e-09
GC_6_311 b_6 NI_6 NS_311 0 2.3094344038707324e-03
GC_6_312 b_6 NI_6 NS_312 0 -6.8959419595272381e-03
GC_6_313 b_6 NI_6 NS_313 0 -3.1008218288504797e-04
GC_6_314 b_6 NI_6 NS_314 0 -1.7661234001045787e-04
GC_6_315 b_6 NI_6 NS_315 0 -1.6942448827637325e-03
GC_6_316 b_6 NI_6 NS_316 0 3.2544013461254665e-03
GC_6_317 b_6 NI_6 NS_317 0 3.6661984993595167e-03
GC_6_318 b_6 NI_6 NS_318 0 1.3253540880233791e-03
GC_6_319 b_6 NI_6 NS_319 0 -4.6074654666422308e-07
GC_6_320 b_6 NI_6 NS_320 0 2.5372496899128906e-07
GC_6_321 b_6 NI_6 NS_321 0 6.3470709897479651e-06
GC_6_322 b_6 NI_6 NS_322 0 -9.0540277348176567e-05
GC_6_323 b_6 NI_6 NS_323 0 3.7450443205582432e-05
GC_6_324 b_6 NI_6 NS_324 0 4.4414663461173087e-04
GC_6_325 b_6 NI_6 NS_325 0 4.7112137980943351e-06
GC_6_326 b_6 NI_6 NS_326 0 5.1400578448751181e-06
GC_6_327 b_6 NI_6 NS_327 0 -4.8732853681098671e-05
GC_6_328 b_6 NI_6 NS_328 0 -5.7866687039609989e-05
GC_6_329 b_6 NI_6 NS_329 0 2.3619909316876917e-07
GC_6_330 b_6 NI_6 NS_330 0 -2.6185082299218427e-07
GC_6_331 b_6 NI_6 NS_331 0 1.0128345599584846e-04
GC_6_332 b_6 NI_6 NS_332 0 4.6775376132098109e-05
GC_6_333 b_6 NI_6 NS_333 0 7.5007951422451201e-06
GC_6_334 b_6 NI_6 NS_334 0 1.6377466269731373e-06
GC_6_335 b_6 NI_6 NS_335 0 5.4979362869252014e-07
GC_6_336 b_6 NI_6 NS_336 0 -5.8021261635319020e-06
GC_6_337 b_6 NI_6 NS_337 0 3.0645650404775252e-04
GC_6_338 b_6 NI_6 NS_338 0 -1.7220681471671930e-04
GC_6_339 b_6 NI_6 NS_339 0 -3.0380137899884827e-05
GC_6_340 b_6 NI_6 NS_340 0 5.3286493165877057e-05
GC_6_341 b_6 NI_6 NS_341 0 5.7403087667870379e-03
GC_6_342 b_6 NI_6 NS_342 0 -4.9676091359682683e-04
GC_6_343 b_6 NI_6 NS_343 0 -3.0287300178094266e-07
GC_6_344 b_6 NI_6 NS_344 0 2.0712740265976221e-09
GC_6_345 b_6 NI_6 NS_345 0 -2.1362631196286922e-03
GC_6_346 b_6 NI_6 NS_346 0 2.0558650617156318e-03
GC_6_347 b_6 NI_6 NS_347 0 -5.6368285425103658e-04
GC_6_348 b_6 NI_6 NS_348 0 1.2106233553992127e-03
GC_6_349 b_6 NI_6 NS_349 0 2.1059602341509274e-03
GC_6_350 b_6 NI_6 NS_350 0 -2.0079011909312629e-03
GC_6_351 b_6 NI_6 NS_351 0 -1.9806786179854935e-03
GC_6_352 b_6 NI_6 NS_352 0 -5.1433388339218119e-04
GC_6_353 b_6 NI_6 NS_353 0 7.1068751683564507e-07
GC_6_354 b_6 NI_6 NS_354 0 2.3213112165553577e-06
GC_6_355 b_6 NI_6 NS_355 0 3.9708326778999624e-06
GC_6_356 b_6 NI_6 NS_356 0 -1.6980380326585424e-05
GC_6_357 b_6 NI_6 NS_357 0 2.1944531493056402e-04
GC_6_358 b_6 NI_6 NS_358 0 1.4707432558985699e-04
GC_6_359 b_6 NI_6 NS_359 0 -7.2273878126489406e-06
GC_6_360 b_6 NI_6 NS_360 0 2.8266324967690821e-06
GC_6_361 b_6 NI_6 NS_361 0 -6.6659900016780409e-05
GC_6_362 b_6 NI_6 NS_362 0 -3.4821924795119211e-05
GC_6_363 b_6 NI_6 NS_363 0 2.5397971200108589e-06
GC_6_364 b_6 NI_6 NS_364 0 -6.3351568824667841e-08
GC_6_365 b_6 NI_6 NS_365 0 -3.9623929312108291e-04
GC_6_366 b_6 NI_6 NS_366 0 2.1414933478213890e-04
GC_6_367 b_6 NI_6 NS_367 0 3.5141890747250070e-06
GC_6_368 b_6 NI_6 NS_368 0 2.5696908440780404e-05
GC_6_369 b_6 NI_6 NS_369 0 -3.9930522672334352e-07
GC_6_370 b_6 NI_6 NS_370 0 1.3819878885708266e-05
GC_6_371 b_6 NI_6 NS_371 0 4.0151958417967575e-04
GC_6_372 b_6 NI_6 NS_372 0 -2.3371863573041222e-04
GC_6_373 b_6 NI_6 NS_373 0 -1.0493955405766366e-05
GC_6_374 b_6 NI_6 NS_374 0 -1.7880258058269762e-05
GC_6_375 b_6 NI_6 NS_375 0 -6.3951134583731676e-03
GC_6_376 b_6 NI_6 NS_376 0 -2.3781867975623855e-05
GC_6_377 b_6 NI_6 NS_377 0 -2.5485819995405096e-06
GC_6_378 b_6 NI_6 NS_378 0 -7.9728793129731629e-10
GC_6_379 b_6 NI_6 NS_379 0 1.5307391215666905e-03
GC_6_380 b_6 NI_6 NS_380 0 -4.4623371408368572e-03
GC_6_381 b_6 NI_6 NS_381 0 -2.2304637285967637e-04
GC_6_382 b_6 NI_6 NS_382 0 7.2350814968276302e-04
GC_6_383 b_6 NI_6 NS_383 0 1.0093195098844062e-03
GC_6_384 b_6 NI_6 NS_384 0 8.9321507959967076e-04
GC_6_385 b_6 NI_6 NS_385 0 1.5186890007362985e-03
GC_6_386 b_6 NI_6 NS_386 0 -6.0196205222927639e-05
GC_6_387 b_6 NI_6 NS_387 0 -1.0877546320154797e-06
GC_6_388 b_6 NI_6 NS_388 0 9.7781376740810116e-07
GC_6_389 b_6 NI_6 NS_389 0 7.2087175992825203e-06
GC_6_390 b_6 NI_6 NS_390 0 -8.7170162695910367e-05
GC_6_391 b_6 NI_6 NS_391 0 2.4865908071693432e-05
GC_6_392 b_6 NI_6 NS_392 0 4.3046784505187404e-04
GC_6_393 b_6 NI_6 NS_393 0 1.0752707990476520e-05
GC_6_394 b_6 NI_6 NS_394 0 1.0506743464341019e-05
GC_6_395 b_6 NI_6 NS_395 0 -7.4276533980518445e-05
GC_6_396 b_6 NI_6 NS_396 0 -9.1464439591981838e-05
GC_6_397 b_6 NI_6 NS_397 0 -2.0937189260242305e-07
GC_6_398 b_6 NI_6 NS_398 0 -3.2000761655897165e-07
GC_6_399 b_6 NI_6 NS_399 0 -1.3885867054658601e-04
GC_6_400 b_6 NI_6 NS_400 0 2.5435660580648914e-04
GC_6_401 b_6 NI_6 NS_401 0 -6.5013093919765549e-07
GC_6_402 b_6 NI_6 NS_402 0 -2.6367857936215684e-06
GC_6_403 b_6 NI_6 NS_403 0 -1.2321075643677266e-07
GC_6_404 b_6 NI_6 NS_404 0 -7.8646786905136415e-06
GC_6_405 b_6 NI_6 NS_405 0 3.1397806596348063e-04
GC_6_406 b_6 NI_6 NS_406 0 -2.3071870277451925e-04
GC_6_407 b_6 NI_6 NS_407 0 -3.2997646857659135e-05
GC_6_408 b_6 NI_6 NS_408 0 5.3916330671465853e-05
GD_6_1 b_6 NI_6 NA_1 0 -3.9477680891773026e-03
GD_6_2 b_6 NI_6 NA_2 0 2.9032617111062697e-03
GD_6_3 b_6 NI_6 NA_3 0 -8.8109985294029924e-03
GD_6_4 b_6 NI_6 NA_4 0 2.3321013501177109e-03
GD_6_5 b_6 NI_6 NA_5 0 -4.0969397186779548e-02
GD_6_6 b_6 NI_6 NA_6 0 -2.6043365196471924e-01
GD_6_7 b_6 NI_6 NA_7 0 -1.5077494731883155e-02
GD_6_8 b_6 NI_6 NA_8 0 -7.2274199774254911e-04
GD_6_9 b_6 NI_6 NA_9 0 -9.8259844448069268e-03
GD_6_10 b_6 NI_6 NA_10 0 1.6658817338809908e-03
GD_6_11 b_6 NI_6 NA_11 0 -4.4612996932750530e-03
GD_6_12 b_6 NI_6 NA_12 0 2.5564032129953848e-03
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 -3.0412030314926554e-03
GC_7_2 b_7 NI_7 NS_2 0 5.6947556121811967e-04
GC_7_3 b_7 NI_7 NS_3 0 -9.6944955066841313e-07
GC_7_4 b_7 NI_7 NS_4 0 -1.1830923747264665e-09
GC_7_5 b_7 NI_7 NS_5 0 1.4261246137030150e-03
GC_7_6 b_7 NI_7 NS_6 0 -3.4967944907216952e-04
GC_7_7 b_7 NI_7 NS_7 0 -7.0604123017308656e-04
GC_7_8 b_7 NI_7 NS_8 0 2.7752911067682398e-04
GC_7_9 b_7 NI_7 NS_9 0 2.1133680062194969e-05
GC_7_10 b_7 NI_7 NS_10 0 1.3191331263275551e-04
GC_7_11 b_7 NI_7 NS_11 0 4.8294650382351941e-04
GC_7_12 b_7 NI_7 NS_12 0 1.3021462013956616e-04
GC_7_13 b_7 NI_7 NS_13 0 4.6795668769138247e-08
GC_7_14 b_7 NI_7 NS_14 0 1.5979265636148717e-06
GC_7_15 b_7 NI_7 NS_15 0 1.5105288262869912e-06
GC_7_16 b_7 NI_7 NS_16 0 -3.7040428070809357e-06
GC_7_17 b_7 NI_7 NS_17 0 1.5909935313607496e-04
GC_7_18 b_7 NI_7 NS_18 0 -4.2454103083045664e-05
GC_7_19 b_7 NI_7 NS_19 0 -1.2405611472817706e-06
GC_7_20 b_7 NI_7 NS_20 0 -7.6111416396099406e-06
GC_7_21 b_7 NI_7 NS_21 0 -8.6255186047320175e-05
GC_7_22 b_7 NI_7 NS_22 0 -8.2379058613708720e-06
GC_7_23 b_7 NI_7 NS_23 0 3.9895789279640266e-07
GC_7_24 b_7 NI_7 NS_24 0 1.4327494400895587e-06
GC_7_25 b_7 NI_7 NS_25 0 -5.5169339231041714e-04
GC_7_26 b_7 NI_7 NS_26 0 2.4925963286568016e-04
GC_7_27 b_7 NI_7 NS_27 0 3.1983861974449841e-05
GC_7_28 b_7 NI_7 NS_28 0 -8.8753281140121233e-06
GC_7_29 b_7 NI_7 NS_29 0 5.6251791663293018e-06
GC_7_30 b_7 NI_7 NS_30 0 -1.1560722833079090e-05
GC_7_31 b_7 NI_7 NS_31 0 6.1009966378419050e-04
GC_7_32 b_7 NI_7 NS_32 0 -1.7156158849538232e-05
GC_7_33 b_7 NI_7 NS_33 0 3.0105783990231258e-06
GC_7_34 b_7 NI_7 NS_34 0 8.8667497954694643e-07
GC_7_35 b_7 NI_7 NS_35 0 6.3021192656896752e-03
GC_7_36 b_7 NI_7 NS_36 0 -4.8523183435758181e-04
GC_7_37 b_7 NI_7 NS_37 0 -2.3563503224703845e-07
GC_7_38 b_7 NI_7 NS_38 0 2.0297667139674028e-09
GC_7_39 b_7 NI_7 NS_39 0 -1.7529292272707401e-03
GC_7_40 b_7 NI_7 NS_40 0 1.9670466786717369e-03
GC_7_41 b_7 NI_7 NS_41 0 -5.9233315903076220e-04
GC_7_42 b_7 NI_7 NS_42 0 8.6220035894382251e-04
GC_7_43 b_7 NI_7 NS_43 0 1.0952545005728620e-03
GC_7_44 b_7 NI_7 NS_44 0 -1.0969412772404679e-03
GC_7_45 b_7 NI_7 NS_45 0 -1.2933335593663785e-03
GC_7_46 b_7 NI_7 NS_46 0 -3.1772190865540670e-04
GC_7_47 b_7 NI_7 NS_47 0 -1.5279832634677631e-06
GC_7_48 b_7 NI_7 NS_48 0 3.3437120450130647e-07
GC_7_49 b_7 NI_7 NS_49 0 5.1384323221686196e-06
GC_7_50 b_7 NI_7 NS_50 0 -1.8057624122574487e-05
GC_7_51 b_7 NI_7 NS_51 0 2.1377371073490179e-04
GC_7_52 b_7 NI_7 NS_52 0 1.5569633027185200e-04
GC_7_53 b_7 NI_7 NS_53 0 -6.8565110892957003e-06
GC_7_54 b_7 NI_7 NS_54 0 5.3984649780299798e-06
GC_7_55 b_7 NI_7 NS_55 0 -9.2285334790373038e-05
GC_7_56 b_7 NI_7 NS_56 0 -5.0608525620140898e-05
GC_7_57 b_7 NI_7 NS_57 0 1.3333682742486236e-06
GC_7_58 b_7 NI_7 NS_58 0 -8.2508048437780410e-07
GC_7_59 b_7 NI_7 NS_59 0 -3.2746501875499076e-04
GC_7_60 b_7 NI_7 NS_60 0 2.0147154469170737e-04
GC_7_61 b_7 NI_7 NS_61 0 -4.8480662356705933e-06
GC_7_62 b_7 NI_7 NS_62 0 2.3607231688729464e-05
GC_7_63 b_7 NI_7 NS_63 0 -4.0408717148428937e-06
GC_7_64 b_7 NI_7 NS_64 0 1.4044851644367170e-05
GC_7_65 b_7 NI_7 NS_65 0 4.2754547028501047e-04
GC_7_66 b_7 NI_7 NS_66 0 -2.1230034161668599e-04
GC_7_67 b_7 NI_7 NS_67 0 -5.7389551729573700e-06
GC_7_68 b_7 NI_7 NS_68 0 -1.5729883527850475e-05
GC_7_69 b_7 NI_7 NS_69 0 -1.2182969463431703e-02
GC_7_70 b_7 NI_7 NS_70 0 1.5127463584190934e-03
GC_7_71 b_7 NI_7 NS_71 0 -3.3241718608319450e-06
GC_7_72 b_7 NI_7 NS_72 0 -2.1976805161879196e-09
GC_7_73 b_7 NI_7 NS_73 0 2.9892911221719117e-03
GC_7_74 b_7 NI_7 NS_74 0 -2.4636886532097505e-03
GC_7_75 b_7 NI_7 NS_75 0 4.8879450687479330e-04
GC_7_76 b_7 NI_7 NS_76 0 -9.6542722386783270e-05
GC_7_77 b_7 NI_7 NS_77 0 -1.0400652308267693e-03
GC_7_78 b_7 NI_7 NS_78 0 -4.3708536237982643e-04
GC_7_79 b_7 NI_7 NS_79 0 1.1709985673143191e-03
GC_7_80 b_7 NI_7 NS_80 0 1.7045205419919911e-04
GC_7_81 b_7 NI_7 NS_81 0 2.9974084387633192e-07
GC_7_82 b_7 NI_7 NS_82 0 1.3651905231572448e-06
GC_7_83 b_7 NI_7 NS_83 0 1.6036026719554953e-06
GC_7_84 b_7 NI_7 NS_84 0 -3.7533199661686696e-06
GC_7_85 b_7 NI_7 NS_85 0 1.6137306341497138e-04
GC_7_86 b_7 NI_7 NS_86 0 -4.7713925001475436e-05
GC_7_87 b_7 NI_7 NS_87 0 -9.3179771460827150e-07
GC_7_88 b_7 NI_7 NS_88 0 -5.3192012001567976e-06
GC_7_89 b_7 NI_7 NS_89 0 -5.6222236355036466e-05
GC_7_90 b_7 NI_7 NS_90 0 -5.3174155503303013e-06
GC_7_91 b_7 NI_7 NS_91 0 2.7875374455515758e-06
GC_7_92 b_7 NI_7 NS_92 0 3.7719158238574910e-06
GC_7_93 b_7 NI_7 NS_93 0 2.2642360559110847e-04
GC_7_94 b_7 NI_7 NS_94 0 1.1810399845972606e-04
GC_7_95 b_7 NI_7 NS_95 0 -3.0719019264778658e-05
GC_7_96 b_7 NI_7 NS_96 0 1.3608512050652233e-05
GC_7_97 b_7 NI_7 NS_97 0 2.4674886334141358e-06
GC_7_98 b_7 NI_7 NS_98 0 -7.8408045845661112e-06
GC_7_99 b_7 NI_7 NS_99 0 5.9446190408749824e-04
GC_7_100 b_7 NI_7 NS_100 0 1.8328742760273315e-05
GC_7_101 b_7 NI_7 NS_101 0 1.8685429442273524e-06
GC_7_102 b_7 NI_7 NS_102 0 8.0899735263990939e-07
GC_7_103 b_7 NI_7 NS_103 0 1.6300902114362272e-02
GC_7_104 b_7 NI_7 NS_104 0 -1.1352095280791335e-03
GC_7_105 b_7 NI_7 NS_105 0 -3.5750731502236731e-07
GC_7_106 b_7 NI_7 NS_106 0 3.7690159332734756e-09
GC_7_107 b_7 NI_7 NS_107 0 -2.7066875603831289e-03
GC_7_108 b_7 NI_7 NS_108 0 5.8402546149941255e-03
GC_7_109 b_7 NI_7 NS_109 0 5.1197853210600310e-04
GC_7_110 b_7 NI_7 NS_110 0 -8.9615446632327711e-04
GC_7_111 b_7 NI_7 NS_111 0 -5.1273461322416209e-03
GC_7_112 b_7 NI_7 NS_112 0 -2.0836614595096479e-03
GC_7_113 b_7 NI_7 NS_113 0 -1.6635040020136973e-03
GC_7_114 b_7 NI_7 NS_114 0 2.1256905395813383e-03
GC_7_115 b_7 NI_7 NS_115 0 -6.3217909495993197e-08
GC_7_116 b_7 NI_7 NS_116 0 -2.7912609971006112e-07
GC_7_117 b_7 NI_7 NS_117 0 5.4974348595560928e-06
GC_7_118 b_7 NI_7 NS_118 0 -1.8741474203053373e-05
GC_7_119 b_7 NI_7 NS_119 0 2.2025717437800625e-04
GC_7_120 b_7 NI_7 NS_120 0 1.5559196205531219e-04
GC_7_121 b_7 NI_7 NS_121 0 -3.2405082461791811e-06
GC_7_122 b_7 NI_7 NS_122 0 4.3866654181432811e-06
GC_7_123 b_7 NI_7 NS_123 0 -6.3858213474351949e-05
GC_7_124 b_7 NI_7 NS_124 0 -3.3516335562008744e-05
GC_7_125 b_7 NI_7 NS_125 0 4.1296702311904974e-06
GC_7_126 b_7 NI_7 NS_126 0 -1.8922747460380279e-06
GC_7_127 b_7 NI_7 NS_127 0 1.3105258968907369e-04
GC_7_128 b_7 NI_7 NS_128 0 5.3620921872703417e-05
GC_7_129 b_7 NI_7 NS_129 0 1.9051505783012243e-06
GC_7_130 b_7 NI_7 NS_130 0 -9.5269217416974014e-06
GC_7_131 b_7 NI_7 NS_131 0 -3.6347725174475549e-06
GC_7_132 b_7 NI_7 NS_132 0 6.5922657014439617e-06
GC_7_133 b_7 NI_7 NS_133 0 4.0826133894212994e-04
GC_7_134 b_7 NI_7 NS_134 0 -1.4713924496800740e-04
GC_7_135 b_7 NI_7 NS_135 0 -6.8246002260244941e-06
GC_7_136 b_7 NI_7 NS_136 0 -1.5527401808320491e-05
GC_7_137 b_7 NI_7 NS_137 0 -2.4578683792133689e-02
GC_7_138 b_7 NI_7 NS_138 0 2.3109324713985473e-03
GC_7_139 b_7 NI_7 NS_139 0 -1.1969288085985311e-05
GC_7_140 b_7 NI_7 NS_140 0 -6.5212986068258466e-09
GC_7_141 b_7 NI_7 NS_141 0 9.9904325170989978e-03
GC_7_142 b_7 NI_7 NS_142 0 -7.1631519529352112e-03
GC_7_143 b_7 NI_7 NS_143 0 8.9129181880669053e-04
GC_7_144 b_7 NI_7 NS_144 0 -5.5497976880868537e-04
GC_7_145 b_7 NI_7 NS_145 0 -2.1589313740661815e-03
GC_7_146 b_7 NI_7 NS_146 0 8.3730779697860662e-04
GC_7_147 b_7 NI_7 NS_147 0 1.8697579183990156e-03
GC_7_148 b_7 NI_7 NS_148 0 2.1874797612346022e-03
GC_7_149 b_7 NI_7 NS_149 0 -9.6504195222339605e-08
GC_7_150 b_7 NI_7 NS_150 0 -3.2649108999113817e-07
GC_7_151 b_7 NI_7 NS_151 0 1.7081423741295994e-06
GC_7_152 b_7 NI_7 NS_152 0 -4.4546909996919903e-06
GC_7_153 b_7 NI_7 NS_153 0 1.5966999074733964e-04
GC_7_154 b_7 NI_7 NS_154 0 -4.2446823709545654e-05
GC_7_155 b_7 NI_7 NS_155 0 -7.7544062900734700e-08
GC_7_156 b_7 NI_7 NS_156 0 -1.4563104737390997e-06
GC_7_157 b_7 NI_7 NS_157 0 -2.0936781085124325e-05
GC_7_158 b_7 NI_7 NS_158 0 1.4234188933379033e-06
GC_7_159 b_7 NI_7 NS_159 0 9.3960745410940893e-07
GC_7_160 b_7 NI_7 NS_160 0 1.2655888658727410e-06
GC_7_161 b_7 NI_7 NS_161 0 8.2956417943038198e-04
GC_7_162 b_7 NI_7 NS_162 0 -1.9269096420187923e-05
GC_7_163 b_7 NI_7 NS_163 0 -8.0481899714629341e-05
GC_7_164 b_7 NI_7 NS_164 0 2.7088140903814880e-05
GC_7_165 b_7 NI_7 NS_165 0 1.0654380499785611e-06
GC_7_166 b_7 NI_7 NS_166 0 -3.4209768063778329e-06
GC_7_167 b_7 NI_7 NS_167 0 6.7614907616212676e-04
GC_7_168 b_7 NI_7 NS_168 0 1.7111328208388719e-05
GC_7_169 b_7 NI_7 NS_169 0 3.6397611861945537e-07
GC_7_170 b_7 NI_7 NS_170 0 1.4601819160563883e-06
GC_7_171 b_7 NI_7 NS_171 0 3.9398691003677246e-02
GC_7_172 b_7 NI_7 NS_172 0 -3.8027458015513216e-03
GC_7_173 b_7 NI_7 NS_173 0 -2.2107981974961209e-07
GC_7_174 b_7 NI_7 NS_174 0 7.6575469703689323e-09
GC_7_175 b_7 NI_7 NS_175 0 -1.2692397775008354e-02
GC_7_176 b_7 NI_7 NS_176 0 1.3989841726815517e-02
GC_7_177 b_7 NI_7 NS_177 0 2.0040860788082073e-03
GC_7_178 b_7 NI_7 NS_178 0 -1.7541345385665788e-03
GC_7_179 b_7 NI_7 NS_179 0 -6.8895800242454400e-03
GC_7_180 b_7 NI_7 NS_180 0 -6.9691634032585719e-03
GC_7_181 b_7 NI_7 NS_181 0 -5.8144427396627195e-03
GC_7_182 b_7 NI_7 NS_182 0 1.5417699163369450e-03
GC_7_183 b_7 NI_7 NS_183 0 1.0895417895338065e-06
GC_7_184 b_7 NI_7 NS_184 0 5.5556074718766602e-07
GC_7_185 b_7 NI_7 NS_185 0 4.8279232122393968e-06
GC_7_186 b_7 NI_7 NS_186 0 -1.8629319594123197e-05
GC_7_187 b_7 NI_7 NS_187 0 2.2422802922418271e-04
GC_7_188 b_7 NI_7 NS_188 0 1.4853378646293393e-04
GC_7_189 b_7 NI_7 NS_189 0 -1.8957992423068588e-06
GC_7_190 b_7 NI_7 NS_190 0 9.9824063271796655e-07
GC_7_191 b_7 NI_7 NS_191 0 -2.5684840989503782e-05
GC_7_192 b_7 NI_7 NS_192 0 -9.5445546021876122e-06
GC_7_193 b_7 NI_7 NS_193 0 2.5020814944428739e-06
GC_7_194 b_7 NI_7 NS_194 0 -3.5815147621036648e-07
GC_7_195 b_7 NI_7 NS_195 0 4.2655454605637779e-04
GC_7_196 b_7 NI_7 NS_196 0 -1.7189299241006606e-04
GC_7_197 b_7 NI_7 NS_197 0 -1.9651569830372679e-06
GC_7_198 b_7 NI_7 NS_198 0 -3.6011901431196111e-05
GC_7_199 b_7 NI_7 NS_199 0 -4.9733150068749976e-06
GC_7_200 b_7 NI_7 NS_200 0 3.4938480413594016e-06
GC_7_201 b_7 NI_7 NS_201 0 4.6661137104767807e-04
GC_7_202 b_7 NI_7 NS_202 0 -2.0891821496363971e-04
GC_7_203 b_7 NI_7 NS_203 0 -8.4037803717594768e-06
GC_7_204 b_7 NI_7 NS_204 0 -1.6195804878853653e-05
GC_7_205 b_7 NI_7 NS_205 0 -2.2105767379430408e-01
GC_7_206 b_7 NI_7 NS_206 0 5.6004957284162757e-02
GC_7_207 b_7 NI_7 NS_207 0 4.0814826571303061e-05
GC_7_208 b_7 NI_7 NS_208 0 -5.8077548940950909e-08
GC_7_209 b_7 NI_7 NS_209 0 8.3862769847962801e-02
GC_7_210 b_7 NI_7 NS_210 0 5.5479028958122069e-03
GC_7_211 b_7 NI_7 NS_211 0 2.7959812303380107e-03
GC_7_212 b_7 NI_7 NS_212 0 1.4194919901821931e-03
GC_7_213 b_7 NI_7 NS_213 0 -1.9881186408531779e-03
GC_7_214 b_7 NI_7 NS_214 0 3.4641552296436574e-03
GC_7_215 b_7 NI_7 NS_215 0 -5.8618435258962426e-03
GC_7_216 b_7 NI_7 NS_216 0 5.9285235059740342e-03
GC_7_217 b_7 NI_7 NS_217 0 2.5030538953189653e-07
GC_7_218 b_7 NI_7 NS_218 0 1.4266328126738940e-06
GC_7_219 b_7 NI_7 NS_219 0 2.6748028730263164e-06
GC_7_220 b_7 NI_7 NS_220 0 -4.1276970986816935e-06
GC_7_221 b_7 NI_7 NS_221 0 1.4812327349713651e-04
GC_7_222 b_7 NI_7 NS_222 0 -4.5917373256396590e-05
GC_7_223 b_7 NI_7 NS_223 0 5.5812821472574181e-07
GC_7_224 b_7 NI_7 NS_224 0 1.2917568486311654e-06
GC_7_225 b_7 NI_7 NS_225 0 2.6437534438817306e-05
GC_7_226 b_7 NI_7 NS_226 0 1.5368590954116895e-05
GC_7_227 b_7 NI_7 NS_227 0 2.8517937460059618e-06
GC_7_228 b_7 NI_7 NS_228 0 8.5522097759554193e-07
GC_7_229 b_7 NI_7 NS_229 0 8.3704442095901331e-04
GC_7_230 b_7 NI_7 NS_230 0 -1.4567804025461854e-04
GC_7_231 b_7 NI_7 NS_231 0 -7.8266303423381715e-05
GC_7_232 b_7 NI_7 NS_232 0 2.2034303164149007e-05
GC_7_233 b_7 NI_7 NS_233 0 -4.1080619306929927e-06
GC_7_234 b_7 NI_7 NS_234 0 4.6061736576720382e-06
GC_7_235 b_7 NI_7 NS_235 0 5.7893465093993761e-04
GC_7_236 b_7 NI_7 NS_236 0 -2.8694311273532228e-05
GC_7_237 b_7 NI_7 NS_237 0 1.9031915522715680e-06
GC_7_238 b_7 NI_7 NS_238 0 1.1072585316905288e-06
GC_7_239 b_7 NI_7 NS_239 0 3.6118853045414165e-02
GC_7_240 b_7 NI_7 NS_240 0 3.2901178109076730e-02
GC_7_241 b_7 NI_7 NS_241 0 1.6608659779673512e-04
GC_7_242 b_7 NI_7 NS_242 0 2.5222102479627659e-07
GC_7_243 b_7 NI_7 NS_243 0 -5.7099385792707520e-02
GC_7_244 b_7 NI_7 NS_244 0 -1.6554041662914010e-02
GC_7_245 b_7 NI_7 NS_245 0 3.0381071847565376e-04
GC_7_246 b_7 NI_7 NS_246 0 2.8396370686485013e-03
GC_7_247 b_7 NI_7 NS_247 0 2.6539842521486499e-03
GC_7_248 b_7 NI_7 NS_248 0 1.8432765990409886e-02
GC_7_249 b_7 NI_7 NS_249 0 1.0450786661727149e-02
GC_7_250 b_7 NI_7 NS_250 0 3.8579154645308291e-03
GC_7_251 b_7 NI_7 NS_251 0 -1.0200232573058210e-06
GC_7_252 b_7 NI_7 NS_252 0 -7.3365615737721665e-07
GC_7_253 b_7 NI_7 NS_253 0 3.5691522700182158e-06
GC_7_254 b_7 NI_7 NS_254 0 -1.9664697103243355e-05
GC_7_255 b_7 NI_7 NS_255 0 2.3864830403772685e-04
GC_7_256 b_7 NI_7 NS_256 0 1.5790963167183969e-04
GC_7_257 b_7 NI_7 NS_257 0 1.6021208006286077e-06
GC_7_258 b_7 NI_7 NS_258 0 1.1959903472291744e-06
GC_7_259 b_7 NI_7 NS_259 0 3.7214412087763496e-05
GC_7_260 b_7 NI_7 NS_260 0 -7.4509706027628245e-06
GC_7_261 b_7 NI_7 NS_261 0 -1.5650600057384704e-06
GC_7_262 b_7 NI_7 NS_262 0 -2.1807384273092135e-06
GC_7_263 b_7 NI_7 NS_263 0 6.2362382787164560e-04
GC_7_264 b_7 NI_7 NS_264 0 -2.4925864212722041e-04
GC_7_265 b_7 NI_7 NS_265 0 -1.9908266407807977e-06
GC_7_266 b_7 NI_7 NS_266 0 -4.5514818561003171e-05
GC_7_267 b_7 NI_7 NS_267 0 -2.9072124866273262e-06
GC_7_268 b_7 NI_7 NS_268 0 -9.4548118162430470e-06
GC_7_269 b_7 NI_7 NS_269 0 5.8460407822737029e-04
GC_7_270 b_7 NI_7 NS_270 0 -6.6855928233880733e-05
GC_7_271 b_7 NI_7 NS_271 0 -1.1291737812030620e-05
GC_7_272 b_7 NI_7 NS_272 0 -1.6930902205911066e-05
GC_7_273 b_7 NI_7 NS_273 0 -1.7778391520302066e-02
GC_7_274 b_7 NI_7 NS_274 0 2.1786079336024991e-03
GC_7_275 b_7 NI_7 NS_275 0 -6.6124705484837135e-06
GC_7_276 b_7 NI_7 NS_276 0 -4.4041428339838611e-09
GC_7_277 b_7 NI_7 NS_277 0 5.5407698558496846e-03
GC_7_278 b_7 NI_7 NS_278 0 -4.5230173731980582e-03
GC_7_279 b_7 NI_7 NS_279 0 4.0038719170724062e-04
GC_7_280 b_7 NI_7 NS_280 0 2.6209851496845389e-04
GC_7_281 b_7 NI_7 NS_281 0 6.1251881775006649e-04
GC_7_282 b_7 NI_7 NS_282 0 6.0960528109209159e-04
GC_7_283 b_7 NI_7 NS_283 0 1.4621434490319682e-03
GC_7_284 b_7 NI_7 NS_284 0 2.9810360270641275e-04
GC_7_285 b_7 NI_7 NS_285 0 -5.0465734478318622e-07
GC_7_286 b_7 NI_7 NS_286 0 -1.6251999825922555e-06
GC_7_287 b_7 NI_7 NS_287 0 1.5745516158433385e-06
GC_7_288 b_7 NI_7 NS_288 0 -3.9815566687363300e-06
GC_7_289 b_7 NI_7 NS_289 0 1.6202374069076617e-04
GC_7_290 b_7 NI_7 NS_290 0 -4.7085097781530384e-05
GC_7_291 b_7 NI_7 NS_291 0 2.3014984815416448e-06
GC_7_292 b_7 NI_7 NS_292 0 6.1542418435430563e-06
GC_7_293 b_7 NI_7 NS_293 0 4.8461287675382141e-05
GC_7_294 b_7 NI_7 NS_294 0 6.6357721651424614e-06
GC_7_295 b_7 NI_7 NS_295 0 2.6422803665982075e-06
GC_7_296 b_7 NI_7 NS_296 0 3.7288709732751735e-06
GC_7_297 b_7 NI_7 NS_297 0 3.6947047039453989e-04
GC_7_298 b_7 NI_7 NS_298 0 -1.2188342342622763e-04
GC_7_299 b_7 NI_7 NS_299 0 -2.3367852352202634e-05
GC_7_300 b_7 NI_7 NS_300 0 -6.6910662785453605e-06
GC_7_301 b_7 NI_7 NS_301 0 -3.1818549239852671e-06
GC_7_302 b_7 NI_7 NS_302 0 7.0909937763915366e-06
GC_7_303 b_7 NI_7 NS_303 0 5.4875940473383977e-04
GC_7_304 b_7 NI_7 NS_304 0 4.0365143832332001e-05
GC_7_305 b_7 NI_7 NS_305 0 9.5606496971545286e-07
GC_7_306 b_7 NI_7 NS_306 0 -3.4755857646609014e-07
GC_7_307 b_7 NI_7 NS_307 0 2.5740500079821961e-02
GC_7_308 b_7 NI_7 NS_308 0 -2.0976068903327599e-03
GC_7_309 b_7 NI_7 NS_309 0 -1.0947919408435835e-06
GC_7_310 b_7 NI_7 NS_310 0 7.2513548591664364e-09
GC_7_311 b_7 NI_7 NS_311 0 -6.9028765993847689e-03
GC_7_312 b_7 NI_7 NS_312 0 1.0506579063186368e-02
GC_7_313 b_7 NI_7 NS_313 0 1.5623150324953307e-03
GC_7_314 b_7 NI_7 NS_314 0 -6.4922338994897186e-04
GC_7_315 b_7 NI_7 NS_315 0 -4.6832293766877493e-03
GC_7_316 b_7 NI_7 NS_316 0 -6.9564974206373972e-03
GC_7_317 b_7 NI_7 NS_317 0 -5.7119223768850166e-03
GC_7_318 b_7 NI_7 NS_318 0 2.4219387619475756e-03
GC_7_319 b_7 NI_7 NS_319 0 1.2990315728960695e-06
GC_7_320 b_7 NI_7 NS_320 0 1.1298257654283665e-06
GC_7_321 b_7 NI_7 NS_321 0 4.9622026277099364e-06
GC_7_322 b_7 NI_7 NS_322 0 -1.9114669066549316e-05
GC_7_323 b_7 NI_7 NS_323 0 2.2449725832379483e-04
GC_7_324 b_7 NI_7 NS_324 0 1.5622514384400267e-04
GC_7_325 b_7 NI_7 NS_325 0 4.7180299343380592e-06
GC_7_326 b_7 NI_7 NS_326 0 -4.1267896311691730e-06
GC_7_327 b_7 NI_7 NS_327 0 5.6541578937594214e-05
GC_7_328 b_7 NI_7 NS_328 0 3.6141683861986508e-05
GC_7_329 b_7 NI_7 NS_329 0 5.6957738103371448e-06
GC_7_330 b_7 NI_7 NS_330 0 -1.4708921991581448e-06
GC_7_331 b_7 NI_7 NS_331 0 1.4100909130500180e-04
GC_7_332 b_7 NI_7 NS_332 0 -1.2193604368578754e-04
GC_7_333 b_7 NI_7 NS_333 0 -5.7452326357799178e-06
GC_7_334 b_7 NI_7 NS_334 0 -1.7327225714343404e-05
GC_7_335 b_7 NI_7 NS_335 0 1.6459941897087785e-06
GC_7_336 b_7 NI_7 NS_336 0 -6.6143337762846285e-06
GC_7_337 b_7 NI_7 NS_337 0 3.3818692100031559e-04
GC_7_338 b_7 NI_7 NS_338 0 -1.6638581928829502e-04
GC_7_339 b_7 NI_7 NS_339 0 -6.5649727651029518e-06
GC_7_340 b_7 NI_7 NS_340 0 -1.5760820030931337e-05
GC_7_341 b_7 NI_7 NS_341 0 -1.2023419092377087e-02
GC_7_342 b_7 NI_7 NS_342 0 1.5260919459704184e-03
GC_7_343 b_7 NI_7 NS_343 0 -3.1104012823549747e-06
GC_7_344 b_7 NI_7 NS_344 0 -2.7309963060117682e-09
GC_7_345 b_7 NI_7 NS_345 0 2.7363513933532945e-03
GC_7_346 b_7 NI_7 NS_346 0 -2.1648117517680580e-03
GC_7_347 b_7 NI_7 NS_347 0 -7.8970066021462066e-04
GC_7_348 b_7 NI_7 NS_348 0 8.0138126679632645e-04
GC_7_349 b_7 NI_7 NS_349 0 2.4482986074664224e-03
GC_7_350 b_7 NI_7 NS_350 0 -5.3758980399439113e-04
GC_7_351 b_7 NI_7 NS_351 0 -4.7796306483866593e-05
GC_7_352 b_7 NI_7 NS_352 0 -5.3654918575454476e-04
GC_7_353 b_7 NI_7 NS_353 0 -1.1099919288308560e-06
GC_7_354 b_7 NI_7 NS_354 0 -2.0123166377973366e-06
GC_7_355 b_7 NI_7 NS_355 0 1.3370501714709121e-06
GC_7_356 b_7 NI_7 NS_356 0 -3.8185050233590836e-06
GC_7_357 b_7 NI_7 NS_357 0 1.5648782207699282e-04
GC_7_358 b_7 NI_7 NS_358 0 -4.4825149571404577e-05
GC_7_359 b_7 NI_7 NS_359 0 1.5539125833697816e-06
GC_7_360 b_7 NI_7 NS_360 0 8.5738736675557685e-06
GC_7_361 b_7 NI_7 NS_361 0 8.4905604113631679e-05
GC_7_362 b_7 NI_7 NS_362 0 6.1729064926317469e-06
GC_7_363 b_7 NI_7 NS_363 0 1.5450320047440889e-07
GC_7_364 b_7 NI_7 NS_364 0 8.5063055174734090e-07
GC_7_365 b_7 NI_7 NS_365 0 -2.4355781583708922e-04
GC_7_366 b_7 NI_7 NS_366 0 -8.8488604710477165e-05
GC_7_367 b_7 NI_7 NS_367 0 4.1292908686097894e-05
GC_7_368 b_7 NI_7 NS_368 0 -3.3063222116587220e-05
GC_7_369 b_7 NI_7 NS_369 0 -5.5267406492114198e-06
GC_7_370 b_7 NI_7 NS_370 0 9.4374254855421016e-06
GC_7_371 b_7 NI_7 NS_371 0 5.3645398236419172e-04
GC_7_372 b_7 NI_7 NS_372 0 1.4628629135243103e-05
GC_7_373 b_7 NI_7 NS_373 0 1.9965236519969796e-06
GC_7_374 b_7 NI_7 NS_374 0 -6.6339708884354423e-07
GC_7_375 b_7 NI_7 NS_375 0 1.3936744846619040e-02
GC_7_376 b_7 NI_7 NS_376 0 -1.2484194231042417e-03
GC_7_377 b_7 NI_7 NS_377 0 2.8352968579886967e-07
GC_7_378 b_7 NI_7 NS_378 0 3.8421647041486327e-09
GC_7_379 b_7 NI_7 NS_379 0 -4.7465211065939681e-03
GC_7_380 b_7 NI_7 NS_380 0 5.5905923155164742e-03
GC_7_381 b_7 NI_7 NS_381 0 -1.3138895257199101e-04
GC_7_382 b_7 NI_7 NS_382 0 1.0235719868745702e-03
GC_7_383 b_7 NI_7 NS_383 0 8.8111154574122648e-04
GC_7_384 b_7 NI_7 NS_384 0 -4.4268491399224149e-03
GC_7_385 b_7 NI_7 NS_385 0 -4.1857698833725867e-03
GC_7_386 b_7 NI_7 NS_386 0 -1.4272711829487507e-05
GC_7_387 b_7 NI_7 NS_387 0 3.1299331269864953e-08
GC_7_388 b_7 NI_7 NS_388 0 1.3833941497988372e-06
GC_7_389 b_7 NI_7 NS_389 0 5.0846045067941040e-06
GC_7_390 b_7 NI_7 NS_390 0 -1.8531650370893533e-05
GC_7_391 b_7 NI_7 NS_391 0 2.1293939324695696e-04
GC_7_392 b_7 NI_7 NS_392 0 1.5751652131911853e-04
GC_7_393 b_7 NI_7 NS_393 0 7.4030530525224811e-06
GC_7_394 b_7 NI_7 NS_394 0 -5.0261408487172666e-06
GC_7_395 b_7 NI_7 NS_395 0 8.8747249632210244e-05
GC_7_396 b_7 NI_7 NS_396 0 5.3004724974302409e-05
GC_7_397 b_7 NI_7 NS_397 0 1.3083430985712266e-06
GC_7_398 b_7 NI_7 NS_398 0 -8.3288329406511509e-07
GC_7_399 b_7 NI_7 NS_399 0 -2.0379438739217038e-04
GC_7_400 b_7 NI_7 NS_400 0 -5.2154924728486936e-05
GC_7_401 b_7 NI_7 NS_401 0 -9.3552807206169868e-06
GC_7_402 b_7 NI_7 NS_402 0 1.1802202570288724e-05
GC_7_403 b_7 NI_7 NS_403 0 4.6625648753280074e-06
GC_7_404 b_7 NI_7 NS_404 0 -1.0818819039668815e-05
GC_7_405 b_7 NI_7 NS_405 0 3.7299569678764152e-04
GC_7_406 b_7 NI_7 NS_406 0 -1.7985701727822235e-04
GC_7_407 b_7 NI_7 NS_407 0 -6.6060902977622797e-06
GC_7_408 b_7 NI_7 NS_408 0 -1.6686381589305360e-05
GD_7_1 b_7 NI_7 NA_1 0 1.8204794536386718e-03
GD_7_2 b_7 NI_7 NA_2 0 -5.3303552334879297e-03
GD_7_3 b_7 NI_7 NA_3 0 7.7119980859052641e-03
GD_7_4 b_7 NI_7 NA_4 0 -7.9128323227508502e-03
GD_7_5 b_7 NI_7 NA_5 0 1.1444631997385078e-02
GD_7_6 b_7 NI_7 NA_6 0 -1.5077496109543840e-02
GD_7_7 b_7 NI_7 NA_7 0 9.8484722417077078e-02
GD_7_8 b_7 NI_7 NA_8 0 -3.9916235302937100e-02
GD_7_9 b_7 NI_7 NA_9 0 5.8062368438598095e-03
GD_7_10 b_7 NI_7 NA_10 0 -9.6183970673708648e-03
GD_7_11 b_7 NI_7 NA_11 0 6.8515445000185927e-03
GD_7_12 b_7 NI_7 NA_12 0 -6.2212602914455692e-03
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 6.4456076645890738e-03
GC_8_2 b_8 NI_8 NS_2 0 -5.3498891881723944e-04
GC_8_3 b_8 NI_8 NS_3 0 -1.5274965368659877e-07
GC_8_4 b_8 NI_8 NS_4 0 1.9703655189379567e-09
GC_8_5 b_8 NI_8 NS_5 0 -1.8570169331086543e-03
GC_8_6 b_8 NI_8 NS_6 0 2.2024766293488461e-03
GC_8_7 b_8 NI_8 NS_7 0 -3.9584143158859214e-04
GC_8_8 b_8 NI_8 NS_8 0 8.9321588500430589e-04
GC_8_9 b_8 NI_8 NS_9 0 9.6371897874081508e-04
GC_8_10 b_8 NI_8 NS_10 0 -1.7581737738040931e-03
GC_8_11 b_8 NI_8 NS_11 0 -1.6761462395052404e-03
GC_8_12 b_8 NI_8 NS_12 0 -1.3762077783835265e-04
GC_8_13 b_8 NI_8 NS_13 0 2.9027668562378198e-07
GC_8_14 b_8 NI_8 NS_14 0 1.3250059386485847e-06
GC_8_15 b_8 NI_8 NS_15 0 4.8630162020058741e-06
GC_8_16 b_8 NI_8 NS_16 0 -1.7947927876948374e-05
GC_8_17 b_8 NI_8 NS_17 0 2.1644136404267250e-04
GC_8_18 b_8 NI_8 NS_18 0 1.5536782882926046e-04
GC_8_19 b_8 NI_8 NS_19 0 -8.1691623886045291e-06
GC_8_20 b_8 NI_8 NS_20 0 1.5866622488752703e-06
GC_8_21 b_8 NI_8 NS_21 0 -8.3115441279932943e-05
GC_8_22 b_8 NI_8 NS_22 0 -4.1380887588794286e-05
GC_8_23 b_8 NI_8 NS_23 0 2.2215012980947801e-06
GC_8_24 b_8 NI_8 NS_24 0 -8.9785716469413241e-08
GC_8_25 b_8 NI_8 NS_25 0 -3.1780949669257331e-04
GC_8_26 b_8 NI_8 NS_26 0 2.2472202059463617e-04
GC_8_27 b_8 NI_8 NS_27 0 1.6263470697112912e-06
GC_8_28 b_8 NI_8 NS_28 0 2.0683364661414751e-05
GC_8_29 b_8 NI_8 NS_29 0 -1.7045417947880502e-06
GC_8_30 b_8 NI_8 NS_30 0 1.2689147437570736e-05
GC_8_31 b_8 NI_8 NS_31 0 4.2602827045606798e-04
GC_8_32 b_8 NI_8 NS_32 0 -2.1085468201233564e-04
GC_8_33 b_8 NI_8 NS_33 0 -1.0779384952600398e-05
GC_8_34 b_8 NI_8 NS_34 0 -1.8806989501244236e-05
GC_8_35 b_8 NI_8 NS_35 0 -5.7896359764916710e-03
GC_8_36 b_8 NI_8 NS_36 0 -2.7497678827253365e-05
GC_8_37 b_8 NI_8 NS_37 0 -2.5204442267890410e-06
GC_8_38 b_8 NI_8 NS_38 0 -7.2602484043715719e-10
GC_8_39 b_8 NI_8 NS_39 0 1.6323978030745000e-03
GC_8_40 b_8 NI_8 NS_40 0 -4.3337499452629378e-03
GC_8_41 b_8 NI_8 NS_41 0 -2.9015476822279662e-04
GC_8_42 b_8 NI_8 NS_42 0 5.8974323784873224e-04
GC_8_43 b_8 NI_8 NS_43 0 7.3788949153355326e-04
GC_8_44 b_8 NI_8 NS_44 0 1.3739484937081068e-03
GC_8_45 b_8 NI_8 NS_45 0 1.7166822533918650e-03
GC_8_46 b_8 NI_8 NS_46 0 -5.7802790704113553e-05
GC_8_47 b_8 NI_8 NS_47 0 -3.0733744962436864e-07
GC_8_48 b_8 NI_8 NS_48 0 6.6872113543893772e-07
GC_8_49 b_8 NI_8 NS_49 0 7.8606297006299040e-06
GC_8_50 b_8 NI_8 NS_50 0 -8.7460138442289485e-05
GC_8_51 b_8 NI_8 NS_51 0 1.9144427434964002e-05
GC_8_52 b_8 NI_8 NS_52 0 4.3309099588595418e-04
GC_8_53 b_8 NI_8 NS_53 0 1.0851084359893508e-05
GC_8_54 b_8 NI_8 NS_54 0 1.3094906853609532e-05
GC_8_55 b_8 NI_8 NS_55 0 -9.0554765558113065e-05
GC_8_56 b_8 NI_8 NS_56 0 -1.0588300230855218e-04
GC_8_57 b_8 NI_8 NS_57 0 -2.7377920546530239e-07
GC_8_58 b_8 NI_8 NS_58 0 -1.4854607445981325e-07
GC_8_59 b_8 NI_8 NS_59 0 -1.2193564975519982e-04
GC_8_60 b_8 NI_8 NS_60 0 2.2194778783686617e-04
GC_8_61 b_8 NI_8 NS_61 0 -3.8811151307633279e-06
GC_8_62 b_8 NI_8 NS_62 0 -1.6252255528859578e-06
GC_8_63 b_8 NI_8 NS_63 0 1.1926461973206792e-07
GC_8_64 b_8 NI_8 NS_64 0 -7.9284300982634729e-06
GC_8_65 b_8 NI_8 NS_65 0 3.2983690331979865e-04
GC_8_66 b_8 NI_8 NS_66 0 -2.2758407669674392e-04
GC_8_67 b_8 NI_8 NS_67 0 -3.3402909825700344e-05
GC_8_68 b_8 NI_8 NS_68 0 5.3566444942571511e-05
GC_8_69 b_8 NI_8 NS_69 0 1.9539864659851826e-02
GC_8_70 b_8 NI_8 NS_70 0 -1.4587579704421615e-03
GC_8_71 b_8 NI_8 NS_71 0 5.0631618782208103e-07
GC_8_72 b_8 NI_8 NS_72 0 3.5449472667069252e-09
GC_8_73 b_8 NI_8 NS_73 0 -2.8896458367441992e-03
GC_8_74 b_8 NI_8 NS_74 0 6.9183056891248115e-03
GC_8_75 b_8 NI_8 NS_75 0 6.4936763760759973e-04
GC_8_76 b_8 NI_8 NS_76 0 -1.0592189977668238e-03
GC_8_77 b_8 NI_8 NS_77 0 -5.9460610678175622e-03
GC_8_78 b_8 NI_8 NS_78 0 -2.6288933151914222e-03
GC_8_79 b_8 NI_8 NS_79 0 -2.2281767729589578e-03
GC_8_80 b_8 NI_8 NS_80 0 2.7254518752580898e-03
GC_8_81 b_8 NI_8 NS_81 0 1.4086371782063429e-06
GC_8_82 b_8 NI_8 NS_82 0 4.8155757420340916e-07
GC_8_83 b_8 NI_8 NS_83 0 4.8716948360453152e-06
GC_8_84 b_8 NI_8 NS_84 0 -1.8248516149753335e-05
GC_8_85 b_8 NI_8 NS_85 0 2.2516092974016796e-04
GC_8_86 b_8 NI_8 NS_86 0 1.5520201546621548e-04
GC_8_87 b_8 NI_8 NS_87 0 -6.1722616680249591e-06
GC_8_88 b_8 NI_8 NS_88 0 6.6588211048036970e-07
GC_8_89 b_8 NI_8 NS_89 0 -4.6945677731341830e-05
GC_8_90 b_8 NI_8 NS_90 0 -2.4503295372884753e-05
GC_8_91 b_8 NI_8 NS_91 0 5.3163391177240232e-06
GC_8_92 b_8 NI_8 NS_92 0 -9.3506105817022857e-07
GC_8_93 b_8 NI_8 NS_93 0 1.3689602797298109e-04
GC_8_94 b_8 NI_8 NS_94 0 5.5135393666544682e-05
GC_8_95 b_8 NI_8 NS_95 0 -3.6746156388078233e-07
GC_8_96 b_8 NI_8 NS_96 0 -1.3497485671449868e-05
GC_8_97 b_8 NI_8 NS_97 0 -1.3785368402654739e-06
GC_8_98 b_8 NI_8 NS_98 0 6.6746579571404860e-06
GC_8_99 b_8 NI_8 NS_99 0 4.0169371199079499e-04
GC_8_100 b_8 NI_8 NS_100 0 -1.4649294196184527e-04
GC_8_101 b_8 NI_8 NS_101 0 -9.3748913337622158e-06
GC_8_102 b_8 NI_8 NS_102 0 -1.7858700645776702e-05
GC_8_103 b_8 NI_8 NS_103 0 -4.9127777750153359e-03
GC_8_104 b_8 NI_8 NS_104 0 -7.5207590786772311e-04
GC_8_105 b_8 NI_8 NS_105 0 -4.5512761827283214e-06
GC_8_106 b_8 NI_8 NS_106 0 -2.4409739690057217e-09
GC_8_107 b_8 NI_8 NS_107 0 2.3205562928772672e-03
GC_8_108 b_8 NI_8 NS_108 0 -6.8635247908530785e-03
GC_8_109 b_8 NI_8 NS_109 0 -3.5597553101852382e-04
GC_8_110 b_8 NI_8 NS_110 0 -2.1653021975204996e-04
GC_8_111 b_8 NI_8 NS_111 0 -1.6737845002869648e-03
GC_8_112 b_8 NI_8 NS_112 0 3.5898850356951874e-03
GC_8_113 b_8 NI_8 NS_113 0 3.7506861466992223e-03
GC_8_114 b_8 NI_8 NS_114 0 1.1601539480015040e-03
GC_8_115 b_8 NI_8 NS_115 0 7.4442193569425017e-08
GC_8_116 b_8 NI_8 NS_116 0 -8.8681900073433979e-08
GC_8_117 b_8 NI_8 NS_117 0 7.4438665282512068e-06
GC_8_118 b_8 NI_8 NS_118 0 -9.0632568619946927e-05
GC_8_119 b_8 NI_8 NS_119 0 2.8998836190743606e-05
GC_8_120 b_8 NI_8 NS_120 0 4.4602407610476658e-04
GC_8_121 b_8 NI_8 NS_121 0 5.6027058431404405e-06
GC_8_122 b_8 NI_8 NS_122 0 6.3752437512517614e-06
GC_8_123 b_8 NI_8 NS_123 0 -6.1282031221498721e-05
GC_8_124 b_8 NI_8 NS_124 0 -6.4161656577257770e-05
GC_8_125 b_8 NI_8 NS_125 0 -1.4468284807546990e-07
GC_8_126 b_8 NI_8 NS_126 0 -1.0445760200833703e-07
GC_8_127 b_8 NI_8 NS_127 0 1.1598003119330362e-04
GC_8_128 b_8 NI_8 NS_128 0 1.2163957626410961e-05
GC_8_129 b_8 NI_8 NS_129 0 4.8641709262714712e-06
GC_8_130 b_8 NI_8 NS_130 0 2.4934865540611719e-06
GC_8_131 b_8 NI_8 NS_131 0 4.2042018630213669e-07
GC_8_132 b_8 NI_8 NS_132 0 -5.8406542509170704e-06
GC_8_133 b_8 NI_8 NS_133 0 3.2454858332802951e-04
GC_8_134 b_8 NI_8 NS_134 0 -1.7111048346205165e-04
GC_8_135 b_8 NI_8 NS_135 0 -3.1502439749098976e-05
GC_8_136 b_8 NI_8 NS_136 0 5.2850961696935429e-05
GC_8_137 b_8 NI_8 NS_137 0 3.8454742911046308e-02
GC_8_138 b_8 NI_8 NS_138 0 -3.7520081276326014e-03
GC_8_139 b_8 NI_8 NS_139 0 -5.5177037901763975e-07
GC_8_140 b_8 NI_8 NS_140 0 7.7762979387534236e-09
GC_8_141 b_8 NI_8 NS_141 0 -1.2629000922412618e-02
GC_8_142 b_8 NI_8 NS_142 0 1.3572289695441414e-02
GC_8_143 b_8 NI_8 NS_143 0 2.0569629791117659e-03
GC_8_144 b_8 NI_8 NS_144 0 -1.6516364327325676e-03
GC_8_145 b_8 NI_8 NS_145 0 -6.5723459303843107e-03
GC_8_146 b_8 NI_8 NS_146 0 -6.8978476261807370e-03
GC_8_147 b_8 NI_8 NS_147 0 -5.7915730630407909e-03
GC_8_148 b_8 NI_8 NS_148 0 1.3642171335044528e-03
GC_8_149 b_8 NI_8 NS_149 0 1.0765546872575650e-06
GC_8_150 b_8 NI_8 NS_150 0 5.5287466452047075e-07
GC_8_151 b_8 NI_8 NS_151 0 5.2734393886361289e-06
GC_8_152 b_8 NI_8 NS_152 0 -1.9056269407794178e-05
GC_8_153 b_8 NI_8 NS_153 0 2.2164006511371685e-04
GC_8_154 b_8 NI_8 NS_154 0 1.5206293087351101e-04
GC_8_155 b_8 NI_8 NS_155 0 -9.7582818370848662e-07
GC_8_156 b_8 NI_8 NS_156 0 -1.0091765632950008e-07
GC_8_157 b_8 NI_8 NS_157 0 -2.8383041093123451e-05
GC_8_158 b_8 NI_8 NS_158 0 -4.3744720341810213e-06
GC_8_159 b_8 NI_8 NS_159 0 2.4953800004499741e-06
GC_8_160 b_8 NI_8 NS_160 0 -3.1052415658028056e-07
GC_8_161 b_8 NI_8 NS_161 0 4.5430660477625145e-04
GC_8_162 b_8 NI_8 NS_162 0 -1.5640574726895101e-04
GC_8_163 b_8 NI_8 NS_163 0 -4.9385753008221439e-06
GC_8_164 b_8 NI_8 NS_164 0 -3.9842778645483427e-05
GC_8_165 b_8 NI_8 NS_165 0 -5.4037811119432640e-06
GC_8_166 b_8 NI_8 NS_166 0 1.8079695164720970e-06
GC_8_167 b_8 NI_8 NS_167 0 4.7145019782791257e-04
GC_8_168 b_8 NI_8 NS_168 0 -2.1130533646028754e-04
GC_8_169 b_8 NI_8 NS_169 0 -8.1755646093271944e-06
GC_8_170 b_8 NI_8 NS_170 0 -1.5839886118406487e-05
GC_8_171 b_8 NI_8 NS_171 0 -3.6774134597637380e-03
GC_8_172 b_8 NI_8 NS_172 0 -2.0338603920770615e-03
GC_8_173 b_8 NI_8 NS_173 0 -1.2217707399416696e-05
GC_8_174 b_8 NI_8 NS_174 0 -6.2795235008564861e-09
GC_8_175 b_8 NI_8 NS_175 0 6.9045378805828485e-03
GC_8_176 b_8 NI_8 NS_176 0 -9.3401850447258628e-03
GC_8_177 b_8 NI_8 NS_177 0 -3.6092172546548282e-04
GC_8_178 b_8 NI_8 NS_178 0 -2.9917291272877375e-04
GC_8_179 b_8 NI_8 NS_179 0 -3.6364347826075023e-03
GC_8_180 b_8 NI_8 NS_180 0 4.8358168571554063e-03
GC_8_181 b_8 NI_8 NS_181 0 3.2294595112594081e-03
GC_8_182 b_8 NI_8 NS_182 0 3.8338758403074448e-03
GC_8_183 b_8 NI_8 NS_183 0 1.9283583218343988e-07
GC_8_184 b_8 NI_8 NS_184 0 -4.0058210102773033e-07
GC_8_185 b_8 NI_8 NS_185 0 6.5086392272841973e-06
GC_8_186 b_8 NI_8 NS_186 0 -8.9957219597691234e-05
GC_8_187 b_8 NI_8 NS_187 0 4.3652196576468300e-05
GC_8_188 b_8 NI_8 NS_188 0 4.4486709211397530e-04
GC_8_189 b_8 NI_8 NS_189 0 3.6744130457657556e-06
GC_8_190 b_8 NI_8 NS_190 0 4.8664914709081460e-06
GC_8_191 b_8 NI_8 NS_191 0 -1.9158460939989660e-05
GC_8_192 b_8 NI_8 NS_192 0 -3.5878297809324474e-05
GC_8_193 b_8 NI_8 NS_193 0 -1.0708906173049717e-07
GC_8_194 b_8 NI_8 NS_194 0 -1.0085259504641648e-06
GC_8_195 b_8 NI_8 NS_195 0 2.5235126883978019e-04
GC_8_196 b_8 NI_8 NS_196 0 -2.0036361622063889e-04
GC_8_197 b_8 NI_8 NS_197 0 1.0238278650083441e-05
GC_8_198 b_8 NI_8 NS_198 0 4.6973424883066097e-06
GC_8_199 b_8 NI_8 NS_199 0 -1.4850963127521040e-06
GC_8_200 b_8 NI_8 NS_200 0 -4.2845935316806036e-06
GC_8_201 b_8 NI_8 NS_201 0 3.6102275207961464e-04
GC_8_202 b_8 NI_8 NS_202 0 -2.1690425479713713e-04
GC_8_203 b_8 NI_8 NS_203 0 -3.3168601671227379e-05
GC_8_204 b_8 NI_8 NS_204 0 6.2037108356079483e-05
GC_8_205 b_8 NI_8 NS_205 0 3.6118852962850438e-02
GC_8_206 b_8 NI_8 NS_206 0 3.2901178112152228e-02
GC_8_207 b_8 NI_8 NS_207 0 1.6608659793221518e-04
GC_8_208 b_8 NI_8 NS_208 0 2.5222102506678524e-07
GC_8_209 b_8 NI_8 NS_209 0 -5.7099385794151053e-02
GC_8_210 b_8 NI_8 NS_210 0 -1.6554041713479978e-02
GC_8_211 b_8 NI_8 NS_211 0 3.0381070531848310e-04
GC_8_212 b_8 NI_8 NS_212 0 2.8396370671535205e-03
GC_8_213 b_8 NI_8 NS_213 0 2.6539842870026329e-03
GC_8_214 b_8 NI_8 NS_214 0 1.8432766053993188e-02
GC_8_215 b_8 NI_8 NS_215 0 1.0450786690501123e-02
GC_8_216 b_8 NI_8 NS_216 0 3.8579154233918944e-03
GC_8_217 b_8 NI_8 NS_217 0 -1.0200232685184101e-06
GC_8_218 b_8 NI_8 NS_218 0 -7.3365617541285520e-07
GC_8_219 b_8 NI_8 NS_219 0 3.5691522214466255e-06
GC_8_220 b_8 NI_8 NS_220 0 -1.9664697145545529e-05
GC_8_221 b_8 NI_8 NS_221 0 2.3864830433269527e-04
GC_8_222 b_8 NI_8 NS_222 0 1.5790963175562437e-04
GC_8_223 b_8 NI_8 NS_223 0 1.6021207569363909e-06
GC_8_224 b_8 NI_8 NS_224 0 1.1959903789237575e-06
GC_8_225 b_8 NI_8 NS_225 0 3.7214412406378002e-05
GC_8_226 b_8 NI_8 NS_226 0 -7.4509705139469417e-06
GC_8_227 b_8 NI_8 NS_227 0 -1.5650598145485269e-06
GC_8_228 b_8 NI_8 NS_228 0 -2.1807381983636893e-06
GC_8_229 b_8 NI_8 NS_229 0 6.2362382960735971e-04
GC_8_230 b_8 NI_8 NS_230 0 -2.4925864231499262e-04
GC_8_231 b_8 NI_8 NS_231 0 -1.9908265988164019e-06
GC_8_232 b_8 NI_8 NS_232 0 -4.5514818697457807e-05
GC_8_233 b_8 NI_8 NS_233 0 -2.9072125484837368e-06
GC_8_234 b_8 NI_8 NS_234 0 -9.4548118729560651e-06
GC_8_235 b_8 NI_8 NS_235 0 5.8460408070400518e-04
GC_8_236 b_8 NI_8 NS_236 0 -6.6855928459623253e-05
GC_8_237 b_8 NI_8 NS_237 0 -1.1291737838780182e-05
GC_8_238 b_8 NI_8 NS_238 0 -1.6930902081775095e-05
GC_8_239 b_8 NI_8 NS_239 0 1.4186169612531234e-02
GC_8_240 b_8 NI_8 NS_240 0 2.9077957569956452e-02
GC_8_241 b_8 NI_8 NS_241 0 6.3260145885409507e-05
GC_8_242 b_8 NI_8 NS_242 0 -7.0302349429072691e-08
GC_8_243 b_8 NI_8 NS_243 0 4.8375953178860946e-02
GC_8_244 b_8 NI_8 NS_244 0 4.1444030144130617e-02
GC_8_245 b_8 NI_8 NS_245 0 -3.5561866211056802e-03
GC_8_246 b_8 NI_8 NS_246 0 6.3624045132632358e-04
GC_8_247 b_8 NI_8 NS_247 0 -1.3982023790296753e-02
GC_8_248 b_8 NI_8 NS_248 0 1.6129242393673554e-02
GC_8_249 b_8 NI_8 NS_249 0 2.1632679823592200e-03
GC_8_250 b_8 NI_8 NS_250 0 6.4643666299310240e-03
GC_8_251 b_8 NI_8 NS_251 0 -1.0670654161999676e-06
GC_8_252 b_8 NI_8 NS_252 0 -2.4843903736671342e-06
GC_8_253 b_8 NI_8 NS_253 0 6.6904913143085878e-06
GC_8_254 b_8 NI_8 NS_254 0 -8.9013375854307296e-05
GC_8_255 b_8 NI_8 NS_255 0 4.1422856004383435e-05
GC_8_256 b_8 NI_8 NS_256 0 4.3668192054273483e-04
GC_8_257 b_8 NI_8 NS_257 0 -3.0670195263489305e-06
GC_8_258 b_8 NI_8 NS_258 0 -3.5305084029557269e-06
GC_8_259 b_8 NI_8 NS_259 0 2.1351123632954012e-05
GC_8_260 b_8 NI_8 NS_260 0 1.7973360850514117e-05
GC_8_261 b_8 NI_8 NS_261 0 -2.5323699486054146e-06
GC_8_262 b_8 NI_8 NS_262 0 -7.5217523573493384e-09
GC_8_263 b_8 NI_8 NS_263 0 3.6709287780821090e-04
GC_8_264 b_8 NI_8 NS_264 0 -2.3123094804842765e-04
GC_8_265 b_8 NI_8 NS_265 0 1.2434679832332849e-05
GC_8_266 b_8 NI_8 NS_266 0 -1.7994206894433577e-06
GC_8_267 b_8 NI_8 NS_267 0 -9.0104168048851485e-07
GC_8_268 b_8 NI_8 NS_268 0 -1.5118155588277276e-06
GC_8_269 b_8 NI_8 NS_269 0 4.3035108766038729e-04
GC_8_270 b_8 NI_8 NS_270 0 -1.4798832571999608e-04
GC_8_271 b_8 NI_8 NS_271 0 -3.5899622661554434e-05
GC_8_272 b_8 NI_8 NS_272 0 6.2104714043591792e-05
GC_8_273 b_8 NI_8 NS_273 0 2.3333371240479146e-02
GC_8_274 b_8 NI_8 NS_274 0 -1.8683240644925571e-03
GC_8_275 b_8 NI_8 NS_275 0 -1.6903885709722657e-06
GC_8_276 b_8 NI_8 NS_276 0 7.3847305185869226e-09
GC_8_277 b_8 NI_8 NS_277 0 -6.9236399939087345e-03
GC_8_278 b_8 NI_8 NS_278 0 9.6263104092905484e-03
GC_8_279 b_8 NI_8 NS_279 0 1.3142812804751954e-03
GC_8_280 b_8 NI_8 NS_280 0 -6.2517992082713352e-04
GC_8_281 b_8 NI_8 NS_281 0 -3.9891724677713495e-03
GC_8_282 b_8 NI_8 NS_282 0 -6.0814156646032992e-03
GC_8_283 b_8 NI_8 NS_283 0 -5.0774928365282627e-03
GC_8_284 b_8 NI_8 NS_284 0 1.6832883684737958e-03
GC_8_285 b_8 NI_8 NS_285 0 -1.3877231366405029e-07
GC_8_286 b_8 NI_8 NS_286 0 2.5534459003025351e-07
GC_8_287 b_8 NI_8 NS_287 0 5.3297151508651062e-06
GC_8_288 b_8 NI_8 NS_288 0 -1.8588382296628635e-05
GC_8_289 b_8 NI_8 NS_289 0 2.2051713991521726e-04
GC_8_290 b_8 NI_8 NS_290 0 1.5578626515140909e-04
GC_8_291 b_8 NI_8 NS_291 0 7.7028315236788311e-06
GC_8_292 b_8 NI_8 NS_292 0 -1.3769447586689752e-06
GC_8_293 b_8 NI_8 NS_293 0 4.1764237660063899e-05
GC_8_294 b_8 NI_8 NS_294 0 3.3482846759840680e-05
GC_8_295 b_8 NI_8 NS_295 0 5.2550725612901560e-06
GC_8_296 b_8 NI_8 NS_296 0 -4.8495826364367126e-07
GC_8_297 b_8 NI_8 NS_297 0 1.3357278495331276e-04
GC_8_298 b_8 NI_8 NS_298 0 -1.4505217208812324e-04
GC_8_299 b_8 NI_8 NS_299 0 2.0200138068096835e-06
GC_8_300 b_8 NI_8 NS_300 0 -1.2605138108088661e-05
GC_8_301 b_8 NI_8 NS_301 0 -6.7586064515833897e-07
GC_8_302 b_8 NI_8 NS_302 0 -8.6496638671949081e-06
GC_8_303 b_8 NI_8 NS_303 0 3.6146974351865382e-04
GC_8_304 b_8 NI_8 NS_304 0 -1.5508511952677252e-04
GC_8_305 b_8 NI_8 NS_305 0 -9.2250633672166022e-06
GC_8_306 b_8 NI_8 NS_306 0 -1.6650536809679033e-05
GC_8_307 b_8 NI_8 NS_307 0 -2.4727892452595596e-03
GC_8_308 b_8 NI_8 NS_308 0 -2.1404410422217607e-03
GC_8_309 b_8 NI_8 NS_309 0 -5.6405347651437646e-06
GC_8_310 b_8 NI_8 NS_310 0 -6.6599211146302139e-09
GC_8_311 b_8 NI_8 NS_311 0 1.8699579157953081e-03
GC_8_312 b_8 NI_8 NS_312 0 -8.0993383605137935e-03
GC_8_313 b_8 NI_8 NS_313 0 9.7895842147925733e-05
GC_8_314 b_8 NI_8 NS_314 0 -1.3612591063429731e-04
GC_8_315 b_8 NI_8 NS_315 0 -2.0319502763059653e-03
GC_8_316 b_8 NI_8 NS_316 0 1.9463855232590068e-03
GC_8_317 b_8 NI_8 NS_317 0 2.6837535182417335e-03
GC_8_318 b_8 NI_8 NS_318 0 2.4381983261298687e-03
GC_8_319 b_8 NI_8 NS_319 0 3.1569007364304178e-07
GC_8_320 b_8 NI_8 NS_320 0 -6.2394638108743093e-07
GC_8_321 b_8 NI_8 NS_321 0 5.8928463405478877e-06
GC_8_322 b_8 NI_8 NS_322 0 -9.1618194597631821e-05
GC_8_323 b_8 NI_8 NS_323 0 4.2514445546303478e-05
GC_8_324 b_8 NI_8 NS_324 0 4.5508237972961076e-04
GC_8_325 b_8 NI_8 NS_325 0 -4.5880732859386333e-06
GC_8_326 b_8 NI_8 NS_326 0 -5.7899136742462364e-06
GC_8_327 b_8 NI_8 NS_327 0 5.7780559868307821e-05
GC_8_328 b_8 NI_8 NS_328 0 5.0883138198675282e-05
GC_8_329 b_8 NI_8 NS_329 0 4.8887380909221559e-07
GC_8_330 b_8 NI_8 NS_330 0 5.5911292369571818e-07
GC_8_331 b_8 NI_8 NS_331 0 1.0136133604081744e-04
GC_8_332 b_8 NI_8 NS_332 0 -9.7926649852804866e-05
GC_8_333 b_8 NI_8 NS_333 0 5.6059825683967160e-06
GC_8_334 b_8 NI_8 NS_334 0 -2.0302080671969748e-06
GC_8_335 b_8 NI_8 NS_335 0 -2.9368586269290154e-07
GC_8_336 b_8 NI_8 NS_336 0 3.5644610582326871e-06
GC_8_337 b_8 NI_8 NS_337 0 2.9850567919678601e-04
GC_8_338 b_8 NI_8 NS_338 0 -1.6051048169958912e-04
GC_8_339 b_8 NI_8 NS_339 0 -3.1201534354432984e-05
GC_8_340 b_8 NI_8 NS_340 0 5.3477379800696382e-05
GC_8_341 b_8 NI_8 NS_341 0 1.0740925978591751e-02
GC_8_342 b_8 NI_8 NS_342 0 -9.6976192700084216e-04
GC_8_343 b_8 NI_8 NS_343 0 -6.2799767332387998e-07
GC_8_344 b_8 NI_8 NS_344 0 4.1451923359120994e-09
GC_8_345 b_8 NI_8 NS_345 0 -4.8261859198392640e-03
GC_8_346 b_8 NI_8 NS_346 0 4.6840554393832064e-03
GC_8_347 b_8 NI_8 NS_347 0 -1.9243514759718078e-04
GC_8_348 b_8 NI_8 NS_348 0 1.3745685530163203e-03
GC_8_349 b_8 NI_8 NS_349 0 2.0442187716053065e-03
GC_8_350 b_8 NI_8 NS_350 0 -4.4549747358375328e-03
GC_8_351 b_8 NI_8 NS_351 0 -4.0090245214969697e-03
GC_8_352 b_8 NI_8 NS_352 0 -6.7731303179064978e-04
GC_8_353 b_8 NI_8 NS_353 0 -1.6709041333259036e-06
GC_8_354 b_8 NI_8 NS_354 0 6.2749941077405259e-07
GC_8_355 b_8 NI_8 NS_355 0 4.6629313642803109e-06
GC_8_356 b_8 NI_8 NS_356 0 -1.7454699684218823e-05
GC_8_357 b_8 NI_8 NS_357 0 2.1287305560809480e-04
GC_8_358 b_8 NI_8 NS_358 0 1.5128574232116808e-04
GC_8_359 b_8 NI_8 NS_359 0 9.3468072412780423e-06
GC_8_360 b_8 NI_8 NS_360 0 -1.5100336834400396e-06
GC_8_361 b_8 NI_8 NS_361 0 7.7831610161082772e-05
GC_8_362 b_8 NI_8 NS_362 0 4.4691204705768574e-05
GC_8_363 b_8 NI_8 NS_363 0 1.4455558528350435e-06
GC_8_364 b_8 NI_8 NS_364 0 -2.6675599472433161e-07
GC_8_365 b_8 NI_8 NS_365 0 -2.2726106566281387e-04
GC_8_366 b_8 NI_8 NS_366 0 -5.7066904325172742e-05
GC_8_367 b_8 NI_8 NS_367 0 4.9703310774054641e-06
GC_8_368 b_8 NI_8 NS_368 0 1.8016233212741194e-05
GC_8_369 b_8 NI_8 NS_369 0 2.6720324289219830e-06
GC_8_370 b_8 NI_8 NS_370 0 -1.1310600498151365e-05
GC_8_371 b_8 NI_8 NS_371 0 3.7933824271754583e-04
GC_8_372 b_8 NI_8 NS_372 0 -1.7766597389534826e-04
GC_8_373 b_8 NI_8 NS_373 0 -1.1701706426603382e-05
GC_8_374 b_8 NI_8 NS_374 0 -1.8821135874550287e-05
GC_8_375 b_8 NI_8 NS_375 0 -4.9772963625904863e-03
GC_8_376 b_8 NI_8 NS_376 0 -1.1266635021507205e-03
GC_8_377 b_8 NI_8 NS_377 0 -2.6341836392848709e-06
GC_8_378 b_8 NI_8 NS_378 0 -3.8357207781905658e-09
GC_8_379 b_8 NI_8 NS_379 0 1.0462676953431353e-03
GC_8_380 b_8 NI_8 NS_380 0 -6.0151277880830202e-03
GC_8_381 b_8 NI_8 NS_381 0 -8.7833602828229240e-05
GC_8_382 b_8 NI_8 NS_382 0 9.4914417440151392e-04
GC_8_383 b_8 NI_8 NS_383 0 1.1864350842801436e-03
GC_8_384 b_8 NI_8 NS_384 0 1.5554323535880288e-04
GC_8_385 b_8 NI_8 NS_385 0 8.2659459613248782e-04
GC_8_386 b_8 NI_8 NS_386 0 5.1629912963909775e-04
GC_8_387 b_8 NI_8 NS_387 0 -2.9638420366674803e-07
GC_8_388 b_8 NI_8 NS_388 0 -2.2021675746224836e-07
GC_8_389 b_8 NI_8 NS_389 0 6.8168004634307266e-06
GC_8_390 b_8 NI_8 NS_390 0 -8.8474630665708886e-05
GC_8_391 b_8 NI_8 NS_391 0 2.8604114632493713e-05
GC_8_392 b_8 NI_8 NS_392 0 4.4299737981713314e-04
GC_8_393 b_8 NI_8 NS_393 0 -1.0363779088422638e-05
GC_8_394 b_8 NI_8 NS_394 0 -1.2493028354860854e-05
GC_8_395 b_8 NI_8 NS_395 0 8.9670276425075985e-05
GC_8_396 b_8 NI_8 NS_396 0 9.7367343027190831e-05
GC_8_397 b_8 NI_8 NS_397 0 -6.5671015184429849e-07
GC_8_398 b_8 NI_8 NS_398 0 6.5978774146717956e-07
GC_8_399 b_8 NI_8 NS_399 0 -8.9565246176924224e-05
GC_8_400 b_8 NI_8 NS_400 0 2.2613766763481564e-05
GC_8_401 b_8 NI_8 NS_401 0 -3.5415333198195460e-06
GC_8_402 b_8 NI_8 NS_402 0 -9.0492559986798801e-06
GC_8_403 b_8 NI_8 NS_403 0 -1.4574059829762385e-07
GC_8_404 b_8 NI_8 NS_404 0 7.3218988395220009e-06
GC_8_405 b_8 NI_8 NS_405 0 3.1925333122234472e-04
GC_8_406 b_8 NI_8 NS_406 0 -2.0400939837737311e-04
GC_8_407 b_8 NI_8 NS_407 0 -3.4234310081067063e-05
GC_8_408 b_8 NI_8 NS_408 0 5.4063726225776720e-05
GD_8_1 b_8 NI_8 NA_1 0 -4.7377929921478962e-03
GD_8_2 b_8 NI_8 NA_2 0 1.6709479412704480e-03
GD_8_3 b_8 NI_8 NA_3 0 -9.8543400229626991e-03
GD_8_4 b_8 NI_8 NA_4 0 1.3409618009834331e-03
GD_8_5 b_8 NI_8 NA_5 0 -1.4684084197946829e-02
GD_8_6 b_8 NI_8 NA_6 0 -7.2274282389396495e-04
GD_8_7 b_8 NI_8 NA_7 0 -3.9916235283360114e-02
GD_8_8 b_8 NI_8 NA_8 0 -2.5906426024993334e-01
GD_8_9 b_8 NI_8 NA_9 0 -8.0982221532315355e-03
GD_8_10 b_8 NI_8 NA_10 0 3.1638889657657323e-03
GD_8_11 b_8 NI_8 NA_11 0 -3.9371620877495178e-03
GD_8_12 b_8 NI_8 NA_12 0 3.6971917478044948e-03
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 4.2780775545272183e-03
GC_9_2 b_9 NI_9 NS_2 0 -2.4442427659941888e-05
GC_9_3 b_9 NI_9 NS_3 0 2.2728663145574589e-07
GC_9_4 b_9 NI_9 NS_4 0 -8.6803302636143215e-10
GC_9_5 b_9 NI_9 NS_5 0 1.6291288436339434e-03
GC_9_6 b_9 NI_9 NS_6 0 1.5105407174463971e-03
GC_9_7 b_9 NI_9 NS_7 0 9.5865247756229076e-04
GC_9_8 b_9 NI_9 NS_8 0 -8.7360007684605479e-05
GC_9_9 b_9 NI_9 NS_9 0 -5.6543793758830870e-03
GC_9_10 b_9 NI_9 NS_10 0 -9.5774035740114189e-04
GC_9_11 b_9 NI_9 NS_11 0 1.4993382979464531e-03
GC_9_12 b_9 NI_9 NS_12 0 2.3679278433225265e-03
GC_9_13 b_9 NI_9 NS_13 0 1.0637146155661194e-05
GC_9_14 b_9 NI_9 NS_14 0 -2.9607302937779836e-06
GC_9_15 b_9 NI_9 NS_15 0 1.2804731223465866e-06
GC_9_16 b_9 NI_9 NS_16 0 -3.5278309073005505e-06
GC_9_17 b_9 NI_9 NS_17 0 1.6382644657371364e-04
GC_9_18 b_9 NI_9 NS_18 0 -4.1962138139153920e-05
GC_9_19 b_9 NI_9 NS_19 0 -4.1065362809078862e-06
GC_9_20 b_9 NI_9 NS_20 0 -1.8042520802119693e-05
GC_9_21 b_9 NI_9 NS_21 0 -2.1791303482005699e-04
GC_9_22 b_9 NI_9 NS_22 0 -1.3664069101907491e-05
GC_9_23 b_9 NI_9 NS_23 0 6.1487119528707730e-08
GC_9_24 b_9 NI_9 NS_24 0 4.3404358231684215e-06
GC_9_25 b_9 NI_9 NS_25 0 -3.4339548016633001e-04
GC_9_26 b_9 NI_9 NS_26 0 4.2457527417561185e-04
GC_9_27 b_9 NI_9 NS_27 0 1.3347172027170953e-05
GC_9_28 b_9 NI_9 NS_28 0 8.9637009519858066e-06
GC_9_29 b_9 NI_9 NS_29 0 5.0120629594039278e-06
GC_9_30 b_9 NI_9 NS_30 0 -2.3884498494576774e-05
GC_9_31 b_9 NI_9 NS_31 0 5.8616815874442795e-04
GC_9_32 b_9 NI_9 NS_32 0 2.9526529362768570e-05
GC_9_33 b_9 NI_9 NS_33 0 2.6951043442772973e-06
GC_9_34 b_9 NI_9 NS_34 0 2.4424423305051336e-07
GC_9_35 b_9 NI_9 NS_35 0 6.2643044338411375e-03
GC_9_36 b_9 NI_9 NS_36 0 -4.6635257792946715e-04
GC_9_37 b_9 NI_9 NS_37 0 5.2644515671030929e-07
GC_9_38 b_9 NI_9 NS_38 0 8.5729666707193798e-10
GC_9_39 b_9 NI_9 NS_39 0 -4.4023379787443546e-04
GC_9_40 b_9 NI_9 NS_40 0 1.4050096387519979e-03
GC_9_41 b_9 NI_9 NS_41 0 7.1670781981928615e-04
GC_9_42 b_9 NI_9 NS_42 0 -1.6614223459408305e-04
GC_9_43 b_9 NI_9 NS_43 0 -3.5734921309564698e-03
GC_9_44 b_9 NI_9 NS_44 0 -1.3823875921051623e-04
GC_9_45 b_9 NI_9 NS_45 0 8.7967974785522042e-04
GC_9_46 b_9 NI_9 NS_46 0 9.8463327370956473e-04
GC_9_47 b_9 NI_9 NS_47 0 -2.1142382917706802e-06
GC_9_48 b_9 NI_9 NS_48 0 1.1689092252731480e-05
GC_9_49 b_9 NI_9 NS_49 0 4.7477588899698154e-06
GC_9_50 b_9 NI_9 NS_50 0 -1.8050486347383198e-05
GC_9_51 b_9 NI_9 NS_51 0 2.1686576670453312e-04
GC_9_52 b_9 NI_9 NS_52 0 1.6156568952420462e-04
GC_9_53 b_9 NI_9 NS_53 0 -1.6486314446421522e-05
GC_9_54 b_9 NI_9 NS_54 0 1.5243506756267160e-05
GC_9_55 b_9 NI_9 NS_55 0 -2.4229882603106408e-04
GC_9_56 b_9 NI_9 NS_56 0 -1.2113166748674599e-04
GC_9_57 b_9 NI_9 NS_57 0 2.0521153412441863e-06
GC_9_58 b_9 NI_9 NS_58 0 -6.6686309101975140e-07
GC_9_59 b_9 NI_9 NS_59 0 -1.3208029747303036e-04
GC_9_60 b_9 NI_9 NS_60 0 3.1764827592439820e-04
GC_9_61 b_9 NI_9 NS_61 0 -6.6161046956599770e-07
GC_9_62 b_9 NI_9 NS_62 0 1.1199387925560263e-05
GC_9_63 b_9 NI_9 NS_63 0 -1.9951507715464563e-06
GC_9_64 b_9 NI_9 NS_64 0 2.3329564648415064e-05
GC_9_65 b_9 NI_9 NS_65 0 4.2464533875462155e-04
GC_9_66 b_9 NI_9 NS_66 0 -1.5506488968340987e-04
GC_9_67 b_9 NI_9 NS_67 0 -7.3055960461463049e-06
GC_9_68 b_9 NI_9 NS_68 0 -1.4769053502513062e-05
GC_9_69 b_9 NI_9 NS_69 0 1.0790907058165228e-03
GC_9_70 b_9 NI_9 NS_70 0 3.6986590112763154e-04
GC_9_71 b_9 NI_9 NS_71 0 -7.4221642894409143e-07
GC_9_72 b_9 NI_9 NS_72 0 -1.1521192543761998e-09
GC_9_73 b_9 NI_9 NS_73 0 2.5188278887038288e-03
GC_9_74 b_9 NI_9 NS_74 0 8.3574233984148969e-04
GC_9_75 b_9 NI_9 NS_75 0 9.4959851458765164e-04
GC_9_76 b_9 NI_9 NS_76 0 -6.6482084209030623e-04
GC_9_77 b_9 NI_9 NS_77 0 -7.3156009102915958e-03
GC_9_78 b_9 NI_9 NS_78 0 -8.6890700298536058e-04
GC_9_79 b_9 NI_9 NS_79 0 2.4824478534353485e-03
GC_9_80 b_9 NI_9 NS_80 0 2.9941125978072227e-03
GC_9_81 b_9 NI_9 NS_81 0 9.5599118241516124e-06
GC_9_82 b_9 NI_9 NS_82 0 -2.8930231610747309e-06
GC_9_83 b_9 NI_9 NS_83 0 1.5618302144910990e-06
GC_9_84 b_9 NI_9 NS_84 0 -3.3663602173853014e-06
GC_9_85 b_9 NI_9 NS_85 0 1.6490364995346094e-04
GC_9_86 b_9 NI_9 NS_86 0 -4.8937686783918421e-05
GC_9_87 b_9 NI_9 NS_87 0 -1.9579643837876413e-06
GC_9_88 b_9 NI_9 NS_88 0 -1.1770668425427888e-05
GC_9_89 b_9 NI_9 NS_89 0 -1.7597065923211671e-04
GC_9_90 b_9 NI_9 NS_90 0 -2.7651143684768436e-06
GC_9_91 b_9 NI_9 NS_91 0 5.2963550282158017e-06
GC_9_92 b_9 NI_9 NS_92 0 1.0703069288018954e-05
GC_9_93 b_9 NI_9 NS_93 0 -4.0449060801955605e-05
GC_9_94 b_9 NI_9 NS_94 0 3.3603200779643830e-04
GC_9_95 b_9 NI_9 NS_95 0 -4.8728451427344663e-06
GC_9_96 b_9 NI_9 NS_96 0 6.8159909850308001e-06
GC_9_97 b_9 NI_9 NS_97 0 3.1009174934411967e-06
GC_9_98 b_9 NI_9 NS_98 0 -1.5270704217327099e-05
GC_9_99 b_9 NI_9 NS_99 0 5.1361891738543278e-04
GC_9_100 b_9 NI_9 NS_100 0 9.9783714717364925e-05
GC_9_101 b_9 NI_9 NS_101 0 2.0115067240257417e-06
GC_9_102 b_9 NI_9 NS_102 0 -1.2198648014672334e-06
GC_9_103 b_9 NI_9 NS_103 0 1.2731602859921955e-02
GC_9_104 b_9 NI_9 NS_104 0 -8.4088922915392863e-04
GC_9_105 b_9 NI_9 NS_105 0 8.3150706751299832e-07
GC_9_106 b_9 NI_9 NS_106 0 1.3529482288401959e-09
GC_9_107 b_9 NI_9 NS_107 0 -2.5330492146754754e-04
GC_9_108 b_9 NI_9 NS_108 0 3.2320868702207964e-03
GC_9_109 b_9 NI_9 NS_109 0 5.3010339492274249e-04
GC_9_110 b_9 NI_9 NS_110 0 -8.1327885327372844e-04
GC_9_111 b_9 NI_9 NS_111 0 -6.6985401008901879e-03
GC_9_112 b_9 NI_9 NS_112 0 2.1814979152690115e-04
GC_9_113 b_9 NI_9 NS_113 0 1.3645734879909875e-03
GC_9_114 b_9 NI_9 NS_114 0 2.5519262947149598e-03
GC_9_115 b_9 NI_9 NS_115 0 -7.8161726757202053e-07
GC_9_116 b_9 NI_9 NS_116 0 8.8972167433004294e-06
GC_9_117 b_9 NI_9 NS_117 0 4.9389978532591491e-06
GC_9_118 b_9 NI_9 NS_118 0 -1.8813917087134590e-05
GC_9_119 b_9 NI_9 NS_119 0 2.2493266510182711e-04
GC_9_120 b_9 NI_9 NS_120 0 1.6206128579177132e-04
GC_9_121 b_9 NI_9 NS_121 0 -6.6593406268269258e-06
GC_9_122 b_9 NI_9 NS_122 0 1.5108013510597318e-05
GC_9_123 b_9 NI_9 NS_123 0 -2.1050272549685286e-04
GC_9_124 b_9 NI_9 NS_124 0 -8.7765546420438381e-05
GC_9_125 b_9 NI_9 NS_125 0 1.0354574132222429e-05
GC_9_126 b_9 NI_9 NS_126 0 -8.1155611209136291e-07
GC_9_127 b_9 NI_9 NS_127 0 3.1102233579865236e-05
GC_9_128 b_9 NI_9 NS_128 0 2.2468720286608772e-04
GC_9_129 b_9 NI_9 NS_129 0 5.2817774961292535e-06
GC_9_130 b_9 NI_9 NS_130 0 2.5308857637583606e-07
GC_9_131 b_9 NI_9 NS_131 0 -1.1577827098867198e-06
GC_9_132 b_9 NI_9 NS_132 0 1.2849329851610081e-05
GC_9_133 b_9 NI_9 NS_133 0 3.6363086952812706e-04
GC_9_134 b_9 NI_9 NS_134 0 -9.4572865299594416e-05
GC_9_135 b_9 NI_9 NS_135 0 -7.6350517370222275e-06
GC_9_136 b_9 NI_9 NS_136 0 -1.5070718298649345e-05
GC_9_137 b_9 NI_9 NS_137 0 -1.1524578734828343e-02
GC_9_138 b_9 NI_9 NS_138 0 1.5028382728781405e-03
GC_9_139 b_9 NI_9 NS_139 0 -3.3155461469337443e-06
GC_9_140 b_9 NI_9 NS_140 0 -2.1612858118715477e-09
GC_9_141 b_9 NI_9 NS_141 0 3.1885439714747468e-03
GC_9_142 b_9 NI_9 NS_142 0 -2.5019624034808242e-03
GC_9_143 b_9 NI_9 NS_143 0 2.4757069382873174e-04
GC_9_144 b_9 NI_9 NS_144 0 -2.7440475035845735e-04
GC_9_145 b_9 NI_9 NS_145 0 -9.9884777829573014e-04
GC_9_146 b_9 NI_9 NS_146 0 4.3453762789786373e-04
GC_9_147 b_9 NI_9 NS_147 0 1.4320858813477312e-03
GC_9_148 b_9 NI_9 NS_148 0 1.3282549803649387e-04
GC_9_149 b_9 NI_9 NS_149 0 -6.3884606475307025e-07
GC_9_150 b_9 NI_9 NS_150 0 3.0385878458642441e-06
GC_9_151 b_9 NI_9 NS_151 0 1.6337265833809756e-06
GC_9_152 b_9 NI_9 NS_152 0 -3.8354230391141444e-06
GC_9_153 b_9 NI_9 NS_153 0 1.6248306422745416e-04
GC_9_154 b_9 NI_9 NS_154 0 -4.7229210106610947e-05
GC_9_155 b_9 NI_9 NS_155 0 2.1173807949400776e-07
GC_9_156 b_9 NI_9 NS_156 0 -3.8697217842517744e-06
GC_9_157 b_9 NI_9 NS_157 0 -4.6869146911311405e-05
GC_9_158 b_9 NI_9 NS_158 0 3.4179083785770844e-06
GC_9_159 b_9 NI_9 NS_159 0 3.1486075900883506e-06
GC_9_160 b_9 NI_9 NS_160 0 4.7800365815910693e-06
GC_9_161 b_9 NI_9 NS_161 0 1.5357999830623397e-04
GC_9_162 b_9 NI_9 NS_162 0 9.4630131856042693e-05
GC_9_163 b_9 NI_9 NS_163 0 -2.5099752708591496e-05
GC_9_164 b_9 NI_9 NS_164 0 2.4893982614809900e-06
GC_9_165 b_9 NI_9 NS_165 0 2.2973685517516310e-06
GC_9_166 b_9 NI_9 NS_166 0 -5.4819244598590039e-06
GC_9_167 b_9 NI_9 NS_167 0 5.8775318416666119e-04
GC_9_168 b_9 NI_9 NS_168 0 -6.3349391282254909e-06
GC_9_169 b_9 NI_9 NS_169 0 1.6267958313119381e-06
GC_9_170 b_9 NI_9 NS_170 0 6.1434608480281431e-07
GC_9_171 b_9 NI_9 NS_171 0 1.9252399606140350e-02
GC_9_172 b_9 NI_9 NS_172 0 -1.4019191907404273e-03
GC_9_173 b_9 NI_9 NS_173 0 2.9704688845700097e-07
GC_9_174 b_9 NI_9 NS_174 0 3.6651279852820646e-09
GC_9_175 b_9 NI_9 NS_175 0 -2.9344176522639394e-03
GC_9_176 b_9 NI_9 NS_176 0 6.9317190015224621e-03
GC_9_177 b_9 NI_9 NS_177 0 4.8453209783057884e-04
GC_9_178 b_9 NI_9 NS_178 0 -9.3438379029201868e-04
GC_9_179 b_9 NI_9 NS_179 0 -5.3627142156728660e-03
GC_9_180 b_9 NI_9 NS_180 0 -2.7018998286908670e-03
GC_9_181 b_9 NI_9 NS_181 0 -2.3571635980292106e-03
GC_9_182 b_9 NI_9 NS_182 0 2.6137203130178824e-03
GC_9_183 b_9 NI_9 NS_183 0 1.7829410510314040e-06
GC_9_184 b_9 NI_9 NS_184 0 1.3392132078428003e-06
GC_9_185 b_9 NI_9 NS_185 0 4.6156931768843070e-06
GC_9_186 b_9 NI_9 NS_186 0 -1.8386300398508250e-05
GC_9_187 b_9 NI_9 NS_187 0 2.2705407254158355e-04
GC_9_188 b_9 NI_9 NS_188 0 1.5334470545011038e-04
GC_9_189 b_9 NI_9 NS_189 0 -5.8952981119383920e-06
GC_9_190 b_9 NI_9 NS_190 0 1.9408004722781840e-06
GC_9_191 b_9 NI_9 NS_191 0 -3.7069794078240588e-05
GC_9_192 b_9 NI_9 NS_192 0 -2.4795825136500876e-05
GC_9_193 b_9 NI_9 NS_193 0 5.8375808628788018e-06
GC_9_194 b_9 NI_9 NS_194 0 -7.1649673785496897e-07
GC_9_195 b_9 NI_9 NS_195 0 5.2722613289450644e-05
GC_9_196 b_9 NI_9 NS_196 0 4.5308805069849958e-05
GC_9_197 b_9 NI_9 NS_197 0 3.5772896482531648e-06
GC_9_198 b_9 NI_9 NS_198 0 -7.1102902331096374e-06
GC_9_199 b_9 NI_9 NS_199 0 -3.9538077180752958e-07
GC_9_200 b_9 NI_9 NS_200 0 8.3386399838414908e-06
GC_9_201 b_9 NI_9 NS_201 0 3.8217129597562747e-04
GC_9_202 b_9 NI_9 NS_202 0 -1.6632278031411952e-04
GC_9_203 b_9 NI_9 NS_203 0 -8.8253403941028880e-06
GC_9_204 b_9 NI_9 NS_204 0 -1.6230668436182587e-05
GC_9_205 b_9 NI_9 NS_205 0 -1.7778392396978135e-02
GC_9_206 b_9 NI_9 NS_206 0 2.1786080156320073e-03
GC_9_207 b_9 NI_9 NS_207 0 -6.6124713816806817e-06
GC_9_208 b_9 NI_9 NS_208 0 -4.4041324219519401e-09
GC_9_209 b_9 NI_9 NS_209 0 5.5407698410552333e-03
GC_9_210 b_9 NI_9 NS_210 0 -4.5230176046346608e-03
GC_9_211 b_9 NI_9 NS_211 0 4.0038716954193739e-04
GC_9_212 b_9 NI_9 NS_212 0 2.6209856052156400e-04
GC_9_213 b_9 NI_9 NS_213 0 6.1251912528365352e-04
GC_9_214 b_9 NI_9 NS_214 0 6.0960535246500644e-04
GC_9_215 b_9 NI_9 NS_215 0 1.4621434656959416e-03
GC_9_216 b_9 NI_9 NS_216 0 2.9810339469136968e-04
GC_9_217 b_9 NI_9 NS_217 0 -5.0465749141283525e-07
GC_9_218 b_9 NI_9 NS_218 0 -1.6252000566394854e-06
GC_9_219 b_9 NI_9 NS_219 0 1.5745516368072425e-06
GC_9_220 b_9 NI_9 NS_220 0 -3.9815566935404295e-06
GC_9_221 b_9 NI_9 NS_221 0 1.6202374061971073e-04
GC_9_222 b_9 NI_9 NS_222 0 -4.7085097607472371e-05
GC_9_223 b_9 NI_9 NS_223 0 2.3014983616224081e-06
GC_9_224 b_9 NI_9 NS_224 0 6.1542417360692755e-06
GC_9_225 b_9 NI_9 NS_225 0 4.8461287883073841e-05
GC_9_226 b_9 NI_9 NS_226 0 6.6357733445691264e-06
GC_9_227 b_9 NI_9 NS_227 0 2.6422803435089483e-06
GC_9_228 b_9 NI_9 NS_228 0 3.7288712982787986e-06
GC_9_229 b_9 NI_9 NS_229 0 3.6947047176775973e-04
GC_9_230 b_9 NI_9 NS_230 0 -1.2188342861389345e-04
GC_9_231 b_9 NI_9 NS_231 0 -2.3367852416987079e-05
GC_9_232 b_9 NI_9 NS_232 0 -6.6910662077826323e-06
GC_9_233 b_9 NI_9 NS_233 0 -3.1818550162020773e-06
GC_9_234 b_9 NI_9 NS_234 0 7.0909938410558783e-06
GC_9_235 b_9 NI_9 NS_235 0 5.4875940916308786e-04
GC_9_236 b_9 NI_9 NS_236 0 4.0365140520212956e-05
GC_9_237 b_9 NI_9 NS_237 0 9.5606490888659279e-07
GC_9_238 b_9 NI_9 NS_238 0 -3.4755849103727580e-07
GC_9_239 b_9 NI_9 NS_239 0 2.3333371255327657e-02
GC_9_240 b_9 NI_9 NS_240 0 -1.8683240537129221e-03
GC_9_241 b_9 NI_9 NS_241 0 -1.6903891289285324e-06
GC_9_242 b_9 NI_9 NS_242 0 7.3847401566364447e-09
GC_9_243 b_9 NI_9 NS_243 0 -6.9236399793582599e-03
GC_9_244 b_9 NI_9 NS_244 0 9.6263104246176005e-03
GC_9_245 b_9 NI_9 NS_245 0 1.3142812808997607e-03
GC_9_246 b_9 NI_9 NS_246 0 -6.2517993043078614e-04
GC_9_247 b_9 NI_9 NS_247 0 -3.9891724978760919e-03
GC_9_248 b_9 NI_9 NS_248 0 -6.0814156405244128e-03
GC_9_249 b_9 NI_9 NS_249 0 -5.0774928238794441e-03
GC_9_250 b_9 NI_9 NS_250 0 1.6832883705821045e-03
GC_9_251 b_9 NI_9 NS_251 0 -1.3877235075463475e-07
GC_9_252 b_9 NI_9 NS_252 0 2.5534457313773685e-07
GC_9_253 b_9 NI_9 NS_253 0 5.3297151853936724e-06
GC_9_254 b_9 NI_9 NS_254 0 -1.8588382272186462e-05
GC_9_255 b_9 NI_9 NS_255 0 2.2051713967598960e-04
GC_9_256 b_9 NI_9 NS_256 0 1.5578626510793809e-04
GC_9_257 b_9 NI_9 NS_257 0 7.7028315653177443e-06
GC_9_258 b_9 NI_9 NS_258 0 -1.3769447394459206e-06
GC_9_259 b_9 NI_9 NS_259 0 4.1764237404032355e-05
GC_9_260 b_9 NI_9 NS_260 0 3.3482846643882425e-05
GC_9_261 b_9 NI_9 NS_261 0 5.2550726062935078e-06
GC_9_262 b_9 NI_9 NS_262 0 -4.8495830144076974e-07
GC_9_263 b_9 NI_9 NS_263 0 1.3357278624331388e-04
GC_9_264 b_9 NI_9 NS_264 0 -1.4505216979168506e-04
GC_9_265 b_9 NI_9 NS_265 0 2.0200145061563221e-06
GC_9_266 b_9 NI_9 NS_266 0 -1.2605138511260858e-05
GC_9_267 b_9 NI_9 NS_267 0 -6.7586095268086359e-07
GC_9_268 b_9 NI_9 NS_268 0 -8.6496641828972453e-06
GC_9_269 b_9 NI_9 NS_269 0 3.6146974513167609e-04
GC_9_270 b_9 NI_9 NS_270 0 -1.5508511978946609e-04
GC_9_271 b_9 NI_9 NS_271 0 -9.2250634479657421e-06
GC_9_272 b_9 NI_9 NS_272 0 -1.6650536788986404e-05
GC_9_273 b_9 NI_9 NS_273 0 -2.3048863481339468e-01
GC_9_274 b_9 NI_9 NS_274 0 5.7061714307863123e-02
GC_9_275 b_9 NI_9 NS_275 0 3.4329105409039437e-05
GC_9_276 b_9 NI_9 NS_276 0 -5.5335773284275802e-08
GC_9_277 b_9 NI_9 NS_277 0 8.5704351786406077e-02
GC_9_278 b_9 NI_9 NS_278 0 1.1006899096108274e-03
GC_9_279 b_9 NI_9 NS_279 0 7.6996340129787473e-04
GC_9_280 b_9 NI_9 NS_280 0 1.5446894754097972e-03
GC_9_281 b_9 NI_9 NS_281 0 2.4816199003943815e-03
GC_9_282 b_9 NI_9 NS_282 0 8.1647583409929503e-03
GC_9_283 b_9 NI_9 NS_283 0 -3.1929164009863770e-03
GC_9_284 b_9 NI_9 NS_284 0 4.2708121744568315e-03
GC_9_285 b_9 NI_9 NS_285 0 -9.1111436692784221e-06
GC_9_286 b_9 NI_9 NS_286 0 3.6845137176112767e-06
GC_9_287 b_9 NI_9 NS_287 0 3.5461322708233099e-06
GC_9_288 b_9 NI_9 NS_288 0 -3.3655670644077820e-06
GC_9_289 b_9 NI_9 NS_289 0 1.4694335562713309e-04
GC_9_290 b_9 NI_9 NS_290 0 -4.9675134018204962e-05
GC_9_291 b_9 NI_9 NS_291 0 6.8159664547574178e-06
GC_9_292 b_9 NI_9 NS_292 0 1.0915593020977576e-05
GC_9_293 b_9 NI_9 NS_293 0 1.4832592169782899e-04
GC_9_294 b_9 NI_9 NS_294 0 3.1629749267591817e-05
GC_9_295 b_9 NI_9 NS_295 0 9.2809979614479875e-06
GC_9_296 b_9 NI_9 NS_296 0 1.1206105756645182e-05
GC_9_297 b_9 NI_9 NS_297 0 1.8465373333338651e-04
GC_9_298 b_9 NI_9 NS_298 0 -2.8691348907043071e-04
GC_9_299 b_9 NI_9 NS_299 0 -8.9496057788501477e-06
GC_9_300 b_9 NI_9 NS_300 0 -7.5888665537806006e-06
GC_9_301 b_9 NI_9 NS_301 0 -8.8243766502381312e-07
GC_9_302 b_9 NI_9 NS_302 0 1.8793088843583391e-05
GC_9_303 b_9 NI_9 NS_303 0 3.5716364424106303e-04
GC_9_304 b_9 NI_9 NS_304 0 1.2243281657072788e-05
GC_9_305 b_9 NI_9 NS_305 0 3.6938511833438500e-06
GC_9_306 b_9 NI_9 NS_306 0 -1.8026678103289338e-06
GC_9_307 b_9 NI_9 NS_307 0 2.6377228646991754e-02
GC_9_308 b_9 NI_9 NS_308 0 3.3943766034111061e-02
GC_9_309 b_9 NI_9 NS_309 0 1.5544087314345057e-04
GC_9_310 b_9 NI_9 NS_310 0 2.7395448244037608e-07
GC_9_311 b_9 NI_9 NS_311 0 -5.7971853057587668e-02
GC_9_312 b_9 NI_9 NS_312 0 -1.9523358955226486e-02
GC_9_313 b_9 NI_9 NS_313 0 -8.5048812575383025e-04
GC_9_314 b_9 NI_9 NS_314 0 4.6890372796694396e-03
GC_9_315 b_9 NI_9 NS_315 0 9.9946671122744662e-03
GC_9_316 b_9 NI_9 NS_316 0 1.7986124303456506e-02
GC_9_317 b_9 NI_9 NS_317 0 1.0158280822908341e-02
GC_9_318 b_9 NI_9 NS_318 0 1.3966072945028358e-03
GC_9_319 b_9 NI_9 NS_319 0 -8.7988267307520834e-07
GC_9_320 b_9 NI_9 NS_320 0 -8.2600730859958384e-06
GC_9_321 b_9 NI_9 NS_321 0 3.2007960053844404e-06
GC_9_322 b_9 NI_9 NS_322 0 -1.8479701984716023e-05
GC_9_323 b_9 NI_9 NS_323 0 2.4269315572997957e-04
GC_9_324 b_9 NI_9 NS_324 0 1.5663785409542139e-04
GC_9_325 b_9 NI_9 NS_325 0 9.0237503976735897e-06
GC_9_326 b_9 NI_9 NS_326 0 -1.2384717387842416e-05
GC_9_327 b_9 NI_9 NS_327 0 2.0385538859530773e-04
GC_9_328 b_9 NI_9 NS_328 0 6.4185898771064120e-05
GC_9_329 b_9 NI_9 NS_329 0 1.2063455855681007e-05
GC_9_330 b_9 NI_9 NS_330 0 -5.6963167609459224e-07
GC_9_331 b_9 NI_9 NS_331 0 1.1620688519430915e-04
GC_9_332 b_9 NI_9 NS_332 0 -2.7952026570698230e-04
GC_9_333 b_9 NI_9 NS_333 0 -3.9324218917187953e-06
GC_9_334 b_9 NI_9 NS_334 0 -1.1295611412713255e-05
GC_9_335 b_9 NI_9 NS_335 0 4.0268231245209534e-07
GC_9_336 b_9 NI_9 NS_336 0 -1.4577434588897148e-05
GC_9_337 b_9 NI_9 NS_337 0 3.6552633615395474e-04
GC_9_338 b_9 NI_9 NS_338 0 -6.4395370567094136e-05
GC_9_339 b_9 NI_9 NS_339 0 -8.6615743575986289e-06
GC_9_340 b_9 NI_9 NS_340 0 -1.5011367952074047e-05
GC_9_341 b_9 NI_9 NS_341 0 -3.3835124596732956e-02
GC_9_342 b_9 NI_9 NS_342 0 3.2816955007957879e-03
GC_9_343 b_9 NI_9 NS_343 0 -1.5878941234393265e-05
GC_9_344 b_9 NI_9 NS_344 0 -5.7011060155701546e-09
GC_9_345 b_9 NI_9 NS_345 0 1.0193799751307124e-02
GC_9_346 b_9 NI_9 NS_346 0 -1.0005631665709626e-02
GC_9_347 b_9 NI_9 NS_347 0 -1.8931606034215422e-03
GC_9_348 b_9 NI_9 NS_348 0 2.3331609590966664e-04
GC_9_349 b_9 NI_9 NS_349 0 5.6460458546476093e-03
GC_9_350 b_9 NI_9 NS_350 0 3.4668903081221491e-03
GC_9_351 b_9 NI_9 NS_351 0 1.8126045338247513e-03
GC_9_352 b_9 NI_9 NS_352 0 -6.0940552833109777e-04
GC_9_353 b_9 NI_9 NS_353 0 -1.1153607347990862e-05
GC_9_354 b_9 NI_9 NS_354 0 2.9591229282834307e-06
GC_9_355 b_9 NI_9 NS_355 0 2.0985250557413684e-06
GC_9_356 b_9 NI_9 NS_356 0 -3.7144259274978780e-06
GC_9_357 b_9 NI_9 NS_357 0 1.5365448567491573e-04
GC_9_358 b_9 NI_9 NS_358 0 -4.4022668830516496e-05
GC_9_359 b_9 NI_9 NS_359 0 5.6750763489808746e-06
GC_9_360 b_9 NI_9 NS_360 0 1.9312491119877673e-05
GC_9_361 b_9 NI_9 NS_361 0 2.1080976830060058e-04
GC_9_362 b_9 NI_9 NS_362 0 1.6100574326974222e-05
GC_9_363 b_9 NI_9 NS_363 0 1.2459252943378358e-06
GC_9_364 b_9 NI_9 NS_364 0 2.9947500136260750e-06
GC_9_365 b_9 NI_9 NS_365 0 1.7957942685104580e-04
GC_9_366 b_9 NI_9 NS_366 0 -3.8393602584723763e-04
GC_9_367 b_9 NI_9 NS_367 0 1.2979329329586175e-05
GC_9_368 b_9 NI_9 NS_368 0 -1.5583482611603187e-05
GC_9_369 b_9 NI_9 NS_369 0 -4.3320602578248556e-06
GC_9_370 b_9 NI_9 NS_370 0 2.3111133528156850e-05
GC_9_371 b_9 NI_9 NS_371 0 4.2270792083167467e-04
GC_9_372 b_9 NI_9 NS_372 0 4.0240119061734892e-05
GC_9_373 b_9 NI_9 NS_373 0 2.6664227608049595e-06
GC_9_374 b_9 NI_9 NS_374 0 -2.1740411229961431e-06
GC_9_375 b_9 NI_9 NS_375 0 2.9656895282391831e-02
GC_9_376 b_9 NI_9 NS_376 0 -3.2240697027102788e-03
GC_9_377 b_9 NI_9 NS_377 0 -3.0243019347554196e-06
GC_9_378 b_9 NI_9 NS_378 0 1.0013019326749722e-08
GC_9_379 b_9 NI_9 NS_379 0 -1.4820438036213773e-02
GC_9_380 b_9 NI_9 NS_380 0 1.1000113964905358e-02
GC_9_381 b_9 NI_9 NS_381 0 7.4272090439269744e-05
GC_9_382 b_9 NI_9 NS_382 0 1.0507078815430245e-03
GC_9_383 b_9 NI_9 NS_383 0 3.9319046178113333e-03
GC_9_384 b_9 NI_9 NS_384 0 -8.2689639627675920e-03
GC_9_385 b_9 NI_9 NS_385 0 -7.9225737943441239e-03
GC_9_386 b_9 NI_9 NS_386 0 -2.3804952810260495e-03
GC_9_387 b_9 NI_9 NS_387 0 1.7230070630720407e-06
GC_9_388 b_9 NI_9 NS_388 0 -9.5635434321006207e-06
GC_9_389 b_9 NI_9 NS_389 0 5.2441221550967882e-06
GC_9_390 b_9 NI_9 NS_390 0 -1.7522146578804036e-05
GC_9_391 b_9 NI_9 NS_391 0 2.1111779376394162e-04
GC_9_392 b_9 NI_9 NS_392 0 1.5544864456888384e-04
GC_9_393 b_9 NI_9 NS_393 0 1.8456680222168503e-05
GC_9_394 b_9 NI_9 NS_394 0 -1.4649661607402191e-05
GC_9_395 b_9 NI_9 NS_395 0 2.3050904767441202e-04
GC_9_396 b_9 NI_9 NS_396 0 1.2623634413957640e-04
GC_9_397 b_9 NI_9 NS_397 0 5.0505520873998884e-06
GC_9_398 b_9 NI_9 NS_398 0 -2.9278728571162569e-07
GC_9_399 b_9 NI_9 NS_399 0 -7.4157371133087616e-05
GC_9_400 b_9 NI_9 NS_400 0 -3.5714707733436617e-04
GC_9_401 b_9 NI_9 NS_401 0 -1.0631053676210192e-05
GC_9_402 b_9 NI_9 NS_402 0 -4.3754644839212874e-07
GC_9_403 b_9 NI_9 NS_403 0 9.2793586555763696e-07
GC_9_404 b_9 NI_9 NS_404 0 -1.9517769450521893e-05
GC_9_405 b_9 NI_9 NS_405 0 2.6513898960768361e-04
GC_9_406 b_9 NI_9 NS_406 0 -2.0076379050513747e-04
GC_9_407 b_9 NI_9 NS_407 0 -6.1723358290226027e-06
GC_9_408 b_9 NI_9 NS_408 0 -1.5741341472034612e-05
GD_9_1 b_9 NI_9 NA_1 0 -3.4471340395326850e-03
GD_9_2 b_9 NI_9 NA_2 0 -5.1900729096658717e-03
GD_9_3 b_9 NI_9 NA_3 0 6.5939034291084212e-04
GD_9_4 b_9 NI_9 NA_4 0 -9.4804162595827721e-03
GD_9_5 b_9 NI_9 NA_5 0 6.3443277963975576e-03
GD_9_6 b_9 NI_9 NA_6 0 -9.8259845682618311e-03
GD_9_7 b_9 NI_9 NA_7 0 5.8062375642934077e-03
GD_9_8 b_9 NI_9 NA_8 0 -8.0982221953389624e-03
GD_9_9 b_9 NI_9 NA_9 0 1.0014380429093206e-01
GD_9_10 b_9 NI_9 NA_10 0 -3.6009240316180254e-02
GD_9_11 b_9 NI_9 NA_11 0 1.6093931511265383e-02
GD_9_12 b_9 NI_9 NA_12 0 -1.0119953228779448e-02
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 4.7345931239919040e-03
GC_10_2 b_10 NI_10 NS_2 0 -3.4366397665360816e-04
GC_10_3 b_10 NI_10 NS_3 0 1.5106549684211601e-07
GC_10_4 b_10 NI_10 NS_4 0 9.4135327202205412e-10
GC_10_5 b_10 NI_10 NS_5 0 -4.3449916255642831e-04
GC_10_6 b_10 NI_10 NS_6 0 8.6125803679138488e-04
GC_10_7 b_10 NI_10 NS_7 0 6.2368403239653804e-04
GC_10_8 b_10 NI_10 NS_8 0 -2.1825012580032105e-04
GC_10_9 b_10 NI_10 NS_9 0 -3.2458430929379754e-03
GC_10_10 b_10 NI_10 NS_10 0 3.0259882412938963e-04
GC_10_11 b_10 NI_10 NS_11 0 1.1838452400879894e-03
GC_10_12 b_10 NI_10 NS_12 0 5.8640913360021984e-04
GC_10_13 b_10 NI_10 NS_13 0 -1.2006608247065487e-06
GC_10_14 b_10 NI_10 NS_14 0 9.7221990239294080e-06
GC_10_15 b_10 NI_10 NS_15 0 5.2673962328645263e-06
GC_10_16 b_10 NI_10 NS_16 0 -1.8464037509674791e-05
GC_10_17 b_10 NI_10 NS_17 0 2.1399819749199186e-04
GC_10_18 b_10 NI_10 NS_18 0 1.5993556892925223e-04
GC_10_19 b_10 NI_10 NS_19 0 -1.3115166425760577e-05
GC_10_20 b_10 NI_10 NS_20 0 1.3797167748628355e-05
GC_10_21 b_10 NI_10 NS_21 0 -2.5483634954047115e-04
GC_10_22 b_10 NI_10 NS_22 0 -1.0341574828507873e-04
GC_10_23 b_10 NI_10 NS_23 0 2.8834983272898978e-06
GC_10_24 b_10 NI_10 NS_24 0 2.4756065937590648e-07
GC_10_25 b_10 NI_10 NS_25 0 -1.1059815474702066e-04
GC_10_26 b_10 NI_10 NS_26 0 3.2429607805637653e-04
GC_10_27 b_10 NI_10 NS_27 0 5.9064427207464875e-06
GC_10_28 b_10 NI_10 NS_28 0 1.2326823047412884e-05
GC_10_29 b_10 NI_10 NS_29 0 -4.9392300185445654e-06
GC_10_30 b_10 NI_10 NS_30 0 1.7366727917652610e-05
GC_10_31 b_10 NI_10 NS_31 0 4.3369367172690768e-04
GC_10_32 b_10 NI_10 NS_32 0 -1.4839602084086006e-04
GC_10_33 b_10 NI_10 NS_33 0 -1.0122545971081957e-05
GC_10_34 b_10 NI_10 NS_34 0 -1.6813558988817324e-05
GC_10_35 b_10 NI_10 NS_35 0 -4.6173019676015606e-04
GC_10_36 b_10 NI_10 NS_36 0 -1.1208627305361846e-04
GC_10_37 b_10 NI_10 NS_37 0 -8.0019625527931700e-07
GC_10_38 b_10 NI_10 NS_38 0 -5.5569558209048363e-10
GC_10_39 b_10 NI_10 NS_39 0 1.5551336522293515e-03
GC_10_40 b_10 NI_10 NS_40 0 -1.5631973634058192e-03
GC_10_41 b_10 NI_10 NS_41 0 2.9645586880369266e-04
GC_10_42 b_10 NI_10 NS_42 0 -4.4836041136607843e-04
GC_10_43 b_10 NI_10 NS_43 0 -2.3601671362829561e-03
GC_10_44 b_10 NI_10 NS_44 0 1.9282171837100876e-03
GC_10_45 b_10 NI_10 NS_45 0 1.8153468150377326e-03
GC_10_46 b_10 NI_10 NS_46 0 3.8370455800140741e-04
GC_10_47 b_10 NI_10 NS_47 0 -1.2365186445302783e-05
GC_10_48 b_10 NI_10 NS_48 0 -2.8898136423095863e-06
GC_10_49 b_10 NI_10 NS_49 0 6.9308393552346285e-06
GC_10_50 b_10 NI_10 NS_50 0 -8.9428339989491975e-05
GC_10_51 b_10 NI_10 NS_51 0 1.7788896003025626e-05
GC_10_52 b_10 NI_10 NS_52 0 4.4732108481862639e-04
GC_10_53 b_10 NI_10 NS_53 0 2.6645754594356438e-05
GC_10_54 b_10 NI_10 NS_54 0 5.5947524041722610e-06
GC_10_55 b_10 NI_10 NS_55 0 -2.4952494131784755e-04
GC_10_56 b_10 NI_10 NS_56 0 -1.7932622736942477e-04
GC_10_57 b_10 NI_10 NS_57 0 -9.2902813779353352e-08
GC_10_58 b_10 NI_10 NS_58 0 2.8214125341276705e-06
GC_10_59 b_10 NI_10 NS_59 0 1.4313752497521666e-05
GC_10_60 b_10 NI_10 NS_60 0 2.3791383102531789e-04
GC_10_61 b_10 NI_10 NS_61 0 6.7360420671779913e-07
GC_10_62 b_10 NI_10 NS_62 0 2.4254125609717691e-06
GC_10_63 b_10 NI_10 NS_63 0 2.2085229880440293e-06
GC_10_64 b_10 NI_10 NS_64 0 -1.3837913943926980e-05
GC_10_65 b_10 NI_10 NS_65 0 3.1315539978905599e-04
GC_10_66 b_10 NI_10 NS_66 0 -2.0751176523839350e-04
GC_10_67 b_10 NI_10 NS_67 0 -3.0450876805000090e-05
GC_10_68 b_10 NI_10 NS_68 0 4.6772907075472424e-05
GC_10_69 b_10 NI_10 NS_69 0 1.2357087775158928e-02
GC_10_70 b_10 NI_10 NS_70 0 -8.3524101144391062e-04
GC_10_71 b_10 NI_10 NS_71 0 7.9833682990120052e-07
GC_10_72 b_10 NI_10 NS_72 0 1.3505754885982753e-09
GC_10_73 b_10 NI_10 NS_73 0 -3.3438272475417116e-04
GC_10_74 b_10 NI_10 NS_74 0 3.1464952091546207e-03
GC_10_75 b_10 NI_10 NS_75 0 5.4102973171624386e-04
GC_10_76 b_10 NI_10 NS_76 0 -8.2844818909817253e-04
GC_10_77 b_10 NI_10 NS_77 0 -6.5662376841553200e-03
GC_10_78 b_10 NI_10 NS_78 0 1.8740072953897104e-04
GC_10_79 b_10 NI_10 NS_79 0 1.2913377266328060e-03
GC_10_80 b_10 NI_10 NS_80 0 2.4130254199949078e-03
GC_10_81 b_10 NI_10 NS_81 0 -5.9102998426158533e-07
GC_10_82 b_10 NI_10 NS_82 0 8.0114927703934715e-06
GC_10_83 b_10 NI_10 NS_83 0 4.9765819209678084e-06
GC_10_84 b_10 NI_10 NS_84 0 -1.8625746570262536e-05
GC_10_85 b_10 NI_10 NS_85 0 2.2553292379757023e-04
GC_10_86 b_10 NI_10 NS_86 0 1.5925064817678270e-04
GC_10_87 b_10 NI_10 NS_87 0 -6.9114932050004536e-06
GC_10_88 b_10 NI_10 NS_88 0 1.1731554699295282e-05
GC_10_89 b_10 NI_10 NS_89 0 -2.0665040990710775e-04
GC_10_90 b_10 NI_10 NS_90 0 -7.2190628965988502e-05
GC_10_91 b_10 NI_10 NS_91 0 1.0482418993598183e-05
GC_10_92 b_10 NI_10 NS_92 0 -4.2889891240142125e-07
GC_10_93 b_10 NI_10 NS_93 0 6.1794823919826840e-05
GC_10_94 b_10 NI_10 NS_94 0 2.3789648061569091e-04
GC_10_95 b_10 NI_10 NS_95 0 2.0787885153740619e-06
GC_10_96 b_10 NI_10 NS_96 0 -3.3484114384450097e-06
GC_10_97 b_10 NI_10 NS_97 0 -1.5157136519148424e-06
GC_10_98 b_10 NI_10 NS_98 0 1.0569425687497188e-05
GC_10_99 b_10 NI_10 NS_99 0 3.6571859213623784e-04
GC_10_100 b_10 NI_10 NS_100 0 -9.1099374630979629e-05
GC_10_101 b_10 NI_10 NS_101 0 -8.1607273804297069e-06
GC_10_102 b_10 NI_10 NS_102 0 -1.6472603830863770e-05
GC_10_103 b_10 NI_10 NS_103 0 1.2332915416069410e-03
GC_10_104 b_10 NI_10 NS_104 0 -4.6498891285266694e-04
GC_10_105 b_10 NI_10 NS_105 0 -9.8632323328785831e-07
GC_10_106 b_10 NI_10 NS_106 0 -1.1653325293524539e-09
GC_10_107 b_10 NI_10 NS_107 0 2.0799342247385748e-03
GC_10_108 b_10 NI_10 NS_108 0 -2.1873212986626167e-03
GC_10_109 b_10 NI_10 NS_109 0 1.8471843080111459e-04
GC_10_110 b_10 NI_10 NS_110 0 -5.2135535402630462e-04
GC_10_111 b_10 NI_10 NS_111 0 -3.6465033491088024e-03
GC_10_112 b_10 NI_10 NS_112 0 2.3603704954216955e-03
GC_10_113 b_10 NI_10 NS_113 0 2.5594549863323501e-03
GC_10_114 b_10 NI_10 NS_114 0 1.3026062354531407e-03
GC_10_115 b_10 NI_10 NS_115 0 -9.6684348706427965e-06
GC_10_116 b_10 NI_10 NS_116 0 -1.9351402809317624e-06
GC_10_117 b_10 NI_10 NS_117 0 6.1010352537726630e-06
GC_10_118 b_10 NI_10 NS_118 0 -9.2664054145529049e-05
GC_10_119 b_10 NI_10 NS_119 0 3.0550624722386510e-05
GC_10_120 b_10 NI_10 NS_120 0 4.6219133516291574e-04
GC_10_121 b_10 NI_10 NS_121 0 2.4328099864403732e-05
GC_10_122 b_10 NI_10 NS_122 0 -3.1911981083693529e-06
GC_10_123 b_10 NI_10 NS_123 0 -2.1045952377661361e-04
GC_10_124 b_10 NI_10 NS_124 0 -1.0665595923016790e-04
GC_10_125 b_10 NI_10 NS_125 0 1.1242573388593096e-06
GC_10_126 b_10 NI_10 NS_126 0 6.6237956703931831e-06
GC_10_127 b_10 NI_10 NS_127 0 8.9366512082654314e-05
GC_10_128 b_10 NI_10 NS_128 0 1.4423243527630290e-04
GC_10_129 b_10 NI_10 NS_129 0 5.0242071570445875e-06
GC_10_130 b_10 NI_10 NS_130 0 2.3546880176338230e-06
GC_10_131 b_10 NI_10 NS_131 0 2.3010161365866188e-06
GC_10_132 b_10 NI_10 NS_132 0 -8.3740559775785090e-06
GC_10_133 b_10 NI_10 NS_133 0 2.6520153753901478e-04
GC_10_134 b_10 NI_10 NS_134 0 -1.5544770678729640e-04
GC_10_135 b_10 NI_10 NS_135 0 -2.8175361977158992e-05
GC_10_136 b_10 NI_10 NS_136 0 4.5776749047949653e-05
GC_10_137 b_10 NI_10 NS_137 0 1.5887108330815573e-02
GC_10_138 b_10 NI_10 NS_138 0 -1.1065483007351897e-03
GC_10_139 b_10 NI_10 NS_139 0 -6.9482761410226685e-07
GC_10_140 b_10 NI_10 NS_140 0 4.0370243047966941e-09
GC_10_141 b_10 NI_10 NS_141 0 -2.6793994926235399e-03
GC_10_142 b_10 NI_10 NS_142 0 5.7506103254746895e-03
GC_10_143 b_10 NI_10 NS_143 0 5.0127015551655282e-04
GC_10_144 b_10 NI_10 NS_144 0 -8.0585931703735071e-04
GC_10_145 b_10 NI_10 NS_145 0 -4.6410356595106518e-03
GC_10_146 b_10 NI_10 NS_146 0 -2.3166589898902133e-03
GC_10_147 b_10 NI_10 NS_147 0 -1.9437663346064768e-03
GC_10_148 b_10 NI_10 NS_148 0 2.0985168268281471e-03
GC_10_149 b_10 NI_10 NS_149 0 -1.3675634831868491e-06
GC_10_150 b_10 NI_10 NS_150 0 -9.4761366413428654e-07
GC_10_151 b_10 NI_10 NS_151 0 5.5591359580563887e-06
GC_10_152 b_10 NI_10 NS_152 0 -1.9042841596820535e-05
GC_10_153 b_10 NI_10 NS_153 0 2.2142554833841984e-04
GC_10_154 b_10 NI_10 NS_154 0 1.5402699193825366e-04
GC_10_155 b_10 NI_10 NS_155 0 -2.8123794958195715e-06
GC_10_156 b_10 NI_10 NS_156 0 1.1745248490257218e-06
GC_10_157 b_10 NI_10 NS_157 0 -5.0332746951517896e-05
GC_10_158 b_10 NI_10 NS_158 0 -1.4751892427487686e-05
GC_10_159 b_10 NI_10 NS_159 0 5.0029522132263445e-06
GC_10_160 b_10 NI_10 NS_160 0 -1.8290711292860468e-06
GC_10_161 b_10 NI_10 NS_161 0 1.1691826845729411e-04
GC_10_162 b_10 NI_10 NS_162 0 8.9643912861467022e-05
GC_10_163 b_10 NI_10 NS_163 0 -3.8140015818317012e-06
GC_10_164 b_10 NI_10 NS_164 0 -1.4295581012425306e-05
GC_10_165 b_10 NI_10 NS_165 0 -3.4180295690205712e-06
GC_10_166 b_10 NI_10 NS_166 0 4.3446193950113452e-06
GC_10_167 b_10 NI_10 NS_167 0 3.8469774508882634e-04
GC_10_168 b_10 NI_10 NS_168 0 -1.6609326385889171e-04
GC_10_169 b_10 NI_10 NS_169 0 -6.4782699861662027e-06
GC_10_170 b_10 NI_10 NS_170 0 -1.5188851905790642e-05
GC_10_171 b_10 NI_10 NS_171 0 -4.9892366871059054e-03
GC_10_172 b_10 NI_10 NS_172 0 -7.7323316954521859e-04
GC_10_173 b_10 NI_10 NS_173 0 -4.5212466708209343e-06
GC_10_174 b_10 NI_10 NS_174 0 -2.5022812634819196e-09
GC_10_175 b_10 NI_10 NS_175 0 2.3094343804283620e-03
GC_10_176 b_10 NI_10 NS_176 0 -6.8959419883895708e-03
GC_10_177 b_10 NI_10 NS_177 0 -3.1008219149799036e-04
GC_10_178 b_10 NI_10 NS_178 0 -1.7661233471079761e-04
GC_10_179 b_10 NI_10 NS_179 0 -1.6942448083445984e-03
GC_10_180 b_10 NI_10 NS_180 0 3.2544013744003186e-03
GC_10_181 b_10 NI_10 NS_181 0 3.6661984838529476e-03
GC_10_182 b_10 NI_10 NS_182 0 1.3253540305185505e-03
GC_10_183 b_10 NI_10 NS_183 0 -4.6074659727810393e-07
GC_10_184 b_10 NI_10 NS_184 0 2.5372489576375721e-07
GC_10_185 b_10 NI_10 NS_185 0 6.3470710057991505e-06
GC_10_186 b_10 NI_10 NS_186 0 -9.0540277353614275e-05
GC_10_187 b_10 NI_10 NS_187 0 3.7450443113809123e-05
GC_10_188 b_10 NI_10 NS_188 0 4.4414663464575443e-04
GC_10_189 b_10 NI_10 NS_189 0 4.7112137710693838e-06
GC_10_190 b_10 NI_10 NS_190 0 5.1400578276550467e-06
GC_10_191 b_10 NI_10 NS_191 0 -4.8732853494422395e-05
GC_10_192 b_10 NI_10 NS_192 0 -5.7866686895742323e-05
GC_10_193 b_10 NI_10 NS_193 0 2.3619918345203137e-07
GC_10_194 b_10 NI_10 NS_194 0 -2.6185085317846270e-07
GC_10_195 b_10 NI_10 NS_195 0 1.0128345871346912e-04
GC_10_196 b_10 NI_10 NS_196 0 4.6775374395906494e-05
GC_10_197 b_10 NI_10 NS_197 0 7.5007950134572985e-06
GC_10_198 b_10 NI_10 NS_198 0 1.6377463980228366e-06
GC_10_199 b_10 NI_10 NS_199 0 5.4979348982295964e-07
GC_10_200 b_10 NI_10 NS_200 0 -5.8021262262659412e-06
GC_10_201 b_10 NI_10 NS_201 0 3.0645650626092628e-04
GC_10_202 b_10 NI_10 NS_202 0 -1.7220681838990776e-04
GC_10_203 b_10 NI_10 NS_203 0 -3.0380137872329849e-05
GC_10_204 b_10 NI_10 NS_204 0 5.3286493388729955e-05
GC_10_205 b_10 NI_10 NS_205 0 2.5740499808455008e-02
GC_10_206 b_10 NI_10 NS_206 0 -2.0976068390319551e-03
GC_10_207 b_10 NI_10 NS_207 0 -1.0947926686529961e-06
GC_10_208 b_10 NI_10 NS_208 0 7.2513647006353288e-09
GC_10_209 b_10 NI_10 NS_209 0 -6.9028765137921222e-03
GC_10_210 b_10 NI_10 NS_210 0 1.0506578882317923e-02
GC_10_211 b_10 NI_10 NS_211 0 1.5623149900318011e-03
GC_10_212 b_10 NI_10 NS_212 0 -6.4922343608729614e-04
GC_10_213 b_10 NI_10 NS_213 0 -4.6832294280894559e-03
GC_10_214 b_10 NI_10 NS_214 0 -6.9564970339168041e-03
GC_10_215 b_10 NI_10 NS_215 0 -5.7119221359228905e-03
GC_10_216 b_10 NI_10 NS_216 0 2.4219386348828180e-03
GC_10_217 b_10 NI_10 NS_217 0 1.2990317485018807e-06
GC_10_218 b_10 NI_10 NS_218 0 1.1298255907733703e-06
GC_10_219 b_10 NI_10 NS_219 0 4.9622026500544225e-06
GC_10_220 b_10 NI_10 NS_220 0 -1.9114669005070678e-05
GC_10_221 b_10 NI_10 NS_221 0 2.2449725805261247e-04
GC_10_222 b_10 NI_10 NS_222 0 1.5622514328248415e-04
GC_10_223 b_10 NI_10 NS_223 0 4.7180300520798724e-06
GC_10_224 b_10 NI_10 NS_224 0 -4.1267896393294258e-06
GC_10_225 b_10 NI_10 NS_225 0 5.6541577842305166e-05
GC_10_226 b_10 NI_10 NS_226 0 3.6141683787426358e-05
GC_10_227 b_10 NI_10 NS_227 0 5.6957737072678015e-06
GC_10_228 b_10 NI_10 NS_228 0 -1.4708920917742760e-06
GC_10_229 b_10 NI_10 NS_229 0 1.4100910704853631e-04
GC_10_230 b_10 NI_10 NS_230 0 -1.2193603396733039e-04
GC_10_231 b_10 NI_10 NS_231 0 -5.7452300006536825e-06
GC_10_232 b_10 NI_10 NS_232 0 -1.7327227106766947e-05
GC_10_233 b_10 NI_10 NS_233 0 1.6459930377928095e-06
GC_10_234 b_10 NI_10 NS_234 0 -6.6143358552455952e-06
GC_10_235 b_10 NI_10 NS_235 0 3.3818693476706408e-04
GC_10_236 b_10 NI_10 NS_236 0 -1.6638582124996141e-04
GC_10_237 b_10 NI_10 NS_237 0 -6.5649728286709330e-06
GC_10_238 b_10 NI_10 NS_238 0 -1.5760819642921875e-05
GC_10_239 b_10 NI_10 NS_239 0 -2.4727893369617627e-03
GC_10_240 b_10 NI_10 NS_240 0 -2.1404410331977335e-03
GC_10_241 b_10 NI_10 NS_241 0 -5.6405352192729703e-06
GC_10_242 b_10 NI_10 NS_242 0 -6.6599108650051501e-09
GC_10_243 b_10 NI_10 NS_243 0 1.8699578800150266e-03
GC_10_244 b_10 NI_10 NS_244 0 -8.0993383538212668e-03
GC_10_245 b_10 NI_10 NS_245 0 9.7895812634545969e-05
GC_10_246 b_10 NI_10 NS_246 0 -1.3612586224815188e-04
GC_10_247 b_10 NI_10 NS_247 0 -2.0319500257450240e-03
GC_10_248 b_10 NI_10 NS_248 0 1.9463854487649116e-03
GC_10_249 b_10 NI_10 NS_249 0 2.6837533926339936e-03
GC_10_250 b_10 NI_10 NS_250 0 2.4381982875422109e-03
GC_10_251 b_10 NI_10 NS_251 0 3.1568987056633983e-07
GC_10_252 b_10 NI_10 NS_252 0 -6.2394653978942625e-07
GC_10_253 b_10 NI_10 NS_253 0 5.8928463131551336e-06
GC_10_254 b_10 NI_10 NS_254 0 -9.1618194588104083e-05
GC_10_255 b_10 NI_10 NS_255 0 4.2514445699956705e-05
GC_10_256 b_10 NI_10 NS_256 0 4.5508237980534309e-04
GC_10_257 b_10 NI_10 NS_257 0 -4.5880733500244905e-06
GC_10_258 b_10 NI_10 NS_258 0 -5.7899137022809619e-06
GC_10_259 b_10 NI_10 NS_259 0 5.7780560422473740e-05
GC_10_260 b_10 NI_10 NS_260 0 5.0883138329369166e-05
GC_10_261 b_10 NI_10 NS_261 0 4.8887372097300904e-07
GC_10_262 b_10 NI_10 NS_262 0 5.5911296280951561e-07
GC_10_263 b_10 NI_10 NS_263 0 1.0136133259106800e-04
GC_10_264 b_10 NI_10 NS_264 0 -9.7926668951334414e-05
GC_10_265 b_10 NI_10 NS_265 0 5.6059793929518219e-06
GC_10_266 b_10 NI_10 NS_266 0 -2.0302088474052469e-06
GC_10_267 b_10 NI_10 NS_267 0 -2.9368644427029732e-07
GC_10_268 b_10 NI_10 NS_268 0 3.5644639060358630e-06
GC_10_269 b_10 NI_10 NS_269 0 2.9850566763966774e-04
GC_10_270 b_10 NI_10 NS_270 0 -1.6051048694514617e-04
GC_10_271 b_10 NI_10 NS_271 0 -3.1201534177001448e-05
GC_10_272 b_10 NI_10 NS_272 0 5.3477379752633964e-05
GC_10_273 b_10 NI_10 NS_273 0 2.6377228271941090e-02
GC_10_274 b_10 NI_10 NS_274 0 3.3943766074286875e-02
GC_10_275 b_10 NI_10 NS_275 0 1.5544087318339345e-04
GC_10_276 b_10 NI_10 NS_276 0 2.7395447777247941e-07
GC_10_277 b_10 NI_10 NS_277 0 -5.7971852989757593e-02
GC_10_278 b_10 NI_10 NS_278 0 -1.9523359206299318e-02
GC_10_279 b_10 NI_10 NS_279 0 -8.5048815360834603e-04
GC_10_280 b_10 NI_10 NS_280 0 4.6890372188612079e-03
GC_10_281 b_10 NI_10 NS_281 0 9.9946669586183871e-03
GC_10_282 b_10 NI_10 NS_282 0 1.7986124688712333e-02
GC_10_283 b_10 NI_10 NS_283 0 1.0158281180582913e-02
GC_10_284 b_10 NI_10 NS_284 0 1.3966071686541261e-03
GC_10_285 b_10 NI_10 NS_285 0 -8.7988262788526464e-07
GC_10_286 b_10 NI_10 NS_286 0 -8.2600733158448406e-06
GC_10_287 b_10 NI_10 NS_287 0 3.2007960603097015e-06
GC_10_288 b_10 NI_10 NS_288 0 -1.8479701988332949e-05
GC_10_289 b_10 NI_10 NS_289 0 2.4269315514052425e-04
GC_10_290 b_10 NI_10 NS_290 0 1.5663785390251144e-04
GC_10_291 b_10 NI_10 NS_291 0 9.0237506555223417e-06
GC_10_292 b_10 NI_10 NS_292 0 -1.2384717643532482e-05
GC_10_293 b_10 NI_10 NS_293 0 2.0385538607106197e-04
GC_10_294 b_10 NI_10 NS_294 0 6.4185900314386488e-05
GC_10_295 b_10 NI_10 NS_295 0 1.2063454803136384e-05
GC_10_296 b_10 NI_10 NS_296 0 -5.6963006190563599e-07
GC_10_297 b_10 NI_10 NS_297 0 1.1620689029274169e-04
GC_10_298 b_10 NI_10 NS_298 0 -2.7952025080104698e-04
GC_10_299 b_10 NI_10 NS_299 0 -3.9324202599231615e-06
GC_10_300 b_10 NI_10 NS_300 0 -1.1295611703611435e-05
GC_10_301 b_10 NI_10 NS_301 0 4.0268286221255260e-07
GC_10_302 b_10 NI_10 NS_302 0 -1.4577435451276860e-05
GC_10_303 b_10 NI_10 NS_303 0 3.6552635051423609e-04
GC_10_304 b_10 NI_10 NS_304 0 -6.4395354237071177e-05
GC_10_305 b_10 NI_10 NS_305 0 -8.6615748972825440e-06
GC_10_306 b_10 NI_10 NS_306 0 -1.5011368059659242e-05
GC_10_307 b_10 NI_10 NS_307 0 8.1970317144409704e-03
GC_10_308 b_10 NI_10 NS_308 0 2.9804063792575788e-02
GC_10_309 b_10 NI_10 NS_309 0 5.6939211370658875e-05
GC_10_310 b_10 NI_10 NS_310 0 -6.6702373421094939e-08
GC_10_311 b_10 NI_10 NS_311 0 5.0849658642520980e-02
GC_10_312 b_10 NI_10 NS_312 0 3.9022555818531604e-02
GC_10_313 b_10 NI_10 NS_313 0 -3.5123161393005010e-03
GC_10_314 b_10 NI_10 NS_314 0 1.4689605439370799e-03
GC_10_315 b_10 NI_10 NS_315 0 -1.3463639240741850e-02
GC_10_316 b_10 NI_10 NS_316 0 1.4700514077886718e-02
GC_10_317 b_10 NI_10 NS_317 0 3.2249608757335736e-03
GC_10_318 b_10 NI_10 NS_318 0 8.1989888242326309e-03
GC_10_319 b_10 NI_10 NS_319 0 9.7612449681455968e-06
GC_10_320 b_10 NI_10 NS_320 0 1.5509577042510849e-07
GC_10_321 b_10 NI_10 NS_321 0 6.5858874161578971e-06
GC_10_322 b_10 NI_10 NS_322 0 -9.0425676207555312e-05
GC_10_323 b_10 NI_10 NS_323 0 2.9482586197004969e-05
GC_10_324 b_10 NI_10 NS_324 0 4.3881175771395007e-04
GC_10_325 b_10 NI_10 NS_325 0 -2.1476610965299978e-05
GC_10_326 b_10 NI_10 NS_326 0 2.5633192458626627e-06
GC_10_327 b_10 NI_10 NS_327 0 1.9183919571674478e-04
GC_10_328 b_10 NI_10 NS_328 0 9.4588595342064434e-05
GC_10_329 b_10 NI_10 NS_329 0 1.6781246825837781e-06
GC_10_330 b_10 NI_10 NS_330 0 2.3973613961046093e-06
GC_10_331 b_10 NI_10 NS_331 0 2.1106697056901323e-05
GC_10_332 b_10 NI_10 NS_332 0 -6.0826236416921145e-05
GC_10_333 b_10 NI_10 NS_333 0 3.8454997355334328e-06
GC_10_334 b_10 NI_10 NS_334 0 -3.1393971382050069e-06
GC_10_335 b_10 NI_10 NS_335 0 5.7218636134590188e-08
GC_10_336 b_10 NI_10 NS_336 0 6.3663951925201986e-06
GC_10_337 b_10 NI_10 NS_337 0 2.0215556275080668e-04
GC_10_338 b_10 NI_10 NS_338 0 -1.3163279188138136e-05
GC_10_339 b_10 NI_10 NS_339 0 -2.8457049269446445e-05
GC_10_340 b_10 NI_10 NS_340 0 4.4374418120277529e-05
GC_10_341 b_10 NI_10 NS_341 0 3.2850472587252835e-02
GC_10_342 b_10 NI_10 NS_342 0 -3.5239937827609255e-03
GC_10_343 b_10 NI_10 NS_343 0 -1.9760090748773960e-06
GC_10_344 b_10 NI_10 NS_344 0 9.6963953625196126e-09
GC_10_345 b_10 NI_10 NS_345 0 -1.5289655212845926e-02
GC_10_346 b_10 NI_10 NS_346 0 1.2292223627691692e-02
GC_10_347 b_10 NI_10 NS_347 0 5.9227433561263335e-05
GC_10_348 b_10 NI_10 NS_348 0 1.1227030362235876e-03
GC_10_349 b_10 NI_10 NS_349 0 3.7337144562585170e-03
GC_10_350 b_10 NI_10 NS_350 0 -9.1134170382652039e-03
GC_10_351 b_10 NI_10 NS_351 0 -8.6972415420631284e-03
GC_10_352 b_10 NI_10 NS_352 0 -1.9939969079513032e-03
GC_10_353 b_10 NI_10 NS_353 0 1.1834787466760915e-07
GC_10_354 b_10 NI_10 NS_354 0 -8.3061522435479074e-06
GC_10_355 b_10 NI_10 NS_355 0 4.0706506375038552e-06
GC_10_356 b_10 NI_10 NS_356 0 -1.7106739370690922e-05
GC_10_357 b_10 NI_10 NS_357 0 2.1829470490025569e-04
GC_10_358 b_10 NI_10 NS_358 0 1.5154613310346712e-04
GC_10_359 b_10 NI_10 NS_359 0 1.5248662207223610e-05
GC_10_360 b_10 NI_10 NS_360 0 -1.5589035678016964e-05
GC_10_361 b_10 NI_10 NS_361 0 2.4540912509815632e-04
GC_10_362 b_10 NI_10 NS_362 0 1.1630279115578611e-04
GC_10_363 b_10 NI_10 NS_363 0 6.7159694219718895e-06
GC_10_364 b_10 NI_10 NS_364 0 1.0255439571914992e-06
GC_10_365 b_10 NI_10 NS_365 0 -1.3236041109646382e-04
GC_10_366 b_10 NI_10 NS_366 0 -3.9484274743345054e-04
GC_10_367 b_10 NI_10 NS_367 0 -3.3181439416489031e-06
GC_10_368 b_10 NI_10 NS_368 0 4.8895768000356011e-06
GC_10_369 b_10 NI_10 NS_369 0 3.8158362948448041e-06
GC_10_370 b_10 NI_10 NS_370 0 -1.5708439489842647e-05
GC_10_371 b_10 NI_10 NS_371 0 2.5429179030867627e-04
GC_10_372 b_10 NI_10 NS_372 0 -2.1880108610291901e-04
GC_10_373 b_10 NI_10 NS_373 0 -8.2383992345027786e-06
GC_10_374 b_10 NI_10 NS_374 0 -1.6537645436218985e-05
GC_10_375 b_10 NI_10 NS_375 0 -1.5709205027216306e-02
GC_10_376 b_10 NI_10 NS_376 0 -1.2852372777193779e-03
GC_10_377 b_10 NI_10 NS_377 0 -1.6948759460277894e-05
GC_10_378 b_10 NI_10 NS_378 0 -4.9324766628217516e-09
GC_10_379 b_10 NI_10 NS_379 0 7.2871525376396219e-03
GC_10_380 b_10 NI_10 NS_380 0 -1.3528681851472690e-02
GC_10_381 b_10 NI_10 NS_381 0 -9.6944396299748293e-04
GC_10_382 b_10 NI_10 NS_382 0 1.6623626014738305e-03
GC_10_383 b_10 NI_10 NS_383 0 2.2776297773858998e-03
GC_10_384 b_10 NI_10 NS_384 0 3.2069839663737888e-03
GC_10_385 b_10 NI_10 NS_385 0 2.7331975090545664e-03
GC_10_386 b_10 NI_10 NS_386 0 2.2195793986139259e-03
GC_10_387 b_10 NI_10 NS_387 0 1.1760832467426582e-05
GC_10_388 b_10 NI_10 NS_388 0 2.9617407590441483e-06
GC_10_389 b_10 NI_10 NS_389 0 7.0112857658020606e-06
GC_10_390 b_10 NI_10 NS_390 0 -8.8599702108795416e-05
GC_10_391 b_10 NI_10 NS_391 0 2.0588917232839076e-05
GC_10_392 b_10 NI_10 NS_392 0 4.3950844927498356e-04
GC_10_393 b_10 NI_10 NS_393 0 -2.5994275150990319e-05
GC_10_394 b_10 NI_10 NS_394 0 -6.1374918738778291e-06
GC_10_395 b_10 NI_10 NS_395 0 2.4842737250354023e-04
GC_10_396 b_10 NI_10 NS_396 0 1.7728963335768831e-04
GC_10_397 b_10 NI_10 NS_397 0 7.4130882161508581e-07
GC_10_398 b_10 NI_10 NS_398 0 1.1002428152899740e-06
GC_10_399 b_10 NI_10 NS_399 0 -8.7761636656888303e-05
GC_10_400 b_10 NI_10 NS_400 0 -1.8930879285145930e-04
GC_10_401 b_10 NI_10 NS_401 0 -4.8544283167664126e-06
GC_10_402 b_10 NI_10 NS_402 0 -5.7048652146901790e-06
GC_10_403 b_10 NI_10 NS_403 0 -2.0432777140302368e-06
GC_10_404 b_10 NI_10 NS_404 0 1.3068856560829426e-05
GC_10_405 b_10 NI_10 NS_405 0 2.4719793390214458e-04
GC_10_406 b_10 NI_10 NS_406 0 -1.3516403589174743e-04
GC_10_407 b_10 NI_10 NS_407 0 -3.0989886099481182e-05
GC_10_408 b_10 NI_10 NS_408 0 4.6298398693814924e-05
GD_10_1 b_10 NI_10 NA_1 0 -3.9608797226965298e-03
GD_10_2 b_10 NI_10 NA_2 0 -1.5923232891671495e-03
GD_10_3 b_10 NI_10 NA_3 0 -8.9344813522449166e-03
GD_10_4 b_10 NI_10 NA_4 0 -3.4066763589321999e-03
GD_10_5 b_10 NI_10 NA_5 0 -7.8366524273498824e-03
GD_10_6 b_10 NI_10 NA_6 0 1.6658818469890895e-03
GD_10_7 b_10 NI_10 NA_7 0 -9.6183972420804727e-03
GD_10_8 b_10 NI_10 NA_8 0 3.1638889255645951e-03
GD_10_9 b_10 NI_10 NA_9 0 -3.6009240211638698e-02
GD_10_10 b_10 NI_10 NA_10 0 -2.5820833543326255e-01
GD_10_11 b_10 NI_10 NA_11 0 -1.1910516112496359e-02
GD_10_12 b_10 NI_10 NA_12 0 7.1021985925394668e-03
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 6.5904971742592180e-03
GC_11_2 b_11 NI_11 NS_2 0 -2.5708654893186010e-04
GC_11_3 b_11 NI_11 NS_3 0 6.0981618186841058e-07
GC_11_4 b_11 NI_11 NS_4 0 -6.1638260617559366e-10
GC_11_5 b_11 NI_11 NS_5 0 1.5645486830453104e-03
GC_11_6 b_11 NI_11 NS_6 0 2.0017579519746522e-03
GC_11_7 b_11 NI_11 NS_7 0 1.8705673153532863e-03
GC_11_8 b_11 NI_11 NS_8 0 -6.5671384922311453e-04
GC_11_9 b_11 NI_11 NS_9 0 -7.8873518083643433e-03
GC_11_10 b_11 NI_11 NS_10 0 -7.2195768597574058e-04
GC_11_11 b_11 NI_11 NS_11 0 1.8083927322584421e-03
GC_11_12 b_11 NI_11 NS_12 0 2.8496919132865585e-03
GC_11_13 b_11 NI_11 NS_13 0 1.2293839369298914e-05
GC_11_14 b_11 NI_11 NS_14 0 -4.0951764691715024e-06
GC_11_15 b_11 NI_11 NS_15 0 1.0123920071657480e-06
GC_11_16 b_11 NI_11 NS_16 0 -3.0941636451086744e-06
GC_11_17 b_11 NI_11 NS_17 0 1.5883069884276292e-04
GC_11_18 b_11 NI_11 NS_18 0 -4.1862824866728754e-05
GC_11_19 b_11 NI_11 NS_19 0 -3.5225833722975277e-06
GC_11_20 b_11 NI_11 NS_20 0 -2.4785541164721773e-05
GC_11_21 b_11 NI_11 NS_21 0 -2.9916783253732242e-04
GC_11_22 b_11 NI_11 NS_22 0 -1.5012626899696225e-05
GC_11_23 b_11 NI_11 NS_23 0 -1.3306432788461077e-06
GC_11_24 b_11 NI_11 NS_24 0 2.2026966864196431e-06
GC_11_25 b_11 NI_11 NS_25 0 -1.7548038587253411e-04
GC_11_26 b_11 NI_11 NS_26 0 4.5531564790149474e-04
GC_11_27 b_11 NI_11 NS_27 0 -1.5540275149495429e-05
GC_11_28 b_11 NI_11 NS_28 0 2.7587095613996364e-05
GC_11_29 b_11 NI_11 NS_29 0 9.3391634303932588e-06
GC_11_30 b_11 NI_11 NS_30 0 -3.1663591433936329e-05
GC_11_31 b_11 NI_11 NS_31 0 6.5652987697573735e-04
GC_11_32 b_11 NI_11 NS_32 0 2.9008193747401563e-05
GC_11_33 b_11 NI_11 NS_33 0 3.5006002612726904e-06
GC_11_34 b_11 NI_11 NS_34 0 7.0858341223378549e-07
GC_11_35 b_11 NI_11 NS_35 0 7.0746105818804365e-03
GC_11_36 b_11 NI_11 NS_36 0 -4.6534114599575214e-04
GC_11_37 b_11 NI_11 NS_37 0 7.9559940484940433e-07
GC_11_38 b_11 NI_11 NS_38 0 2.7002132704761320e-10
GC_11_39 b_11 NI_11 NS_39 0 5.8202986621402235e-04
GC_11_40 b_11 NI_11 NS_40 0 1.6089618682722238e-03
GC_11_41 b_11 NI_11 NS_41 0 1.4710534523524805e-03
GC_11_42 b_11 NI_11 NS_42 0 -1.3561543085244549e-03
GC_11_43 b_11 NI_11 NS_43 0 -6.8784178760176173e-03
GC_11_44 b_11 NI_11 NS_44 0 6.8762023651887751e-04
GC_11_45 b_11 NI_11 NS_45 0 1.7513870352558717e-03
GC_11_46 b_11 NI_11 NS_46 0 2.1300727286511141e-03
GC_11_47 b_11 NI_11 NS_47 0 -1.2009232082002195e-06
GC_11_48 b_11 NI_11 NS_48 0 1.2906686835087843e-05
GC_11_49 b_11 NI_11 NS_49 0 3.9210508218762630e-06
GC_11_50 b_11 NI_11 NS_50 0 -1.6465800029986685e-05
GC_11_51 b_11 NI_11 NS_51 0 2.1124397652342756e-04
GC_11_52 b_11 NI_11 NS_52 0 1.5297127814358904e-04
GC_11_53 b_11 NI_11 NS_53 0 -2.4085320669994810e-05
GC_11_54 b_11 NI_11 NS_54 0 1.7724139081842514e-05
GC_11_55 b_11 NI_11 NS_55 0 -3.2648902583783931e-04
GC_11_56 b_11 NI_11 NS_56 0 -1.6305721302213347e-04
GC_11_57 b_11 NI_11 NS_57 0 1.3021069813360914e-07
GC_11_58 b_11 NI_11 NS_58 0 -3.6100417652829220e-07
GC_11_59 b_11 NI_11 NS_59 0 5.9196555678334759e-06
GC_11_60 b_11 NI_11 NS_60 0 3.7180673820558599e-04
GC_11_61 b_11 NI_11 NS_61 0 2.0490350413728704e-06
GC_11_62 b_11 NI_11 NS_62 0 -2.2602763477617131e-06
GC_11_63 b_11 NI_11 NS_63 0 -7.6497676581617920e-06
GC_11_64 b_11 NI_11 NS_64 0 3.1776634880725590e-05
GC_11_65 b_11 NI_11 NS_65 0 4.8282708954547441e-04
GC_11_66 b_11 NI_11 NS_66 0 -1.4040043120083711e-04
GC_11_67 b_11 NI_11 NS_67 0 -9.6615549012573673e-06
GC_11_68 b_11 NI_11 NS_68 0 -1.6431034758061317e-05
GC_11_69 b_11 NI_11 NS_69 0 4.7652830814229755e-03
GC_11_70 b_11 NI_11 NS_70 0 -3.6921529843050613e-05
GC_11_71 b_11 NI_11 NS_71 0 2.5169131650066477e-07
GC_11_72 b_11 NI_11 NS_72 0 -8.9160760708988326e-10
GC_11_73 b_11 NI_11 NS_73 0 1.7124161087228513e-03
GC_11_74 b_11 NI_11 NS_74 0 1.5475804069780682e-03
GC_11_75 b_11 NI_11 NS_75 0 7.4430420975781203e-04
GC_11_76 b_11 NI_11 NS_76 0 -1.6023165108241982e-04
GC_11_77 b_11 NI_11 NS_77 0 -5.5314504006866412e-03
GC_11_78 b_11 NI_11 NS_78 0 -4.4655616227984399e-04
GC_11_79 b_11 NI_11 NS_79 0 1.6138149360579385e-03
GC_11_80 b_11 NI_11 NS_80 0 2.2938448178103014e-03
GC_11_81 b_11 NI_11 NS_81 0 1.0323274818931940e-05
GC_11_82 b_11 NI_11 NS_82 0 -3.6656011193678495e-06
GC_11_83 b_11 NI_11 NS_83 0 1.0985199168819868e-06
GC_11_84 b_11 NI_11 NS_84 0 -3.3395124958954973e-06
GC_11_85 b_11 NI_11 NS_85 0 1.6102097134514830e-04
GC_11_86 b_11 NI_11 NS_86 0 -4.5218442348266320e-05
GC_11_87 b_11 NI_11 NS_87 0 -3.1585125545714931e-06
GC_11_88 b_11 NI_11 NS_88 0 -1.6482095671275182e-05
GC_11_89 b_11 NI_11 NS_89 0 -2.0490222586878616e-04
GC_11_90 b_11 NI_11 NS_90 0 -4.3169639021589365e-06
GC_11_91 b_11 NI_11 NS_91 0 4.0857885049895718e-07
GC_11_92 b_11 NI_11 NS_92 0 4.2656654597150523e-06
GC_11_93 b_11 NI_11 NS_93 0 -3.9050386395179509e-04
GC_11_94 b_11 NI_11 NS_94 0 4.0661316947696036e-04
GC_11_95 b_11 NI_11 NS_95 0 1.9145331847226602e-05
GC_11_96 b_11 NI_11 NS_96 0 -1.9537011475473159e-06
GC_11_97 b_11 NI_11 NS_97 0 4.3210311732329511e-06
GC_11_98 b_11 NI_11 NS_98 0 -2.1205016069143586e-05
GC_11_99 b_11 NI_11 NS_99 0 5.8047115429727889e-04
GC_11_100 b_11 NI_11 NS_100 0 2.7934966805040774e-05
GC_11_101 b_11 NI_11 NS_101 0 2.9211800834105284e-06
GC_11_102 b_11 NI_11 NS_102 0 2.0872312884100151e-07
GC_11_103 b_11 NI_11 NS_103 0 3.9364551925647768e-03
GC_11_104 b_11 NI_11 NS_104 0 -2.9699663310858558e-04
GC_11_105 b_11 NI_11 NS_105 0 2.1277166764066754e-08
GC_11_106 b_11 NI_11 NS_106 0 1.0071886551888427e-09
GC_11_107 b_11 NI_11 NS_107 0 -6.0188150510479476e-04
GC_11_108 b_11 NI_11 NS_108 0 6.3457881057924642e-04
GC_11_109 b_11 NI_11 NS_109 0 5.9730461051647884e-04
GC_11_110 b_11 NI_11 NS_110 0 -1.8891702578264371e-05
GC_11_111 b_11 NI_11 NS_111 0 -2.6175296706305497e-03
GC_11_112 b_11 NI_11 NS_112 0 1.4294197263675279e-04
GC_11_113 b_11 NI_11 NS_113 0 1.0967122916278288e-03
GC_11_114 b_11 NI_11 NS_114 0 3.2349916497159177e-04
GC_11_115 b_11 NI_11 NS_115 0 -1.1429475455863845e-06
GC_11_116 b_11 NI_11 NS_116 0 1.0601000513358398e-05
GC_11_117 b_11 NI_11 NS_117 0 4.6084306948697177e-06
GC_11_118 b_11 NI_11 NS_118 0 -1.7489066520044106e-05
GC_11_119 b_11 NI_11 NS_119 0 2.1443605039431403e-04
GC_11_120 b_11 NI_11 NS_120 0 1.5572073092174309e-04
GC_11_121 b_11 NI_11 NS_121 0 -1.2547827020403254e-05
GC_11_122 b_11 NI_11 NS_122 0 1.6348273337184345e-05
GC_11_123 b_11 NI_11 NS_123 0 -2.4668937816388451e-04
GC_11_124 b_11 NI_11 NS_124 0 -1.0716621240105062e-04
GC_11_125 b_11 NI_11 NS_125 0 2.8564354845742988e-06
GC_11_126 b_11 NI_11 NS_126 0 -1.6180605501619011e-07
GC_11_127 b_11 NI_11 NS_127 0 -1.5020941112582089e-04
GC_11_128 b_11 NI_11 NS_128 0 3.2792650767531371e-04
GC_11_129 b_11 NI_11 NS_129 0 3.9939787971405451e-06
GC_11_130 b_11 NI_11 NS_130 0 1.2466440144833831e-05
GC_11_131 b_11 NI_11 NS_131 0 -4.2364877186023545e-06
GC_11_132 b_11 NI_11 NS_132 0 1.8937067454884047e-05
GC_11_133 b_11 NI_11 NS_133 0 4.2604238851028342e-04
GC_11_134 b_11 NI_11 NS_134 0 -1.5478300459843185e-04
GC_11_135 b_11 NI_11 NS_135 0 -9.7361844389681194e-06
GC_11_136 b_11 NI_11 NS_136 0 -1.6103565636454414e-05
GC_11_137 b_11 NI_11 NS_137 0 -2.8622044608859493e-03
GC_11_138 b_11 NI_11 NS_138 0 5.8851188567024158e-04
GC_11_139 b_11 NI_11 NS_139 0 -1.0298726390181808e-06
GC_11_140 b_11 NI_11 NS_140 0 -1.2010063910683944e-09
GC_11_141 b_11 NI_11 NS_141 0 1.5323549843585045e-03
GC_11_142 b_11 NI_11 NS_142 0 -4.5396929986005273e-04
GC_11_143 b_11 NI_11 NS_143 0 -1.0401353605748234e-03
GC_11_144 b_11 NI_11 NS_144 0 5.4146745787973180e-05
GC_11_145 b_11 NI_11 NS_145 0 3.3884510805422437e-04
GC_11_146 b_11 NI_11 NS_146 0 1.1008711520298349e-03
GC_11_147 b_11 NI_11 NS_147 0 6.7206486523692540e-04
GC_11_148 b_11 NI_11 NS_148 0 -1.1552602301880997e-04
GC_11_149 b_11 NI_11 NS_149 0 -9.2189463411264345e-07
GC_11_150 b_11 NI_11 NS_150 0 3.4633231089203190e-06
GC_11_151 b_11 NI_11 NS_151 0 1.4049618668629127e-06
GC_11_152 b_11 NI_11 NS_152 0 -3.6180745173334891e-06
GC_11_153 b_11 NI_11 NS_153 0 1.5695188764615104e-04
GC_11_154 b_11 NI_11 NS_154 0 -4.4913647878615782e-05
GC_11_155 b_11 NI_11 NS_155 0 3.7329361723161207e-07
GC_11_156 b_11 NI_11 NS_156 0 -4.8331645594830735e-06
GC_11_157 b_11 NI_11 NS_157 0 -6.8575192157057857e-05
GC_11_158 b_11 NI_11 NS_158 0 7.6708143858736326e-06
GC_11_159 b_11 NI_11 NS_159 0 6.6535559048027262e-07
GC_11_160 b_11 NI_11 NS_160 0 1.7916857623663641e-06
GC_11_161 b_11 NI_11 NS_161 0 -6.1779647875208387e-04
GC_11_162 b_11 NI_11 NS_162 0 2.1697441979672745e-04
GC_11_163 b_11 NI_11 NS_163 0 4.0716318355684318e-05
GC_11_164 b_11 NI_11 NS_164 0 -2.3436320996607686e-05
GC_11_165 b_11 NI_11 NS_165 0 4.5511189338773960e-06
GC_11_166 b_11 NI_11 NS_166 0 -6.9727957931297484e-06
GC_11_167 b_11 NI_11 NS_167 0 5.9902869043770791e-04
GC_11_168 b_11 NI_11 NS_168 0 -4.6277914776284931e-05
GC_11_169 b_11 NI_11 NS_169 0 2.9055004477589648e-06
GC_11_170 b_11 NI_11 NS_170 0 6.8394009621211600e-07
GC_11_171 b_11 NI_11 NS_171 0 5.7403212039234359e-03
GC_11_172 b_11 NI_11 NS_172 0 -4.9676224184750620e-04
GC_11_173 b_11 NI_11 NS_173 0 -3.0285971987339069e-07
GC_11_174 b_11 NI_11 NS_174 0 2.0709799517999618e-09
GC_11_175 b_11 NI_11 NS_175 0 -2.1362638642202516e-03
GC_11_176 b_11 NI_11 NS_176 0 2.0558687567760062e-03
GC_11_177 b_11 NI_11 NS_177 0 -5.6368257837554562e-04
GC_11_178 b_11 NI_11 NS_178 0 1.2106229108160645e-03
GC_11_179 b_11 NI_11 NS_179 0 2.1059573345629280e-03
GC_11_180 b_11 NI_11 NS_180 0 -2.0079026854109235e-03
GC_11_181 b_11 NI_11 NS_181 0 -1.9806799138105129e-03
GC_11_182 b_11 NI_11 NS_182 0 -5.1433192851249002e-04
GC_11_183 b_11 NI_11 NS_183 0 7.1068816970838688e-07
GC_11_184 b_11 NI_11 NS_184 0 2.3213113989950085e-06
GC_11_185 b_11 NI_11 NS_185 0 3.9708329136103656e-06
GC_11_186 b_11 NI_11 NS_186 0 -1.6980381064575673e-05
GC_11_187 b_11 NI_11 NS_187 0 2.1944531383214974e-04
GC_11_188 b_11 NI_11 NS_188 0 1.4707433161083487e-04
GC_11_189 b_11 NI_11 NS_189 0 -7.2273881048286486e-06
GC_11_190 b_11 NI_11 NS_190 0 2.8266319700110507e-06
GC_11_191 b_11 NI_11 NS_191 0 -6.6659895958017901e-05
GC_11_192 b_11 NI_11 NS_192 0 -3.4821920500270080e-05
GC_11_193 b_11 NI_11 NS_193 0 2.5397973616791483e-06
GC_11_194 b_11 NI_11 NS_194 0 -6.3352157634170958e-08
GC_11_195 b_11 NI_11 NS_195 0 -3.9623932305397246e-04
GC_11_196 b_11 NI_11 NS_196 0 2.1414936205330684e-04
GC_11_197 b_11 NI_11 NS_197 0 3.5141898799756159e-06
GC_11_198 b_11 NI_11 NS_198 0 2.5696910121500275e-05
GC_11_199 b_11 NI_11 NS_199 0 -3.9930421683831875e-07
GC_11_200 b_11 NI_11 NS_200 0 1.3819879835150695e-05
GC_11_201 b_11 NI_11 NS_201 0 4.0151954294154955e-04
GC_11_202 b_11 NI_11 NS_202 0 -2.3371861775782135e-04
GC_11_203 b_11 NI_11 NS_203 0 -1.0493955086723401e-05
GC_11_204 b_11 NI_11 NS_204 0 -1.7880258885812424e-05
GC_11_205 b_11 NI_11 NS_205 0 -1.2023412524613657e-02
GC_11_206 b_11 NI_11 NS_206 0 1.5260909726964860e-03
GC_11_207 b_11 NI_11 NS_207 0 -3.1103879496602479e-06
GC_11_208 b_11 NI_11 NS_208 0 -2.7311491549456816e-09
GC_11_209 b_11 NI_11 NS_209 0 2.7363500911700613e-03
GC_11_210 b_11 NI_11 NS_210 0 -2.1648095732052335e-03
GC_11_211 b_11 NI_11 NS_211 0 -7.8970034570543580e-04
GC_11_212 b_11 NI_11 NS_212 0 8.0138119715785275e-04
GC_11_213 b_11 NI_11 NS_213 0 2.4482977022492768e-03
GC_11_214 b_11 NI_11 NS_214 0 -5.3759162611108433e-04
GC_11_215 b_11 NI_11 NS_215 0 -4.7797753794446699e-05
GC_11_216 b_11 NI_11 NS_216 0 -5.3654849055087214e-04
GC_11_217 b_11 NI_11 NS_217 0 -1.1099915592061889e-06
GC_11_218 b_11 NI_11 NS_218 0 -2.0123160353280910e-06
GC_11_219 b_11 NI_11 NS_219 0 1.3370505208517884e-06
GC_11_220 b_11 NI_11 NS_220 0 -3.8185054380926480e-06
GC_11_221 b_11 NI_11 NS_221 0 1.5648781969091562e-04
GC_11_222 b_11 NI_11 NS_222 0 -4.4825145726379293e-05
GC_11_223 b_11 NI_11 NS_223 0 1.5539122479999530e-06
GC_11_224 b_11 NI_11 NS_224 0 8.5738731593666525e-06
GC_11_225 b_11 NI_11 NS_225 0 8.4905606969111773e-05
GC_11_226 b_11 NI_11 NS_226 0 6.1729117055171494e-06
GC_11_227 b_11 NI_11 NS_227 0 1.5450380397723871e-07
GC_11_228 b_11 NI_11 NS_228 0 8.5063051690902433e-07
GC_11_229 b_11 NI_11 NS_229 0 -2.4355784047680183e-04
GC_11_230 b_11 NI_11 NS_230 0 -8.8488600017971354e-05
GC_11_231 b_11 NI_11 NS_231 0 4.1292908549286610e-05
GC_11_232 b_11 NI_11 NS_232 0 -3.3063221425079361e-05
GC_11_233 b_11 NI_11 NS_233 0 -5.5267407429947569e-06
GC_11_234 b_11 NI_11 NS_234 0 9.4374261515540724e-06
GC_11_235 b_11 NI_11 NS_235 0 5.3645395308599066e-04
GC_11_236 b_11 NI_11 NS_236 0 1.4628619089776525e-05
GC_11_237 b_11 NI_11 NS_237 0 1.9965241991125924e-06
GC_11_238 b_11 NI_11 NS_238 0 -6.6339729036827784e-07
GC_11_239 b_11 NI_11 NS_239 0 1.0740932060516932e-02
GC_11_240 b_11 NI_11 NS_240 0 -9.6976288621372555e-04
GC_11_241 b_11 NI_11 NS_241 0 -6.2798410600020054e-07
GC_11_242 b_11 NI_11 NS_242 0 4.1450453344662773e-09
GC_11_243 b_11 NI_11 NS_243 0 -4.8261873414535746e-03
GC_11_244 b_11 NI_11 NS_244 0 4.6840574959655830e-03
GC_11_245 b_11 NI_11 NS_245 0 -1.9243484202241447e-04
GC_11_246 b_11 NI_11 NS_246 0 1.3745685368306241e-03
GC_11_247 b_11 NI_11 NS_247 0 2.0442181541639325e-03
GC_11_248 b_11 NI_11 NS_248 0 -4.4549766255966364e-03
GC_11_249 b_11 NI_11 NS_249 0 -4.0090260290626513e-03
GC_11_250 b_11 NI_11 NS_250 0 -6.7731249001654580e-04
GC_11_251 b_11 NI_11 NS_251 0 -1.6709039471237483e-06
GC_11_252 b_11 NI_11 NS_252 0 6.2749989653182146e-07
GC_11_253 b_11 NI_11 NS_253 0 4.6629318501588797e-06
GC_11_254 b_11 NI_11 NS_254 0 -1.7454700038141407e-05
GC_11_255 b_11 NI_11 NS_255 0 2.1287305228318986e-04
GC_11_256 b_11 NI_11 NS_256 0 1.5128574594756072e-04
GC_11_257 b_11 NI_11 NS_257 0 9.3468071513204006e-06
GC_11_258 b_11 NI_11 NS_258 0 -1.5100342071812882e-06
GC_11_259 b_11 NI_11 NS_259 0 7.7831611439755266e-05
GC_11_260 b_11 NI_11 NS_260 0 4.4691209663383202e-05
GC_11_261 b_11 NI_11 NS_261 0 1.4455564211186945e-06
GC_11_262 b_11 NI_11 NS_262 0 -2.6675626652074775e-07
GC_11_263 b_11 NI_11 NS_263 0 -2.2726109504053179e-04
GC_11_264 b_11 NI_11 NS_264 0 -5.7066907307492150e-05
GC_11_265 b_11 NI_11 NS_265 0 4.9703305959138357e-06
GC_11_266 b_11 NI_11 NS_266 0 1.8016234396344570e-05
GC_11_267 b_11 NI_11 NS_267 0 2.6720323390104067e-06
GC_11_268 b_11 NI_11 NS_268 0 -1.1310599518461368e-05
GC_11_269 b_11 NI_11 NS_269 0 3.7933821088176155e-04
GC_11_270 b_11 NI_11 NS_270 0 -1.7766598710550568e-04
GC_11_271 b_11 NI_11 NS_271 0 -1.1701705813337291e-05
GC_11_272 b_11 NI_11 NS_272 0 -1.8821136104863797e-05
GC_11_273 b_11 NI_11 NS_273 0 -3.3835127070151613e-02
GC_11_274 b_11 NI_11 NS_274 0 3.2816952524806638e-03
GC_11_275 b_11 NI_11 NS_275 0 -1.5878931873327682e-05
GC_11_276 b_11 NI_11 NS_276 0 -5.7011516637311961e-09
GC_11_277 b_11 NI_11 NS_277 0 1.0193798057749618e-02
GC_11_278 b_11 NI_11 NS_278 0 -1.0005632062877839e-02
GC_11_279 b_11 NI_11 NS_279 0 -1.8931606119316250e-03
GC_11_280 b_11 NI_11 NS_280 0 2.3331662916374504e-04
GC_11_281 b_11 NI_11 NS_281 0 5.6460487629264589e-03
GC_11_282 b_11 NI_11 NS_282 0 3.4668890174292828e-03
GC_11_283 b_11 NI_11 NS_283 0 1.8126030643520726e-03
GC_11_284 b_11 NI_11 NS_284 0 -6.0940695179018589e-04
GC_11_285 b_11 NI_11 NS_285 0 -1.1153608351667405e-05
GC_11_286 b_11 NI_11 NS_286 0 2.9591228839482261e-06
GC_11_287 b_11 NI_11 NS_287 0 2.0985253836974496e-06
GC_11_288 b_11 NI_11 NS_288 0 -3.7144259370389897e-06
GC_11_289 b_11 NI_11 NS_289 0 1.5365448238209486e-04
GC_11_290 b_11 NI_11 NS_290 0 -4.4022668050939518e-05
GC_11_291 b_11 NI_11 NS_291 0 5.6750764129017924e-06
GC_11_292 b_11 NI_11 NS_292 0 1.9312490393457342e-05
GC_11_293 b_11 NI_11 NS_293 0 2.1080976723294480e-04
GC_11_294 b_11 NI_11 NS_294 0 1.6100580521359033e-05
GC_11_295 b_11 NI_11 NS_295 0 1.2459259441288702e-06
GC_11_296 b_11 NI_11 NS_296 0 2.9947500544197611e-06
GC_11_297 b_11 NI_11 NS_297 0 1.7957942733314377e-04
GC_11_298 b_11 NI_11 NS_298 0 -3.8393613595189192e-04
GC_11_299 b_11 NI_11 NS_299 0 1.2979314814191741e-05
GC_11_300 b_11 NI_11 NS_300 0 -1.5583491129384082e-05
GC_11_301 b_11 NI_11 NS_301 0 -4.3320671731046821e-06
GC_11_302 b_11 NI_11 NS_302 0 2.3111144697108292e-05
GC_11_303 b_11 NI_11 NS_303 0 4.2270787522050786e-04
GC_11_304 b_11 NI_11 NS_304 0 4.0240050294477466e-05
GC_11_305 b_11 NI_11 NS_305 0 2.6664246026282233e-06
GC_11_306 b_11 NI_11 NS_306 0 -2.1740416778806806e-06
GC_11_307 b_11 NI_11 NS_307 0 3.2850475390866787e-02
GC_11_308 b_11 NI_11 NS_308 0 -3.5239944320197849e-03
GC_11_309 b_11 NI_11 NS_309 0 -1.9759978112809740e-06
GC_11_310 b_11 NI_11 NS_310 0 9.6963504096010097e-09
GC_11_311 b_11 NI_11 NS_311 0 -1.5289656551483845e-02
GC_11_312 b_11 NI_11 NS_312 0 1.2292224700810895e-02
GC_11_313 b_11 NI_11 NS_313 0 5.9227679670577924e-05
GC_11_314 b_11 NI_11 NS_314 0 1.1227030856325911e-03
GC_11_315 b_11 NI_11 NS_315 0 3.7337145323375802e-03
GC_11_316 b_11 NI_11 NS_316 0 -9.1134184512235220e-03
GC_11_317 b_11 NI_11 NS_317 0 -8.6972426872503460e-03
GC_11_318 b_11 NI_11 NS_318 0 -1.9939969921796644e-03
GC_11_319 b_11 NI_11 NS_319 0 1.1834780476771154e-07
GC_11_320 b_11 NI_11 NS_320 0 -8.3061519722165440e-06
GC_11_321 b_11 NI_11 NS_321 0 4.0706510436770074e-06
GC_11_322 b_11 NI_11 NS_322 0 -1.7106739543639383e-05
GC_11_323 b_11 NI_11 NS_323 0 2.1829470173642077e-04
GC_11_324 b_11 NI_11 NS_324 0 1.5154613525815105e-04
GC_11_325 b_11 NI_11 NS_325 0 1.5248662223839422e-05
GC_11_326 b_11 NI_11 NS_326 0 -1.5589036163283982e-05
GC_11_327 b_11 NI_11 NS_327 0 2.4540912514571918e-04
GC_11_328 b_11 NI_11 NS_328 0 1.1630279609413247e-04
GC_11_329 b_11 NI_11 NS_329 0 6.7159703415845616e-06
GC_11_330 b_11 NI_11 NS_330 0 1.0255440187206238e-06
GC_11_331 b_11 NI_11 NS_331 0 -1.3236042633016116e-04
GC_11_332 b_11 NI_11 NS_332 0 -3.9484275098406059e-04
GC_11_333 b_11 NI_11 NS_333 0 -3.3181442890401266e-06
GC_11_334 b_11 NI_11 NS_334 0 4.8895776114243075e-06
GC_11_335 b_11 NI_11 NS_335 0 3.8158365488448764e-06
GC_11_336 b_11 NI_11 NS_336 0 -1.5708438936134302e-05
GC_11_337 b_11 NI_11 NS_337 0 2.5429178663090237e-04
GC_11_338 b_11 NI_11 NS_338 0 -2.1880110305506347e-04
GC_11_339 b_11 NI_11 NS_339 0 -8.2384009046678529e-06
GC_11_340 b_11 NI_11 NS_340 0 -1.6537645220364260e-05
GC_11_341 b_11 NI_11 NS_341 0 -2.3531005745253064e-01
GC_11_342 b_11 NI_11 NS_342 0 5.7440312415981673e-02
GC_11_343 b_11 NI_11 NS_343 0 3.4376134557584744e-05
GC_11_344 b_11 NI_11 NS_344 0 -5.6713874126097491e-08
GC_11_345 b_11 NI_11 NS_345 0 8.4103777509869526e-02
GC_11_346 b_11 NI_11 NS_346 0 2.2117925755600807e-03
GC_11_347 b_11 NI_11 NS_347 0 1.7692062312993823e-04
GC_11_348 b_11 NI_11 NS_348 0 1.9540138399147806e-03
GC_11_349 b_11 NI_11 NS_349 0 7.0788049812392619e-03
GC_11_350 b_11 NI_11 NS_350 0 5.4727467570125973e-03
GC_11_351 b_11 NI_11 NS_351 0 -6.9549309008340096e-03
GC_11_352 b_11 NI_11 NS_352 0 2.3420266372967376e-03
GC_11_353 b_11 NI_11 NS_353 0 -1.2805167854405243e-05
GC_11_354 b_11 NI_11 NS_354 0 5.7609506984891091e-06
GC_11_355 b_11 NI_11 NS_355 0 2.7150205528544257e-06
GC_11_356 b_11 NI_11 NS_356 0 -3.4746330676413788e-06
GC_11_357 b_11 NI_11 NS_357 0 1.3913562285804585e-04
GC_11_358 b_11 NI_11 NS_358 0 -4.2204037778942299e-05
GC_11_359 b_11 NI_11 NS_359 0 4.6147042592834133e-06
GC_11_360 b_11 NI_11 NS_360 0 2.6100950783461522e-05
GC_11_361 b_11 NI_11 NS_361 0 2.9878849416394872e-04
GC_11_362 b_11 NI_11 NS_362 0 3.0709503922879302e-05
GC_11_363 b_11 NI_11 NS_363 0 2.3839696790709053e-06
GC_11_364 b_11 NI_11 NS_364 0 -7.5475175179684969e-08
GC_11_365 b_11 NI_11 NS_365 0 6.7694978781016220e-04
GC_11_366 b_11 NI_11 NS_366 0 -6.8505704035459389e-04
GC_11_367 b_11 NI_11 NS_367 0 -2.0963496218396894e-05
GC_11_368 b_11 NI_11 NS_368 0 4.6281569141492279e-06
GC_11_369 b_11 NI_11 NS_369 0 -1.1647776640134387e-05
GC_11_370 b_11 NI_11 NS_370 0 3.4055353255788897e-05
GC_11_371 b_11 NI_11 NS_371 0 3.3517041446496666e-04
GC_11_372 b_11 NI_11 NS_372 0 -1.8977860195205547e-05
GC_11_373 b_11 NI_11 NS_373 0 5.2506341605314484e-06
GC_11_374 b_11 NI_11 NS_374 0 -2.5610915676791306e-06
GC_11_375 b_11 NI_11 NS_375 0 3.2724706258644029e-02
GC_11_376 b_11 NI_11 NS_376 0 3.2736866451345700e-02
GC_11_377 b_11 NI_11 NS_377 0 1.6523826391137434e-04
GC_11_378 b_11 NI_11 NS_378 0 2.5349383293241769e-07
GC_11_379 b_11 NI_11 NS_379 0 -6.0934733057427908e-02
GC_11_380 b_11 NI_11 NS_380 0 -1.7132987174366700e-02
GC_11_381 b_11 NI_11 NS_381 0 -1.7899288550700544e-03
GC_11_382 b_11 NI_11 NS_382 0 4.8602801592216140e-03
GC_11_383 b_11 NI_11 NS_383 0 1.2185135287179637e-02
GC_11_384 b_11 NI_11 NS_384 0 1.6811852628881130e-02
GC_11_385 b_11 NI_11 NS_385 0 7.1137388361608000e-03
GC_11_386 b_11 NI_11 NS_386 0 8.1970615233297985e-05
GC_11_387 b_11 NI_11 NS_387 0 -5.2197828031974734e-07
GC_11_388 b_11 NI_11 NS_388 0 -1.3005900105788046e-05
GC_11_389 b_11 NI_11 NS_389 0 2.7206797921878804e-06
GC_11_390 b_11 NI_11 NS_390 0 -1.7277000711605512e-05
GC_11_391 b_11 NI_11 NS_391 0 2.2114793525987856e-04
GC_11_392 b_11 NI_11 NS_392 0 1.5871324659615267e-04
GC_11_393 b_11 NI_11 NS_393 0 2.4015035143101963e-05
GC_11_394 b_11 NI_11 NS_394 0 -1.4432352217034474e-05
GC_11_395 b_11 NI_11 NS_395 0 3.3597212254563231e-04
GC_11_396 b_11 NI_11 NS_396 0 1.4568791189526007e-04
GC_11_397 b_11 NI_11 NS_397 0 -1.2531814801653733e-06
GC_11_398 b_11 NI_11 NS_398 0 -9.3013107855436504e-07
GC_11_399 b_11 NI_11 NS_399 0 3.7106916885653056e-04
GC_11_400 b_11 NI_11 NS_400 0 -6.4126372716687586e-04
GC_11_401 b_11 NI_11 NS_401 0 -3.8412966732137480e-06
GC_11_402 b_11 NI_11 NS_402 0 -2.4749017461650801e-05
GC_11_403 b_11 NI_11 NS_403 0 3.2526383287192302e-06
GC_11_404 b_11 NI_11 NS_404 0 -3.4178724922346622e-05
GC_11_405 b_11 NI_11 NS_405 0 4.2186431390820399e-04
GC_11_406 b_11 NI_11 NS_406 0 -5.1895124895972440e-05
GC_11_407 b_11 NI_11 NS_407 0 -1.1686949289103079e-05
GC_11_408 b_11 NI_11 NS_408 0 -1.7937695238829897e-05
GD_11_1 b_11 NI_11 NA_1 0 -5.1252094069501901e-03
GD_11_2 b_11 NI_11 NA_2 0 -4.8175277143955525e-03
GD_11_3 b_11 NI_11 NA_3 0 -4.2636986075969968e-03
GD_11_4 b_11 NI_11 NA_4 0 -3.4892434087148917e-03
GD_11_5 b_11 NI_11 NA_5 0 1.2181903169224703e-03
GD_11_6 b_11 NI_11 NA_6 0 -4.4613088143037978e-03
GD_11_7 b_11 NI_11 NA_7 0 6.8515421669424386e-03
GD_11_8 b_11 NI_11 NA_8 0 -3.9371638264554384e-03
GD_11_9 b_11 NI_11 NA_9 0 1.6093936552799858e-02
GD_11_10 b_11 NI_11 NA_10 0 -1.1910514918679158e-02
GD_11_11 b_11 NI_11 NA_11 0 1.0795451869903004e-01
GD_11_12 b_11 NI_11 NA_12 0 -3.5191575883040283e-02
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 7.0918497914602471e-03
GC_12_2 b_12 NI_12 NS_2 0 -4.6171629817053843e-04
GC_12_3 b_12 NI_12 NS_3 0 7.8399023967037056e-07
GC_12_4 b_12 NI_12 NS_4 0 2.7793517231239117e-10
GC_12_5 b_12 NI_12 NS_5 0 5.9929371947466353e-04
GC_12_6 b_12 NI_12 NS_6 0 1.5791892094341856e-03
GC_12_7 b_12 NI_12 NS_7 0 1.3769530191934712e-03
GC_12_8 b_12 NI_12 NS_8 0 -1.3596435477110879e-03
GC_12_9 b_12 NI_12 NS_9 0 -6.7299577014755816e-03
GC_12_10 b_12 NI_12 NS_10 0 8.7059485289296668e-04
GC_12_11 b_12 NI_12 NS_11 0 1.7678503908029207e-03
GC_12_12 b_12 NI_12 NS_12 0 2.0430373666466676e-03
GC_12_13 b_12 NI_12 NS_13 0 -2.0298651939313861e-06
GC_12_14 b_12 NI_12 NS_14 0 1.1883912769448550e-05
GC_12_15 b_12 NI_12 NS_15 0 4.7055760862836707e-06
GC_12_16 b_12 NI_12 NS_16 0 -1.7366820363344177e-05
GC_12_17 b_12 NI_12 NS_17 0 2.0850591213509532e-04
GC_12_18 b_12 NI_12 NS_18 0 1.5751373054571040e-04
GC_12_19 b_12 NI_12 NS_19 0 -2.2776422390340912e-05
GC_12_20 b_12 NI_12 NS_20 0 1.5281476060992603e-05
GC_12_21 b_12 NI_12 NS_21 0 -3.2850132382824209e-04
GC_12_22 b_12 NI_12 NS_22 0 -1.5665465045767377e-04
GC_12_23 b_12 NI_12 NS_23 0 3.0793834868926044e-07
GC_12_24 b_12 NI_12 NS_24 0 -2.2371736507970293e-07
GC_12_25 b_12 NI_12 NS_25 0 -5.0290843723953911e-06
GC_12_26 b_12 NI_12 NS_26 0 3.5547550321884713e-04
GC_12_27 b_12 NI_12 NS_27 0 5.4551211707487873e-06
GC_12_28 b_12 NI_12 NS_28 0 2.1525782159090576e-06
GC_12_29 b_12 NI_12 NS_29 0 -7.4406691866509952e-06
GC_12_30 b_12 NI_12 NS_30 0 2.9076698573710994e-05
GC_12_31 b_12 NI_12 NS_31 0 4.8737385208360315e-04
GC_12_32 b_12 NI_12 NS_32 0 -1.4037010353227191e-04
GC_12_33 b_12 NI_12 NS_33 0 -9.8137158137936701e-06
GC_12_34 b_12 NI_12 NS_34 0 -1.7335114430768381e-05
GC_12_35 b_12 NI_12 NS_35 0 2.4230028956626986e-03
GC_12_36 b_12 NI_12 NS_36 0 -9.8387394385423250e-05
GC_12_37 b_12 NI_12 NS_37 0 -4.3917260008279619e-07
GC_12_38 b_12 NI_12 NS_38 0 -2.3815598289238033e-10
GC_12_39 b_12 NI_12 NS_39 0 1.9634674238368064e-03
GC_12_40 b_12 NI_12 NS_40 0 -3.3509769770803769e-04
GC_12_41 b_12 NI_12 NS_41 0 5.4668619928719287e-04
GC_12_42 b_12 NI_12 NS_42 0 -1.2699747383749160e-03
GC_12_43 b_12 NI_12 NS_43 0 -4.6180391593397671e-03
GC_12_44 b_12 NI_12 NS_44 0 2.4918450674381639e-03
GC_12_45 b_12 NI_12 NS_45 0 2.2235333647192259e-03
GC_12_46 b_12 NI_12 NS_46 0 1.4004592264383613e-03
GC_12_47 b_12 NI_12 NS_47 0 -1.4840252846836711e-05
GC_12_48 b_12 NI_12 NS_48 0 -5.1143433184959633e-06
GC_12_49 b_12 NI_12 NS_49 0 7.9411390260710906e-06
GC_12_50 b_12 NI_12 NS_50 0 -8.5623186820538819e-05
GC_12_51 b_12 NI_12 NS_51 0 5.9387466143540643e-06
GC_12_52 b_12 NI_12 NS_52 0 4.2775704370299990e-04
GC_12_53 b_12 NI_12 NS_53 0 3.8912321862454498e-05
GC_12_54 b_12 NI_12 NS_54 0 2.2642833621339910e-05
GC_12_55 b_12 NI_12 NS_55 0 -3.2645315917656048e-04
GC_12_56 b_12 NI_12 NS_56 0 -3.0819342936092887e-04
GC_12_57 b_12 NI_12 NS_57 0 1.8762505659429799e-08
GC_12_58 b_12 NI_12 NS_58 0 1.7867139890528043e-07
GC_12_59 b_12 NI_12 NS_59 0 7.5346669631508439e-05
GC_12_60 b_12 NI_12 NS_60 0 2.4783109832974523e-04
GC_12_61 b_12 NI_12 NS_61 0 4.4739639551544536e-06
GC_12_62 b_12 NI_12 NS_62 0 1.0116694842117591e-05
GC_12_63 b_12 NI_12 NS_63 0 1.3524359338736486e-06
GC_12_64 b_12 NI_12 NS_64 0 -2.3185503376281683e-05
GC_12_65 b_12 NI_12 NS_65 0 3.3336077469771043e-04
GC_12_66 b_12 NI_12 NS_66 0 -2.1080813336662890e-04
GC_12_67 b_12 NI_12 NS_67 0 -3.2992078424257538e-05
GC_12_68 b_12 NI_12 NS_68 0 4.6785746304139202e-05
GC_12_69 b_12 NI_12 NS_69 0 5.6565104888912001e-03
GC_12_70 b_12 NI_12 NS_70 0 -4.4119117057139334e-04
GC_12_71 b_12 NI_12 NS_71 0 4.6096157655606291e-07
GC_12_72 b_12 NI_12 NS_72 0 8.8242390044361049e-10
GC_12_73 b_12 NI_12 NS_73 0 -5.8577913087898303e-04
GC_12_74 b_12 NI_12 NS_74 0 1.2278740208574656e-03
GC_12_75 b_12 NI_12 NS_75 0 5.9221013806723009e-04
GC_12_76 b_12 NI_12 NS_76 0 -6.7902228745398790e-05
GC_12_77 b_12 NI_12 NS_77 0 -2.9555051291182987e-03
GC_12_78 b_12 NI_12 NS_78 0 -1.1020655528962630e-04
GC_12_79 b_12 NI_12 NS_79 0 7.6426852890754864e-04
GC_12_80 b_12 NI_12 NS_80 0 6.6649185605493404e-04
GC_12_81 b_12 NI_12 NS_81 0 -2.4629469468153632e-06
GC_12_82 b_12 NI_12 NS_82 0 1.0671816327320843e-05
GC_12_83 b_12 NI_12 NS_83 0 4.8800840654196127e-06
GC_12_84 b_12 NI_12 NS_84 0 -1.7866073773009926e-05
GC_12_85 b_12 NI_12 NS_85 0 2.1554385567010970e-04
GC_12_86 b_12 NI_12 NS_86 0 1.5960848162302740e-04
GC_12_87 b_12 NI_12 NS_87 0 -1.4650885929117881e-05
GC_12_88 b_12 NI_12 NS_88 0 1.1245295656762322e-05
GC_12_89 b_12 NI_12 NS_89 0 -2.3255592555264308e-04
GC_12_90 b_12 NI_12 NS_90 0 -9.8410689871078193e-05
GC_12_91 b_12 NI_12 NS_91 0 2.5120254351309516e-06
GC_12_92 b_12 NI_12 NS_92 0 -5.6360477849433305e-07
GC_12_93 b_12 NI_12 NS_93 0 -1.5371760836781006e-04
GC_12_94 b_12 NI_12 NS_94 0 3.2102337311738229e-04
GC_12_95 b_12 NI_12 NS_95 0 -4.5645635694412994e-07
GC_12_96 b_12 NI_12 NS_96 0 1.2225113852424451e-05
GC_12_97 b_12 NI_12 NS_97 0 -1.5482956223918301e-06
GC_12_98 b_12 NI_12 NS_98 0 1.9004479383174351e-05
GC_12_99 b_12 NI_12 NS_99 0 4.2222587460466910e-04
GC_12_100 b_12 NI_12 NS_100 0 -1.5487110847158155e-04
GC_12_101 b_12 NI_12 NS_101 0 -7.6611114955227126e-06
GC_12_102 b_12 NI_12 NS_102 0 -1.6383417264958292e-05
GC_12_103 b_12 NI_12 NS_103 0 -7.1107541204436654e-04
GC_12_104 b_12 NI_12 NS_104 0 -1.0886741671459968e-04
GC_12_105 b_12 NI_12 NS_105 0 -8.1091816754327505e-07
GC_12_106 b_12 NI_12 NS_106 0 -5.8896374352250936e-10
GC_12_107 b_12 NI_12 NS_107 0 1.5100183848132207e-03
GC_12_108 b_12 NI_12 NS_108 0 -1.5895073923755376e-03
GC_12_109 b_12 NI_12 NS_109 0 3.5732116400193320e-04
GC_12_110 b_12 NI_12 NS_110 0 -4.0707445912455099e-04
GC_12_111 b_12 NI_12 NS_111 0 -2.3298841524700647e-03
GC_12_112 b_12 NI_12 NS_112 0 1.6988277554911273e-03
GC_12_113 b_12 NI_12 NS_113 0 1.7485515571815527e-03
GC_12_114 b_12 NI_12 NS_114 0 3.8653449281827974e-04
GC_12_115 b_12 NI_12 NS_115 0 -1.2185526670873028e-05
GC_12_116 b_12 NI_12 NS_116 0 -3.3252706034112958e-06
GC_12_117 b_12 NI_12 NS_117 0 7.3132799415179013e-06
GC_12_118 b_12 NI_12 NS_118 0 -8.9166320993637764e-05
GC_12_119 b_12 NI_12 NS_119 0 1.5646765883131196e-05
GC_12_120 b_12 NI_12 NS_120 0 4.4586684816458777e-04
GC_12_121 b_12 NI_12 NS_121 0 2.7022162808638414e-05
GC_12_122 b_12 NI_12 NS_122 0 4.4550584721133170e-06
GC_12_123 b_12 NI_12 NS_123 0 -2.4050569016618225e-04
GC_12_124 b_12 NI_12 NS_124 0 -1.7353534191056046e-04
GC_12_125 b_12 NI_12 NS_125 0 -1.3726810061776088e-07
GC_12_126 b_12 NI_12 NS_126 0 2.5285102613826860e-06
GC_12_127 b_12 NI_12 NS_127 0 3.6206565532477183e-06
GC_12_128 b_12 NI_12 NS_128 0 2.5996820071154722e-04
GC_12_129 b_12 NI_12 NS_129 0 3.1493560595960116e-06
GC_12_130 b_12 NI_12 NS_130 0 1.6102220818290540e-06
GC_12_131 b_12 NI_12 NS_131 0 1.7946365295986384e-06
GC_12_132 b_12 NI_12 NS_132 0 -1.3999347707322027e-05
GC_12_133 b_12 NI_12 NS_133 0 3.1093345948536919e-04
GC_12_134 b_12 NI_12 NS_134 0 -2.0352139483486499e-04
GC_12_135 b_12 NI_12 NS_135 0 -3.1096404437801461e-05
GC_12_136 b_12 NI_12 NS_136 0 4.6536347840627337e-05
GC_12_137 b_12 NI_12 NS_137 0 5.4021915109088809e-03
GC_12_138 b_12 NI_12 NS_138 0 -4.3347041531720585e-04
GC_12_139 b_12 NI_12 NS_139 0 -4.7316388994856155e-07
GC_12_140 b_12 NI_12 NS_140 0 2.1518604563602693e-09
GC_12_141 b_12 NI_12 NS_141 0 -1.9034798304654976e-03
GC_12_142 b_12 NI_12 NS_142 0 1.7235837900078158e-03
GC_12_143 b_12 NI_12 NS_143 0 -7.6963967366949293e-04
GC_12_144 b_12 NI_12 NS_144 0 9.4718963763853797e-04
GC_12_145 b_12 NI_12 NS_145 0 1.9703905496639214e-03
GC_12_146 b_12 NI_12 NS_146 0 -1.0335461861524765e-03
GC_12_147 b_12 NI_12 NS_147 0 -1.4931659050930631e-03
GC_12_148 b_12 NI_12 NS_148 0 -7.1921904121939617e-04
GC_12_149 b_12 NI_12 NS_149 0 -3.1306277256056093e-06
GC_12_150 b_12 NI_12 NS_150 0 -9.4461694871495806e-07
GC_12_151 b_12 NI_12 NS_151 0 5.4250483145182997e-06
GC_12_152 b_12 NI_12 NS_152 0 -1.8420696429615884e-05
GC_12_153 b_12 NI_12 NS_153 0 2.1202949840831053e-04
GC_12_154 b_12 NI_12 NS_154 0 1.5543282000323919e-04
GC_12_155 b_12 NI_12 NS_155 0 -4.1713394816652230e-06
GC_12_156 b_12 NI_12 NS_156 0 1.2719169810938734e-06
GC_12_157 b_12 NI_12 NS_157 0 -7.8345093850077865e-05
GC_12_158 b_12 NI_12 NS_158 0 -2.1931706819699464e-05
GC_12_159 b_12 NI_12 NS_159 0 1.6913556323487986e-06
GC_12_160 b_12 NI_12 NS_160 0 -7.6928567921969549e-07
GC_12_161 b_12 NI_12 NS_161 0 -3.4506707819707626e-04
GC_12_162 b_12 NI_12 NS_162 0 2.2281254495658061e-04
GC_12_163 b_12 NI_12 NS_163 0 -8.3649277327889862e-06
GC_12_164 b_12 NI_12 NS_164 0 2.0621718487104089e-05
GC_12_165 b_12 NI_12 NS_165 0 -3.2667030722376924e-06
GC_12_166 b_12 NI_12 NS_166 0 9.6005345501586721e-06
GC_12_167 b_12 NI_12 NS_167 0 4.1271426934801113e-04
GC_12_168 b_12 NI_12 NS_168 0 -2.3123692117707617e-04
GC_12_169 b_12 NI_12 NS_169 0 -5.5405070964848976e-06
GC_12_170 b_12 NI_12 NS_170 0 -1.5541171684278643e-05
GC_12_171 b_12 NI_12 NS_171 0 -6.3951021741088312e-03
GC_12_172 b_12 NI_12 NS_172 0 -2.3783108151938688e-05
GC_12_173 b_12 NI_12 NS_173 0 -2.5485691726449258e-06
GC_12_174 b_12 NI_12 NS_174 0 -7.9759324360269189e-10
GC_12_175 b_12 NI_12 NS_175 0 1.5307383227665251e-03
GC_12_176 b_12 NI_12 NS_176 0 -4.4623337415699406e-03
GC_12_177 b_12 NI_12 NS_177 0 -2.2304610618305369e-04
GC_12_178 b_12 NI_12 NS_178 0 7.2350779701030310e-04
GC_12_179 b_12 NI_12 NS_179 0 1.0093170567694312e-03
GC_12_180 b_12 NI_12 NS_180 0 8.9321352094758706e-04
GC_12_181 b_12 NI_12 NS_181 0 1.5186876505331936e-03
GC_12_182 b_12 NI_12 NS_182 0 -6.0194469681754589e-05
GC_12_183 b_12 NI_12 NS_183 0 -1.0877541359814826e-06
GC_12_184 b_12 NI_12 NS_184 0 9.7781402829674724e-07
GC_12_185 b_12 NI_12 NS_185 0 7.2087177239118294e-06
GC_12_186 b_12 NI_12 NS_186 0 -8.7170163146132448e-05
GC_12_187 b_12 NI_12 NS_187 0 2.4865907211427475e-05
GC_12_188 b_12 NI_12 NS_188 0 4.3046785004867362e-04
GC_12_189 b_12 NI_12 NS_189 0 1.0752707601450207e-05
GC_12_190 b_12 NI_12 NS_190 0 1.0506743129900463e-05
GC_12_191 b_12 NI_12 NS_191 0 -7.4276529153277488e-05
GC_12_192 b_12 NI_12 NS_192 0 -9.1464436208432362e-05
GC_12_193 b_12 NI_12 NS_193 0 -2.0937102532120052e-07
GC_12_194 b_12 NI_12 NS_194 0 -3.2000860858210709e-07
GC_12_195 b_12 NI_12 NS_195 0 -1.3885870299092652e-04
GC_12_196 b_12 NI_12 NS_196 0 2.5435662702331198e-04
GC_12_197 b_12 NI_12 NS_197 0 -6.5013013106614582e-07
GC_12_198 b_12 NI_12 NS_198 0 -2.6367835736132276e-06
GC_12_199 b_12 NI_12 NS_199 0 -1.2320950719266049e-07
GC_12_200 b_12 NI_12 NS_200 0 -7.8646778842242478e-06
GC_12_201 b_12 NI_12 NS_201 0 3.1397802795283533e-04
GC_12_202 b_12 NI_12 NS_202 0 -2.3071869344332851e-04
GC_12_203 b_12 NI_12 NS_203 0 -3.2997646825010636e-05
GC_12_204 b_12 NI_12 NS_204 0 5.3916329890326607e-05
GC_12_205 b_12 NI_12 NS_205 0 1.3936750548694690e-02
GC_12_206 b_12 NI_12 NS_206 0 -1.2484203547880716e-03
GC_12_207 b_12 NI_12 NS_207 0 2.8354314945840004e-07
GC_12_208 b_12 NI_12 NS_208 0 3.8420151946958098e-09
GC_12_209 b_12 NI_12 NS_209 0 -4.7465225610172244e-03
GC_12_210 b_12 NI_12 NS_210 0 5.5905942338339452e-03
GC_12_211 b_12 NI_12 NS_211 0 -1.3138867824258335e-04
GC_12_212 b_12 NI_12 NS_212 0 1.0235720043542968e-03
GC_12_213 b_12 NI_12 NS_213 0 8.8111113064689300e-04
GC_12_214 b_12 NI_12 NS_214 0 -4.4268509474025761e-03
GC_12_215 b_12 NI_12 NS_215 0 -4.1857713582038594e-03
GC_12_216 b_12 NI_12 NS_216 0 -1.4272309606988831e-05
GC_12_217 b_12 NI_12 NS_217 0 3.1299454465437259e-08
GC_12_218 b_12 NI_12 NS_218 0 1.3833946973820873e-06
GC_12_219 b_12 NI_12 NS_219 0 5.0846050248910007e-06
GC_12_220 b_12 NI_12 NS_220 0 -1.8531650726133757e-05
GC_12_221 b_12 NI_12 NS_221 0 2.1293938965086229e-04
GC_12_222 b_12 NI_12 NS_222 0 1.5751652486226171e-04
GC_12_223 b_12 NI_12 NS_223 0 7.4030530031346945e-06
GC_12_224 b_12 NI_12 NS_224 0 -5.0261413861836046e-06
GC_12_225 b_12 NI_12 NS_225 0 8.8747250471163256e-05
GC_12_226 b_12 NI_12 NS_226 0 5.3004730174246515e-05
GC_12_227 b_12 NI_12 NS_227 0 1.3083437171332484e-06
GC_12_228 b_12 NI_12 NS_228 0 -8.3288338959608503e-07
GC_12_229 b_12 NI_12 NS_229 0 -2.0379441753783241e-04
GC_12_230 b_12 NI_12 NS_230 0 -5.2154931435704433e-05
GC_12_231 b_12 NI_12 NS_231 0 -9.3552815655733701e-06
GC_12_232 b_12 NI_12 NS_232 0 1.1802204564078875e-05
GC_12_233 b_12 NI_12 NS_233 0 4.6625653576242680e-06
GC_12_234 b_12 NI_12 NS_234 0 -1.0818817826878400e-05
GC_12_235 b_12 NI_12 NS_235 0 3.7299566824070001e-04
GC_12_236 b_12 NI_12 NS_236 0 -1.7985703097944040e-04
GC_12_237 b_12 NI_12 NS_237 0 -6.6060896338987326e-06
GC_12_238 b_12 NI_12 NS_238 0 -1.6686381850653957e-05
GC_12_239 b_12 NI_12 NS_239 0 -4.9772910896456538e-03
GC_12_240 b_12 NI_12 NS_240 0 -1.1266643529689640e-03
GC_12_241 b_12 NI_12 NS_241 0 -2.6341708700385613e-06
GC_12_242 b_12 NI_12 NS_242 0 -3.8358654127033019e-09
GC_12_243 b_12 NI_12 NS_243 0 1.0462664272477969e-03
GC_12_244 b_12 NI_12 NS_244 0 -6.0151260514778801e-03
GC_12_245 b_12 NI_12 NS_245 0 -8.7833336302619973e-05
GC_12_246 b_12 NI_12 NS_246 0 9.4914415164105807e-04
GC_12_247 b_12 NI_12 NS_247 0 1.1864345172459760e-03
GC_12_248 b_12 NI_12 NS_248 0 1.5554165197538314e-04
GC_12_249 b_12 NI_12 NS_249 0 8.2659335499771366e-04
GC_12_250 b_12 NI_12 NS_250 0 5.1629955730622776e-04
GC_12_251 b_12 NI_12 NS_251 0 -2.9638396104115540e-07
GC_12_252 b_12 NI_12 NS_252 0 -2.2021630740161471e-07
GC_12_253 b_12 NI_12 NS_253 0 6.8168008497221241e-06
GC_12_254 b_12 NI_12 NS_254 0 -8.8474630890139616e-05
GC_12_255 b_12 NI_12 NS_255 0 2.8604111530207097e-05
GC_12_256 b_12 NI_12 NS_256 0 4.4299738249024807e-04
GC_12_257 b_12 NI_12 NS_257 0 -1.0363779117260595e-05
GC_12_258 b_12 NI_12 NS_258 0 -1.2493028772536341e-05
GC_12_259 b_12 NI_12 NS_259 0 8.9670277202776697e-05
GC_12_260 b_12 NI_12 NS_260 0 9.7367347326795842e-05
GC_12_261 b_12 NI_12 NS_261 0 -6.5670960725981244e-07
GC_12_262 b_12 NI_12 NS_262 0 6.5978772479396110e-07
GC_12_263 b_12 NI_12 NS_263 0 -8.9565272280627041e-05
GC_12_264 b_12 NI_12 NS_264 0 2.2613767600273246e-05
GC_12_265 b_12 NI_12 NS_265 0 -3.5415336241131986e-06
GC_12_266 b_12 NI_12 NS_266 0 -9.0492543711766060e-06
GC_12_267 b_12 NI_12 NS_267 0 -1.4574007693618493e-07
GC_12_268 b_12 NI_12 NS_268 0 7.3218997594901718e-06
GC_12_269 b_12 NI_12 NS_269 0 3.1925330957455536e-04
GC_12_270 b_12 NI_12 NS_270 0 -2.0400940367125214e-04
GC_12_271 b_12 NI_12 NS_271 0 -3.4234310094000023e-05
GC_12_272 b_12 NI_12 NS_272 0 5.4063725607148064e-05
GC_12_273 b_12 NI_12 NS_273 0 2.9656910325822527e-02
GC_12_274 b_12 NI_12 NS_274 0 -3.2240710615324564e-03
GC_12_275 b_12 NI_12 NS_275 0 -3.0242884577545581e-06
GC_12_276 b_12 NI_12 NS_276 0 1.0012975955410279e-08
GC_12_277 b_12 NI_12 NS_277 0 -1.4820437656735495e-02
GC_12_278 b_12 NI_12 NS_278 0 1.1000118134645156e-02
GC_12_279 b_12 NI_12 NS_279 0 7.4272684059373717e-05
GC_12_280 b_12 NI_12 NS_280 0 1.0507069708176921e-03
GC_12_281 b_12 NI_12 NS_281 0 3.9318983208203578e-03
GC_12_282 b_12 NI_12 NS_282 0 -8.2689653683234027e-03
GC_12_283 b_12 NI_12 NS_283 0 -7.9225737659077995e-03
GC_12_284 b_12 NI_12 NS_284 0 -2.3804916213319336e-03
GC_12_285 b_12 NI_12 NS_285 0 1.7230085691224870e-06
GC_12_286 b_12 NI_12 NS_286 0 -9.5635417741211182e-06
GC_12_287 b_12 NI_12 NS_287 0 5.2441220113645213e-06
GC_12_288 b_12 NI_12 NS_288 0 -1.7522146783344789e-05
GC_12_289 b_12 NI_12 NS_289 0 2.1111779570685791e-04
GC_12_290 b_12 NI_12 NS_290 0 1.5544864654285930e-04
GC_12_291 b_12 NI_12 NS_291 0 1.8456679960384097e-05
GC_12_292 b_12 NI_12 NS_292 0 -1.4649661224851075e-05
GC_12_293 b_12 NI_12 NS_293 0 2.3050905121949503e-04
GC_12_294 b_12 NI_12 NS_294 0 1.2623634044912910e-04
GC_12_295 b_12 NI_12 NS_295 0 5.0505510521077014e-06
GC_12_296 b_12 NI_12 NS_296 0 -2.9278756998618038e-07
GC_12_297 b_12 NI_12 NS_297 0 -7.4157463101595878e-05
GC_12_298 b_12 NI_12 NS_298 0 -3.5714688593890977e-04
GC_12_299 b_12 NI_12 NS_299 0 -1.0631028954115732e-05
GC_12_300 b_12 NI_12 NS_300 0 -4.3752481927563254e-07
GC_12_301 b_12 NI_12 NS_301 0 9.2794980912119219e-07
GC_12_302 b_12 NI_12 NS_302 0 -1.9517784016937868e-05
GC_12_303 b_12 NI_12 NS_303 0 2.6513899405992530e-04
GC_12_304 b_12 NI_12 NS_304 0 -2.0076366107916042e-04
GC_12_305 b_12 NI_12 NS_305 0 -6.1723377981796085e-06
GC_12_306 b_12 NI_12 NS_306 0 -1.5741342079358015e-05
GC_12_307 b_12 NI_12 NS_307 0 -1.5709202977264216e-02
GC_12_308 b_12 NI_12 NS_308 0 -1.2852377346699497e-03
GC_12_309 b_12 NI_12 NS_309 0 -1.6948749949338027e-05
GC_12_310 b_12 NI_12 NS_310 0 -4.9325201096850420e-09
GC_12_311 b_12 NI_12 NS_311 0 7.2871517503671187e-03
GC_12_312 b_12 NI_12 NS_312 0 -1.3528681160454930e-02
GC_12_313 b_12 NI_12 NS_313 0 -9.6944374512814577e-04
GC_12_314 b_12 NI_12 NS_314 0 1.6623626397277984e-03
GC_12_315 b_12 NI_12 NS_315 0 2.2776295521392486e-03
GC_12_316 b_12 NI_12 NS_316 0 3.2069828681123942e-03
GC_12_317 b_12 NI_12 NS_317 0 2.7331968758511497e-03
GC_12_318 b_12 NI_12 NS_318 0 2.2195795937111650e-03
GC_12_319 b_12 NI_12 NS_319 0 1.1760832703476865e-05
GC_12_320 b_12 NI_12 NS_320 0 2.9617409166189521e-06
GC_12_321 b_12 NI_12 NS_321 0 7.0112858347957106e-06
GC_12_322 b_12 NI_12 NS_322 0 -8.8599702107063959e-05
GC_12_323 b_12 NI_12 NS_323 0 2.0588916038624325e-05
GC_12_324 b_12 NI_12 NS_324 0 4.3950844952571713e-04
GC_12_325 b_12 NI_12 NS_325 0 -2.5994275149227010e-05
GC_12_326 b_12 NI_12 NS_326 0 -6.1374918495775940e-06
GC_12_327 b_12 NI_12 NS_327 0 2.4842737211969889e-04
GC_12_328 b_12 NI_12 NS_328 0 1.7728963419060391e-04
GC_12_329 b_12 NI_12 NS_329 0 7.4130893792789666e-07
GC_12_330 b_12 NI_12 NS_330 0 1.1002428071542538e-06
GC_12_331 b_12 NI_12 NS_331 0 -8.7761661771038036e-05
GC_12_332 b_12 NI_12 NS_332 0 -1.8930878958226804e-04
GC_12_333 b_12 NI_12 NS_333 0 -4.8544284757692293e-06
GC_12_334 b_12 NI_12 NS_334 0 -5.7048634552030375e-06
GC_12_335 b_12 NI_12 NS_335 0 -2.0432769362112074e-06
GC_12_336 b_12 NI_12 NS_336 0 1.3068857642177785e-05
GC_12_337 b_12 NI_12 NS_337 0 2.4719791746856141e-04
GC_12_338 b_12 NI_12 NS_338 0 -1.3516402708012762e-04
GC_12_339 b_12 NI_12 NS_339 0 -3.0989886279489757e-05
GC_12_340 b_12 NI_12 NS_340 0 4.6298397489286863e-05
GC_12_341 b_12 NI_12 NS_341 0 3.2724712848655073e-02
GC_12_342 b_12 NI_12 NS_342 0 3.2736865829842872e-02
GC_12_343 b_12 NI_12 NS_343 0 1.6523826842596316e-04
GC_12_344 b_12 NI_12 NS_344 0 2.5349385201451214e-07
GC_12_345 b_12 NI_12 NS_345 0 -6.0934733235492505e-02
GC_12_346 b_12 NI_12 NS_346 0 -1.7132985253020181e-02
GC_12_347 b_12 NI_12 NS_347 0 -1.7899288486096245e-03
GC_12_348 b_12 NI_12 NS_348 0 4.8602799554595339e-03
GC_12_349 b_12 NI_12 NS_349 0 1.2185134042684244e-02
GC_12_350 b_12 NI_12 NS_350 0 1.6811852108492429e-02
GC_12_351 b_12 NI_12 NS_351 0 7.1137381325896256e-03
GC_12_352 b_12 NI_12 NS_352 0 8.1971668483051511e-05
GC_12_353 b_12 NI_12 NS_353 0 -5.2197829980936962e-07
GC_12_354 b_12 NI_12 NS_354 0 -1.3005900083568962e-05
GC_12_355 b_12 NI_12 NS_355 0 2.7206797507700593e-06
GC_12_356 b_12 NI_12 NS_356 0 -1.7277001032917340e-05
GC_12_357 b_12 NI_12 NS_357 0 2.2114793591013112e-04
GC_12_358 b_12 NI_12 NS_358 0 1.5871324948177104e-04
GC_12_359 b_12 NI_12 NS_359 0 2.4015034757781868e-05
GC_12_360 b_12 NI_12 NS_360 0 -1.4432352317698314e-05
GC_12_361 b_12 NI_12 NS_361 0 3.3597212679355279e-04
GC_12_362 b_12 NI_12 NS_362 0 1.4568791291196109e-04
GC_12_363 b_12 NI_12 NS_363 0 -1.2531813364834015e-06
GC_12_364 b_12 NI_12 NS_364 0 -9.3013173451061838e-07
GC_12_365 b_12 NI_12 NS_365 0 3.7106916007323469e-04
GC_12_366 b_12 NI_12 NS_366 0 -6.4126373706166592e-04
GC_12_367 b_12 NI_12 NS_367 0 -3.8412984249672822e-06
GC_12_368 b_12 NI_12 NS_368 0 -2.4749018005479831e-05
GC_12_369 b_12 NI_12 NS_369 0 3.2526367684450603e-06
GC_12_370 b_12 NI_12 NS_370 0 -3.4178723602264679e-05
GC_12_371 b_12 NI_12 NS_371 0 4.2186427370161328e-04
GC_12_372 b_12 NI_12 NS_372 0 -5.1895135702768504e-05
GC_12_373 b_12 NI_12 NS_373 0 -1.1686946616027080e-05
GC_12_374 b_12 NI_12 NS_374 0 -1.7937694350618287e-05
GC_12_375 b_12 NI_12 NS_375 0 4.2201837536707254e-03
GC_12_376 b_12 NI_12 NS_376 0 2.9204513907572730e-02
GC_12_377 b_12 NI_12 NS_377 0 5.8739838230819135e-05
GC_12_378 b_12 NI_12 NS_378 0 -7.0229537413896974e-08
GC_12_379 b_12 NI_12 NS_379 0 4.8322536494817853e-02
GC_12_380 b_12 NI_12 NS_380 0 3.6908801395367744e-02
GC_12_381 b_12 NI_12 NS_381 0 -4.6968298894514956e-03
GC_12_382 b_12 NI_12 NS_382 0 2.5557764748820396e-03
GC_12_383 b_12 NI_12 NS_383 0 -7.2918034652796320e-03
GC_12_384 b_12 NI_12 NS_384 0 1.5060047268266220e-02
GC_12_385 b_12 NI_12 NS_385 0 1.0981764362058026e-03
GC_12_386 b_12 NI_12 NS_386 0 4.7287169266712788e-03
GC_12_387 b_12 NI_12 NS_387 0 1.2811237967185636e-05
GC_12_388 b_12 NI_12 NS_388 0 2.6464103517361870e-06
GC_12_389 b_12 NI_12 NS_389 0 7.3338745377910708e-06
GC_12_390 b_12 NI_12 NS_390 0 -8.5275195054598544e-05
GC_12_391 b_12 NI_12 NS_391 0 1.1345850783583701e-05
GC_12_392 b_12 NI_12 NS_392 0 4.2586114593162961e-04
GC_12_393 b_12 NI_12 NS_393 0 -3.7496538317018099e-05
GC_12_394 b_12 NI_12 NS_394 0 -2.1913383555818310e-05
GC_12_395 b_12 NI_12 NS_395 0 3.2373882268205655e-04
GC_12_396 b_12 NI_12 NS_396 0 3.0002357458530047e-04
GC_12_397 b_12 NI_12 NS_397 0 -2.8234443462946003e-06
GC_12_398 b_12 NI_12 NS_398 0 1.5860362933572922e-06
GC_12_399 b_12 NI_12 NS_399 0 1.5265579516734497e-04
GC_12_400 b_12 NI_12 NS_400 0 -4.2565284157939585e-04
GC_12_401 b_12 NI_12 NS_401 0 -3.9169688855094544e-06
GC_12_402 b_12 NI_12 NS_402 0 -8.9382001199418510e-06
GC_12_403 b_12 NI_12 NS_403 0 -2.7669257818435537e-06
GC_12_404 b_12 NI_12 NS_404 0 1.8944329863211846e-05
GC_12_405 b_12 NI_12 NS_405 0 3.4993096041980139e-04
GC_12_406 b_12 NI_12 NS_406 0 -8.3943082752623187e-05
GC_12_407 b_12 NI_12 NS_407 0 -3.6053520230202817e-05
GC_12_408 b_12 NI_12 NS_408 0 4.6757704612185648e-05
GD_12_1 b_12 NI_12 NA_1 0 -5.0035970948097003e-03
GD_12_2 b_12 NI_12 NA_2 0 -3.5936837648275631e-03
GD_12_3 b_12 NI_12 NA_3 0 -4.7388169087013658e-03
GD_12_4 b_12 NI_12 NA_4 0 -1.1463015675026299e-03
GD_12_5 b_12 NI_12 NA_5 0 -4.6948962146504602e-03
GD_12_6 b_12 NI_12 NA_6 0 2.5563951663638454e-03
GD_12_7 b_12 NI_12 NA_7 0 -6.2212618473697816e-03
GD_12_8 b_12 NI_12 NA_8 0 3.6971902711345583e-03
GD_12_9 b_12 NI_12 NA_9 0 -1.0119964535331044e-02
GD_12_10 b_12 NI_12 NA_10 0 7.1021990973039791e-03
GD_12_11 b_12 NI_12 NA_11 0 -3.5191581735794647e-02
GD_12_12 b_12 NI_12 NA_12 0 -2.5228578540554830e-01
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 3.4256132957802641e+00
GS_1_1 0 NS_1 NA_1 0 1.5251913417194629e+00
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 8.6582773449483081e+00
GS_2_1 0 NS_2 NA_1 0 1.5251913417194629e+00
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 3.1453339577953656e+01
GS_3_1 0 NS_3 NA_1 0 1.5251913417194629e+00
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 1.2483716714088728e+03
GS_4_1 0 NS_4 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 9.5700292143510275e+00
RS_6 NS_6 0 9.5700292143510275e+00
GL_5 0 NS_5 NS_6 0 1.4040628101439498e-01
GL_6 0 NS_6 NS_5 0 -1.4040628101439498e-01
GS_5_1 0 NS_5 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 4.0462967855885069e+01
RS_8 NS_8 0 4.0462967855885061e+01
GL_7 0 NS_7 NS_8 0 2.6673201695183885e-01
GL_8 0 NS_8 NS_7 0 -2.6673201695183885e-01
GS_7_1 0 NS_7 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 1.9059070407967361e+01
RS_10 NS_10 0 1.9059070407967358e+01
GL_9 0 NS_9 NS_10 0 2.4185814461526237e-01
GL_10 0 NS_10 NS_9 0 -2.4185814461526237e-01
GS_9_1 0 NS_9 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 1.7666316379915560e+01
RS_12 NS_12 0 1.7666316379915564e+01
GL_11 0 NS_11 NS_12 0 1.9702615210896449e-01
GL_12 0 NS_12 NS_11 0 -1.9702615210896449e-01
GS_11_1 0 NS_11 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 3.4591856087420081e+02
RS_14 NS_14 0 3.4591856087420081e+02
GL_13 0 NS_13 NS_14 0 2.4170685235821462e-01
GL_14 0 NS_14 NS_13 0 -2.4170685235821462e-01
GS_13_1 0 NS_13 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 3.4257938362763537e+02
RS_16 NS_16 0 3.4257938362763537e+02
GL_15 0 NS_15 NS_16 0 1.4255159266867465e-01
GL_16 0 NS_16 NS_15 0 -1.4255159266867465e-01
GS_15_1 0 NS_15 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 1.0126954757407573e+02
RS_18 NS_18 0 1.0126954757407573e+02
GL_17 0 NS_17 NS_18 0 1.4356554078688363e-01
GL_18 0 NS_18 NS_17 0 -1.4356554078688363e-01
GS_17_1 0 NS_17 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 3.5335368091933424e+02
RS_20 NS_20 0 3.5335368091933418e+02
GL_19 0 NS_19 NS_20 0 1.6640381409742028e-01
GL_20 0 NS_20 NS_19 0 -1.6640381409742028e-01
GS_19_1 0 NS_19 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 1.1172419684791065e+02
RS_22 NS_22 0 1.1172419684791066e+02
GL_21 0 NS_21 NS_22 0 1.6662138407694810e-01
GL_22 0 NS_22 NS_21 0 -1.6662138407694810e-01
GS_21_1 0 NS_21 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 2.3124949155545121e+02
RS_24 NS_24 0 2.3124949155545121e+02
GL_23 0 NS_23 NS_24 0 1.8384390380970300e-01
GL_24 0 NS_24 NS_23 0 -1.8384390380970300e-01
GS_23_1 0 NS_23 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 8.6778721170894016e+01
RS_26 NS_26 0 8.6778721170894002e+01
GL_25 0 NS_25 NS_26 0 2.2562932600183958e-01
GL_26 0 NS_26 NS_25 0 -2.2562932600183958e-01
GS_25_1 0 NS_25 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 3.2996671012988776e+02
RS_28 NS_28 0 3.2996671012988776e+02
GL_27 0 NS_27 NS_28 0 2.2283373301463522e-01
GL_28 0 NS_28 NS_27 0 -2.2283373301463522e-01
GS_27_1 0 NS_27 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 3.9174610175015977e+02
RS_30 NS_30 0 3.9174610175015977e+02
GL_29 0 NS_29 NS_30 0 2.1918798560265801e-01
GL_30 0 NS_30 NS_29 0 -2.1918798560265801e-01
GS_29_1 0 NS_29 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 7.1523254667023437e+01
RS_32 NS_32 0 7.1523254667023451e+01
GL_31 0 NS_31 NS_32 0 2.0613705597202187e-01
GL_32 0 NS_32 NS_31 0 -2.0613705597202187e-01
GS_31_1 0 NS_31 NA_1 0 1.5251913417194629e+00
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 3.4487804113693971e+02
RS_34 NS_34 0 3.4487804113693966e+02
GL_33 0 NS_33 NS_34 0 2.0650350471279413e-01
GL_34 0 NS_34 NS_33 0 -2.0650350471279413e-01
GS_33_1 0 NS_33 NA_1 0 1.5251913417194629e+00
*
* Real pole n. 35
CS_35 NS_35 0 9.9999999999999998e-13
RS_35 NS_35 0 3.4256132957802641e+00
GS_35_2 0 NS_35 NA_2 0 1.5251913417194629e+00
*
* Real pole n. 36
CS_36 NS_36 0 9.9999999999999998e-13
RS_36 NS_36 0 8.6582773449483081e+00
GS_36_2 0 NS_36 NA_2 0 1.5251913417194629e+00
*
* Real pole n. 37
CS_37 NS_37 0 9.9999999999999998e-13
RS_37 NS_37 0 3.1453339577953656e+01
GS_37_2 0 NS_37 NA_2 0 1.5251913417194629e+00
*
* Real pole n. 38
CS_38 NS_38 0 9.9999999999999998e-13
RS_38 NS_38 0 1.2483716714088728e+03
GS_38_2 0 NS_38 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 9.5700292143510275e+00
RS_40 NS_40 0 9.5700292143510275e+00
GL_39 0 NS_39 NS_40 0 1.4040628101439498e-01
GL_40 0 NS_40 NS_39 0 -1.4040628101439498e-01
GS_39_2 0 NS_39 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 4.0462967855885069e+01
RS_42 NS_42 0 4.0462967855885061e+01
GL_41 0 NS_41 NS_42 0 2.6673201695183885e-01
GL_42 0 NS_42 NS_41 0 -2.6673201695183885e-01
GS_41_2 0 NS_41 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 1.9059070407967361e+01
RS_44 NS_44 0 1.9059070407967358e+01
GL_43 0 NS_43 NS_44 0 2.4185814461526237e-01
GL_44 0 NS_44 NS_43 0 -2.4185814461526237e-01
GS_43_2 0 NS_43 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 1.7666316379915560e+01
RS_46 NS_46 0 1.7666316379915564e+01
GL_45 0 NS_45 NS_46 0 1.9702615210896449e-01
GL_46 0 NS_46 NS_45 0 -1.9702615210896449e-01
GS_45_2 0 NS_45 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 3.4591856087420081e+02
RS_48 NS_48 0 3.4591856087420081e+02
GL_47 0 NS_47 NS_48 0 2.4170685235821462e-01
GL_48 0 NS_48 NS_47 0 -2.4170685235821462e-01
GS_47_2 0 NS_47 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 3.4257938362763537e+02
RS_50 NS_50 0 3.4257938362763537e+02
GL_49 0 NS_49 NS_50 0 1.4255159266867465e-01
GL_50 0 NS_50 NS_49 0 -1.4255159266867465e-01
GS_49_2 0 NS_49 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 1.0126954757407573e+02
RS_52 NS_52 0 1.0126954757407573e+02
GL_51 0 NS_51 NS_52 0 1.4356554078688363e-01
GL_52 0 NS_52 NS_51 0 -1.4356554078688363e-01
GS_51_2 0 NS_51 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 3.5335368091933424e+02
RS_54 NS_54 0 3.5335368091933418e+02
GL_53 0 NS_53 NS_54 0 1.6640381409742028e-01
GL_54 0 NS_54 NS_53 0 -1.6640381409742028e-01
GS_53_2 0 NS_53 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 1.1172419684791065e+02
RS_56 NS_56 0 1.1172419684791066e+02
GL_55 0 NS_55 NS_56 0 1.6662138407694810e-01
GL_56 0 NS_56 NS_55 0 -1.6662138407694810e-01
GS_55_2 0 NS_55 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 2.3124949155545121e+02
RS_58 NS_58 0 2.3124949155545121e+02
GL_57 0 NS_57 NS_58 0 1.8384390380970300e-01
GL_58 0 NS_58 NS_57 0 -1.8384390380970300e-01
GS_57_2 0 NS_57 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 8.6778721170894016e+01
RS_60 NS_60 0 8.6778721170894002e+01
GL_59 0 NS_59 NS_60 0 2.2562932600183958e-01
GL_60 0 NS_60 NS_59 0 -2.2562932600183958e-01
GS_59_2 0 NS_59 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 3.2996671012988776e+02
RS_62 NS_62 0 3.2996671012988776e+02
GL_61 0 NS_61 NS_62 0 2.2283373301463522e-01
GL_62 0 NS_62 NS_61 0 -2.2283373301463522e-01
GS_61_2 0 NS_61 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 3.9174610175015977e+02
RS_64 NS_64 0 3.9174610175015977e+02
GL_63 0 NS_63 NS_64 0 2.1918798560265801e-01
GL_64 0 NS_64 NS_63 0 -2.1918798560265801e-01
GS_63_2 0 NS_63 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 7.1523254667023437e+01
RS_66 NS_66 0 7.1523254667023451e+01
GL_65 0 NS_65 NS_66 0 2.0613705597202187e-01
GL_66 0 NS_66 NS_65 0 -2.0613705597202187e-01
GS_65_2 0 NS_65 NA_2 0 1.5251913417194629e+00
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 3.4487804113693971e+02
RS_68 NS_68 0 3.4487804113693966e+02
GL_67 0 NS_67 NS_68 0 2.0650350471279413e-01
GL_68 0 NS_68 NS_67 0 -2.0650350471279413e-01
GS_67_2 0 NS_67 NA_2 0 1.5251913417194629e+00
*
* Real pole n. 69
CS_69 NS_69 0 9.9999999999999998e-13
RS_69 NS_69 0 3.4256132957802641e+00
GS_69_3 0 NS_69 NA_3 0 1.5251913417194629e+00
*
* Real pole n. 70
CS_70 NS_70 0 9.9999999999999998e-13
RS_70 NS_70 0 8.6582773449483081e+00
GS_70_3 0 NS_70 NA_3 0 1.5251913417194629e+00
*
* Real pole n. 71
CS_71 NS_71 0 9.9999999999999998e-13
RS_71 NS_71 0 3.1453339577953656e+01
GS_71_3 0 NS_71 NA_3 0 1.5251913417194629e+00
*
* Real pole n. 72
CS_72 NS_72 0 9.9999999999999998e-13
RS_72 NS_72 0 1.2483716714088728e+03
GS_72_3 0 NS_72 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 9.5700292143510275e+00
RS_74 NS_74 0 9.5700292143510275e+00
GL_73 0 NS_73 NS_74 0 1.4040628101439498e-01
GL_74 0 NS_74 NS_73 0 -1.4040628101439498e-01
GS_73_3 0 NS_73 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 4.0462967855885069e+01
RS_76 NS_76 0 4.0462967855885061e+01
GL_75 0 NS_75 NS_76 0 2.6673201695183885e-01
GL_76 0 NS_76 NS_75 0 -2.6673201695183885e-01
GS_75_3 0 NS_75 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 1.9059070407967361e+01
RS_78 NS_78 0 1.9059070407967358e+01
GL_77 0 NS_77 NS_78 0 2.4185814461526237e-01
GL_78 0 NS_78 NS_77 0 -2.4185814461526237e-01
GS_77_3 0 NS_77 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 1.7666316379915560e+01
RS_80 NS_80 0 1.7666316379915564e+01
GL_79 0 NS_79 NS_80 0 1.9702615210896449e-01
GL_80 0 NS_80 NS_79 0 -1.9702615210896449e-01
GS_79_3 0 NS_79 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 3.4591856087420081e+02
RS_82 NS_82 0 3.4591856087420081e+02
GL_81 0 NS_81 NS_82 0 2.4170685235821462e-01
GL_82 0 NS_82 NS_81 0 -2.4170685235821462e-01
GS_81_3 0 NS_81 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 3.4257938362763537e+02
RS_84 NS_84 0 3.4257938362763537e+02
GL_83 0 NS_83 NS_84 0 1.4255159266867465e-01
GL_84 0 NS_84 NS_83 0 -1.4255159266867465e-01
GS_83_3 0 NS_83 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 1.0126954757407573e+02
RS_86 NS_86 0 1.0126954757407573e+02
GL_85 0 NS_85 NS_86 0 1.4356554078688363e-01
GL_86 0 NS_86 NS_85 0 -1.4356554078688363e-01
GS_85_3 0 NS_85 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 3.5335368091933424e+02
RS_88 NS_88 0 3.5335368091933418e+02
GL_87 0 NS_87 NS_88 0 1.6640381409742028e-01
GL_88 0 NS_88 NS_87 0 -1.6640381409742028e-01
GS_87_3 0 NS_87 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 1.1172419684791065e+02
RS_90 NS_90 0 1.1172419684791066e+02
GL_89 0 NS_89 NS_90 0 1.6662138407694810e-01
GL_90 0 NS_90 NS_89 0 -1.6662138407694810e-01
GS_89_3 0 NS_89 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 2.3124949155545121e+02
RS_92 NS_92 0 2.3124949155545121e+02
GL_91 0 NS_91 NS_92 0 1.8384390380970300e-01
GL_92 0 NS_92 NS_91 0 -1.8384390380970300e-01
GS_91_3 0 NS_91 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 8.6778721170894016e+01
RS_94 NS_94 0 8.6778721170894002e+01
GL_93 0 NS_93 NS_94 0 2.2562932600183958e-01
GL_94 0 NS_94 NS_93 0 -2.2562932600183958e-01
GS_93_3 0 NS_93 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 3.2996671012988776e+02
RS_96 NS_96 0 3.2996671012988776e+02
GL_95 0 NS_95 NS_96 0 2.2283373301463522e-01
GL_96 0 NS_96 NS_95 0 -2.2283373301463522e-01
GS_95_3 0 NS_95 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 3.9174610175015977e+02
RS_98 NS_98 0 3.9174610175015977e+02
GL_97 0 NS_97 NS_98 0 2.1918798560265801e-01
GL_98 0 NS_98 NS_97 0 -2.1918798560265801e-01
GS_97_3 0 NS_97 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 7.1523254667023437e+01
RS_100 NS_100 0 7.1523254667023451e+01
GL_99 0 NS_99 NS_100 0 2.0613705597202187e-01
GL_100 0 NS_100 NS_99 0 -2.0613705597202187e-01
GS_99_3 0 NS_99 NA_3 0 1.5251913417194629e+00
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 3.4487804113693971e+02
RS_102 NS_102 0 3.4487804113693966e+02
GL_101 0 NS_101 NS_102 0 2.0650350471279413e-01
GL_102 0 NS_102 NS_101 0 -2.0650350471279413e-01
GS_101_3 0 NS_101 NA_3 0 1.5251913417194629e+00
*
* Real pole n. 103
CS_103 NS_103 0 9.9999999999999998e-13
RS_103 NS_103 0 3.4256132957802641e+00
GS_103_4 0 NS_103 NA_4 0 1.5251913417194629e+00
*
* Real pole n. 104
CS_104 NS_104 0 9.9999999999999998e-13
RS_104 NS_104 0 8.6582773449483081e+00
GS_104_4 0 NS_104 NA_4 0 1.5251913417194629e+00
*
* Real pole n. 105
CS_105 NS_105 0 9.9999999999999998e-13
RS_105 NS_105 0 3.1453339577953656e+01
GS_105_4 0 NS_105 NA_4 0 1.5251913417194629e+00
*
* Real pole n. 106
CS_106 NS_106 0 9.9999999999999998e-13
RS_106 NS_106 0 1.2483716714088728e+03
GS_106_4 0 NS_106 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 9.5700292143510275e+00
RS_108 NS_108 0 9.5700292143510275e+00
GL_107 0 NS_107 NS_108 0 1.4040628101439498e-01
GL_108 0 NS_108 NS_107 0 -1.4040628101439498e-01
GS_107_4 0 NS_107 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 4.0462967855885069e+01
RS_110 NS_110 0 4.0462967855885061e+01
GL_109 0 NS_109 NS_110 0 2.6673201695183885e-01
GL_110 0 NS_110 NS_109 0 -2.6673201695183885e-01
GS_109_4 0 NS_109 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 1.9059070407967361e+01
RS_112 NS_112 0 1.9059070407967358e+01
GL_111 0 NS_111 NS_112 0 2.4185814461526237e-01
GL_112 0 NS_112 NS_111 0 -2.4185814461526237e-01
GS_111_4 0 NS_111 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 1.7666316379915560e+01
RS_114 NS_114 0 1.7666316379915564e+01
GL_113 0 NS_113 NS_114 0 1.9702615210896449e-01
GL_114 0 NS_114 NS_113 0 -1.9702615210896449e-01
GS_113_4 0 NS_113 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 3.4591856087420081e+02
RS_116 NS_116 0 3.4591856087420081e+02
GL_115 0 NS_115 NS_116 0 2.4170685235821462e-01
GL_116 0 NS_116 NS_115 0 -2.4170685235821462e-01
GS_115_4 0 NS_115 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 3.4257938362763537e+02
RS_118 NS_118 0 3.4257938362763537e+02
GL_117 0 NS_117 NS_118 0 1.4255159266867465e-01
GL_118 0 NS_118 NS_117 0 -1.4255159266867465e-01
GS_117_4 0 NS_117 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 1.0126954757407573e+02
RS_120 NS_120 0 1.0126954757407573e+02
GL_119 0 NS_119 NS_120 0 1.4356554078688363e-01
GL_120 0 NS_120 NS_119 0 -1.4356554078688363e-01
GS_119_4 0 NS_119 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 3.5335368091933424e+02
RS_122 NS_122 0 3.5335368091933418e+02
GL_121 0 NS_121 NS_122 0 1.6640381409742028e-01
GL_122 0 NS_122 NS_121 0 -1.6640381409742028e-01
GS_121_4 0 NS_121 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 1.1172419684791065e+02
RS_124 NS_124 0 1.1172419684791066e+02
GL_123 0 NS_123 NS_124 0 1.6662138407694810e-01
GL_124 0 NS_124 NS_123 0 -1.6662138407694810e-01
GS_123_4 0 NS_123 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 2.3124949155545121e+02
RS_126 NS_126 0 2.3124949155545121e+02
GL_125 0 NS_125 NS_126 0 1.8384390380970300e-01
GL_126 0 NS_126 NS_125 0 -1.8384390380970300e-01
GS_125_4 0 NS_125 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 8.6778721170894016e+01
RS_128 NS_128 0 8.6778721170894002e+01
GL_127 0 NS_127 NS_128 0 2.2562932600183958e-01
GL_128 0 NS_128 NS_127 0 -2.2562932600183958e-01
GS_127_4 0 NS_127 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 3.2996671012988776e+02
RS_130 NS_130 0 3.2996671012988776e+02
GL_129 0 NS_129 NS_130 0 2.2283373301463522e-01
GL_130 0 NS_130 NS_129 0 -2.2283373301463522e-01
GS_129_4 0 NS_129 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 3.9174610175015977e+02
RS_132 NS_132 0 3.9174610175015977e+02
GL_131 0 NS_131 NS_132 0 2.1918798560265801e-01
GL_132 0 NS_132 NS_131 0 -2.1918798560265801e-01
GS_131_4 0 NS_131 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 133/134
CS_133 NS_133 0 9.9999999999999998e-13
CS_134 NS_134 0 9.9999999999999998e-13
RS_133 NS_133 0 7.1523254667023437e+01
RS_134 NS_134 0 7.1523254667023451e+01
GL_133 0 NS_133 NS_134 0 2.0613705597202187e-01
GL_134 0 NS_134 NS_133 0 -2.0613705597202187e-01
GS_133_4 0 NS_133 NA_4 0 1.5251913417194629e+00
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 3.4487804113693971e+02
RS_136 NS_136 0 3.4487804113693966e+02
GL_135 0 NS_135 NS_136 0 2.0650350471279413e-01
GL_136 0 NS_136 NS_135 0 -2.0650350471279413e-01
GS_135_4 0 NS_135 NA_4 0 1.5251913417194629e+00
*
* Real pole n. 137
CS_137 NS_137 0 9.9999999999999998e-13
RS_137 NS_137 0 3.4256132957802641e+00
GS_137_5 0 NS_137 NA_5 0 1.5251913417194629e+00
*
* Real pole n. 138
CS_138 NS_138 0 9.9999999999999998e-13
RS_138 NS_138 0 8.6582773449483081e+00
GS_138_5 0 NS_138 NA_5 0 1.5251913417194629e+00
*
* Real pole n. 139
CS_139 NS_139 0 9.9999999999999998e-13
RS_139 NS_139 0 3.1453339577953656e+01
GS_139_5 0 NS_139 NA_5 0 1.5251913417194629e+00
*
* Real pole n. 140
CS_140 NS_140 0 9.9999999999999998e-13
RS_140 NS_140 0 1.2483716714088728e+03
GS_140_5 0 NS_140 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 9.5700292143510275e+00
RS_142 NS_142 0 9.5700292143510275e+00
GL_141 0 NS_141 NS_142 0 1.4040628101439498e-01
GL_142 0 NS_142 NS_141 0 -1.4040628101439498e-01
GS_141_5 0 NS_141 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 4.0462967855885069e+01
RS_144 NS_144 0 4.0462967855885061e+01
GL_143 0 NS_143 NS_144 0 2.6673201695183885e-01
GL_144 0 NS_144 NS_143 0 -2.6673201695183885e-01
GS_143_5 0 NS_143 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 1.9059070407967361e+01
RS_146 NS_146 0 1.9059070407967358e+01
GL_145 0 NS_145 NS_146 0 2.4185814461526237e-01
GL_146 0 NS_146 NS_145 0 -2.4185814461526237e-01
GS_145_5 0 NS_145 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 1.7666316379915560e+01
RS_148 NS_148 0 1.7666316379915564e+01
GL_147 0 NS_147 NS_148 0 1.9702615210896449e-01
GL_148 0 NS_148 NS_147 0 -1.9702615210896449e-01
GS_147_5 0 NS_147 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 3.4591856087420081e+02
RS_150 NS_150 0 3.4591856087420081e+02
GL_149 0 NS_149 NS_150 0 2.4170685235821462e-01
GL_150 0 NS_150 NS_149 0 -2.4170685235821462e-01
GS_149_5 0 NS_149 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 3.4257938362763537e+02
RS_152 NS_152 0 3.4257938362763537e+02
GL_151 0 NS_151 NS_152 0 1.4255159266867465e-01
GL_152 0 NS_152 NS_151 0 -1.4255159266867465e-01
GS_151_5 0 NS_151 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 1.0126954757407573e+02
RS_154 NS_154 0 1.0126954757407573e+02
GL_153 0 NS_153 NS_154 0 1.4356554078688363e-01
GL_154 0 NS_154 NS_153 0 -1.4356554078688363e-01
GS_153_5 0 NS_153 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 3.5335368091933424e+02
RS_156 NS_156 0 3.5335368091933418e+02
GL_155 0 NS_155 NS_156 0 1.6640381409742028e-01
GL_156 0 NS_156 NS_155 0 -1.6640381409742028e-01
GS_155_5 0 NS_155 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 1.1172419684791065e+02
RS_158 NS_158 0 1.1172419684791066e+02
GL_157 0 NS_157 NS_158 0 1.6662138407694810e-01
GL_158 0 NS_158 NS_157 0 -1.6662138407694810e-01
GS_157_5 0 NS_157 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 2.3124949155545121e+02
RS_160 NS_160 0 2.3124949155545121e+02
GL_159 0 NS_159 NS_160 0 1.8384390380970300e-01
GL_160 0 NS_160 NS_159 0 -1.8384390380970300e-01
GS_159_5 0 NS_159 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 8.6778721170894016e+01
RS_162 NS_162 0 8.6778721170894002e+01
GL_161 0 NS_161 NS_162 0 2.2562932600183958e-01
GL_162 0 NS_162 NS_161 0 -2.2562932600183958e-01
GS_161_5 0 NS_161 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 163/164
CS_163 NS_163 0 9.9999999999999998e-13
CS_164 NS_164 0 9.9999999999999998e-13
RS_163 NS_163 0 3.2996671012988776e+02
RS_164 NS_164 0 3.2996671012988776e+02
GL_163 0 NS_163 NS_164 0 2.2283373301463522e-01
GL_164 0 NS_164 NS_163 0 -2.2283373301463522e-01
GS_163_5 0 NS_163 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 3.9174610175015977e+02
RS_166 NS_166 0 3.9174610175015977e+02
GL_165 0 NS_165 NS_166 0 2.1918798560265801e-01
GL_166 0 NS_166 NS_165 0 -2.1918798560265801e-01
GS_165_5 0 NS_165 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 7.1523254667023437e+01
RS_168 NS_168 0 7.1523254667023451e+01
GL_167 0 NS_167 NS_168 0 2.0613705597202187e-01
GL_168 0 NS_168 NS_167 0 -2.0613705597202187e-01
GS_167_5 0 NS_167 NA_5 0 1.5251913417194629e+00
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 3.4487804113693971e+02
RS_170 NS_170 0 3.4487804113693966e+02
GL_169 0 NS_169 NS_170 0 2.0650350471279413e-01
GL_170 0 NS_170 NS_169 0 -2.0650350471279413e-01
GS_169_5 0 NS_169 NA_5 0 1.5251913417194629e+00
*
* Real pole n. 171
CS_171 NS_171 0 9.9999999999999998e-13
RS_171 NS_171 0 3.4256132957802641e+00
GS_171_6 0 NS_171 NA_6 0 1.5251913417194629e+00
*
* Real pole n. 172
CS_172 NS_172 0 9.9999999999999998e-13
RS_172 NS_172 0 8.6582773449483081e+00
GS_172_6 0 NS_172 NA_6 0 1.5251913417194629e+00
*
* Real pole n. 173
CS_173 NS_173 0 9.9999999999999998e-13
RS_173 NS_173 0 3.1453339577953656e+01
GS_173_6 0 NS_173 NA_6 0 1.5251913417194629e+00
*
* Real pole n. 174
CS_174 NS_174 0 9.9999999999999998e-13
RS_174 NS_174 0 1.2483716714088728e+03
GS_174_6 0 NS_174 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 9.5700292143510275e+00
RS_176 NS_176 0 9.5700292143510275e+00
GL_175 0 NS_175 NS_176 0 1.4040628101439498e-01
GL_176 0 NS_176 NS_175 0 -1.4040628101439498e-01
GS_175_6 0 NS_175 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 4.0462967855885069e+01
RS_178 NS_178 0 4.0462967855885061e+01
GL_177 0 NS_177 NS_178 0 2.6673201695183885e-01
GL_178 0 NS_178 NS_177 0 -2.6673201695183885e-01
GS_177_6 0 NS_177 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 1.9059070407967361e+01
RS_180 NS_180 0 1.9059070407967358e+01
GL_179 0 NS_179 NS_180 0 2.4185814461526237e-01
GL_180 0 NS_180 NS_179 0 -2.4185814461526237e-01
GS_179_6 0 NS_179 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 181/182
CS_181 NS_181 0 9.9999999999999998e-13
CS_182 NS_182 0 9.9999999999999998e-13
RS_181 NS_181 0 1.7666316379915560e+01
RS_182 NS_182 0 1.7666316379915564e+01
GL_181 0 NS_181 NS_182 0 1.9702615210896449e-01
GL_182 0 NS_182 NS_181 0 -1.9702615210896449e-01
GS_181_6 0 NS_181 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 183/184
CS_183 NS_183 0 9.9999999999999998e-13
CS_184 NS_184 0 9.9999999999999998e-13
RS_183 NS_183 0 3.4591856087420081e+02
RS_184 NS_184 0 3.4591856087420081e+02
GL_183 0 NS_183 NS_184 0 2.4170685235821462e-01
GL_184 0 NS_184 NS_183 0 -2.4170685235821462e-01
GS_183_6 0 NS_183 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 3.4257938362763537e+02
RS_186 NS_186 0 3.4257938362763537e+02
GL_185 0 NS_185 NS_186 0 1.4255159266867465e-01
GL_186 0 NS_186 NS_185 0 -1.4255159266867465e-01
GS_185_6 0 NS_185 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 1.0126954757407573e+02
RS_188 NS_188 0 1.0126954757407573e+02
GL_187 0 NS_187 NS_188 0 1.4356554078688363e-01
GL_188 0 NS_188 NS_187 0 -1.4356554078688363e-01
GS_187_6 0 NS_187 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 3.5335368091933424e+02
RS_190 NS_190 0 3.5335368091933418e+02
GL_189 0 NS_189 NS_190 0 1.6640381409742028e-01
GL_190 0 NS_190 NS_189 0 -1.6640381409742028e-01
GS_189_6 0 NS_189 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 1.1172419684791065e+02
RS_192 NS_192 0 1.1172419684791066e+02
GL_191 0 NS_191 NS_192 0 1.6662138407694810e-01
GL_192 0 NS_192 NS_191 0 -1.6662138407694810e-01
GS_191_6 0 NS_191 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 2.3124949155545121e+02
RS_194 NS_194 0 2.3124949155545121e+02
GL_193 0 NS_193 NS_194 0 1.8384390380970300e-01
GL_194 0 NS_194 NS_193 0 -1.8384390380970300e-01
GS_193_6 0 NS_193 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 8.6778721170894016e+01
RS_196 NS_196 0 8.6778721170894002e+01
GL_195 0 NS_195 NS_196 0 2.2562932600183958e-01
GL_196 0 NS_196 NS_195 0 -2.2562932600183958e-01
GS_195_6 0 NS_195 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 3.2996671012988776e+02
RS_198 NS_198 0 3.2996671012988776e+02
GL_197 0 NS_197 NS_198 0 2.2283373301463522e-01
GL_198 0 NS_198 NS_197 0 -2.2283373301463522e-01
GS_197_6 0 NS_197 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 3.9174610175015977e+02
RS_200 NS_200 0 3.9174610175015977e+02
GL_199 0 NS_199 NS_200 0 2.1918798560265801e-01
GL_200 0 NS_200 NS_199 0 -2.1918798560265801e-01
GS_199_6 0 NS_199 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 201/202
CS_201 NS_201 0 9.9999999999999998e-13
CS_202 NS_202 0 9.9999999999999998e-13
RS_201 NS_201 0 7.1523254667023437e+01
RS_202 NS_202 0 7.1523254667023451e+01
GL_201 0 NS_201 NS_202 0 2.0613705597202187e-01
GL_202 0 NS_202 NS_201 0 -2.0613705597202187e-01
GS_201_6 0 NS_201 NA_6 0 1.5251913417194629e+00
*
* Complex pair n. 203/204
CS_203 NS_203 0 9.9999999999999998e-13
CS_204 NS_204 0 9.9999999999999998e-13
RS_203 NS_203 0 3.4487804113693971e+02
RS_204 NS_204 0 3.4487804113693966e+02
GL_203 0 NS_203 NS_204 0 2.0650350471279413e-01
GL_204 0 NS_204 NS_203 0 -2.0650350471279413e-01
GS_203_6 0 NS_203 NA_6 0 1.5251913417194629e+00
*
* Real pole n. 205
CS_205 NS_205 0 9.9999999999999998e-13
RS_205 NS_205 0 3.4256132957802641e+00
GS_205_7 0 NS_205 NA_7 0 1.5251913417194629e+00
*
* Real pole n. 206
CS_206 NS_206 0 9.9999999999999998e-13
RS_206 NS_206 0 8.6582773449483081e+00
GS_206_7 0 NS_206 NA_7 0 1.5251913417194629e+00
*
* Real pole n. 207
CS_207 NS_207 0 9.9999999999999998e-13
RS_207 NS_207 0 3.1453339577953656e+01
GS_207_7 0 NS_207 NA_7 0 1.5251913417194629e+00
*
* Real pole n. 208
CS_208 NS_208 0 9.9999999999999998e-13
RS_208 NS_208 0 1.2483716714088728e+03
GS_208_7 0 NS_208 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 9.5700292143510275e+00
RS_210 NS_210 0 9.5700292143510275e+00
GL_209 0 NS_209 NS_210 0 1.4040628101439498e-01
GL_210 0 NS_210 NS_209 0 -1.4040628101439498e-01
GS_209_7 0 NS_209 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 4.0462967855885069e+01
RS_212 NS_212 0 4.0462967855885061e+01
GL_211 0 NS_211 NS_212 0 2.6673201695183885e-01
GL_212 0 NS_212 NS_211 0 -2.6673201695183885e-01
GS_211_7 0 NS_211 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 1.9059070407967361e+01
RS_214 NS_214 0 1.9059070407967358e+01
GL_213 0 NS_213 NS_214 0 2.4185814461526237e-01
GL_214 0 NS_214 NS_213 0 -2.4185814461526237e-01
GS_213_7 0 NS_213 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 1.7666316379915560e+01
RS_216 NS_216 0 1.7666316379915564e+01
GL_215 0 NS_215 NS_216 0 1.9702615210896449e-01
GL_216 0 NS_216 NS_215 0 -1.9702615210896449e-01
GS_215_7 0 NS_215 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 3.4591856087420081e+02
RS_218 NS_218 0 3.4591856087420081e+02
GL_217 0 NS_217 NS_218 0 2.4170685235821462e-01
GL_218 0 NS_218 NS_217 0 -2.4170685235821462e-01
GS_217_7 0 NS_217 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 3.4257938362763537e+02
RS_220 NS_220 0 3.4257938362763537e+02
GL_219 0 NS_219 NS_220 0 1.4255159266867465e-01
GL_220 0 NS_220 NS_219 0 -1.4255159266867465e-01
GS_219_7 0 NS_219 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 221/222
CS_221 NS_221 0 9.9999999999999998e-13
CS_222 NS_222 0 9.9999999999999998e-13
RS_221 NS_221 0 1.0126954757407573e+02
RS_222 NS_222 0 1.0126954757407573e+02
GL_221 0 NS_221 NS_222 0 1.4356554078688363e-01
GL_222 0 NS_222 NS_221 0 -1.4356554078688363e-01
GS_221_7 0 NS_221 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 223/224
CS_223 NS_223 0 9.9999999999999998e-13
CS_224 NS_224 0 9.9999999999999998e-13
RS_223 NS_223 0 3.5335368091933424e+02
RS_224 NS_224 0 3.5335368091933418e+02
GL_223 0 NS_223 NS_224 0 1.6640381409742028e-01
GL_224 0 NS_224 NS_223 0 -1.6640381409742028e-01
GS_223_7 0 NS_223 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 225/226
CS_225 NS_225 0 9.9999999999999998e-13
CS_226 NS_226 0 9.9999999999999998e-13
RS_225 NS_225 0 1.1172419684791065e+02
RS_226 NS_226 0 1.1172419684791066e+02
GL_225 0 NS_225 NS_226 0 1.6662138407694810e-01
GL_226 0 NS_226 NS_225 0 -1.6662138407694810e-01
GS_225_7 0 NS_225 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 2.3124949155545121e+02
RS_228 NS_228 0 2.3124949155545121e+02
GL_227 0 NS_227 NS_228 0 1.8384390380970300e-01
GL_228 0 NS_228 NS_227 0 -1.8384390380970300e-01
GS_227_7 0 NS_227 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 229/230
CS_229 NS_229 0 9.9999999999999998e-13
CS_230 NS_230 0 9.9999999999999998e-13
RS_229 NS_229 0 8.6778721170894016e+01
RS_230 NS_230 0 8.6778721170894002e+01
GL_229 0 NS_229 NS_230 0 2.2562932600183958e-01
GL_230 0 NS_230 NS_229 0 -2.2562932600183958e-01
GS_229_7 0 NS_229 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 3.2996671012988776e+02
RS_232 NS_232 0 3.2996671012988776e+02
GL_231 0 NS_231 NS_232 0 2.2283373301463522e-01
GL_232 0 NS_232 NS_231 0 -2.2283373301463522e-01
GS_231_7 0 NS_231 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 3.9174610175015977e+02
RS_234 NS_234 0 3.9174610175015977e+02
GL_233 0 NS_233 NS_234 0 2.1918798560265801e-01
GL_234 0 NS_234 NS_233 0 -2.1918798560265801e-01
GS_233_7 0 NS_233 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 7.1523254667023437e+01
RS_236 NS_236 0 7.1523254667023451e+01
GL_235 0 NS_235 NS_236 0 2.0613705597202187e-01
GL_236 0 NS_236 NS_235 0 -2.0613705597202187e-01
GS_235_7 0 NS_235 NA_7 0 1.5251913417194629e+00
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 3.4487804113693971e+02
RS_238 NS_238 0 3.4487804113693966e+02
GL_237 0 NS_237 NS_238 0 2.0650350471279413e-01
GL_238 0 NS_238 NS_237 0 -2.0650350471279413e-01
GS_237_7 0 NS_237 NA_7 0 1.5251913417194629e+00
*
* Real pole n. 239
CS_239 NS_239 0 9.9999999999999998e-13
RS_239 NS_239 0 3.4256132957802641e+00
GS_239_8 0 NS_239 NA_8 0 1.5251913417194629e+00
*
* Real pole n. 240
CS_240 NS_240 0 9.9999999999999998e-13
RS_240 NS_240 0 8.6582773449483081e+00
GS_240_8 0 NS_240 NA_8 0 1.5251913417194629e+00
*
* Real pole n. 241
CS_241 NS_241 0 9.9999999999999998e-13
RS_241 NS_241 0 3.1453339577953656e+01
GS_241_8 0 NS_241 NA_8 0 1.5251913417194629e+00
*
* Real pole n. 242
CS_242 NS_242 0 9.9999999999999998e-13
RS_242 NS_242 0 1.2483716714088728e+03
GS_242_8 0 NS_242 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 243/244
CS_243 NS_243 0 9.9999999999999998e-13
CS_244 NS_244 0 9.9999999999999998e-13
RS_243 NS_243 0 9.5700292143510275e+00
RS_244 NS_244 0 9.5700292143510275e+00
GL_243 0 NS_243 NS_244 0 1.4040628101439498e-01
GL_244 0 NS_244 NS_243 0 -1.4040628101439498e-01
GS_243_8 0 NS_243 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 245/246
CS_245 NS_245 0 9.9999999999999998e-13
CS_246 NS_246 0 9.9999999999999998e-13
RS_245 NS_245 0 4.0462967855885069e+01
RS_246 NS_246 0 4.0462967855885061e+01
GL_245 0 NS_245 NS_246 0 2.6673201695183885e-01
GL_246 0 NS_246 NS_245 0 -2.6673201695183885e-01
GS_245_8 0 NS_245 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 247/248
CS_247 NS_247 0 9.9999999999999998e-13
CS_248 NS_248 0 9.9999999999999998e-13
RS_247 NS_247 0 1.9059070407967361e+01
RS_248 NS_248 0 1.9059070407967358e+01
GL_247 0 NS_247 NS_248 0 2.4185814461526237e-01
GL_248 0 NS_248 NS_247 0 -2.4185814461526237e-01
GS_247_8 0 NS_247 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 249/250
CS_249 NS_249 0 9.9999999999999998e-13
CS_250 NS_250 0 9.9999999999999998e-13
RS_249 NS_249 0 1.7666316379915560e+01
RS_250 NS_250 0 1.7666316379915564e+01
GL_249 0 NS_249 NS_250 0 1.9702615210896449e-01
GL_250 0 NS_250 NS_249 0 -1.9702615210896449e-01
GS_249_8 0 NS_249 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 251/252
CS_251 NS_251 0 9.9999999999999998e-13
CS_252 NS_252 0 9.9999999999999998e-13
RS_251 NS_251 0 3.4591856087420081e+02
RS_252 NS_252 0 3.4591856087420081e+02
GL_251 0 NS_251 NS_252 0 2.4170685235821462e-01
GL_252 0 NS_252 NS_251 0 -2.4170685235821462e-01
GS_251_8 0 NS_251 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 253/254
CS_253 NS_253 0 9.9999999999999998e-13
CS_254 NS_254 0 9.9999999999999998e-13
RS_253 NS_253 0 3.4257938362763537e+02
RS_254 NS_254 0 3.4257938362763537e+02
GL_253 0 NS_253 NS_254 0 1.4255159266867465e-01
GL_254 0 NS_254 NS_253 0 -1.4255159266867465e-01
GS_253_8 0 NS_253 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 255/256
CS_255 NS_255 0 9.9999999999999998e-13
CS_256 NS_256 0 9.9999999999999998e-13
RS_255 NS_255 0 1.0126954757407573e+02
RS_256 NS_256 0 1.0126954757407573e+02
GL_255 0 NS_255 NS_256 0 1.4356554078688363e-01
GL_256 0 NS_256 NS_255 0 -1.4356554078688363e-01
GS_255_8 0 NS_255 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 257/258
CS_257 NS_257 0 9.9999999999999998e-13
CS_258 NS_258 0 9.9999999999999998e-13
RS_257 NS_257 0 3.5335368091933424e+02
RS_258 NS_258 0 3.5335368091933418e+02
GL_257 0 NS_257 NS_258 0 1.6640381409742028e-01
GL_258 0 NS_258 NS_257 0 -1.6640381409742028e-01
GS_257_8 0 NS_257 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 259/260
CS_259 NS_259 0 9.9999999999999998e-13
CS_260 NS_260 0 9.9999999999999998e-13
RS_259 NS_259 0 1.1172419684791065e+02
RS_260 NS_260 0 1.1172419684791066e+02
GL_259 0 NS_259 NS_260 0 1.6662138407694810e-01
GL_260 0 NS_260 NS_259 0 -1.6662138407694810e-01
GS_259_8 0 NS_259 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 261/262
CS_261 NS_261 0 9.9999999999999998e-13
CS_262 NS_262 0 9.9999999999999998e-13
RS_261 NS_261 0 2.3124949155545121e+02
RS_262 NS_262 0 2.3124949155545121e+02
GL_261 0 NS_261 NS_262 0 1.8384390380970300e-01
GL_262 0 NS_262 NS_261 0 -1.8384390380970300e-01
GS_261_8 0 NS_261 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 263/264
CS_263 NS_263 0 9.9999999999999998e-13
CS_264 NS_264 0 9.9999999999999998e-13
RS_263 NS_263 0 8.6778721170894016e+01
RS_264 NS_264 0 8.6778721170894002e+01
GL_263 0 NS_263 NS_264 0 2.2562932600183958e-01
GL_264 0 NS_264 NS_263 0 -2.2562932600183958e-01
GS_263_8 0 NS_263 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 265/266
CS_265 NS_265 0 9.9999999999999998e-13
CS_266 NS_266 0 9.9999999999999998e-13
RS_265 NS_265 0 3.2996671012988776e+02
RS_266 NS_266 0 3.2996671012988776e+02
GL_265 0 NS_265 NS_266 0 2.2283373301463522e-01
GL_266 0 NS_266 NS_265 0 -2.2283373301463522e-01
GS_265_8 0 NS_265 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 267/268
CS_267 NS_267 0 9.9999999999999998e-13
CS_268 NS_268 0 9.9999999999999998e-13
RS_267 NS_267 0 3.9174610175015977e+02
RS_268 NS_268 0 3.9174610175015977e+02
GL_267 0 NS_267 NS_268 0 2.1918798560265801e-01
GL_268 0 NS_268 NS_267 0 -2.1918798560265801e-01
GS_267_8 0 NS_267 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 269/270
CS_269 NS_269 0 9.9999999999999998e-13
CS_270 NS_270 0 9.9999999999999998e-13
RS_269 NS_269 0 7.1523254667023437e+01
RS_270 NS_270 0 7.1523254667023451e+01
GL_269 0 NS_269 NS_270 0 2.0613705597202187e-01
GL_270 0 NS_270 NS_269 0 -2.0613705597202187e-01
GS_269_8 0 NS_269 NA_8 0 1.5251913417194629e+00
*
* Complex pair n. 271/272
CS_271 NS_271 0 9.9999999999999998e-13
CS_272 NS_272 0 9.9999999999999998e-13
RS_271 NS_271 0 3.4487804113693971e+02
RS_272 NS_272 0 3.4487804113693966e+02
GL_271 0 NS_271 NS_272 0 2.0650350471279413e-01
GL_272 0 NS_272 NS_271 0 -2.0650350471279413e-01
GS_271_8 0 NS_271 NA_8 0 1.5251913417194629e+00
*
* Real pole n. 273
CS_273 NS_273 0 9.9999999999999998e-13
RS_273 NS_273 0 3.4256132957802641e+00
GS_273_9 0 NS_273 NA_9 0 1.5251913417194629e+00
*
* Real pole n. 274
CS_274 NS_274 0 9.9999999999999998e-13
RS_274 NS_274 0 8.6582773449483081e+00
GS_274_9 0 NS_274 NA_9 0 1.5251913417194629e+00
*
* Real pole n. 275
CS_275 NS_275 0 9.9999999999999998e-13
RS_275 NS_275 0 3.1453339577953656e+01
GS_275_9 0 NS_275 NA_9 0 1.5251913417194629e+00
*
* Real pole n. 276
CS_276 NS_276 0 9.9999999999999998e-13
RS_276 NS_276 0 1.2483716714088728e+03
GS_276_9 0 NS_276 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 277/278
CS_277 NS_277 0 9.9999999999999998e-13
CS_278 NS_278 0 9.9999999999999998e-13
RS_277 NS_277 0 9.5700292143510275e+00
RS_278 NS_278 0 9.5700292143510275e+00
GL_277 0 NS_277 NS_278 0 1.4040628101439498e-01
GL_278 0 NS_278 NS_277 0 -1.4040628101439498e-01
GS_277_9 0 NS_277 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 279/280
CS_279 NS_279 0 9.9999999999999998e-13
CS_280 NS_280 0 9.9999999999999998e-13
RS_279 NS_279 0 4.0462967855885069e+01
RS_280 NS_280 0 4.0462967855885061e+01
GL_279 0 NS_279 NS_280 0 2.6673201695183885e-01
GL_280 0 NS_280 NS_279 0 -2.6673201695183885e-01
GS_279_9 0 NS_279 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 281/282
CS_281 NS_281 0 9.9999999999999998e-13
CS_282 NS_282 0 9.9999999999999998e-13
RS_281 NS_281 0 1.9059070407967361e+01
RS_282 NS_282 0 1.9059070407967358e+01
GL_281 0 NS_281 NS_282 0 2.4185814461526237e-01
GL_282 0 NS_282 NS_281 0 -2.4185814461526237e-01
GS_281_9 0 NS_281 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 283/284
CS_283 NS_283 0 9.9999999999999998e-13
CS_284 NS_284 0 9.9999999999999998e-13
RS_283 NS_283 0 1.7666316379915560e+01
RS_284 NS_284 0 1.7666316379915564e+01
GL_283 0 NS_283 NS_284 0 1.9702615210896449e-01
GL_284 0 NS_284 NS_283 0 -1.9702615210896449e-01
GS_283_9 0 NS_283 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 285/286
CS_285 NS_285 0 9.9999999999999998e-13
CS_286 NS_286 0 9.9999999999999998e-13
RS_285 NS_285 0 3.4591856087420081e+02
RS_286 NS_286 0 3.4591856087420081e+02
GL_285 0 NS_285 NS_286 0 2.4170685235821462e-01
GL_286 0 NS_286 NS_285 0 -2.4170685235821462e-01
GS_285_9 0 NS_285 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 287/288
CS_287 NS_287 0 9.9999999999999998e-13
CS_288 NS_288 0 9.9999999999999998e-13
RS_287 NS_287 0 3.4257938362763537e+02
RS_288 NS_288 0 3.4257938362763537e+02
GL_287 0 NS_287 NS_288 0 1.4255159266867465e-01
GL_288 0 NS_288 NS_287 0 -1.4255159266867465e-01
GS_287_9 0 NS_287 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 289/290
CS_289 NS_289 0 9.9999999999999998e-13
CS_290 NS_290 0 9.9999999999999998e-13
RS_289 NS_289 0 1.0126954757407573e+02
RS_290 NS_290 0 1.0126954757407573e+02
GL_289 0 NS_289 NS_290 0 1.4356554078688363e-01
GL_290 0 NS_290 NS_289 0 -1.4356554078688363e-01
GS_289_9 0 NS_289 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 291/292
CS_291 NS_291 0 9.9999999999999998e-13
CS_292 NS_292 0 9.9999999999999998e-13
RS_291 NS_291 0 3.5335368091933424e+02
RS_292 NS_292 0 3.5335368091933418e+02
GL_291 0 NS_291 NS_292 0 1.6640381409742028e-01
GL_292 0 NS_292 NS_291 0 -1.6640381409742028e-01
GS_291_9 0 NS_291 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 293/294
CS_293 NS_293 0 9.9999999999999998e-13
CS_294 NS_294 0 9.9999999999999998e-13
RS_293 NS_293 0 1.1172419684791065e+02
RS_294 NS_294 0 1.1172419684791066e+02
GL_293 0 NS_293 NS_294 0 1.6662138407694810e-01
GL_294 0 NS_294 NS_293 0 -1.6662138407694810e-01
GS_293_9 0 NS_293 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 295/296
CS_295 NS_295 0 9.9999999999999998e-13
CS_296 NS_296 0 9.9999999999999998e-13
RS_295 NS_295 0 2.3124949155545121e+02
RS_296 NS_296 0 2.3124949155545121e+02
GL_295 0 NS_295 NS_296 0 1.8384390380970300e-01
GL_296 0 NS_296 NS_295 0 -1.8384390380970300e-01
GS_295_9 0 NS_295 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 297/298
CS_297 NS_297 0 9.9999999999999998e-13
CS_298 NS_298 0 9.9999999999999998e-13
RS_297 NS_297 0 8.6778721170894016e+01
RS_298 NS_298 0 8.6778721170894002e+01
GL_297 0 NS_297 NS_298 0 2.2562932600183958e-01
GL_298 0 NS_298 NS_297 0 -2.2562932600183958e-01
GS_297_9 0 NS_297 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 299/300
CS_299 NS_299 0 9.9999999999999998e-13
CS_300 NS_300 0 9.9999999999999998e-13
RS_299 NS_299 0 3.2996671012988776e+02
RS_300 NS_300 0 3.2996671012988776e+02
GL_299 0 NS_299 NS_300 0 2.2283373301463522e-01
GL_300 0 NS_300 NS_299 0 -2.2283373301463522e-01
GS_299_9 0 NS_299 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 301/302
CS_301 NS_301 0 9.9999999999999998e-13
CS_302 NS_302 0 9.9999999999999998e-13
RS_301 NS_301 0 3.9174610175015977e+02
RS_302 NS_302 0 3.9174610175015977e+02
GL_301 0 NS_301 NS_302 0 2.1918798560265801e-01
GL_302 0 NS_302 NS_301 0 -2.1918798560265801e-01
GS_301_9 0 NS_301 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 303/304
CS_303 NS_303 0 9.9999999999999998e-13
CS_304 NS_304 0 9.9999999999999998e-13
RS_303 NS_303 0 7.1523254667023437e+01
RS_304 NS_304 0 7.1523254667023451e+01
GL_303 0 NS_303 NS_304 0 2.0613705597202187e-01
GL_304 0 NS_304 NS_303 0 -2.0613705597202187e-01
GS_303_9 0 NS_303 NA_9 0 1.5251913417194629e+00
*
* Complex pair n. 305/306
CS_305 NS_305 0 9.9999999999999998e-13
CS_306 NS_306 0 9.9999999999999998e-13
RS_305 NS_305 0 3.4487804113693971e+02
RS_306 NS_306 0 3.4487804113693966e+02
GL_305 0 NS_305 NS_306 0 2.0650350471279413e-01
GL_306 0 NS_306 NS_305 0 -2.0650350471279413e-01
GS_305_9 0 NS_305 NA_9 0 1.5251913417194629e+00
*
* Real pole n. 307
CS_307 NS_307 0 9.9999999999999998e-13
RS_307 NS_307 0 3.4256132957802641e+00
GS_307_10 0 NS_307 NA_10 0 1.5251913417194629e+00
*
* Real pole n. 308
CS_308 NS_308 0 9.9999999999999998e-13
RS_308 NS_308 0 8.6582773449483081e+00
GS_308_10 0 NS_308 NA_10 0 1.5251913417194629e+00
*
* Real pole n. 309
CS_309 NS_309 0 9.9999999999999998e-13
RS_309 NS_309 0 3.1453339577953656e+01
GS_309_10 0 NS_309 NA_10 0 1.5251913417194629e+00
*
* Real pole n. 310
CS_310 NS_310 0 9.9999999999999998e-13
RS_310 NS_310 0 1.2483716714088728e+03
GS_310_10 0 NS_310 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 311/312
CS_311 NS_311 0 9.9999999999999998e-13
CS_312 NS_312 0 9.9999999999999998e-13
RS_311 NS_311 0 9.5700292143510275e+00
RS_312 NS_312 0 9.5700292143510275e+00
GL_311 0 NS_311 NS_312 0 1.4040628101439498e-01
GL_312 0 NS_312 NS_311 0 -1.4040628101439498e-01
GS_311_10 0 NS_311 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 313/314
CS_313 NS_313 0 9.9999999999999998e-13
CS_314 NS_314 0 9.9999999999999998e-13
RS_313 NS_313 0 4.0462967855885069e+01
RS_314 NS_314 0 4.0462967855885061e+01
GL_313 0 NS_313 NS_314 0 2.6673201695183885e-01
GL_314 0 NS_314 NS_313 0 -2.6673201695183885e-01
GS_313_10 0 NS_313 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 315/316
CS_315 NS_315 0 9.9999999999999998e-13
CS_316 NS_316 0 9.9999999999999998e-13
RS_315 NS_315 0 1.9059070407967361e+01
RS_316 NS_316 0 1.9059070407967358e+01
GL_315 0 NS_315 NS_316 0 2.4185814461526237e-01
GL_316 0 NS_316 NS_315 0 -2.4185814461526237e-01
GS_315_10 0 NS_315 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 317/318
CS_317 NS_317 0 9.9999999999999998e-13
CS_318 NS_318 0 9.9999999999999998e-13
RS_317 NS_317 0 1.7666316379915560e+01
RS_318 NS_318 0 1.7666316379915564e+01
GL_317 0 NS_317 NS_318 0 1.9702615210896449e-01
GL_318 0 NS_318 NS_317 0 -1.9702615210896449e-01
GS_317_10 0 NS_317 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 319/320
CS_319 NS_319 0 9.9999999999999998e-13
CS_320 NS_320 0 9.9999999999999998e-13
RS_319 NS_319 0 3.4591856087420081e+02
RS_320 NS_320 0 3.4591856087420081e+02
GL_319 0 NS_319 NS_320 0 2.4170685235821462e-01
GL_320 0 NS_320 NS_319 0 -2.4170685235821462e-01
GS_319_10 0 NS_319 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 321/322
CS_321 NS_321 0 9.9999999999999998e-13
CS_322 NS_322 0 9.9999999999999998e-13
RS_321 NS_321 0 3.4257938362763537e+02
RS_322 NS_322 0 3.4257938362763537e+02
GL_321 0 NS_321 NS_322 0 1.4255159266867465e-01
GL_322 0 NS_322 NS_321 0 -1.4255159266867465e-01
GS_321_10 0 NS_321 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 323/324
CS_323 NS_323 0 9.9999999999999998e-13
CS_324 NS_324 0 9.9999999999999998e-13
RS_323 NS_323 0 1.0126954757407573e+02
RS_324 NS_324 0 1.0126954757407573e+02
GL_323 0 NS_323 NS_324 0 1.4356554078688363e-01
GL_324 0 NS_324 NS_323 0 -1.4356554078688363e-01
GS_323_10 0 NS_323 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 325/326
CS_325 NS_325 0 9.9999999999999998e-13
CS_326 NS_326 0 9.9999999999999998e-13
RS_325 NS_325 0 3.5335368091933424e+02
RS_326 NS_326 0 3.5335368091933418e+02
GL_325 0 NS_325 NS_326 0 1.6640381409742028e-01
GL_326 0 NS_326 NS_325 0 -1.6640381409742028e-01
GS_325_10 0 NS_325 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 327/328
CS_327 NS_327 0 9.9999999999999998e-13
CS_328 NS_328 0 9.9999999999999998e-13
RS_327 NS_327 0 1.1172419684791065e+02
RS_328 NS_328 0 1.1172419684791066e+02
GL_327 0 NS_327 NS_328 0 1.6662138407694810e-01
GL_328 0 NS_328 NS_327 0 -1.6662138407694810e-01
GS_327_10 0 NS_327 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 329/330
CS_329 NS_329 0 9.9999999999999998e-13
CS_330 NS_330 0 9.9999999999999998e-13
RS_329 NS_329 0 2.3124949155545121e+02
RS_330 NS_330 0 2.3124949155545121e+02
GL_329 0 NS_329 NS_330 0 1.8384390380970300e-01
GL_330 0 NS_330 NS_329 0 -1.8384390380970300e-01
GS_329_10 0 NS_329 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 331/332
CS_331 NS_331 0 9.9999999999999998e-13
CS_332 NS_332 0 9.9999999999999998e-13
RS_331 NS_331 0 8.6778721170894016e+01
RS_332 NS_332 0 8.6778721170894002e+01
GL_331 0 NS_331 NS_332 0 2.2562932600183958e-01
GL_332 0 NS_332 NS_331 0 -2.2562932600183958e-01
GS_331_10 0 NS_331 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 333/334
CS_333 NS_333 0 9.9999999999999998e-13
CS_334 NS_334 0 9.9999999999999998e-13
RS_333 NS_333 0 3.2996671012988776e+02
RS_334 NS_334 0 3.2996671012988776e+02
GL_333 0 NS_333 NS_334 0 2.2283373301463522e-01
GL_334 0 NS_334 NS_333 0 -2.2283373301463522e-01
GS_333_10 0 NS_333 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 335/336
CS_335 NS_335 0 9.9999999999999998e-13
CS_336 NS_336 0 9.9999999999999998e-13
RS_335 NS_335 0 3.9174610175015977e+02
RS_336 NS_336 0 3.9174610175015977e+02
GL_335 0 NS_335 NS_336 0 2.1918798560265801e-01
GL_336 0 NS_336 NS_335 0 -2.1918798560265801e-01
GS_335_10 0 NS_335 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 337/338
CS_337 NS_337 0 9.9999999999999998e-13
CS_338 NS_338 0 9.9999999999999998e-13
RS_337 NS_337 0 7.1523254667023437e+01
RS_338 NS_338 0 7.1523254667023451e+01
GL_337 0 NS_337 NS_338 0 2.0613705597202187e-01
GL_338 0 NS_338 NS_337 0 -2.0613705597202187e-01
GS_337_10 0 NS_337 NA_10 0 1.5251913417194629e+00
*
* Complex pair n. 339/340
CS_339 NS_339 0 9.9999999999999998e-13
CS_340 NS_340 0 9.9999999999999998e-13
RS_339 NS_339 0 3.4487804113693971e+02
RS_340 NS_340 0 3.4487804113693966e+02
GL_339 0 NS_339 NS_340 0 2.0650350471279413e-01
GL_340 0 NS_340 NS_339 0 -2.0650350471279413e-01
GS_339_10 0 NS_339 NA_10 0 1.5251913417194629e+00
*
* Real pole n. 341
CS_341 NS_341 0 9.9999999999999998e-13
RS_341 NS_341 0 3.4256132957802641e+00
GS_341_11 0 NS_341 NA_11 0 1.5251913417194629e+00
*
* Real pole n. 342
CS_342 NS_342 0 9.9999999999999998e-13
RS_342 NS_342 0 8.6582773449483081e+00
GS_342_11 0 NS_342 NA_11 0 1.5251913417194629e+00
*
* Real pole n. 343
CS_343 NS_343 0 9.9999999999999998e-13
RS_343 NS_343 0 3.1453339577953656e+01
GS_343_11 0 NS_343 NA_11 0 1.5251913417194629e+00
*
* Real pole n. 344
CS_344 NS_344 0 9.9999999999999998e-13
RS_344 NS_344 0 1.2483716714088728e+03
GS_344_11 0 NS_344 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 345/346
CS_345 NS_345 0 9.9999999999999998e-13
CS_346 NS_346 0 9.9999999999999998e-13
RS_345 NS_345 0 9.5700292143510275e+00
RS_346 NS_346 0 9.5700292143510275e+00
GL_345 0 NS_345 NS_346 0 1.4040628101439498e-01
GL_346 0 NS_346 NS_345 0 -1.4040628101439498e-01
GS_345_11 0 NS_345 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 347/348
CS_347 NS_347 0 9.9999999999999998e-13
CS_348 NS_348 0 9.9999999999999998e-13
RS_347 NS_347 0 4.0462967855885069e+01
RS_348 NS_348 0 4.0462967855885061e+01
GL_347 0 NS_347 NS_348 0 2.6673201695183885e-01
GL_348 0 NS_348 NS_347 0 -2.6673201695183885e-01
GS_347_11 0 NS_347 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 349/350
CS_349 NS_349 0 9.9999999999999998e-13
CS_350 NS_350 0 9.9999999999999998e-13
RS_349 NS_349 0 1.9059070407967361e+01
RS_350 NS_350 0 1.9059070407967358e+01
GL_349 0 NS_349 NS_350 0 2.4185814461526237e-01
GL_350 0 NS_350 NS_349 0 -2.4185814461526237e-01
GS_349_11 0 NS_349 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 351/352
CS_351 NS_351 0 9.9999999999999998e-13
CS_352 NS_352 0 9.9999999999999998e-13
RS_351 NS_351 0 1.7666316379915560e+01
RS_352 NS_352 0 1.7666316379915564e+01
GL_351 0 NS_351 NS_352 0 1.9702615210896449e-01
GL_352 0 NS_352 NS_351 0 -1.9702615210896449e-01
GS_351_11 0 NS_351 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 353/354
CS_353 NS_353 0 9.9999999999999998e-13
CS_354 NS_354 0 9.9999999999999998e-13
RS_353 NS_353 0 3.4591856087420081e+02
RS_354 NS_354 0 3.4591856087420081e+02
GL_353 0 NS_353 NS_354 0 2.4170685235821462e-01
GL_354 0 NS_354 NS_353 0 -2.4170685235821462e-01
GS_353_11 0 NS_353 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 355/356
CS_355 NS_355 0 9.9999999999999998e-13
CS_356 NS_356 0 9.9999999999999998e-13
RS_355 NS_355 0 3.4257938362763537e+02
RS_356 NS_356 0 3.4257938362763537e+02
GL_355 0 NS_355 NS_356 0 1.4255159266867465e-01
GL_356 0 NS_356 NS_355 0 -1.4255159266867465e-01
GS_355_11 0 NS_355 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 357/358
CS_357 NS_357 0 9.9999999999999998e-13
CS_358 NS_358 0 9.9999999999999998e-13
RS_357 NS_357 0 1.0126954757407573e+02
RS_358 NS_358 0 1.0126954757407573e+02
GL_357 0 NS_357 NS_358 0 1.4356554078688363e-01
GL_358 0 NS_358 NS_357 0 -1.4356554078688363e-01
GS_357_11 0 NS_357 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 359/360
CS_359 NS_359 0 9.9999999999999998e-13
CS_360 NS_360 0 9.9999999999999998e-13
RS_359 NS_359 0 3.5335368091933424e+02
RS_360 NS_360 0 3.5335368091933418e+02
GL_359 0 NS_359 NS_360 0 1.6640381409742028e-01
GL_360 0 NS_360 NS_359 0 -1.6640381409742028e-01
GS_359_11 0 NS_359 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 361/362
CS_361 NS_361 0 9.9999999999999998e-13
CS_362 NS_362 0 9.9999999999999998e-13
RS_361 NS_361 0 1.1172419684791065e+02
RS_362 NS_362 0 1.1172419684791066e+02
GL_361 0 NS_361 NS_362 0 1.6662138407694810e-01
GL_362 0 NS_362 NS_361 0 -1.6662138407694810e-01
GS_361_11 0 NS_361 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 363/364
CS_363 NS_363 0 9.9999999999999998e-13
CS_364 NS_364 0 9.9999999999999998e-13
RS_363 NS_363 0 2.3124949155545121e+02
RS_364 NS_364 0 2.3124949155545121e+02
GL_363 0 NS_363 NS_364 0 1.8384390380970300e-01
GL_364 0 NS_364 NS_363 0 -1.8384390380970300e-01
GS_363_11 0 NS_363 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 365/366
CS_365 NS_365 0 9.9999999999999998e-13
CS_366 NS_366 0 9.9999999999999998e-13
RS_365 NS_365 0 8.6778721170894016e+01
RS_366 NS_366 0 8.6778721170894002e+01
GL_365 0 NS_365 NS_366 0 2.2562932600183958e-01
GL_366 0 NS_366 NS_365 0 -2.2562932600183958e-01
GS_365_11 0 NS_365 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 367/368
CS_367 NS_367 0 9.9999999999999998e-13
CS_368 NS_368 0 9.9999999999999998e-13
RS_367 NS_367 0 3.2996671012988776e+02
RS_368 NS_368 0 3.2996671012988776e+02
GL_367 0 NS_367 NS_368 0 2.2283373301463522e-01
GL_368 0 NS_368 NS_367 0 -2.2283373301463522e-01
GS_367_11 0 NS_367 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 369/370
CS_369 NS_369 0 9.9999999999999998e-13
CS_370 NS_370 0 9.9999999999999998e-13
RS_369 NS_369 0 3.9174610175015977e+02
RS_370 NS_370 0 3.9174610175015977e+02
GL_369 0 NS_369 NS_370 0 2.1918798560265801e-01
GL_370 0 NS_370 NS_369 0 -2.1918798560265801e-01
GS_369_11 0 NS_369 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 371/372
CS_371 NS_371 0 9.9999999999999998e-13
CS_372 NS_372 0 9.9999999999999998e-13
RS_371 NS_371 0 7.1523254667023437e+01
RS_372 NS_372 0 7.1523254667023451e+01
GL_371 0 NS_371 NS_372 0 2.0613705597202187e-01
GL_372 0 NS_372 NS_371 0 -2.0613705597202187e-01
GS_371_11 0 NS_371 NA_11 0 1.5251913417194629e+00
*
* Complex pair n. 373/374
CS_373 NS_373 0 9.9999999999999998e-13
CS_374 NS_374 0 9.9999999999999998e-13
RS_373 NS_373 0 3.4487804113693971e+02
RS_374 NS_374 0 3.4487804113693966e+02
GL_373 0 NS_373 NS_374 0 2.0650350471279413e-01
GL_374 0 NS_374 NS_373 0 -2.0650350471279413e-01
GS_373_11 0 NS_373 NA_11 0 1.5251913417194629e+00
*
* Real pole n. 375
CS_375 NS_375 0 9.9999999999999998e-13
RS_375 NS_375 0 3.4256132957802641e+00
GS_375_12 0 NS_375 NA_12 0 1.5251913417194629e+00
*
* Real pole n. 376
CS_376 NS_376 0 9.9999999999999998e-13
RS_376 NS_376 0 8.6582773449483081e+00
GS_376_12 0 NS_376 NA_12 0 1.5251913417194629e+00
*
* Real pole n. 377
CS_377 NS_377 0 9.9999999999999998e-13
RS_377 NS_377 0 3.1453339577953656e+01
GS_377_12 0 NS_377 NA_12 0 1.5251913417194629e+00
*
* Real pole n. 378
CS_378 NS_378 0 9.9999999999999998e-13
RS_378 NS_378 0 1.2483716714088728e+03
GS_378_12 0 NS_378 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 379/380
CS_379 NS_379 0 9.9999999999999998e-13
CS_380 NS_380 0 9.9999999999999998e-13
RS_379 NS_379 0 9.5700292143510275e+00
RS_380 NS_380 0 9.5700292143510275e+00
GL_379 0 NS_379 NS_380 0 1.4040628101439498e-01
GL_380 0 NS_380 NS_379 0 -1.4040628101439498e-01
GS_379_12 0 NS_379 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 381/382
CS_381 NS_381 0 9.9999999999999998e-13
CS_382 NS_382 0 9.9999999999999998e-13
RS_381 NS_381 0 4.0462967855885069e+01
RS_382 NS_382 0 4.0462967855885061e+01
GL_381 0 NS_381 NS_382 0 2.6673201695183885e-01
GL_382 0 NS_382 NS_381 0 -2.6673201695183885e-01
GS_381_12 0 NS_381 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 383/384
CS_383 NS_383 0 9.9999999999999998e-13
CS_384 NS_384 0 9.9999999999999998e-13
RS_383 NS_383 0 1.9059070407967361e+01
RS_384 NS_384 0 1.9059070407967358e+01
GL_383 0 NS_383 NS_384 0 2.4185814461526237e-01
GL_384 0 NS_384 NS_383 0 -2.4185814461526237e-01
GS_383_12 0 NS_383 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 385/386
CS_385 NS_385 0 9.9999999999999998e-13
CS_386 NS_386 0 9.9999999999999998e-13
RS_385 NS_385 0 1.7666316379915560e+01
RS_386 NS_386 0 1.7666316379915564e+01
GL_385 0 NS_385 NS_386 0 1.9702615210896449e-01
GL_386 0 NS_386 NS_385 0 -1.9702615210896449e-01
GS_385_12 0 NS_385 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 387/388
CS_387 NS_387 0 9.9999999999999998e-13
CS_388 NS_388 0 9.9999999999999998e-13
RS_387 NS_387 0 3.4591856087420081e+02
RS_388 NS_388 0 3.4591856087420081e+02
GL_387 0 NS_387 NS_388 0 2.4170685235821462e-01
GL_388 0 NS_388 NS_387 0 -2.4170685235821462e-01
GS_387_12 0 NS_387 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 389/390
CS_389 NS_389 0 9.9999999999999998e-13
CS_390 NS_390 0 9.9999999999999998e-13
RS_389 NS_389 0 3.4257938362763537e+02
RS_390 NS_390 0 3.4257938362763537e+02
GL_389 0 NS_389 NS_390 0 1.4255159266867465e-01
GL_390 0 NS_390 NS_389 0 -1.4255159266867465e-01
GS_389_12 0 NS_389 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 391/392
CS_391 NS_391 0 9.9999999999999998e-13
CS_392 NS_392 0 9.9999999999999998e-13
RS_391 NS_391 0 1.0126954757407573e+02
RS_392 NS_392 0 1.0126954757407573e+02
GL_391 0 NS_391 NS_392 0 1.4356554078688363e-01
GL_392 0 NS_392 NS_391 0 -1.4356554078688363e-01
GS_391_12 0 NS_391 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 393/394
CS_393 NS_393 0 9.9999999999999998e-13
CS_394 NS_394 0 9.9999999999999998e-13
RS_393 NS_393 0 3.5335368091933424e+02
RS_394 NS_394 0 3.5335368091933418e+02
GL_393 0 NS_393 NS_394 0 1.6640381409742028e-01
GL_394 0 NS_394 NS_393 0 -1.6640381409742028e-01
GS_393_12 0 NS_393 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 395/396
CS_395 NS_395 0 9.9999999999999998e-13
CS_396 NS_396 0 9.9999999999999998e-13
RS_395 NS_395 0 1.1172419684791065e+02
RS_396 NS_396 0 1.1172419684791066e+02
GL_395 0 NS_395 NS_396 0 1.6662138407694810e-01
GL_396 0 NS_396 NS_395 0 -1.6662138407694810e-01
GS_395_12 0 NS_395 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 397/398
CS_397 NS_397 0 9.9999999999999998e-13
CS_398 NS_398 0 9.9999999999999998e-13
RS_397 NS_397 0 2.3124949155545121e+02
RS_398 NS_398 0 2.3124949155545121e+02
GL_397 0 NS_397 NS_398 0 1.8384390380970300e-01
GL_398 0 NS_398 NS_397 0 -1.8384390380970300e-01
GS_397_12 0 NS_397 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 399/400
CS_399 NS_399 0 9.9999999999999998e-13
CS_400 NS_400 0 9.9999999999999998e-13
RS_399 NS_399 0 8.6778721170894016e+01
RS_400 NS_400 0 8.6778721170894002e+01
GL_399 0 NS_399 NS_400 0 2.2562932600183958e-01
GL_400 0 NS_400 NS_399 0 -2.2562932600183958e-01
GS_399_12 0 NS_399 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 401/402
CS_401 NS_401 0 9.9999999999999998e-13
CS_402 NS_402 0 9.9999999999999998e-13
RS_401 NS_401 0 3.2996671012988776e+02
RS_402 NS_402 0 3.2996671012988776e+02
GL_401 0 NS_401 NS_402 0 2.2283373301463522e-01
GL_402 0 NS_402 NS_401 0 -2.2283373301463522e-01
GS_401_12 0 NS_401 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 403/404
CS_403 NS_403 0 9.9999999999999998e-13
CS_404 NS_404 0 9.9999999999999998e-13
RS_403 NS_403 0 3.9174610175015977e+02
RS_404 NS_404 0 3.9174610175015977e+02
GL_403 0 NS_403 NS_404 0 2.1918798560265801e-01
GL_404 0 NS_404 NS_403 0 -2.1918798560265801e-01
GS_403_12 0 NS_403 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 405/406
CS_405 NS_405 0 9.9999999999999998e-13
CS_406 NS_406 0 9.9999999999999998e-13
RS_405 NS_405 0 7.1523254667023437e+01
RS_406 NS_406 0 7.1523254667023451e+01
GL_405 0 NS_405 NS_406 0 2.0613705597202187e-01
GL_406 0 NS_406 NS_405 0 -2.0613705597202187e-01
GS_405_12 0 NS_405 NA_12 0 1.5251913417194629e+00
*
* Complex pair n. 407/408
CS_407 NS_407 0 9.9999999999999998e-13
CS_408 NS_408 0 9.9999999999999998e-13
RS_407 NS_407 0 3.4487804113693971e+02
RS_408 NS_408 0 3.4487804113693966e+02
GL_407 0 NS_407 NS_408 0 2.0650350471279413e-01
GL_408 0 NS_408 NS_407 0 -2.0650350471279413e-01
GS_407_12 0 NS_407 NA_12 0 1.5251913417194629e+00
*
******************************


.ends
*******************
* End of subcircuit
*******************
