**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [32 16 160] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_15_PCB_wire_2p0inch_lowloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 -1.5530868320838243e-02
GC_1_2 b_1 NI_1 NS_2 0 6.4872575665921759e-09
GC_1_3 b_1 NI_1 NS_3 0 -1.0780988234711904e-06
GC_1_4 b_1 NI_1 NS_4 0 -2.3175274109547209e-05
GC_1_5 b_1 NI_1 NS_5 0 3.3380760479897011e-04
GC_1_6 b_1 NI_1 NS_6 0 -2.0548502423846943e-04
GC_1_7 b_1 NI_1 NS_7 0 -1.5862582242396779e-03
GC_1_8 b_1 NI_1 NS_8 0 -2.3361772915297539e-03
GC_1_9 b_1 NI_1 NS_9 0 -6.3216355249708312e-05
GC_1_10 b_1 NI_1 NS_10 0 4.3863825431021452e-03
GC_1_11 b_1 NI_1 NS_11 0 1.5399048802873965e-03
GC_1_12 b_1 NI_1 NS_12 0 -5.9456443665761643e-03
GC_1_13 b_1 NI_1 NS_13 0 -4.9710137030512013e-03
GC_1_14 b_1 NI_1 NS_14 0 6.5658943387613905e-03
GC_1_15 b_1 NI_1 NS_15 0 1.1033049601678431e-03
GC_1_16 b_1 NI_1 NS_16 0 -4.8869713796920514e-04
GC_1_17 b_1 NI_1 NS_17 0 2.8351211271457162e-03
GC_1_18 b_1 NI_1 NS_18 0 2.3742295355822000e-03
GC_1_19 b_1 NI_1 NS_19 0 -4.4219508017686055e-03
GC_1_20 b_1 NI_1 NS_20 0 -1.3476668926753999e-02
GC_1_21 b_1 NI_1 NS_21 0 1.7485551924605149e-03
GC_1_22 b_1 NI_1 NS_22 0 1.7702185490222219e-02
GC_1_23 b_1 NI_1 NS_23 0 9.8282594327939506e-03
GC_1_24 b_1 NI_1 NS_24 0 -2.3328386621705678e-03
GC_1_25 b_1 NI_1 NS_25 0 -1.3062251318156934e-02
GC_1_26 b_1 NI_1 NS_26 0 2.3406843805529850e-03
GC_1_27 b_1 NI_1 NS_27 0 9.2233753890635928e-03
GC_1_28 b_1 NI_1 NS_28 0 1.9112827881353725e-03
GC_1_29 b_1 NI_1 NS_29 0 -1.7997095998237785e-02
GC_1_30 b_1 NI_1 NS_30 0 -6.3439019430810931e-03
GC_1_31 b_1 NI_1 NS_31 0 1.5754262105909664e-02
GC_1_32 b_1 NI_1 NS_32 0 6.4095337182158265e-03
GC_1_33 b_1 NI_1 NS_33 0 8.1027183200185933e-03
GC_1_34 b_1 NI_1 NS_34 0 -4.2190611020470909e-03
GC_1_35 b_1 NI_1 NS_35 0 -7.4948915553305255e-03
GC_1_36 b_1 NI_1 NS_36 0 2.0941339334177456e-03
GC_1_37 b_1 NI_1 NS_37 0 6.7044800415873382e-03
GC_1_38 b_1 NI_1 NS_38 0 -2.7628606905911201e-03
GC_1_39 b_1 NI_1 NS_39 0 -6.5432407834931589e-03
GC_1_40 b_1 NI_1 NS_40 0 2.9299446522590418e-03
GC_1_41 b_1 NI_1 NS_41 0 7.6773806179844545e-03
GC_1_42 b_1 NI_1 NS_42 0 4.6375265103133659e-04
GC_1_43 b_1 NI_1 NS_43 0 -9.3401575977007986e-03
GC_1_44 b_1 NI_1 NS_44 0 -5.1079553032413339e-03
GC_1_45 b_1 NI_1 NS_45 0 6.8551899767938839e-03
GC_1_46 b_1 NI_1 NS_46 0 4.0869854575189728e-03
GC_1_47 b_1 NI_1 NS_47 0 -3.8349360358261721e-04
GC_1_48 b_1 NI_1 NS_48 0 -9.2299662211745308e-04
GC_1_49 b_1 NI_1 NS_49 0 5.6963375693309939e-03
GC_1_50 b_1 NI_1 NS_50 0 -1.3852990128853365e-03
GC_1_51 b_1 NI_1 NS_51 0 -9.1011041743308107e-03
GC_1_52 b_1 NI_1 NS_52 0 -1.2296019020133515e-03
GC_1_53 b_1 NI_1 NS_53 0 6.0201772757163541e-03
GC_1_54 b_1 NI_1 NS_54 0 7.1817299147957552e-04
GC_1_55 b_1 NI_1 NS_55 0 -2.6199046907131019e-03
GC_1_56 b_1 NI_1 NS_56 0 2.4600285323131296e-04
GC_1_57 b_1 NI_1 NS_57 0 6.7218299050604150e-03
GC_1_58 b_1 NI_1 NS_58 0 -2.2667453976548519e-03
GC_1_59 b_1 NI_1 NS_59 0 -9.2254204622592706e-03
GC_1_60 b_1 NI_1 NS_60 0 1.5046090677211855e-03
GC_1_61 b_1 NI_1 NS_61 0 5.7525390025044230e-03
GC_1_62 b_1 NI_1 NS_62 0 -1.5177985015858960e-03
GC_1_63 b_1 NI_1 NS_63 0 -3.2852539079676300e-03
GC_1_64 b_1 NI_1 NS_64 0 2.3899132658382464e-03
GC_1_65 b_1 NI_1 NS_65 0 7.2874270495532573e-03
GC_1_66 b_1 NI_1 NS_66 0 -4.1034629640531823e-03
GC_1_67 b_1 NI_1 NS_67 0 -8.5232791386866749e-03
GC_1_68 b_1 NI_1 NS_68 0 4.1574394236145321e-03
GC_1_69 b_1 NI_1 NS_69 0 4.8370647226197933e-03
GC_1_70 b_1 NI_1 NS_70 0 -3.8866667833394701e-03
GC_1_71 b_1 NI_1 NS_71 0 -2.3786687275308563e-03
GC_1_72 b_1 NI_1 NS_72 0 4.7281088504797049e-03
GC_1_73 b_1 NI_1 NS_73 0 7.0803230103499417e-03
GC_1_74 b_1 NI_1 NS_74 0 -7.3558602091558295e-03
GC_1_75 b_1 NI_1 NS_75 0 -7.0931612742462652e-03
GC_1_76 b_1 NI_1 NS_76 0 6.8359962682758889e-03
GC_1_77 b_1 NI_1 NS_77 0 1.6811451238135050e-03
GC_1_78 b_1 NI_1 NS_78 0 -5.3216376516710146e-03
GC_1_79 b_1 NI_1 NS_79 0 5.9853529083191549e-04
GC_1_80 b_1 NI_1 NS_80 0 5.4496392043413486e-03
GC_1_81 b_1 NI_1 NS_81 0 -4.1282353587319472e-09
GC_1_82 b_1 NI_1 NS_82 0 -1.3976314252426336e-08
GC_1_83 b_1 NI_1 NS_83 0 2.7262643674317863e-03
GC_1_84 b_1 NI_1 NS_84 0 -8.5984900355557184e-03
GC_1_85 b_1 NI_1 NS_85 0 8.7601828765636824e-04
GC_1_86 b_1 NI_1 NS_86 0 -3.4431550566540047e-03
GC_1_87 b_1 NI_1 NS_87 0 6.3792143208043345e-04
GC_1_88 b_1 NI_1 NS_88 0 4.0228569547314606e-03
GC_1_89 b_1 NI_1 NS_89 0 2.1875522053167217e-03
GC_1_90 b_1 NI_1 NS_90 0 -8.1664821177311279e-03
GC_1_91 b_1 NI_1 NS_91 0 -3.4772864743811858e-03
GC_1_92 b_1 NI_1 NS_92 0 6.9937177099685536e-03
GC_1_93 b_1 NI_1 NS_93 0 -8.5503727188456809e-08
GC_1_94 b_1 NI_1 NS_94 0 -3.1420283073468535e-07
GC_1_95 b_1 NI_1 NS_95 0 -7.9941562802591133e-03
GC_1_96 b_1 NI_1 NS_96 0 5.3784297957891530e-03
GC_1_97 b_1 NI_1 NS_97 0 4.1818213559482662e-03
GC_1_98 b_1 NI_1 NS_98 0 -6.8548439330208032e-03
GC_1_99 b_1 NI_1 NS_99 0 5.3337133193831028e-03
GC_1_100 b_1 NI_1 NS_100 0 7.4258455792823932e-04
GC_1_101 b_1 NI_1 NS_101 0 -2.3535039763461197e-03
GC_1_102 b_1 NI_1 NS_102 0 6.8399075503825088e-03
GC_1_103 b_1 NI_1 NS_103 0 -1.4841908740739218e-03
GC_1_104 b_1 NI_1 NS_104 0 -4.2255112512419053e-03
GC_1_105 b_1 NI_1 NS_105 0 2.3638870734323035e-03
GC_1_106 b_1 NI_1 NS_106 0 5.0284973543175621e-03
GC_1_107 b_1 NI_1 NS_107 0 -1.9828423531963631e-03
GC_1_108 b_1 NI_1 NS_108 0 -8.9598437406871855e-03
GC_1_109 b_1 NI_1 NS_109 0 -1.1185495614699415e-02
GC_1_110 b_1 NI_1 NS_110 0 8.4594985314924632e-09
GC_1_111 b_1 NI_1 NS_111 0 9.8721878574552315e-07
GC_1_112 b_1 NI_1 NS_112 0 3.6199507015198418e-05
GC_1_113 b_1 NI_1 NS_113 0 4.3663018799460314e-03
GC_1_114 b_1 NI_1 NS_114 0 -3.4896621214979850e-03
GC_1_115 b_1 NI_1 NS_115 0 -3.7149213676674854e-03
GC_1_116 b_1 NI_1 NS_116 0 6.2509196129706714e-03
GC_1_117 b_1 NI_1 NS_117 0 -8.7863564569121231e-03
GC_1_118 b_1 NI_1 NS_118 0 -5.9490008506655860e-03
GC_1_119 b_1 NI_1 NS_119 0 9.1761685703224041e-03
GC_1_120 b_1 NI_1 NS_120 0 -5.9808724636429634e-03
GC_1_121 b_1 NI_1 NS_121 0 7.1653427149210242e-03
GC_1_122 b_1 NI_1 NS_122 0 1.1911619516633998e-02
GC_1_123 b_1 NI_1 NS_123 0 -4.2323502246248085e-03
GC_1_124 b_1 NI_1 NS_124 0 -1.1251731311410942e-03
GC_1_125 b_1 NI_1 NS_125 0 -8.8793814729324506e-03
GC_1_126 b_1 NI_1 NS_126 0 -4.5103774349622287e-04
GC_1_127 b_1 NI_1 NS_127 0 1.4527713310507191e-02
GC_1_128 b_1 NI_1 NS_128 0 -1.0355588691760466e-02
GC_1_129 b_1 NI_1 NS_129 0 1.6511395596738761e-02
GC_1_130 b_1 NI_1 NS_130 0 4.0489387043224747e-03
GC_1_131 b_1 NI_1 NS_131 0 -1.1485124336039657e-02
GC_1_132 b_1 NI_1 NS_132 0 -1.9361413256017900e-04
GC_1_133 b_1 NI_1 NS_133 0 -1.6607752081580419e-02
GC_1_134 b_1 NI_1 NS_134 0 -4.4552719964303947e-02
GC_1_135 b_1 NI_1 NS_135 0 1.0667471159289860e-02
GC_1_136 b_1 NI_1 NS_136 0 1.0870824200981976e-03
GC_1_137 b_1 NI_1 NS_137 0 -4.8262935568841779e-02
GC_1_138 b_1 NI_1 NS_138 0 1.1004758939664946e-02
GC_1_139 b_1 NI_1 NS_139 0 -1.0464750686436750e-02
GC_1_140 b_1 NI_1 NS_140 0 5.4279500905995829e-04
GC_1_141 b_1 NI_1 NS_141 0 9.7653630224749845e-03
GC_1_142 b_1 NI_1 NS_142 0 -6.1129099939059861e-04
GC_1_143 b_1 NI_1 NS_143 0 4.5934330574465667e-03
GC_1_144 b_1 NI_1 NS_144 0 2.4194429108418045e-02
GC_1_145 b_1 NI_1 NS_145 0 -1.0736736005889072e-02
GC_1_146 b_1 NI_1 NS_146 0 1.9986342864633717e-03
GC_1_147 b_1 NI_1 NS_147 0 -8.4713022982081110e-03
GC_1_148 b_1 NI_1 NS_148 0 -1.3526361329873744e-02
GC_1_149 b_1 NI_1 NS_149 0 1.0155212753688383e-02
GC_1_150 b_1 NI_1 NS_150 0 9.6273264187683358e-04
GC_1_151 b_1 NI_1 NS_151 0 -1.9169421790722910e-02
GC_1_152 b_1 NI_1 NS_152 0 2.8673863620290875e-02
GC_1_153 b_1 NI_1 NS_153 0 -9.6256415308615742e-03
GC_1_154 b_1 NI_1 NS_154 0 -9.4348281783413900e-04
GC_1_155 b_1 NI_1 NS_155 0 1.8844348159612382e-03
GC_1_156 b_1 NI_1 NS_156 0 -1.3764795551416162e-03
GC_1_157 b_1 NI_1 NS_157 0 9.4635462038030783e-03
GC_1_158 b_1 NI_1 NS_158 0 -2.5486095653160916e-04
GC_1_159 b_1 NI_1 NS_159 0 -1.6535192238852274e-04
GC_1_160 b_1 NI_1 NS_160 0 3.0293306931723211e-02
GC_1_161 b_1 NI_1 NS_161 0 -8.5338138707214319e-03
GC_1_162 b_1 NI_1 NS_162 0 1.7750635776358370e-04
GC_1_163 b_1 NI_1 NS_163 0 2.1345417843923240e-04
GC_1_164 b_1 NI_1 NS_164 0 -5.4660289948873907e-03
GC_1_165 b_1 NI_1 NS_165 0 1.0030295563258294e-02
GC_1_166 b_1 NI_1 NS_166 0 -3.4496677366391461e-04
GC_1_167 b_1 NI_1 NS_167 0 8.9347318283640609e-03
GC_1_168 b_1 NI_1 NS_168 0 2.6406163893342806e-02
GC_1_169 b_1 NI_1 NS_169 0 -8.3546165129830003e-03
GC_1_170 b_1 NI_1 NS_170 0 1.4014782426117504e-03
GC_1_171 b_1 NI_1 NS_171 0 -2.5783437829380155e-03
GC_1_172 b_1 NI_1 NS_172 0 -7.3352780822781840e-03
GC_1_173 b_1 NI_1 NS_173 0 1.0543947028944893e-02
GC_1_174 b_1 NI_1 NS_174 0 -8.2792607460328448e-04
GC_1_175 b_1 NI_1 NS_175 0 1.4465695980430154e-02
GC_1_176 b_1 NI_1 NS_176 0 1.9992681054547944e-02
GC_1_177 b_1 NI_1 NS_177 0 -8.2668415347023697e-03
GC_1_178 b_1 NI_1 NS_178 0 2.9582407908293790e-03
GC_1_179 b_1 NI_1 NS_179 0 -5.5757286531069620e-03
GC_1_180 b_1 NI_1 NS_180 0 -6.9085960741767285e-03
GC_1_181 b_1 NI_1 NS_181 0 1.1230556732160281e-02
GC_1_182 b_1 NI_1 NS_182 0 -1.3725284458290360e-03
GC_1_183 b_1 NI_1 NS_183 0 1.5750291698828071e-02
GC_1_184 b_1 NI_1 NS_184 0 1.2967900121577171e-02
GC_1_185 b_1 NI_1 NS_185 0 -7.1659122868756022e-03
GC_1_186 b_1 NI_1 NS_186 0 5.1305973072879934e-03
GC_1_187 b_1 NI_1 NS_187 0 -6.8667080635905894e-03
GC_1_188 b_1 NI_1 NS_188 0 -4.8393413396225380e-03
GC_1_189 b_1 NI_1 NS_189 0 5.3089322140956139e-09
GC_1_190 b_1 NI_1 NS_190 0 4.4273821506169640e-08
GC_1_191 b_1 NI_1 NS_191 0 1.2002193839018226e-02
GC_1_192 b_1 NI_1 NS_192 0 -2.5686804852326946e-03
GC_1_193 b_1 NI_1 NS_193 0 -5.2367617774666036e-03
GC_1_194 b_1 NI_1 NS_194 0 4.7118170466739729e-03
GC_1_195 b_1 NI_1 NS_195 0 -6.1526719493275187e-03
GC_1_196 b_1 NI_1 NS_196 0 -4.3194220595839375e-03
GC_1_197 b_1 NI_1 NS_197 0 1.1768583380166451e-02
GC_1_198 b_1 NI_1 NS_198 0 -3.7146184684677531e-03
GC_1_199 b_1 NI_1 NS_199 0 1.3012626394160634e-02
GC_1_200 b_1 NI_1 NS_200 0 9.4653980218875437e-03
GC_1_201 b_1 NI_1 NS_201 0 3.9556714058173220e-06
GC_1_202 b_1 NI_1 NS_202 0 -9.4250490833158713e-07
GC_1_203 b_1 NI_1 NS_203 0 1.6124340760127556e-02
GC_1_204 b_1 NI_1 NS_204 0 1.6774826305275950e-02
GC_1_205 b_1 NI_1 NS_205 0 1.2055184277835789e-02
GC_1_206 b_1 NI_1 NS_206 0 -2.4727536272118817e-03
GC_1_207 b_1 NI_1 NS_207 0 -8.3469685278654195e-03
GC_1_208 b_1 NI_1 NS_208 0 8.5427575741755114e-05
GC_1_209 b_1 NI_1 NS_209 0 1.1349985592678913e-02
GC_1_210 b_1 NI_1 NS_210 0 7.3343055724884518e-03
GC_1_211 b_1 NI_1 NS_211 0 -4.6479092981493398e-03
GC_1_212 b_1 NI_1 NS_212 0 7.3635995051594128e-03
GC_1_213 b_1 NI_1 NS_213 0 -8.0750686747775059e-03
GC_1_214 b_1 NI_1 NS_214 0 -3.7254234632548367e-03
GC_1_215 b_1 NI_1 NS_215 0 1.5991408214089314e-02
GC_1_216 b_1 NI_1 NS_216 0 -7.7330117492573425e-03
GC_1_217 b_1 NI_1 NS_217 0 1.1804733745049464e-03
GC_1_218 b_1 NI_1 NS_218 0 -3.5559930485178238e-09
GC_1_219 b_1 NI_1 NS_219 0 -4.8002576637136509e-08
GC_1_220 b_1 NI_1 NS_220 0 -3.4752160399439619e-06
GC_1_221 b_1 NI_1 NS_221 0 -3.6812594757275628e-04
GC_1_222 b_1 NI_1 NS_222 0 1.3598225816639000e-04
GC_1_223 b_1 NI_1 NS_223 0 1.1297229767084471e-03
GC_1_224 b_1 NI_1 NS_224 0 1.9432473214890582e-03
GC_1_225 b_1 NI_1 NS_225 0 -6.5058842661985843e-05
GC_1_226 b_1 NI_1 NS_226 0 -3.4937471195339541e-03
GC_1_227 b_1 NI_1 NS_227 0 -1.5644007735436589e-03
GC_1_228 b_1 NI_1 NS_228 0 5.0906039829275102e-03
GC_1_229 b_1 NI_1 NS_229 0 4.2533992673209750e-03
GC_1_230 b_1 NI_1 NS_230 0 -4.9938033603221530e-03
GC_1_231 b_1 NI_1 NS_231 0 -1.0085547515915304e-03
GC_1_232 b_1 NI_1 NS_232 0 5.6397878144831700e-04
GC_1_233 b_1 NI_1 NS_233 0 -2.0807515163003471e-03
GC_1_234 b_1 NI_1 NS_234 0 -1.8633117440015107e-03
GC_1_235 b_1 NI_1 NS_235 0 3.6454397795403167e-03
GC_1_236 b_1 NI_1 NS_236 0 1.1647366929176957e-02
GC_1_237 b_1 NI_1 NS_237 0 -8.9814148338303388e-04
GC_1_238 b_1 NI_1 NS_238 0 -1.4854322540288489e-02
GC_1_239 b_1 NI_1 NS_239 0 -8.1235361417816496e-03
GC_1_240 b_1 NI_1 NS_240 0 1.9196061451794422e-03
GC_1_241 b_1 NI_1 NS_241 0 1.1263056429606252e-02
GC_1_242 b_1 NI_1 NS_242 0 -1.8122318450235300e-03
GC_1_243 b_1 NI_1 NS_243 0 -7.5672718808769040e-03
GC_1_244 b_1 NI_1 NS_244 0 -1.6811818298721004e-03
GC_1_245 b_1 NI_1 NS_245 0 1.5281711114847187e-02
GC_1_246 b_1 NI_1 NS_246 0 5.3008448916442436e-03
GC_1_247 b_1 NI_1 NS_247 0 -1.3082856900665159e-02
GC_1_248 b_1 NI_1 NS_248 0 -5.4612973817835704e-03
GC_1_249 b_1 NI_1 NS_249 0 -6.6370717900765160e-03
GC_1_250 b_1 NI_1 NS_250 0 3.4566939005134067e-03
GC_1_251 b_1 NI_1 NS_251 0 6.3616039747960516e-03
GC_1_252 b_1 NI_1 NS_252 0 -1.8793243513729383e-03
GC_1_253 b_1 NI_1 NS_253 0 -5.4737176493986966e-03
GC_1_254 b_1 NI_1 NS_254 0 2.1830271446640101e-03
GC_1_255 b_1 NI_1 NS_255 0 5.3937683821950614e-03
GC_1_256 b_1 NI_1 NS_256 0 -2.6324374313278702e-03
GC_1_257 b_1 NI_1 NS_257 0 -6.3064546623561903e-03
GC_1_258 b_1 NI_1 NS_258 0 -4.8381472945087140e-04
GC_1_259 b_1 NI_1 NS_259 0 7.6452800881850677e-03
GC_1_260 b_1 NI_1 NS_260 0 3.6298731666400646e-03
GC_1_261 b_1 NI_1 NS_261 0 -5.8336241539701213e-03
GC_1_262 b_1 NI_1 NS_262 0 -3.4645948161415611e-03
GC_1_263 b_1 NI_1 NS_263 0 2.9620036015146848e-04
GC_1_264 b_1 NI_1 NS_264 0 5.5810466178821355e-04
GC_1_265 b_1 NI_1 NS_265 0 -4.9270628226813070e-03
GC_1_266 b_1 NI_1 NS_266 0 8.9219828341239921e-04
GC_1_267 b_1 NI_1 NS_267 0 6.2063416474648731e-03
GC_1_268 b_1 NI_1 NS_268 0 6.8827499107644216e-04
GC_1_269 b_1 NI_1 NS_269 0 -5.3209621295614677e-03
GC_1_270 b_1 NI_1 NS_270 0 -4.8418936150818444e-04
GC_1_271 b_1 NI_1 NS_271 0 1.5503327192988130e-03
GC_1_272 b_1 NI_1 NS_272 0 -4.3207881492277861e-05
GC_1_273 b_1 NI_1 NS_273 0 -6.0223328276230517e-03
GC_1_274 b_1 NI_1 NS_274 0 1.9232412392108302e-03
GC_1_275 b_1 NI_1 NS_275 0 6.2616666873382427e-03
GC_1_276 b_1 NI_1 NS_276 0 2.1736210789949600e-04
GC_1_277 b_1 NI_1 NS_277 0 -5.0591984903880808e-03
GC_1_278 b_1 NI_1 NS_278 0 1.7016163938226461e-03
GC_1_279 b_1 NI_1 NS_279 0 2.4884732765862003e-03
GC_1_280 b_1 NI_1 NS_280 0 -9.5765139707198153e-04
GC_1_281 b_1 NI_1 NS_281 0 -6.5329629510427513e-03
GC_1_282 b_1 NI_1 NS_282 0 3.8846376443299195e-03
GC_1_283 b_1 NI_1 NS_283 0 7.4932677132106915e-03
GC_1_284 b_1 NI_1 NS_284 0 -1.0960274181880257e-03
GC_1_285 b_1 NI_1 NS_285 0 -3.9851190199831433e-03
GC_1_286 b_1 NI_1 NS_286 0 4.0409800028668062e-03
GC_1_287 b_1 NI_1 NS_287 0 2.8633260163856747e-03
GC_1_288 b_1 NI_1 NS_288 0 -3.0534889789912601e-03
GC_1_289 b_1 NI_1 NS_289 0 -6.0227292275259279e-03
GC_1_290 b_1 NI_1 NS_290 0 7.2373892460004278e-03
GC_1_291 b_1 NI_1 NS_291 0 7.9897111890509329e-03
GC_1_292 b_1 NI_1 NS_292 0 -4.8114595196128854e-03
GC_1_293 b_1 NI_1 NS_293 0 -5.3741900546798915e-04
GC_1_294 b_1 NI_1 NS_294 0 5.0204728210163059e-03
GC_1_295 b_1 NI_1 NS_295 0 2.4825551854831666e-04
GC_1_296 b_1 NI_1 NS_296 0 -4.7581976244320361e-03
GC_1_297 b_1 NI_1 NS_297 0 1.8109240231550959e-09
GC_1_298 b_1 NI_1 NS_298 0 3.2744953923182652e-09
GC_1_299 b_1 NI_1 NS_299 0 -1.4271962547646496e-03
GC_1_300 b_1 NI_1 NS_300 0 7.8707399680795799e-03
GC_1_301 b_1 NI_1 NS_301 0 -1.7997930773597581e-04
GC_1_302 b_1 NI_1 NS_302 0 3.0272441090316983e-03
GC_1_303 b_1 NI_1 NS_303 0 -1.3038553838673966e-04
GC_1_304 b_1 NI_1 NS_304 0 -3.3753037112221030e-03
GC_1_305 b_1 NI_1 NS_305 0 -8.7631252230381095e-04
GC_1_306 b_1 NI_1 NS_306 0 7.5304828374334011e-03
GC_1_307 b_1 NI_1 NS_307 0 3.7888078333932545e-03
GC_1_308 b_1 NI_1 NS_308 0 -6.1574210772036677e-03
GC_1_309 b_1 NI_1 NS_309 0 8.6236228961298154e-08
GC_1_310 b_1 NI_1 NS_310 0 -3.5294047735957657e-07
GC_1_311 b_1 NI_1 NS_311 0 6.7186801411306118e-03
GC_1_312 b_1 NI_1 NS_312 0 -5.3194116322398920e-03
GC_1_313 b_1 NI_1 NS_313 0 -2.6111716281401859e-03
GC_1_314 b_1 NI_1 NS_314 0 6.0542407326549530e-03
GC_1_315 b_1 NI_1 NS_315 0 -4.2922714918651019e-03
GC_1_316 b_1 NI_1 NS_316 0 1.4429424497219179e-05
GC_1_317 b_1 NI_1 NS_317 0 2.7173890707778872e-03
GC_1_318 b_1 NI_1 NS_318 0 -6.2040229563888119e-03
GC_1_319 b_1 NI_1 NS_319 0 2.0957200636999899e-03
GC_1_320 b_1 NI_1 NS_320 0 3.2562724999328769e-03
GC_1_321 b_1 NI_1 NS_321 0 -1.9700344229512056e-03
GC_1_322 b_1 NI_1 NS_322 0 -4.4205369357727051e-03
GC_1_323 b_1 NI_1 NS_323 0 2.8640861854579832e-03
GC_1_324 b_1 NI_1 NS_324 0 8.0083630618385405e-03
GC_1_325 b_1 NI_1 NS_325 0 -3.3036180970061630e-03
GC_1_326 b_1 NI_1 NS_326 0 1.8493832823042814e-09
GC_1_327 b_1 NI_1 NS_327 0 5.6032189490553142e-08
GC_1_328 b_1 NI_1 NS_328 0 1.8929692725188575e-06
GC_1_329 b_1 NI_1 NS_329 0 -9.1167737507262552e-05
GC_1_330 b_1 NI_1 NS_330 0 -5.7737685755106589e-05
GC_1_331 b_1 NI_1 NS_331 0 -1.2657732161165509e-03
GC_1_332 b_1 NI_1 NS_332 0 -2.9559335222127485e-04
GC_1_333 b_1 NI_1 NS_333 0 -1.6792127366473328e-03
GC_1_334 b_1 NI_1 NS_334 0 2.6464981006143404e-03
GC_1_335 b_1 NI_1 NS_335 0 5.1121264532543831e-04
GC_1_336 b_1 NI_1 NS_336 0 5.4276095823366883e-03
GC_1_337 b_1 NI_1 NS_337 0 7.1034902512452829e-03
GC_1_338 b_1 NI_1 NS_338 0 6.3629125422538530e-04
GC_1_339 b_1 NI_1 NS_339 0 6.4433103890677032e-04
GC_1_340 b_1 NI_1 NS_340 0 -6.6091960340223046e-04
GC_1_341 b_1 NI_1 NS_341 0 1.0576976596943556e-03
GC_1_342 b_1 NI_1 NS_342 0 1.5711389936581806e-03
GC_1_343 b_1 NI_1 NS_343 0 1.2687515823413766e-02
GC_1_344 b_1 NI_1 NS_344 0 1.3123211174097885e-02
GC_1_345 b_1 NI_1 NS_345 0 8.7187952794639690e-03
GC_1_346 b_1 NI_1 NS_346 0 -2.0392082089599209e-02
GC_1_347 b_1 NI_1 NS_347 0 8.3891008500467240e-03
GC_1_348 b_1 NI_1 NS_348 0 -2.9045265237153104e-03
GC_1_349 b_1 NI_1 NS_349 0 -1.2701292149288671e-02
GC_1_350 b_1 NI_1 NS_350 0 -3.8806700451772272e-02
GC_1_351 b_1 NI_1 NS_351 0 -7.2523394833819413e-03
GC_1_352 b_1 NI_1 NS_352 0 -2.1332749821331193e-03
GC_1_353 b_1 NI_1 NS_353 0 -5.2307202159103720e-02
GC_1_354 b_1 NI_1 NS_354 0 -1.7936179688050891e-03
GC_1_355 b_1 NI_1 NS_355 0 1.4914415692729588e-02
GC_1_356 b_1 NI_1 NS_356 0 8.6735776565941818e-03
GC_1_357 b_1 NI_1 NS_357 0 -5.9233536256804520e-03
GC_1_358 b_1 NI_1 NS_358 0 5.0044967075035304e-03
GC_1_359 b_1 NI_1 NS_359 0 8.3724176331088241e-03
GC_1_360 b_1 NI_1 NS_360 0 1.1688364625441145e-02
GC_1_361 b_1 NI_1 NS_361 0 4.5592636104997064e-03
GC_1_362 b_1 NI_1 NS_362 0 -2.9327401719611169e-03
GC_1_363 b_1 NI_1 NS_363 0 -7.8986725967775898e-03
GC_1_364 b_1 NI_1 NS_364 0 -8.1490644575003997e-03
GC_1_365 b_1 NI_1 NS_365 0 -5.6808136133521380e-03
GC_1_366 b_1 NI_1 NS_366 0 -6.1281014119028861e-04
GC_1_367 b_1 NI_1 NS_367 0 -1.8070849967427711e-02
GC_1_368 b_1 NI_1 NS_368 0 1.3578963955423523e-02
GC_1_369 b_1 NI_1 NS_369 0 4.7069862003012121e-03
GC_1_370 b_1 NI_1 NS_370 0 4.3794387117467972e-03
GC_1_371 b_1 NI_1 NS_371 0 6.5015855106825436e-04
GC_1_372 b_1 NI_1 NS_372 0 -1.0995439862358935e-04
GC_1_373 b_1 NI_1 NS_373 0 -3.7963997069979001e-03
GC_1_374 b_1 NI_1 NS_374 0 8.8498808111762170e-04
GC_1_375 b_1 NI_1 NS_375 0 -1.1178294264516547e-03
GC_1_376 b_1 NI_1 NS_376 0 1.6699687298610138e-02
GC_1_377 b_1 NI_1 NS_377 0 4.4472802791198692e-03
GC_1_378 b_1 NI_1 NS_378 0 7.0796476542593016e-04
GC_1_379 b_1 NI_1 NS_379 0 -5.1995788484028973e-04
GC_1_380 b_1 NI_1 NS_380 0 -2.2477510619071791e-03
GC_1_381 b_1 NI_1 NS_381 0 -4.9864554978103744e-03
GC_1_382 b_1 NI_1 NS_382 0 2.1108871156513566e-03
GC_1_383 b_1 NI_1 NS_383 0 7.3425260061966155e-03
GC_1_384 b_1 NI_1 NS_384 0 1.4345854400172163e-02
GC_1_385 b_1 NI_1 NS_385 0 4.1872272047987135e-03
GC_1_386 b_1 NI_1 NS_386 0 -1.6838581706049060e-03
GC_1_387 b_1 NI_1 NS_387 0 -3.3981246702574270e-03
GC_1_388 b_1 NI_1 NS_388 0 -2.1006230765289861e-03
GC_1_389 b_1 NI_1 NS_389 0 -5.4204251691831132e-03
GC_1_390 b_1 NI_1 NS_390 0 4.3817243703984732e-03
GC_1_391 b_1 NI_1 NS_391 0 1.3196871817556671e-02
GC_1_392 b_1 NI_1 NS_392 0 8.4333056515530601e-03
GC_1_393 b_1 NI_1 NS_393 0 2.8324335572192925e-03
GC_1_394 b_1 NI_1 NS_394 0 -4.1306068389809075e-03
GC_1_395 b_1 NI_1 NS_395 0 -5.3207874912403665e-03
GC_1_396 b_1 NI_1 NS_396 0 1.1381584327498882e-03
GC_1_397 b_1 NI_1 NS_397 0 -4.4310212147721613e-03
GC_1_398 b_1 NI_1 NS_398 0 8.3104301777177716e-03
GC_1_399 b_1 NI_1 NS_399 0 1.4612784269093021e-02
GC_1_400 b_1 NI_1 NS_400 0 -4.6824610784193819e-04
GC_1_401 b_1 NI_1 NS_401 0 -1.1845326137263396e-03
GC_1_402 b_1 NI_1 NS_402 0 -4.5473896403316902e-03
GC_1_403 b_1 NI_1 NS_403 0 -2.2825677872358348e-03
GC_1_404 b_1 NI_1 NS_404 0 4.3832552638568200e-03
GC_1_405 b_1 NI_1 NS_405 0 1.3569666870060944e-10
GC_1_406 b_1 NI_1 NS_406 0 -1.5466154844224288e-09
GC_1_407 b_1 NI_1 NS_407 0 1.4460253040254922e-03
GC_1_408 b_1 NI_1 NS_408 0 8.2165469656936378e-03
GC_1_409 b_1 NI_1 NS_409 0 -8.7895049051729126e-04
GC_1_410 b_1 NI_1 NS_410 0 -2.2072123281508820e-03
GC_1_411 b_1 NI_1 NS_411 0 -1.4679135720377459e-03
GC_1_412 b_1 NI_1 NS_412 0 2.7519863067537076e-03
GC_1_413 b_1 NI_1 NS_413 0 1.7320139993817166e-03
GC_1_414 b_1 NI_1 NS_414 0 7.6059327053470934e-03
GC_1_415 b_1 NI_1 NS_415 0 7.5874085871717612e-03
GC_1_416 b_1 NI_1 NS_416 0 -3.8276817774250647e-03
GC_1_417 b_1 NI_1 NS_417 0 -5.2100997192587115e-08
GC_1_418 b_1 NI_1 NS_418 0 -2.0817378738744386e-08
GC_1_419 b_1 NI_1 NS_419 0 1.1391243329432347e-02
GC_1_420 b_1 NI_1 NS_420 0 4.4700330913975492e-03
GC_1_421 b_1 NI_1 NS_421 0 -8.6185050907439315e-04
GC_1_422 b_1 NI_1 NS_422 0 6.4916225478167267e-03
GC_1_423 b_1 NI_1 NS_423 0 3.6263738388922751e-03
GC_1_424 b_1 NI_1 NS_424 0 4.0710469182203346e-04
GC_1_425 b_1 NI_1 NS_425 0 6.0525110463776222e-03
GC_1_426 b_1 NI_1 NS_426 0 -4.6635397551543318e-03
GC_1_427 b_1 NI_1 NS_427 0 -3.3929751263156800e-03
GC_1_428 b_1 NI_1 NS_428 0 -1.3533957775770016e-03
GC_1_429 b_1 NI_1 NS_429 0 1.1237978222521250e-04
GC_1_430 b_1 NI_1 NS_430 0 4.4958002947645768e-03
GC_1_431 b_1 NI_1 NS_431 0 7.2795568486024665e-03
GC_1_432 b_1 NI_1 NS_432 0 5.5305047819474576e-03
GC_1_433 b_1 NI_1 NS_433 0 -5.4772840353252395e-05
GC_1_434 b_1 NI_1 NS_434 0 -6.9629493660689059e-12
GC_1_435 b_1 NI_1 NS_435 0 -2.0817913073277382e-10
GC_1_436 b_1 NI_1 NS_436 0 9.8206142046700071e-09
GC_1_437 b_1 NI_1 NS_437 0 5.4129955292066444e-07
GC_1_438 b_1 NI_1 NS_438 0 4.9187588029370276e-08
GC_1_439 b_1 NI_1 NS_439 0 2.9069067458616369e-06
GC_1_440 b_1 NI_1 NS_440 0 -1.4984891738552250e-06
GC_1_441 b_1 NI_1 NS_441 0 -3.1925349829530730e-06
GC_1_442 b_1 NI_1 NS_442 0 -2.5905348778030764e-06
GC_1_443 b_1 NI_1 NS_443 0 4.5917106882760407e-06
GC_1_444 b_1 NI_1 NS_444 0 -3.9820007571934454e-07
GC_1_445 b_1 NI_1 NS_445 0 -7.4318681196242337e-06
GC_1_446 b_1 NI_1 NS_446 0 -7.4641162171818488e-06
GC_1_447 b_1 NI_1 NS_447 0 -2.5846965145825013e-07
GC_1_448 b_1 NI_1 NS_448 0 -1.3549726256211494e-06
GC_1_449 b_1 NI_1 NS_449 0 -5.8670258840623926e-06
GC_1_450 b_1 NI_1 NS_450 0 2.4876411449981935e-06
GC_1_451 b_1 NI_1 NS_451 0 5.2138885635375731e-06
GC_1_452 b_1 NI_1 NS_452 0 -5.0558572957784690e-06
GC_1_453 b_1 NI_1 NS_453 0 -1.6625735785244108e-05
GC_1_454 b_1 NI_1 NS_454 0 5.0766173677375648e-06
GC_1_455 b_1 NI_1 NS_455 0 -1.1389054013052338e-06
GC_1_456 b_1 NI_1 NS_456 0 7.5150225455479287e-06
GC_1_457 b_1 NI_1 NS_457 0 -6.5962450746383150e-06
GC_1_458 b_1 NI_1 NS_458 0 -4.0226074186359979e-06
GC_1_459 b_1 NI_1 NS_459 0 -3.2518604166616544e-06
GC_1_460 b_1 NI_1 NS_460 0 8.3354887816037049e-06
GC_1_461 b_1 NI_1 NS_461 0 -1.2792488618460939e-06
GC_1_462 b_1 NI_1 NS_462 0 -4.0909172896885417e-06
GC_1_463 b_1 NI_1 NS_463 0 -3.9771513962304930e-06
GC_1_464 b_1 NI_1 NS_464 0 1.1475667014148861e-05
GC_1_465 b_1 NI_1 NS_465 0 -1.4782030867609544e-08
GC_1_466 b_1 NI_1 NS_466 0 7.6669268298814251e-06
GC_1_467 b_1 NI_1 NS_467 0 -3.6189376815193057e-06
GC_1_468 b_1 NI_1 NS_468 0 1.4618091075125581e-06
GC_1_469 b_1 NI_1 NS_469 0 -3.4651561561141648e-07
GC_1_470 b_1 NI_1 NS_470 0 8.4080178673610159e-06
GC_1_471 b_1 NI_1 NS_471 0 -5.5944437275723413e-07
GC_1_472 b_1 NI_1 NS_472 0 2.1381467042673498e-06
GC_1_473 b_1 NI_1 NS_473 0 -2.2883709878372640e-06
GC_1_474 b_1 NI_1 NS_474 0 8.4915537092422419e-06
GC_1_475 b_1 NI_1 NS_475 0 7.3273065644404286e-07
GC_1_476 b_1 NI_1 NS_476 0 9.9252259814584731e-06
GC_1_477 b_1 NI_1 NS_477 0 -7.0096485539198338e-07
GC_1_478 b_1 NI_1 NS_478 0 8.9537433388867552e-06
GC_1_479 b_1 NI_1 NS_479 0 -1.2260743868631067e-06
GC_1_480 b_1 NI_1 NS_480 0 4.0765952034157057e-06
GC_1_481 b_1 NI_1 NS_481 0 1.3021507699096236e-06
GC_1_482 b_1 NI_1 NS_482 0 1.2333188024695548e-05
GC_1_483 b_1 NI_1 NS_483 0 1.8798613691079439e-05
GC_1_484 b_1 NI_1 NS_484 0 1.7017274528297146e-05
GC_1_485 b_1 NI_1 NS_485 0 5.0479536326908199e-06
GC_1_486 b_1 NI_1 NS_486 0 7.8839364786011346e-06
GC_1_487 b_1 NI_1 NS_487 0 1.0389989159431335e-05
GC_1_488 b_1 NI_1 NS_488 0 3.8923637340305840e-06
GC_1_489 b_1 NI_1 NS_489 0 6.8759108838637096e-06
GC_1_490 b_1 NI_1 NS_490 0 1.1069323299168399e-05
GC_1_491 b_1 NI_1 NS_491 0 3.3658577748727632e-05
GC_1_492 b_1 NI_1 NS_492 0 -6.2040451214914010e-06
GC_1_493 b_1 NI_1 NS_493 0 8.2351360411225469e-06
GC_1_494 b_1 NI_1 NS_494 0 3.4806556416421720e-06
GC_1_495 b_1 NI_1 NS_495 0 1.2053460491717584e-05
GC_1_496 b_1 NI_1 NS_496 0 -1.0358836552357092e-05
GC_1_497 b_1 NI_1 NS_497 0 1.0858559158242454e-05
GC_1_498 b_1 NI_1 NS_498 0 6.5736101397806447e-06
GC_1_499 b_1 NI_1 NS_499 0 1.7121023107778326e-05
GC_1_500 b_1 NI_1 NS_500 0 -3.0993300016099915e-05
GC_1_501 b_1 NI_1 NS_501 0 8.1831185883472392e-06
GC_1_502 b_1 NI_1 NS_502 0 -2.9223709966197651e-06
GC_1_503 b_1 NI_1 NS_503 0 -3.1852000490213911e-06
GC_1_504 b_1 NI_1 NS_504 0 -1.6372769537781413e-05
GC_1_505 b_1 NI_1 NS_505 0 1.1876730430073047e-05
GC_1_506 b_1 NI_1 NS_506 0 -1.5556620866584189e-06
GC_1_507 b_1 NI_1 NS_507 0 -1.2637533144655237e-05
GC_1_508 b_1 NI_1 NS_508 0 -2.5277365582997518e-05
GC_1_509 b_1 NI_1 NS_509 0 -1.0768097498238817e-07
GC_1_510 b_1 NI_1 NS_510 0 -6.6428261759649856e-06
GC_1_511 b_1 NI_1 NS_511 0 -9.5779958853537360e-06
GC_1_512 b_1 NI_1 NS_512 0 -2.6885576400152161e-06
GC_1_513 b_1 NI_1 NS_513 0 1.0207142841859829e-10
GC_1_514 b_1 NI_1 NS_514 0 4.5675821797114163e-11
GC_1_515 b_1 NI_1 NS_515 0 1.5500864030618115e-06
GC_1_516 b_1 NI_1 NS_516 0 -4.7010659178518667e-06
GC_1_517 b_1 NI_1 NS_517 0 -1.3389449281339345e-06
GC_1_518 b_1 NI_1 NS_518 0 -1.3668614643132152e-06
GC_1_519 b_1 NI_1 NS_519 0 -4.8399314334380905e-06
GC_1_520 b_1 NI_1 NS_520 0 -1.0276602184978542e-06
GC_1_521 b_1 NI_1 NS_521 0 -1.0646411062857677e-06
GC_1_522 b_1 NI_1 NS_522 0 -2.7378264897269780e-06
GC_1_523 b_1 NI_1 NS_523 0 -9.9890614961940441e-06
GC_1_524 b_1 NI_1 NS_524 0 -4.1192122924894110e-06
GC_1_525 b_1 NI_1 NS_525 0 6.6959739397162805e-09
GC_1_526 b_1 NI_1 NS_526 0 5.4073953858017388e-09
GC_1_527 b_1 NI_1 NS_527 0 1.7777235253457072e-06
GC_1_528 b_1 NI_1 NS_528 0 4.4395358542096964e-07
GC_1_529 b_1 NI_1 NS_529 0 -1.5869735788636677e-06
GC_1_530 b_1 NI_1 NS_530 0 3.2264934738449072e-06
GC_1_531 b_1 NI_1 NS_531 0 -8.2721064458509379e-07
GC_1_532 b_1 NI_1 NS_532 0 6.9325933769457430e-07
GC_1_533 b_1 NI_1 NS_533 0 -7.6673739082868226e-06
GC_1_534 b_1 NI_1 NS_534 0 4.7218363040188629e-07
GC_1_535 b_1 NI_1 NS_535 0 -2.2070929496261079e-06
GC_1_536 b_1 NI_1 NS_536 0 1.9527358661088228e-06
GC_1_537 b_1 NI_1 NS_537 0 -2.0870473420942245e-06
GC_1_538 b_1 NI_1 NS_538 0 1.9632477567105223e-06
GC_1_539 b_1 NI_1 NS_539 0 1.2949329871419346e-06
GC_1_540 b_1 NI_1 NS_540 0 2.8398322222945939e-06
GC_1_541 b_1 NI_1 NS_541 0 -1.5264428399970240e-04
GC_1_542 b_1 NI_1 NS_542 0 3.6649132892898950e-11
GC_1_543 b_1 NI_1 NS_543 0 1.8928590922149661e-11
GC_1_544 b_1 NI_1 NS_544 0 9.3054076807431039e-10
GC_1_545 b_1 NI_1 NS_545 0 -2.3228676044917988e-06
GC_1_546 b_1 NI_1 NS_546 0 -1.6428464482290505e-06
GC_1_547 b_1 NI_1 NS_547 0 1.4316065188687036e-06
GC_1_548 b_1 NI_1 NS_548 0 3.8987525939732385e-06
GC_1_549 b_1 NI_1 NS_549 0 3.0058947704748358e-06
GC_1_550 b_1 NI_1 NS_550 0 5.4030088564441270e-06
GC_1_551 b_1 NI_1 NS_551 0 5.4598824609792475e-06
GC_1_552 b_1 NI_1 NS_552 0 -8.4815335176039264e-06
GC_1_553 b_1 NI_1 NS_553 0 -2.3143021991359662e-06
GC_1_554 b_1 NI_1 NS_554 0 -1.2723713125522872e-05
GC_1_555 b_1 NI_1 NS_555 0 -3.7422815479914989e-06
GC_1_556 b_1 NI_1 NS_556 0 2.7239280806643890e-06
GC_1_557 b_1 NI_1 NS_557 0 4.5151374665530798e-06
GC_1_558 b_1 NI_1 NS_558 0 1.5308267084965942e-06
GC_1_559 b_1 NI_1 NS_559 0 8.7546974060670150e-06
GC_1_560 b_1 NI_1 NS_560 0 -3.8479490037179314e-05
GC_1_561 b_1 NI_1 NS_561 0 -4.3264671443631738e-05
GC_1_562 b_1 NI_1 NS_562 0 -1.4454744379327977e-06
GC_1_563 b_1 NI_1 NS_563 0 -1.4749717205410142e-05
GC_1_564 b_1 NI_1 NS_564 0 -8.4842945954629639e-06
GC_1_565 b_1 NI_1 NS_565 0 -7.0816462319778944e-05
GC_1_566 b_1 NI_1 NS_566 0 7.5582598455229229e-05
GC_1_567 b_1 NI_1 NS_567 0 4.8530274531807275e-06
GC_1_568 b_1 NI_1 NS_568 0 1.3247865580993275e-05
GC_1_569 b_1 NI_1 NS_569 0 6.5374369184357010e-05
GC_1_570 b_1 NI_1 NS_570 0 1.2308042481895385e-04
GC_1_571 b_1 NI_1 NS_571 0 -1.3621919957046133e-07
GC_1_572 b_1 NI_1 NS_572 0 -3.7823808583904314e-05
GC_1_573 b_1 NI_1 NS_573 0 1.6963590097517820e-05
GC_1_574 b_1 NI_1 NS_574 0 4.3619938108783868e-06
GC_1_575 b_1 NI_1 NS_575 0 2.5306794315928710e-05
GC_1_576 b_1 NI_1 NS_576 0 -3.1224053636926455e-05
GC_1_577 b_1 NI_1 NS_577 0 -8.6239860494983006e-06
GC_1_578 b_1 NI_1 NS_578 0 -2.7323210456153975e-06
GC_1_579 b_1 NI_1 NS_579 0 -8.1953044485731331e-06
GC_1_580 b_1 NI_1 NS_580 0 2.4464548376856204e-05
GC_1_581 b_1 NI_1 NS_581 0 6.0407838915878882e-06
GC_1_582 b_1 NI_1 NS_582 0 8.5945639768612187e-06
GC_1_583 b_1 NI_1 NS_583 0 5.7640726660439236e-05
GC_1_584 b_1 NI_1 NS_584 0 2.4091623802097210e-05
GC_1_585 b_1 NI_1 NS_585 0 3.6450330993384114e-06
GC_1_586 b_1 NI_1 NS_586 0 -1.2427359565397291e-05
GC_1_587 b_1 NI_1 NS_587 0 -7.2829865777896872e-08
GC_1_588 b_1 NI_1 NS_588 0 -1.3777667482690573e-06
GC_1_589 b_1 NI_1 NS_589 0 7.2151138915891430e-06
GC_1_590 b_1 NI_1 NS_590 0 2.9209468974009380e-06
GC_1_591 b_1 NI_1 NS_591 0 4.2720192042089456e-05
GC_1_592 b_1 NI_1 NS_592 0 -1.9006948602793728e-05
GC_1_593 b_1 NI_1 NS_593 0 -2.4852095675016650e-06
GC_1_594 b_1 NI_1 NS_594 0 -7.7713965379320601e-06
GC_1_595 b_1 NI_1 NS_595 0 -2.8170144077133781e-06
GC_1_596 b_1 NI_1 NS_596 0 1.1098406511235079e-06
GC_1_597 b_1 NI_1 NS_597 0 9.8836296878130054e-06
GC_1_598 b_1 NI_1 NS_598 0 2.6879758237826445e-06
GC_1_599 b_1 NI_1 NS_599 0 2.2660734469142287e-05
GC_1_600 b_1 NI_1 NS_600 0 -3.3266526713047401e-05
GC_1_601 b_1 NI_1 NS_601 0 -5.7339970441297675e-06
GC_1_602 b_1 NI_1 NS_602 0 -4.2993067218084699e-06
GC_1_603 b_1 NI_1 NS_603 0 -8.7801679880195232e-07
GC_1_604 b_1 NI_1 NS_604 0 4.2822877570003244e-06
GC_1_605 b_1 NI_1 NS_605 0 1.2543454714744512e-05
GC_1_606 b_1 NI_1 NS_606 0 -1.7546384261439789e-07
GC_1_607 b_1 NI_1 NS_607 0 6.1365687914324302e-07
GC_1_608 b_1 NI_1 NS_608 0 -3.3004228705351794e-05
GC_1_609 b_1 NI_1 NS_609 0 -6.9295573805267525e-06
GC_1_610 b_1 NI_1 NS_610 0 3.5363856915814961e-07
GC_1_611 b_1 NI_1 NS_611 0 3.8626268484334861e-06
GC_1_612 b_1 NI_1 NS_612 0 3.5637321733248592e-06
GC_1_613 b_1 NI_1 NS_613 0 1.4168106270637756e-05
GC_1_614 b_1 NI_1 NS_614 0 -6.6370175193129667e-06
GC_1_615 b_1 NI_1 NS_615 0 -1.5560866986288483e-05
GC_1_616 b_1 NI_1 NS_616 0 -1.9131989493466493e-05
GC_1_617 b_1 NI_1 NS_617 0 -2.9829588374360874e-06
GC_1_618 b_1 NI_1 NS_618 0 5.0701561833278959e-06
GC_1_619 b_1 NI_1 NS_619 0 4.2041649275303831e-06
GC_1_620 b_1 NI_1 NS_620 0 -1.9026015325060855e-06
GC_1_621 b_1 NI_1 NS_621 0 -2.7722790310416844e-11
GC_1_622 b_1 NI_1 NS_622 0 5.4084110262601355e-12
GC_1_623 b_1 NI_1 NS_623 0 4.8943388946700578e-06
GC_1_624 b_1 NI_1 NS_624 0 -1.1671181898417512e-05
GC_1_625 b_1 NI_1 NS_625 0 -5.0226833666976024e-07
GC_1_626 b_1 NI_1 NS_626 0 2.7925780467032050e-06
GC_1_627 b_1 NI_1 NS_627 0 2.3625598514337450e-06
GC_1_628 b_1 NI_1 NS_628 0 -1.5932478386881160e-06
GC_1_629 b_1 NI_1 NS_629 0 2.1702787462610420e-06
GC_1_630 b_1 NI_1 NS_630 0 -9.8796191162116970e-06
GC_1_631 b_1 NI_1 NS_631 0 -1.0601745811140070e-05
GC_1_632 b_1 NI_1 NS_632 0 -3.5479047838036458e-06
GC_1_633 b_1 NI_1 NS_633 0 -2.2615837183871249e-10
GC_1_634 b_1 NI_1 NS_634 0 4.2333550538492704e-10
GC_1_635 b_1 NI_1 NS_635 0 -9.1524849094126705e-06
GC_1_636 b_1 NI_1 NS_636 0 -5.6556656184864412e-06
GC_1_637 b_1 NI_1 NS_637 0 2.0113014697140588e-06
GC_1_638 b_1 NI_1 NS_638 0 -6.6968795823165202e-06
GC_1_639 b_1 NI_1 NS_639 0 -3.3581444652303078e-06
GC_1_640 b_1 NI_1 NS_640 0 -1.8350860972418478e-07
GC_1_641 b_1 NI_1 NS_641 0 -8.5821482899103483e-06
GC_1_642 b_1 NI_1 NS_642 0 5.9050997224498942e-07
GC_1_643 b_1 NI_1 NS_643 0 2.6252784674000122e-06
GC_1_644 b_1 NI_1 NS_644 0 2.8290986360157644e-06
GC_1_645 b_1 NI_1 NS_645 0 1.0192405471127688e-06
GC_1_646 b_1 NI_1 NS_646 0 -3.7248629659019981e-06
GC_1_647 b_1 NI_1 NS_647 0 -5.3998861493844549e-06
GC_1_648 b_1 NI_1 NS_648 0 -4.2209465551541440e-06
GC_1_649 b_1 NI_1 NS_649 0 4.7667634991338681e-05
GC_1_650 b_1 NI_1 NS_650 0 7.4776847031506445e-12
GC_1_651 b_1 NI_1 NS_651 0 -1.8812256119375492e-11
GC_1_652 b_1 NI_1 NS_652 0 9.9179838164105649e-10
GC_1_653 b_1 NI_1 NS_653 0 -6.5157794694004389e-08
GC_1_654 b_1 NI_1 NS_654 0 2.4828598365694043e-07
GC_1_655 b_1 NI_1 NS_655 0 2.2372320514292207e-07
GC_1_656 b_1 NI_1 NS_656 0 4.0478127486981010e-07
GC_1_657 b_1 NI_1 NS_657 0 -1.7409002867060431e-07
GC_1_658 b_1 NI_1 NS_658 0 2.7593251513154737e-07
GC_1_659 b_1 NI_1 NS_659 0 7.2779076971384783e-07
GC_1_660 b_1 NI_1 NS_660 0 1.4717948094694481e-06
GC_1_661 b_1 NI_1 NS_661 0 1.0335880791094407e-06
GC_1_662 b_1 NI_1 NS_662 0 -4.2692968700297716e-07
GC_1_663 b_1 NI_1 NS_663 0 3.0382920003609948e-07
GC_1_664 b_1 NI_1 NS_664 0 9.1841908444365410e-07
GC_1_665 b_1 NI_1 NS_665 0 7.7986142233585933e-07
GC_1_666 b_1 NI_1 NS_666 0 -3.1608329173884109e-07
GC_1_667 b_1 NI_1 NS_667 0 4.3388026286861650e-06
GC_1_668 b_1 NI_1 NS_668 0 1.5030455980821885e-06
GC_1_669 b_1 NI_1 NS_669 0 -1.5184037606617087e-06
GC_1_670 b_1 NI_1 NS_670 0 -3.5718097889197916e-06
GC_1_671 b_1 NI_1 NS_671 0 2.4364831324376439e-07
GC_1_672 b_1 NI_1 NS_672 0 1.5787640687712293e-06
GC_1_673 b_1 NI_1 NS_673 0 3.1022177414005644e-06
GC_1_674 b_1 NI_1 NS_674 0 -4.6733355510217803e-06
GC_1_675 b_1 NI_1 NS_675 0 -7.4687476832322560e-07
GC_1_676 b_1 NI_1 NS_676 0 5.6934744772133024e-07
GC_1_677 b_1 NI_1 NS_677 0 5.7285804675535073e-06
GC_1_678 b_1 NI_1 NS_678 0 -5.7347848856970326e-06
GC_1_679 b_1 NI_1 NS_679 0 -3.3214859807985778e-06
GC_1_680 b_1 NI_1 NS_680 0 1.7576634704131742e-06
GC_1_681 b_1 NI_1 NS_681 0 8.8321672371989189e-07
GC_1_682 b_1 NI_1 NS_682 0 1.2580676808604446e-06
GC_1_683 b_1 NI_1 NS_683 0 1.6925156656259456e-06
GC_1_684 b_1 NI_1 NS_684 0 -4.0851793469377355e-06
GC_1_685 b_1 NI_1 NS_685 0 6.1027164515327597e-07
GC_1_686 b_1 NI_1 NS_686 0 2.1452821416541284e-07
GC_1_687 b_1 NI_1 NS_687 0 2.5203339336950535e-07
GC_1_688 b_1 NI_1 NS_688 0 -4.0638363195331192e-06
GC_1_689 b_1 NI_1 NS_689 0 -1.5631455390921308e-07
GC_1_690 b_1 NI_1 NS_690 0 1.7770660228377965e-07
GC_1_691 b_1 NI_1 NS_691 0 4.7896809045742640e-06
GC_1_692 b_1 NI_1 NS_692 0 -6.3217698546668245e-06
GC_1_693 b_1 NI_1 NS_693 0 -1.7965573454654146e-06
GC_1_694 b_1 NI_1 NS_694 0 -1.3136933530981270e-06
GC_1_695 b_1 NI_1 NS_695 0 1.3999546725855262e-06
GC_1_696 b_1 NI_1 NS_696 0 -1.1893440076757560e-06
GC_1_697 b_1 NI_1 NS_697 0 4.3391057721770385e-07
GC_1_698 b_1 NI_1 NS_698 0 -2.1052476083066785e-06
GC_1_699 b_1 NI_1 NS_699 0 -1.3418245259665670e-06
GC_1_700 b_1 NI_1 NS_700 0 -1.1874133880432384e-05
GC_1_701 b_1 NI_1 NS_701 0 -2.2438004868045952e-06
GC_1_702 b_1 NI_1 NS_702 0 -1.7319021713360125e-06
GC_1_703 b_1 NI_1 NS_703 0 -2.3535060375479365e-06
GC_1_704 b_1 NI_1 NS_704 0 -4.0395593952659807e-06
GC_1_705 b_1 NI_1 NS_705 0 -1.4505098359950838e-06
GC_1_706 b_1 NI_1 NS_706 0 -2.4379033461916955e-06
GC_1_707 b_1 NI_1 NS_707 0 -1.0686776496428313e-05
GC_1_708 b_1 NI_1 NS_708 0 -7.2206330999653853e-06
GC_1_709 b_1 NI_1 NS_709 0 -3.1790011754201251e-06
GC_1_710 b_1 NI_1 NS_710 0 -8.7765696002126754e-07
GC_1_711 b_1 NI_1 NS_711 0 -5.7557878621449920e-06
GC_1_712 b_1 NI_1 NS_712 0 -4.1572972767071986e-07
GC_1_713 b_1 NI_1 NS_713 0 -3.1006027440169650e-06
GC_1_714 b_1 NI_1 NS_714 0 -1.7564435173153082e-06
GC_1_715 b_1 NI_1 NS_715 0 -1.0631077550859850e-05
GC_1_716 b_1 NI_1 NS_716 0 3.2969265906245892e-06
GC_1_717 b_1 NI_1 NS_717 0 -3.6194761454602404e-06
GC_1_718 b_1 NI_1 NS_718 0 8.1861921741097109e-07
GC_1_719 b_1 NI_1 NS_719 0 -2.8825399718510349e-06
GC_1_720 b_1 NI_1 NS_720 0 3.9154070853532000e-06
GC_1_721 b_1 NI_1 NS_721 0 -4.3323126070155919e-06
GC_1_722 b_1 NI_1 NS_722 0 1.7065222683208521e-07
GC_1_723 b_1 NI_1 NS_723 0 -1.8686337116389320e-06
GC_1_724 b_1 NI_1 NS_724 0 7.2154273629241074e-06
GC_1_725 b_1 NI_1 NS_725 0 -1.5642574239963418e-06
GC_1_726 b_1 NI_1 NS_726 0 2.7942572187065192e-06
GC_1_727 b_1 NI_1 NS_727 0 9.2411099653240610e-07
GC_1_728 b_1 NI_1 NS_728 0 1.8150576312827812e-06
GC_1_729 b_1 NI_1 NS_729 0 -3.0215515435431412e-11
GC_1_730 b_1 NI_1 NS_730 0 -3.9734318930103948e-12
GC_1_731 b_1 NI_1 NS_731 0 -1.7144585895151410e-06
GC_1_732 b_1 NI_1 NS_732 0 2.1408166849345804e-06
GC_1_733 b_1 NI_1 NS_733 0 -3.2467234438535779e-07
GC_1_734 b_1 NI_1 NS_734 0 1.0491055714752952e-06
GC_1_735 b_1 NI_1 NS_735 0 1.4393954742628979e-07
GC_1_736 b_1 NI_1 NS_736 0 6.2162096391356932e-07
GC_1_737 b_1 NI_1 NS_737 0 -1.0469794411795822e-06
GC_1_738 b_1 NI_1 NS_738 0 1.2713193986409870e-06
GC_1_739 b_1 NI_1 NS_739 0 9.7964306394159268e-07
GC_1_740 b_1 NI_1 NS_740 0 1.8202535954245332e-06
GC_1_741 b_1 NI_1 NS_741 0 -1.5166092265821539e-09
GC_1_742 b_1 NI_1 NS_742 0 -7.8069310747819796e-10
GC_1_743 b_1 NI_1 NS_743 0 -4.8493308084957737e-07
GC_1_744 b_1 NI_1 NS_744 0 -2.7294746177595716e-08
GC_1_745 b_1 NI_1 NS_745 0 -3.1063970948731694e-07
GC_1_746 b_1 NI_1 NS_746 0 1.7482714071519435e-07
GC_1_747 b_1 NI_1 NS_747 0 -5.5091839441355379e-07
GC_1_748 b_1 NI_1 NS_748 0 1.5193413497055865e-07
GC_1_749 b_1 NI_1 NS_749 0 6.6426777512670208e-07
GC_1_750 b_1 NI_1 NS_750 0 8.1167777933365757e-07
GC_1_751 b_1 NI_1 NS_751 0 2.1767291504337169e-07
GC_1_752 b_1 NI_1 NS_752 0 6.9613027546740794e-07
GC_1_753 b_1 NI_1 NS_753 0 1.1062267534101281e-08
GC_1_754 b_1 NI_1 NS_754 0 -1.3787266932550285e-07
GC_1_755 b_1 NI_1 NS_755 0 -3.4802849371124018e-07
GC_1_756 b_1 NI_1 NS_756 0 2.9432595917684435e-07
GC_1_757 b_1 NI_1 NS_757 0 -8.9925218205147572e-05
GC_1_758 b_1 NI_1 NS_758 0 3.3207625557556248e-12
GC_1_759 b_1 NI_1 NS_759 0 -4.3129003689820412e-11
GC_1_760 b_1 NI_1 NS_760 0 3.0190931034018415e-10
GC_1_761 b_1 NI_1 NS_761 0 -1.5707265267596847e-06
GC_1_762 b_1 NI_1 NS_762 0 -1.5515335302063219e-06
GC_1_763 b_1 NI_1 NS_763 0 9.5011175720599756e-07
GC_1_764 b_1 NI_1 NS_764 0 7.0859701891566132e-07
GC_1_765 b_1 NI_1 NS_765 0 -2.7109494107501498e-06
GC_1_766 b_1 NI_1 NS_766 0 3.0183023951932276e-06
GC_1_767 b_1 NI_1 NS_767 0 -3.0631388585999040e-06
GC_1_768 b_1 NI_1 NS_768 0 -2.5681884249631681e-06
GC_1_769 b_1 NI_1 NS_769 0 1.4917484025306431e-06
GC_1_770 b_1 NI_1 NS_770 0 8.4629974694011571e-08
GC_1_771 b_1 NI_1 NS_771 0 -1.6569930217449169e-06
GC_1_772 b_1 NI_1 NS_772 0 1.7806143435866220e-06
GC_1_773 b_1 NI_1 NS_773 0 8.7351129920769035e-07
GC_1_774 b_1 NI_1 NS_774 0 4.1342415306663632e-06
GC_1_775 b_1 NI_1 NS_775 0 -4.3581737167262901e-06
GC_1_776 b_1 NI_1 NS_776 0 -1.9912127016043016e-06
GC_1_777 b_1 NI_1 NS_777 0 2.4348167028846871e-06
GC_1_778 b_1 NI_1 NS_778 0 -1.8849460000042840e-06
GC_1_779 b_1 NI_1 NS_779 0 -1.1509994185373718e-06
GC_1_780 b_1 NI_1 NS_780 0 3.2760381443478099e-06
GC_1_781 b_1 NI_1 NS_781 0 -8.2168140607561578e-06
GC_1_782 b_1 NI_1 NS_782 0 1.1138773600274359e-05
GC_1_783 b_1 NI_1 NS_783 0 1.2480494970484499e-06
GC_1_784 b_1 NI_1 NS_784 0 -1.6722613313027214e-06
GC_1_785 b_1 NI_1 NS_785 0 9.8795491316207918e-06
GC_1_786 b_1 NI_1 NS_786 0 1.7077773348590559e-05
GC_1_787 b_1 NI_1 NS_787 0 -6.7062994411341483e-07
GC_1_788 b_1 NI_1 NS_788 0 -4.6941500700339070e-07
GC_1_789 b_1 NI_1 NS_789 0 4.0634322347752696e-07
GC_1_790 b_1 NI_1 NS_790 0 -1.3870388681266231e-06
GC_1_791 b_1 NI_1 NS_791 0 6.8974701929178973e-06
GC_1_792 b_1 NI_1 NS_792 0 -1.5804453785663486e-07
GC_1_793 b_1 NI_1 NS_793 0 7.1137389270233561e-07
GC_1_794 b_1 NI_1 NS_794 0 3.0107782934626998e-06
GC_1_795 b_1 NI_1 NS_795 0 5.0117254369979543e-07
GC_1_796 b_1 NI_1 NS_796 0 2.8944367233467796e-06
GC_1_797 b_1 NI_1 NS_797 0 1.1551647547769495e-06
GC_1_798 b_1 NI_1 NS_798 0 -1.4201288575311080e-06
GC_1_799 b_1 NI_1 NS_799 0 9.2615675512690635e-06
GC_1_800 b_1 NI_1 NS_800 0 5.1119747715524988e-06
GC_1_801 b_1 NI_1 NS_801 0 5.5745192723926379e-07
GC_1_802 b_1 NI_1 NS_802 0 1.1628103680073571e-06
GC_1_803 b_1 NI_1 NS_803 0 4.5595296073938857e-08
GC_1_804 b_1 NI_1 NS_804 0 4.6106330260977726e-07
GC_1_805 b_1 NI_1 NS_805 0 1.2710016590994916e-06
GC_1_806 b_1 NI_1 NS_806 0 -8.4419654567064095e-07
GC_1_807 b_1 NI_1 NS_807 0 9.0349216768769687e-06
GC_1_808 b_1 NI_1 NS_808 0 7.0642340918690939e-07
GC_1_809 b_1 NI_1 NS_809 0 8.3856357416351601e-07
GC_1_810 b_1 NI_1 NS_810 0 1.4664570219485881e-06
GC_1_811 b_1 NI_1 NS_811 0 1.0338784039119723e-06
GC_1_812 b_1 NI_1 NS_812 0 6.2486556908687612e-07
GC_1_813 b_1 NI_1 NS_813 0 1.3512321882111644e-06
GC_1_814 b_1 NI_1 NS_814 0 -9.4049600124989625e-07
GC_1_815 b_1 NI_1 NS_815 0 7.9401962162716770e-06
GC_1_816 b_1 NI_1 NS_816 0 -2.0574255574874029e-06
GC_1_817 b_1 NI_1 NS_817 0 1.1774919014089991e-06
GC_1_818 b_1 NI_1 NS_818 0 1.5557241980196506e-06
GC_1_819 b_1 NI_1 NS_819 0 1.6144528239301847e-06
GC_1_820 b_1 NI_1 NS_820 0 -2.1447501936533188e-07
GC_1_821 b_1 NI_1 NS_821 0 1.3152865803807315e-06
GC_1_822 b_1 NI_1 NS_822 0 -9.8120137166388306e-07
GC_1_823 b_1 NI_1 NS_823 0 5.8097408795829562e-06
GC_1_824 b_1 NI_1 NS_824 0 -3.8285001544996836e-06
GC_1_825 b_1 NI_1 NS_825 0 1.8107800533624054e-06
GC_1_826 b_1 NI_1 NS_826 0 1.4375733721327862e-06
GC_1_827 b_1 NI_1 NS_827 0 1.1299057172966509e-06
GC_1_828 b_1 NI_1 NS_828 0 -1.3882960270743553e-06
GC_1_829 b_1 NI_1 NS_829 0 1.4160198575808448e-06
GC_1_830 b_1 NI_1 NS_830 0 -1.0986934170320665e-06
GC_1_831 b_1 NI_1 NS_831 0 2.9955759506803834e-06
GC_1_832 b_1 NI_1 NS_832 0 -4.1669900521497758e-06
GC_1_833 b_1 NI_1 NS_833 0 2.2265267681847416e-06
GC_1_834 b_1 NI_1 NS_834 0 3.1296075911807403e-07
GC_1_835 b_1 NI_1 NS_835 0 -3.0639582407511614e-07
GC_1_836 b_1 NI_1 NS_836 0 -1.1888589103381794e-06
GC_1_837 b_1 NI_1 NS_837 0 2.5432726302652474e-11
GC_1_838 b_1 NI_1 NS_838 0 -4.1105493673853196e-11
GC_1_839 b_1 NI_1 NS_839 0 8.0940359984332026e-07
GC_1_840 b_1 NI_1 NS_840 0 -1.5691568120885569e-06
GC_1_841 b_1 NI_1 NS_841 0 1.2651505112856283e-06
GC_1_842 b_1 NI_1 NS_842 0 2.2094626122462969e-07
GC_1_843 b_1 NI_1 NS_843 0 1.6270340230431924e-07
GC_1_844 b_1 NI_1 NS_844 0 -5.4918503451125140e-07
GC_1_845 b_1 NI_1 NS_845 0 5.5453548516204060e-07
GC_1_846 b_1 NI_1 NS_846 0 -8.6155696530668564e-07
GC_1_847 b_1 NI_1 NS_847 0 1.3101228494516593e-06
GC_1_848 b_1 NI_1 NS_848 0 -2.0776542728331350e-06
GC_1_849 b_1 NI_1 NS_849 0 4.9004241369849262e-10
GC_1_850 b_1 NI_1 NS_850 0 -1.2286555862142567e-09
GC_1_851 b_1 NI_1 NS_851 0 5.5269638593774206e-07
GC_1_852 b_1 NI_1 NS_852 0 -8.6347743980987401e-07
GC_1_853 b_1 NI_1 NS_853 0 7.1657274256928223e-07
GC_1_854 b_1 NI_1 NS_854 0 -9.5174166386364863e-07
GC_1_855 b_1 NI_1 NS_855 0 9.1484538066207609e-08
GC_1_856 b_1 NI_1 NS_856 0 4.9336706704217216e-08
GC_1_857 b_1 NI_1 NS_857 0 1.3737763923271597e-06
GC_1_858 b_1 NI_1 NS_858 0 -1.2452371583956394e-06
GC_1_859 b_1 NI_1 NS_859 0 1.6627830383908924e-06
GC_1_860 b_1 NI_1 NS_860 0 -3.1746340877092975e-07
GC_1_861 b_1 NI_1 NS_861 0 -2.3880342496467442e-07
GC_1_862 b_1 NI_1 NS_862 0 -7.4467008822728145e-07
GC_1_863 b_1 NI_1 NS_863 0 7.3885048364507687e-07
GC_1_864 b_1 NI_1 NS_864 0 2.9287444171229083e-07
GC_1_865 b_1 NI_1 NS_865 0 8.5353704786034774e-06
GC_1_866 b_1 NI_1 NS_866 0 3.7657752912963307e-12
GC_1_867 b_1 NI_1 NS_867 0 -7.8556109733805345e-11
GC_1_868 b_1 NI_1 NS_868 0 2.5472491386882807e-09
GC_1_869 b_1 NI_1 NS_869 0 1.5490998360342992e-08
GC_1_870 b_1 NI_1 NS_870 0 -8.4748465221595510e-08
GC_1_871 b_1 NI_1 NS_871 0 -2.4892840412059719e-07
GC_1_872 b_1 NI_1 NS_872 0 2.7099898489506464e-07
GC_1_873 b_1 NI_1 NS_873 0 7.4290249282271744e-07
GC_1_874 b_1 NI_1 NS_874 0 -2.8388534064636949e-07
GC_1_875 b_1 NI_1 NS_875 0 -9.6871931849573971e-07
GC_1_876 b_1 NI_1 NS_876 0 -2.3710760025017572e-07
GC_1_877 b_1 NI_1 NS_877 0 1.0260920997630067e-06
GC_1_878 b_1 NI_1 NS_878 0 4.0158045599157042e-07
GC_1_879 b_1 NI_1 NS_879 0 -1.2037285122812623e-07
GC_1_880 b_1 NI_1 NS_880 0 -2.7297917785933942e-07
GC_1_881 b_1 NI_1 NS_881 0 1.1063206438297356e-07
GC_1_882 b_1 NI_1 NS_882 0 -5.1161000512560247e-07
GC_1_883 b_1 NI_1 NS_883 0 -2.0841507820502348e-06
GC_1_884 b_1 NI_1 NS_884 0 8.6187378256231683e-07
GC_1_885 b_1 NI_1 NS_885 0 2.4334047634897882e-06
GC_1_886 b_1 NI_1 NS_886 0 -6.0600261081495405e-07
GC_1_887 b_1 NI_1 NS_887 0 -6.6287061715896148e-07
GC_1_888 b_1 NI_1 NS_888 0 -1.3976071837878993e-06
GC_1_889 b_1 NI_1 NS_889 0 4.2935321629221941e-07
GC_1_890 b_1 NI_1 NS_890 0 1.8452584788722363e-06
GC_1_891 b_1 NI_1 NS_891 0 -3.0162630897667337e-08
GC_1_892 b_1 NI_1 NS_892 0 -1.3237443853160071e-06
GC_1_893 b_1 NI_1 NS_893 0 -6.3111958696000754e-07
GC_1_894 b_1 NI_1 NS_894 0 2.5911444250920180e-06
GC_1_895 b_1 NI_1 NS_895 0 4.5382319377295665e-07
GC_1_896 b_1 NI_1 NS_896 0 -2.2434945526742737e-06
GC_1_897 b_1 NI_1 NS_897 0 -7.9908825013216038e-07
GC_1_898 b_1 NI_1 NS_898 0 -9.3142313348879862e-07
GC_1_899 b_1 NI_1 NS_899 0 3.6009685934546090e-07
GC_1_900 b_1 NI_1 NS_900 0 9.1166050762694868e-07
GC_1_901 b_1 NI_1 NS_901 0 -5.5608512820496737e-07
GC_1_902 b_1 NI_1 NS_902 0 -7.2540373613622828e-07
GC_1_903 b_1 NI_1 NS_903 0 4.7741247983444003e-07
GC_1_904 b_1 NI_1 NS_904 0 7.3899243510952519e-07
GC_1_905 b_1 NI_1 NS_905 0 -1.7328930081318513e-07
GC_1_906 b_1 NI_1 NS_906 0 -8.7767195832874048e-07
GC_1_907 b_1 NI_1 NS_907 0 -3.3590695840111846e-07
GC_1_908 b_1 NI_1 NS_908 0 1.1576097202956247e-06
GC_1_909 b_1 NI_1 NS_909 0 2.5415456978741553e-07
GC_1_910 b_1 NI_1 NS_910 0 -8.4414343334111457e-07
GC_1_911 b_1 NI_1 NS_911 0 -6.4136843093424200e-08
GC_1_912 b_1 NI_1 NS_912 0 6.7380930122215642e-08
GC_1_913 b_1 NI_1 NS_913 0 -2.5853731692925395e-07
GC_1_914 b_1 NI_1 NS_914 0 -5.4962236780302718e-07
GC_1_915 b_1 NI_1 NS_915 0 1.8909250177901109e-07
GC_1_916 b_1 NI_1 NS_916 0 7.1453978311692792e-07
GC_1_917 b_1 NI_1 NS_917 0 -7.9753109727658355e-08
GC_1_918 b_1 NI_1 NS_918 0 -6.3559753890320041e-07
GC_1_919 b_1 NI_1 NS_919 0 1.0309073472571145e-07
GC_1_920 b_1 NI_1 NS_920 0 1.0288950249206237e-07
GC_1_921 b_1 NI_1 NS_921 0 -2.8962126646388242e-07
GC_1_922 b_1 NI_1 NS_922 0 -5.9366754294072890e-07
GC_1_923 b_1 NI_1 NS_923 0 1.6267762729444982e-07
GC_1_924 b_1 NI_1 NS_924 0 2.2629276864260377e-07
GC_1_925 b_1 NI_1 NS_925 0 -2.5661155074527880e-07
GC_1_926 b_1 NI_1 NS_926 0 -5.0830119398613699e-07
GC_1_927 b_1 NI_1 NS_927 0 4.8280332271699601e-08
GC_1_928 b_1 NI_1 NS_928 0 -5.1510551616284063e-08
GC_1_929 b_1 NI_1 NS_929 0 -3.6755844250471756e-07
GC_1_930 b_1 NI_1 NS_930 0 -5.5772108541198000e-07
GC_1_931 b_1 NI_1 NS_931 0 -2.3473065062353649e-07
GC_1_932 b_1 NI_1 NS_932 0 1.8283346331071063e-08
GC_1_933 b_1 NI_1 NS_933 0 -4.3348905959049046e-07
GC_1_934 b_1 NI_1 NS_934 0 -3.4064034261615779e-07
GC_1_935 b_1 NI_1 NS_935 0 -1.2461953039811282e-07
GC_1_936 b_1 NI_1 NS_936 0 1.5315607277837712e-08
GC_1_937 b_1 NI_1 NS_937 0 -5.6246383803517942e-07
GC_1_938 b_1 NI_1 NS_938 0 -4.3868109994738859e-07
GC_1_939 b_1 NI_1 NS_939 0 -3.1884355297299377e-07
GC_1_940 b_1 NI_1 NS_940 0 3.1347599290200543e-07
GC_1_941 b_1 NI_1 NS_941 0 -4.9949265410241812e-07
GC_1_942 b_1 NI_1 NS_942 0 3.7092917034455550e-08
GC_1_943 b_1 NI_1 NS_943 0 -1.1552467529369592e-08
GC_1_944 b_1 NI_1 NS_944 0 6.1370300827156978e-08
GC_1_945 b_1 NI_1 NS_945 0 -3.2703367488811547e-12
GC_1_946 b_1 NI_1 NS_946 0 3.1967953928322777e-12
GC_1_947 b_1 NI_1 NS_947 0 -5.7559168021636518e-07
GC_1_948 b_1 NI_1 NS_948 0 4.6740712153220262e-08
GC_1_949 b_1 NI_1 NS_949 0 -2.8964967534768721e-07
GC_1_950 b_1 NI_1 NS_950 0 1.1772139308035727e-07
GC_1_951 b_1 NI_1 NS_951 0 -6.5538444078424600e-09
GC_1_952 b_1 NI_1 NS_952 0 -6.9121947230200931e-08
GC_1_953 b_1 NI_1 NS_953 0 -6.5992732953559318e-07
GC_1_954 b_1 NI_1 NS_954 0 1.4030097782343075e-07
GC_1_955 b_1 NI_1 NS_955 0 2.8354681568748672e-08
GC_1_956 b_1 NI_1 NS_956 0 1.2330387136638975e-07
GC_1_957 b_1 NI_1 NS_957 0 -6.1638206232475730e-11
GC_1_958 b_1 NI_1 NS_958 0 1.2851368970855106e-10
GC_1_959 b_1 NI_1 NS_959 0 -3.4587946766461037e-08
GC_1_960 b_1 NI_1 NS_960 0 1.9625703786221989e-07
GC_1_961 b_1 NI_1 NS_961 0 -3.6686776912860957e-07
GC_1_962 b_1 NI_1 NS_962 0 -4.3787044899047150e-08
GC_1_963 b_1 NI_1 NS_963 0 -1.8653371176012126e-07
GC_1_964 b_1 NI_1 NS_964 0 -2.5483585216431299e-09
GC_1_965 b_1 NI_1 NS_965 0 1.9191386457617091e-07
GC_1_966 b_1 NI_1 NS_966 0 8.0894692172215104e-08
GC_1_967 b_1 NI_1 NS_967 0 -2.6556150651858720e-07
GC_1_968 b_1 NI_1 NS_968 0 3.1336803412570797e-07
GC_1_969 b_1 NI_1 NS_969 0 1.2476999947103999e-07
GC_1_970 b_1 NI_1 NS_970 0 -1.4419553004833362e-07
GC_1_971 b_1 NI_1 NS_971 0 -5.7833744075171485e-08
GC_1_972 b_1 NI_1 NS_972 0 2.3865274337292768e-07
GC_1_973 b_1 NI_1 NS_973 0 -6.4269038241641059e-05
GC_1_974 b_1 NI_1 NS_974 0 3.5608521625298994e-12
GC_1_975 b_1 NI_1 NS_975 0 5.0181476394742783e-11
GC_1_976 b_1 NI_1 NS_976 0 -1.5818265741576425e-09
GC_1_977 b_1 NI_1 NS_977 0 -1.0723769641530345e-06
GC_1_978 b_1 NI_1 NS_978 0 -1.0588520054610921e-06
GC_1_979 b_1 NI_1 NS_979 0 4.0966175197751305e-07
GC_1_980 b_1 NI_1 NS_980 0 3.5701210772589777e-07
GC_1_981 b_1 NI_1 NS_981 0 -2.2606186537331619e-06
GC_1_982 b_1 NI_1 NS_982 0 2.1080723331958036e-06
GC_1_983 b_1 NI_1 NS_983 0 -2.5321040691744948e-06
GC_1_984 b_1 NI_1 NS_984 0 -1.2387515780846197e-06
GC_1_985 b_1 NI_1 NS_985 0 1.3985056993313348e-06
GC_1_986 b_1 NI_1 NS_986 0 9.9855289668105375e-07
GC_1_987 b_1 NI_1 NS_987 0 -1.1234344727136966e-06
GC_1_988 b_1 NI_1 NS_988 0 1.3407166885449851e-06
GC_1_989 b_1 NI_1 NS_989 0 7.2717974126498260e-07
GC_1_990 b_1 NI_1 NS_990 0 3.0410653348924909e-06
GC_1_991 b_1 NI_1 NS_991 0 -2.8465248643829942e-06
GC_1_992 b_1 NI_1 NS_992 0 4.7256440585627649e-07
GC_1_993 b_1 NI_1 NS_993 0 3.6884688834901371e-06
GC_1_994 b_1 NI_1 NS_994 0 -2.0179785706712499e-06
GC_1_995 b_1 NI_1 NS_995 0 -1.8787145445275323e-07
GC_1_996 b_1 NI_1 NS_996 0 2.5631993848328373e-06
GC_1_997 b_1 NI_1 NS_997 0 -4.0642674639875062e-06
GC_1_998 b_1 NI_1 NS_998 0 4.8363350279059956e-06
GC_1_999 b_1 NI_1 NS_999 0 6.4243858154821154e-07
GC_1_1000 b_1 NI_1 NS_1000 0 -1.5864518387114428e-06
GC_1_1001 b_1 NI_1 NS_1001 0 4.6100806243305420e-06
GC_1_1002 b_1 NI_1 NS_1002 0 9.9431511941856787e-06
GC_1_1003 b_1 NI_1 NS_1003 0 -1.1102489666352662e-07
GC_1_1004 b_1 NI_1 NS_1004 0 5.2377246277050100e-07
GC_1_1005 b_1 NI_1 NS_1005 0 -6.3324620518550039e-09
GC_1_1006 b_1 NI_1 NS_1006 0 -7.8556093714293333e-07
GC_1_1007 b_1 NI_1 NS_1007 0 5.3518716461257863e-06
GC_1_1008 b_1 NI_1 NS_1008 0 4.9529632629283703e-07
GC_1_1009 b_1 NI_1 NS_1009 0 8.4638501459824202e-07
GC_1_1010 b_1 NI_1 NS_1010 0 1.9176019784654787e-06
GC_1_1011 b_1 NI_1 NS_1011 0 3.0815075464149169e-08
GC_1_1012 b_1 NI_1 NS_1012 0 1.1332192727145922e-06
GC_1_1013 b_1 NI_1 NS_1013 0 5.8507493873317939e-07
GC_1_1014 b_1 NI_1 NS_1014 0 -1.1108406342547111e-06
GC_1_1015 b_1 NI_1 NS_1015 0 5.8253763756870823e-06
GC_1_1016 b_1 NI_1 NS_1016 0 4.0748099123876920e-06
GC_1_1017 b_1 NI_1 NS_1017 0 6.0627635993518846e-07
GC_1_1018 b_1 NI_1 NS_1018 0 8.5952665164444521e-07
GC_1_1019 b_1 NI_1 NS_1019 0 1.9691886629190546e-07
GC_1_1020 b_1 NI_1 NS_1020 0 2.4098448075952537e-07
GC_1_1021 b_1 NI_1 NS_1021 0 8.4525701275576515e-07
GC_1_1022 b_1 NI_1 NS_1022 0 -6.7216150114709542e-07
GC_1_1023 b_1 NI_1 NS_1023 0 6.6650755007442849e-06
GC_1_1024 b_1 NI_1 NS_1024 0 7.5449820014682551e-07
GC_1_1025 b_1 NI_1 NS_1025 0 7.7455390263945930e-07
GC_1_1026 b_1 NI_1 NS_1026 0 7.4913651464199227e-07
GC_1_1027 b_1 NI_1 NS_1027 0 6.6483843612190144e-07
GC_1_1028 b_1 NI_1 NS_1028 0 -6.6191831018346201e-08
GC_1_1029 b_1 NI_1 NS_1029 0 8.7154980323628372e-07
GC_1_1030 b_1 NI_1 NS_1030 0 -6.4038365874910943e-07
GC_1_1031 b_1 NI_1 NS_1031 0 5.7752120754334234e-06
GC_1_1032 b_1 NI_1 NS_1032 0 -1.5909564992807787e-06
GC_1_1033 b_1 NI_1 NS_1033 0 8.2383600998361142e-07
GC_1_1034 b_1 NI_1 NS_1034 0 5.6703551462648707e-07
GC_1_1035 b_1 NI_1 NS_1035 0 6.2585199809882424e-07
GC_1_1036 b_1 NI_1 NS_1036 0 -5.5331547324779851e-07
GC_1_1037 b_1 NI_1 NS_1037 0 9.3777565358804005e-07
GC_1_1038 b_1 NI_1 NS_1038 0 -4.4580725816626415e-07
GC_1_1039 b_1 NI_1 NS_1039 0 3.9036532139444350e-06
GC_1_1040 b_1 NI_1 NS_1040 0 -2.9907073926661119e-06
GC_1_1041 b_1 NI_1 NS_1041 0 8.9571182224548302e-07
GC_1_1042 b_1 NI_1 NS_1042 0 3.2737751524085106e-07
GC_1_1043 b_1 NI_1 NS_1043 0 2.1610738223718206e-07
GC_1_1044 b_1 NI_1 NS_1044 0 -7.9556802750517936e-07
GC_1_1045 b_1 NI_1 NS_1045 0 1.1598915171262582e-06
GC_1_1046 b_1 NI_1 NS_1046 0 -3.2475159023610365e-07
GC_1_1047 b_1 NI_1 NS_1047 0 1.6774682826949600e-06
GC_1_1048 b_1 NI_1 NS_1048 0 -3.0902005039372228e-06
GC_1_1049 b_1 NI_1 NS_1049 0 7.9113447536958361e-07
GC_1_1050 b_1 NI_1 NS_1050 0 -1.0639016447596902e-07
GC_1_1051 b_1 NI_1 NS_1051 0 -1.9701914479953946e-07
GC_1_1052 b_1 NI_1 NS_1052 0 -4.0861200597093092e-07
GC_1_1053 b_1 NI_1 NS_1053 0 8.5880951507782980e-12
GC_1_1054 b_1 NI_1 NS_1054 0 -1.5730327612410231e-11
GC_1_1055 b_1 NI_1 NS_1055 0 8.3871767630788946e-07
GC_1_1056 b_1 NI_1 NS_1056 0 -5.9378006517672573e-07
GC_1_1057 b_1 NI_1 NS_1057 0 4.9464417176392867e-07
GC_1_1058 b_1 NI_1 NS_1058 0 -3.5991788841252947e-08
GC_1_1059 b_1 NI_1 NS_1059 0 1.7011718931362604e-08
GC_1_1060 b_1 NI_1 NS_1060 0 -8.9110505216608295e-08
GC_1_1061 b_1 NI_1 NS_1061 0 5.2142187953855885e-07
GC_1_1062 b_1 NI_1 NS_1062 0 -1.7665126343983346e-08
GC_1_1063 b_1 NI_1 NS_1063 0 7.0517929069376941e-07
GC_1_1064 b_1 NI_1 NS_1064 0 -1.5613971828937544e-06
GC_1_1065 b_1 NI_1 NS_1065 0 4.0969158122779004e-10
GC_1_1066 b_1 NI_1 NS_1066 0 -5.8070646204711723e-10
GC_1_1067 b_1 NI_1 NS_1067 0 1.0099580412046372e-06
GC_1_1068 b_1 NI_1 NS_1068 0 -2.7386484742794206e-07
GC_1_1069 b_1 NI_1 NS_1069 0 3.5400824713411028e-07
GC_1_1070 b_1 NI_1 NS_1070 0 -1.7369715843651193e-07
GC_1_1071 b_1 NI_1 NS_1071 0 2.5492777521074502e-07
GC_1_1072 b_1 NI_1 NS_1072 0 2.6554610617675391e-08
GC_1_1073 b_1 NI_1 NS_1073 0 1.0857964010502795e-06
GC_1_1074 b_1 NI_1 NS_1074 0 -1.1750256139168005e-06
GC_1_1075 b_1 NI_1 NS_1075 0 6.5375796995367926e-07
GC_1_1076 b_1 NI_1 NS_1076 0 -3.3455195392977169e-07
GC_1_1077 b_1 NI_1 NS_1077 0 -2.1221517820184706e-07
GC_1_1078 b_1 NI_1 NS_1078 0 -9.8558751132562085e-08
GC_1_1079 b_1 NI_1 NS_1079 0 7.5732237739999659e-07
GC_1_1080 b_1 NI_1 NS_1080 0 3.2283825784083746e-07
GC_1_1081 b_1 NI_1 NS_1081 0 1.0245384258995773e-05
GC_1_1082 b_1 NI_1 NS_1082 0 -4.7958088227125739e-12
GC_1_1083 b_1 NI_1 NS_1083 0 1.0352297964230360e-11
GC_1_1084 b_1 NI_1 NS_1084 0 3.7845454076365777e-10
GC_1_1085 b_1 NI_1 NS_1085 0 1.3513077173965740e-07
GC_1_1086 b_1 NI_1 NS_1086 0 1.0761870573568796e-07
GC_1_1087 b_1 NI_1 NS_1087 0 7.2008562286728628e-07
GC_1_1088 b_1 NI_1 NS_1088 0 -1.8726845596581332e-07
GC_1_1089 b_1 NI_1 NS_1089 0 -5.9812718062634980e-07
GC_1_1090 b_1 NI_1 NS_1090 0 -3.6307219401307903e-07
GC_1_1091 b_1 NI_1 NS_1091 0 1.3990038660999155e-06
GC_1_1092 b_1 NI_1 NS_1092 0 3.2530787826127925e-07
GC_1_1093 b_1 NI_1 NS_1093 0 -9.9970735240279225e-07
GC_1_1094 b_1 NI_1 NS_1094 0 -1.7789827642819512e-06
GC_1_1095 b_1 NI_1 NS_1095 0 2.5546176889479215e-07
GC_1_1096 b_1 NI_1 NS_1096 0 -5.4933497040031238e-09
GC_1_1097 b_1 NI_1 NS_1097 0 -8.7355628960942563e-07
GC_1_1098 b_1 NI_1 NS_1098 0 9.7895470201604934e-08
GC_1_1099 b_1 NI_1 NS_1099 0 2.5713369721440631e-06
GC_1_1100 b_1 NI_1 NS_1100 0 -1.1144100002988219e-06
GC_1_1101 b_1 NI_1 NS_1101 0 -3.9893102937372838e-06
GC_1_1102 b_1 NI_1 NS_1102 0 -2.3993361286701073e-07
GC_1_1103 b_1 NI_1 NS_1103 0 1.2124338328002744e-08
GC_1_1104 b_1 NI_1 NS_1104 0 1.6053661122360611e-06
GC_1_1105 b_1 NI_1 NS_1105 0 -8.3049225972147176e-07
GC_1_1106 b_1 NI_1 NS_1106 0 -2.6088805033676240e-06
GC_1_1107 b_1 NI_1 NS_1107 0 -7.8261942813012342e-07
GC_1_1108 b_1 NI_1 NS_1108 0 1.4932796656384996e-06
GC_1_1109 b_1 NI_1 NS_1109 0 5.8169597730079314e-07
GC_1_1110 b_1 NI_1 NS_1110 0 -3.0275529235370791e-06
GC_1_1111 b_1 NI_1 NS_1111 0 -1.4470915337603056e-06
GC_1_1112 b_1 NI_1 NS_1112 0 2.5662113529757830e-06
GC_1_1113 b_1 NI_1 NS_1113 0 2.3925451555009972e-07
GC_1_1114 b_1 NI_1 NS_1114 0 1.2705007888989326e-06
GC_1_1115 b_1 NI_1 NS_1115 0 -6.9734458799339679e-07
GC_1_1116 b_1 NI_1 NS_1116 0 -1.1693047771733218e-06
GC_1_1117 b_1 NI_1 NS_1117 0 -5.8085651812399973e-08
GC_1_1118 b_1 NI_1 NS_1118 0 1.0861713571512818e-06
GC_1_1119 b_1 NI_1 NS_1119 0 -6.5279035323089893e-07
GC_1_1120 b_1 NI_1 NS_1120 0 -7.6713130307013621e-07
GC_1_1121 b_1 NI_1 NS_1121 0 -5.1252978975319072e-07
GC_1_1122 b_1 NI_1 NS_1122 0 1.1060675790626693e-06
GC_1_1123 b_1 NI_1 NS_1123 0 4.4999149023627219e-08
GC_1_1124 b_1 NI_1 NS_1124 0 -8.8827900048031637e-07
GC_1_1125 b_1 NI_1 NS_1125 0 -9.1171396552981851e-07
GC_1_1126 b_1 NI_1 NS_1126 0 1.0678813358339161e-06
GC_1_1127 b_1 NI_1 NS_1127 0 -1.1158379113938508e-07
GC_1_1128 b_1 NI_1 NS_1128 0 7.9073211351303828e-09
GC_1_1129 b_1 NI_1 NS_1129 0 -3.3925154958139826e-07
GC_1_1130 b_1 NI_1 NS_1130 0 1.0187616704955964e-06
GC_1_1131 b_1 NI_1 NS_1131 0 -9.8166434745908840e-08
GC_1_1132 b_1 NI_1 NS_1132 0 1.1223307960179983e-07
GC_1_1133 b_1 NI_1 NS_1133 0 -3.0039653171284692e-07
GC_1_1134 b_1 NI_1 NS_1134 0 1.0059098942816963e-06
GC_1_1135 b_1 NI_1 NS_1135 0 8.0883136640991456e-08
GC_1_1136 b_1 NI_1 NS_1136 0 1.6439747255968547e-07
GC_1_1137 b_1 NI_1 NS_1137 0 -7.9044592831957276e-08
GC_1_1138 b_1 NI_1 NS_1138 0 1.1304481134805368e-06
GC_1_1139 b_1 NI_1 NS_1139 0 7.8461453791312786e-07
GC_1_1140 b_1 NI_1 NS_1140 0 -9.7570838628202824e-09
GC_1_1141 b_1 NI_1 NS_1141 0 8.4840800416579579e-08
GC_1_1142 b_1 NI_1 NS_1142 0 8.2101370411799943e-07
GC_1_1143 b_1 NI_1 NS_1143 0 3.1724421151258472e-07
GC_1_1144 b_1 NI_1 NS_1144 0 -1.9309458351938130e-07
GC_1_1145 b_1 NI_1 NS_1145 0 1.9072402901890414e-07
GC_1_1146 b_1 NI_1 NS_1146 0 1.0069310086911574e-06
GC_1_1147 b_1 NI_1 NS_1147 0 7.9530340488118118e-07
GC_1_1148 b_1 NI_1 NS_1148 0 -8.1778182733392566e-07
GC_1_1149 b_1 NI_1 NS_1149 0 3.2998208114682366e-07
GC_1_1150 b_1 NI_1 NS_1150 0 5.3262081600105107e-07
GC_1_1151 b_1 NI_1 NS_1151 0 -5.5953898156054471e-09
GC_1_1152 b_1 NI_1 NS_1152 0 -5.5296153982669502e-07
GC_1_1153 b_1 NI_1 NS_1153 0 4.5645165259472984e-07
GC_1_1154 b_1 NI_1 NS_1154 0 7.5300520758601643e-07
GC_1_1155 b_1 NI_1 NS_1155 0 -9.7862811646997938e-09
GC_1_1156 b_1 NI_1 NS_1156 0 -1.1013781191883387e-06
GC_1_1157 b_1 NI_1 NS_1157 0 3.1840056913741531e-07
GC_1_1158 b_1 NI_1 NS_1158 0 1.0305578398258949e-07
GC_1_1159 b_1 NI_1 NS_1159 0 -3.9308071966558556e-07
GC_1_1160 b_1 NI_1 NS_1160 0 -2.5353168797515727e-07
GC_1_1161 b_1 NI_1 NS_1161 0 1.4514794153999483e-12
GC_1_1162 b_1 NI_1 NS_1162 0 3.4002756789709351e-12
GC_1_1163 b_1 NI_1 NS_1163 0 3.9031458344833592e-07
GC_1_1164 b_1 NI_1 NS_1164 0 2.2952284883585700e-07
GC_1_1165 b_1 NI_1 NS_1165 0 1.1980142620547435e-07
GC_1_1166 b_1 NI_1 NS_1166 0 3.5452839185948235e-08
GC_1_1167 b_1 NI_1 NS_1167 0 -2.7884429390230538e-07
GC_1_1168 b_1 NI_1 NS_1168 0 -1.0897418319043582e-07
GC_1_1169 b_1 NI_1 NS_1169 0 3.2155756646742162e-07
GC_1_1170 b_1 NI_1 NS_1170 0 6.8216948095005443e-08
GC_1_1171 b_1 NI_1 NS_1171 0 -3.5584815978295839e-07
GC_1_1172 b_1 NI_1 NS_1172 0 -4.5135914814990749e-07
GC_1_1173 b_1 NI_1 NS_1173 0 -1.0584673380418352e-11
GC_1_1174 b_1 NI_1 NS_1174 0 3.2224626933249412e-10
GC_1_1175 b_1 NI_1 NS_1175 0 1.8885751843225794e-07
GC_1_1176 b_1 NI_1 NS_1176 0 -1.9033778301479452e-07
GC_1_1177 b_1 NI_1 NS_1177 0 -7.7180591096607714e-08
GC_1_1178 b_1 NI_1 NS_1178 0 3.9129238311383908e-07
GC_1_1179 b_1 NI_1 NS_1179 0 -1.7579625661375933e-07
GC_1_1180 b_1 NI_1 NS_1180 0 6.2408373933475997e-08
GC_1_1181 b_1 NI_1 NS_1181 0 -5.3348761012331053e-07
GC_1_1182 b_1 NI_1 NS_1182 0 -2.6042276811469348e-07
GC_1_1183 b_1 NI_1 NS_1183 0 5.9192917077450809e-08
GC_1_1184 b_1 NI_1 NS_1184 0 2.3074546667381306e-08
GC_1_1185 b_1 NI_1 NS_1185 0 -3.6617434570277031e-07
GC_1_1186 b_1 NI_1 NS_1186 0 6.6095492751868394e-08
GC_1_1187 b_1 NI_1 NS_1187 0 1.0697299763773797e-07
GC_1_1188 b_1 NI_1 NS_1188 0 3.2656865005653597e-07
GC_1_1189 b_1 NI_1 NS_1189 0 -2.9911173221486412e-05
GC_1_1190 b_1 NI_1 NS_1190 0 1.1048095222991891e-11
GC_1_1191 b_1 NI_1 NS_1191 0 -3.3938009146698972e-11
GC_1_1192 b_1 NI_1 NS_1192 0 2.1481827751444802e-10
GC_1_1193 b_1 NI_1 NS_1193 0 -4.0868868596511456e-07
GC_1_1194 b_1 NI_1 NS_1194 0 -2.7774318382853672e-07
GC_1_1195 b_1 NI_1 NS_1195 0 -1.0550522727598482e-07
GC_1_1196 b_1 NI_1 NS_1196 0 5.6498322822733933e-07
GC_1_1197 b_1 NI_1 NS_1197 0 2.3968371355330480e-07
GC_1_1198 b_1 NI_1 NS_1198 0 1.4051815282390979e-06
GC_1_1199 b_1 NI_1 NS_1199 0 1.1112307900128348e-06
GC_1_1200 b_1 NI_1 NS_1200 0 -3.7354356343831171e-07
GC_1_1201 b_1 NI_1 NS_1201 0 6.7789713601926417e-07
GC_1_1202 b_1 NI_1 NS_1202 0 -2.0311511425906303e-06
GC_1_1203 b_1 NI_1 NS_1203 0 -6.4633694267672091e-07
GC_1_1204 b_1 NI_1 NS_1204 0 2.8079878975699909e-07
GC_1_1205 b_1 NI_1 NS_1205 0 1.0005713576656666e-06
GC_1_1206 b_1 NI_1 NS_1206 0 6.6401102228363034e-07
GC_1_1207 b_1 NI_1 NS_1207 0 3.8996102973396283e-06
GC_1_1208 b_1 NI_1 NS_1208 0 -3.7317995213882810e-06
GC_1_1209 b_1 NI_1 NS_1209 0 -5.6020120952779304e-06
GC_1_1210 b_1 NI_1 NS_1210 0 -3.8667562489040379e-06
GC_1_1211 b_1 NI_1 NS_1211 0 -9.1897851751228860e-07
GC_1_1212 b_1 NI_1 NS_1212 0 -2.0469352376524306e-06
GC_1_1213 b_1 NI_1 NS_1213 0 -1.3607677665812100e-05
GC_1_1214 b_1 NI_1 NS_1214 0 5.3832308047003920e-06
GC_1_1215 b_1 NI_1 NS_1215 0 -5.4034698902712382e-07
GC_1_1216 b_1 NI_1 NS_1216 0 1.8948093686571101e-06
GC_1_1217 b_1 NI_1 NS_1217 0 7.8102993007884422e-07
GC_1_1218 b_1 NI_1 NS_1218 0 1.9317333584848843e-05
GC_1_1219 b_1 NI_1 NS_1219 0 2.7701902439919061e-06
GC_1_1220 b_1 NI_1 NS_1220 0 -4.5964451452450741e-06
GC_1_1221 b_1 NI_1 NS_1221 0 1.4650388630184302e-06
GC_1_1222 b_1 NI_1 NS_1222 0 1.7125873321931918e-06
GC_1_1223 b_1 NI_1 NS_1223 0 5.3187257311558065e-06
GC_1_1224 b_1 NI_1 NS_1224 0 -2.2434162855938697e-06
GC_1_1225 b_1 NI_1 NS_1225 0 -4.1230591487114323e-07
GC_1_1226 b_1 NI_1 NS_1226 0 -8.1329299385298727e-07
GC_1_1227 b_1 NI_1 NS_1227 0 -2.0580543104909368e-06
GC_1_1228 b_1 NI_1 NS_1228 0 2.3269572623047236e-06
GC_1_1229 b_1 NI_1 NS_1229 0 -3.1363925527938227e-08
GC_1_1230 b_1 NI_1 NS_1230 0 1.2404837727111551e-06
GC_1_1231 b_1 NI_1 NS_1231 0 5.2823865452015492e-06
GC_1_1232 b_1 NI_1 NS_1232 0 5.9487399826125207e-06
GC_1_1233 b_1 NI_1 NS_1233 0 1.4530432179488947e-06
GC_1_1234 b_1 NI_1 NS_1234 0 -1.0228754785201235e-06
GC_1_1235 b_1 NI_1 NS_1235 0 1.1373691227615444e-07
GC_1_1236 b_1 NI_1 NS_1236 0 -4.7316172236600780e-08
GC_1_1237 b_1 NI_1 NS_1237 0 5.0717305568391269e-07
GC_1_1238 b_1 NI_1 NS_1238 0 7.4710388460798672e-07
GC_1_1239 b_1 NI_1 NS_1239 0 6.0612473921484193e-06
GC_1_1240 b_1 NI_1 NS_1240 0 4.9609619779223550e-07
GC_1_1241 b_1 NI_1 NS_1241 0 5.5847156366506730e-07
GC_1_1242 b_1 NI_1 NS_1242 0 -8.6793796623137918e-07
GC_1_1243 b_1 NI_1 NS_1243 0 -1.2620910365202743e-07
GC_1_1244 b_1 NI_1 NS_1244 0 -3.6195021437154026e-08
GC_1_1245 b_1 NI_1 NS_1245 0 6.7933683595153924e-07
GC_1_1246 b_1 NI_1 NS_1246 0 8.5069430376643199e-07
GC_1_1247 b_1 NI_1 NS_1247 0 4.7901354514244203e-06
GC_1_1248 b_1 NI_1 NS_1248 0 -1.9393599982243997e-06
GC_1_1249 b_1 NI_1 NS_1249 0 1.3625256888869693e-07
GC_1_1250 b_1 NI_1 NS_1250 0 -7.2246347539931699e-07
GC_1_1251 b_1 NI_1 NS_1251 0 -1.2136751048157018e-07
GC_1_1252 b_1 NI_1 NS_1252 0 1.4889523479760242e-07
GC_1_1253 b_1 NI_1 NS_1253 0 9.4361099694093632e-07
GC_1_1254 b_1 NI_1 NS_1254 0 7.7800960061430492e-07
GC_1_1255 b_1 NI_1 NS_1255 0 2.7633735593720279e-06
GC_1_1256 b_1 NI_1 NS_1256 0 -3.0197974279882405e-06
GC_1_1257 b_1 NI_1 NS_1257 0 -1.0372492258419068e-07
GC_1_1258 b_1 NI_1 NS_1258 0 -4.8471760937194680e-07
GC_1_1259 b_1 NI_1 NS_1259 0 8.9033616067031618e-08
GC_1_1260 b_1 NI_1 NS_1260 0 2.0201010749836439e-07
GC_1_1261 b_1 NI_1 NS_1261 0 1.3142772270252366e-06
GC_1_1262 b_1 NI_1 NS_1262 0 5.1190794733927497e-07
GC_1_1263 b_1 NI_1 NS_1263 0 6.6544744168990564e-07
GC_1_1264 b_1 NI_1 NS_1264 0 -2.7719631488754048e-06
GC_1_1265 b_1 NI_1 NS_1265 0 -1.6530856232657801e-07
GC_1_1266 b_1 NI_1 NS_1266 0 -1.3965319059630030e-07
GC_1_1267 b_1 NI_1 NS_1267 0 2.2791482261247256e-07
GC_1_1268 b_1 NI_1 NS_1268 0 2.3002434380403737e-08
GC_1_1269 b_1 NI_1 NS_1269 0 1.6157122814673357e-12
GC_1_1270 b_1 NI_1 NS_1270 0 -6.1868902060857049e-12
GC_1_1271 b_1 NI_1 NS_1271 0 9.8141681624976042e-07
GC_1_1272 b_1 NI_1 NS_1272 0 -2.6421942871623969e-07
GC_1_1273 b_1 NI_1 NS_1273 0 -2.6951628682238875e-08
GC_1_1274 b_1 NI_1 NS_1274 0 4.9063544491580503e-08
GC_1_1275 b_1 NI_1 NS_1275 0 2.6324992063835156e-07
GC_1_1276 b_1 NI_1 NS_1276 0 1.1274450322268854e-08
GC_1_1277 b_1 NI_1 NS_1277 0 8.3346126065193629e-07
GC_1_1278 b_1 NI_1 NS_1278 0 -1.5917988203912892e-07
GC_1_1279 b_1 NI_1 NS_1279 0 -6.3278673529717265e-08
GC_1_1280 b_1 NI_1 NS_1280 0 -1.0953391574476952e-06
GC_1_1281 b_1 NI_1 NS_1281 0 7.6569319932331943e-11
GC_1_1282 b_1 NI_1 NS_1282 0 -1.9331137282387902e-10
GC_1_1283 b_1 NI_1 NS_1283 0 6.8054859570820136e-07
GC_1_1284 b_1 NI_1 NS_1284 0 -4.3046071152271011e-07
GC_1_1285 b_1 NI_1 NS_1285 0 4.2750306682817931e-07
GC_1_1286 b_1 NI_1 NS_1286 0 1.6125223086140207e-07
GC_1_1287 b_1 NI_1 NS_1287 0 1.4001448397266218e-07
GC_1_1288 b_1 NI_1 NS_1288 0 -8.2569469654814434e-08
GC_1_1289 b_1 NI_1 NS_1289 0 -1.4342639763531244e-07
GC_1_1290 b_1 NI_1 NS_1290 0 -6.7675448163170973e-07
GC_1_1291 b_1 NI_1 NS_1291 0 2.4259608520321782e-08
GC_1_1292 b_1 NI_1 NS_1292 0 2.3629843032300946e-07
GC_1_1293 b_1 NI_1 NS_1293 0 3.3308558588913117e-07
GC_1_1294 b_1 NI_1 NS_1294 0 -5.5341378354054465e-08
GC_1_1295 b_1 NI_1 NS_1295 0 4.0226660260479828e-07
GC_1_1296 b_1 NI_1 NS_1296 0 2.2651278872068571e-07
GD_1_1 b_1 NI_1 NA_1 0 -1.0697627826309073e-02
GD_1_2 b_1 NI_1 NA_2 0 -4.9158964730094904e-03
GD_1_3 b_1 NI_1 NA_3 0 1.0616253486384260e-02
GD_1_4 b_1 NI_1 NA_4 0 -1.1524190468082207e-03
GD_1_5 b_1 NI_1 NA_5 0 3.5826265727156722e-06
GD_1_6 b_1 NI_1 NA_6 0 1.9212508464231526e-05
GD_1_7 b_1 NI_1 NA_7 0 -2.6048129114249810e-06
GD_1_8 b_1 NI_1 NA_8 0 1.1368434537201947e-05
GD_1_9 b_1 NI_1 NA_9 0 -1.1492068523045698e-06
GD_1_10 b_1 NI_1 NA_10 0 8.8077108006292936e-06
GD_1_11 b_1 NI_1 NA_11 0 -2.2825702197041068e-06
GD_1_12 b_1 NI_1 NA_12 0 3.3590104558761906e-06
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 -1.1185318891512081e-02
GC_2_2 b_2 NI_2 NS_2 0 8.4594325180498540e-09
GC_2_3 b_2 NI_2 NS_3 0 9.8721911449637860e-07
GC_2_4 b_2 NI_2 NS_4 0 3.6199500522715448e-05
GC_2_5 b_2 NI_2 NS_5 0 4.3662906184767291e-03
GC_2_6 b_2 NI_2 NS_6 0 -3.4896484639602974e-03
GC_2_7 b_2 NI_2 NS_7 0 -3.7149072093813004e-03
GC_2_8 b_2 NI_2 NS_8 0 6.2509116279174529e-03
GC_2_9 b_2 NI_2 NS_9 0 -8.7863139627084967e-03
GC_2_10 b_2 NI_2 NS_10 0 -5.9489736257098969e-03
GC_2_11 b_2 NI_2 NS_11 0 9.1761805401024219e-03
GC_2_12 b_2 NI_2 NS_12 0 -5.9808508445949524e-03
GC_2_13 b_2 NI_2 NS_13 0 7.1653533573038638e-03
GC_2_14 b_2 NI_2 NS_14 0 1.1911536903754466e-02
GC_2_15 b_2 NI_2 NS_15 0 -4.2323327784051703e-03
GC_2_16 b_2 NI_2 NS_16 0 -1.1251853986173305e-03
GC_2_17 b_2 NI_2 NS_17 0 -8.8793668752458720e-03
GC_2_18 b_2 NI_2 NS_18 0 -4.5104620536031380e-04
GC_2_19 b_2 NI_2 NS_19 0 1.4527757661353691e-02
GC_2_20 b_2 NI_2 NS_20 0 -1.0355614600562044e-02
GC_2_21 b_2 NI_2 NS_21 0 1.6511274776936972e-02
GC_2_22 b_2 NI_2 NS_22 0 4.0488525528743439e-03
GC_2_23 b_2 NI_2 NS_23 0 -1.1485097255967780e-02
GC_2_24 b_2 NI_2 NS_24 0 -1.9365690960972148e-04
GC_2_25 b_2 NI_2 NS_25 0 -1.6607936563914096e-02
GC_2_26 b_2 NI_2 NS_26 0 -4.4552656828734681e-02
GC_2_27 b_2 NI_2 NS_27 0 1.0667427531020028e-02
GC_2_28 b_2 NI_2 NS_28 0 1.0871078766845174e-03
GC_2_29 b_2 NI_2 NS_29 0 -4.8262950733012719e-02
GC_2_30 b_2 NI_2 NS_30 0 1.1004975277486844e-02
GC_2_31 b_2 NI_2 NS_31 0 -1.0464671151952881e-02
GC_2_32 b_2 NI_2 NS_32 0 5.4274164938456827e-04
GC_2_33 b_2 NI_2 NS_33 0 9.7653643368533008e-03
GC_2_34 b_2 NI_2 NS_34 0 -6.1125784264771119e-04
GC_2_35 b_2 NI_2 NS_35 0 4.5934996371976835e-03
GC_2_36 b_2 NI_2 NS_36 0 2.4194364075232778e-02
GC_2_37 b_2 NI_2 NS_37 0 -1.0736724410978921e-02
GC_2_38 b_2 NI_2 NS_38 0 1.9986022318733503e-03
GC_2_39 b_2 NI_2 NS_39 0 -8.4713467636975369e-03
GC_2_40 b_2 NI_2 NS_40 0 -1.3526340808323538e-02
GC_2_41 b_2 NI_2 NS_41 0 1.0155188700111641e-02
GC_2_42 b_2 NI_2 NS_42 0 9.6274536043311281e-04
GC_2_43 b_2 NI_2 NS_43 0 -1.9169400150860594e-02
GC_2_44 b_2 NI_2 NS_44 0 2.8673901252024691e-02
GC_2_45 b_2 NI_2 NS_45 0 -9.6256171620100212e-03
GC_2_46 b_2 NI_2 NS_46 0 -9.4348245151263592e-04
GC_2_47 b_2 NI_2 NS_47 0 1.8844293453739965e-03
GC_2_48 b_2 NI_2 NS_48 0 -1.3764768671320940e-03
GC_2_49 b_2 NI_2 NS_49 0 9.4635363229341758e-03
GC_2_50 b_2 NI_2 NS_50 0 -2.5484226415299741e-04
GC_2_51 b_2 NI_2 NS_51 0 -1.6528682610979169e-04
GC_2_52 b_2 NI_2 NS_52 0 3.0293323953774674e-02
GC_2_53 b_2 NI_2 NS_53 0 -8.5337896249960479e-03
GC_2_54 b_2 NI_2 NS_54 0 1.7749901864751438e-04
GC_2_55 b_2 NI_2 NS_55 0 2.1346942673064573e-04
GC_2_56 b_2 NI_2 NS_56 0 -5.4660291853263513e-03
GC_2_57 b_2 NI_2 NS_57 0 1.0030308692266938e-02
GC_2_58 b_2 NI_2 NS_58 0 -3.4495594413518998e-04
GC_2_59 b_2 NI_2 NS_59 0 8.9348009028942348e-03
GC_2_60 b_2 NI_2 NS_60 0 2.6406081591113115e-02
GC_2_61 b_2 NI_2 NS_61 0 -8.3546045890684987e-03
GC_2_62 b_2 NI_2 NS_62 0 1.4014497012807940e-03
GC_2_63 b_2 NI_2 NS_63 0 -2.5783542028017452e-03
GC_2_64 b_2 NI_2 NS_64 0 -7.3353097824526625e-03
GC_2_65 b_2 NI_2 NS_65 0 1.0543963545994026e-02
GC_2_66 b_2 NI_2 NS_66 0 -8.2794516716442430e-04
GC_2_67 b_2 NI_2 NS_67 0 1.4465628170017118e-02
GC_2_68 b_2 NI_2 NS_68 0 1.9992578331510708e-02
GC_2_69 b_2 NI_2 NS_69 0 -8.2668756533445954e-03
GC_2_70 b_2 NI_2 NS_70 0 2.9582064059229226e-03
GC_2_71 b_2 NI_2 NS_71 0 -5.5757831722139661e-03
GC_2_72 b_2 NI_2 NS_72 0 -6.9085585185648642e-03
GC_2_73 b_2 NI_2 NS_73 0 1.1230526618477061e-02
GC_2_74 b_2 NI_2 NS_74 0 -1.3725314730132663e-03
GC_2_75 b_2 NI_2 NS_75 0 1.5750266787679469e-02
GC_2_76 b_2 NI_2 NS_76 0 1.2967936069378167e-02
GC_2_77 b_2 NI_2 NS_77 0 -7.1659245948872720e-03
GC_2_78 b_2 NI_2 NS_78 0 5.1306113575499031e-03
GC_2_79 b_2 NI_2 NS_79 0 -6.8666967512978150e-03
GC_2_80 b_2 NI_2 NS_80 0 -4.8393269801176083e-03
GC_2_81 b_2 NI_2 NS_81 0 5.3070768232975490e-09
GC_2_82 b_2 NI_2 NS_82 0 4.4270319074752177e-08
GC_2_83 b_2 NI_2 NS_83 0 1.2002194279759631e-02
GC_2_84 b_2 NI_2 NS_84 0 -2.5686812797779961e-03
GC_2_85 b_2 NI_2 NS_85 0 -5.2367715071774566e-03
GC_2_86 b_2 NI_2 NS_86 0 4.7118183221642219e-03
GC_2_87 b_2 NI_2 NS_87 0 -6.1526759348403291e-03
GC_2_88 b_2 NI_2 NS_88 0 -4.3194122054824712e-03
GC_2_89 b_2 NI_2 NS_89 0 1.1768574648813541e-02
GC_2_90 b_2 NI_2 NS_90 0 -3.7146151958965443e-03
GC_2_91 b_2 NI_2 NS_91 0 1.3012614294512937e-02
GC_2_92 b_2 NI_2 NS_92 0 9.4653951069011699e-03
GC_2_93 b_2 NI_2 NS_93 0 3.9556699659738697e-06
GC_2_94 b_2 NI_2 NS_94 0 -9.4249279161021384e-07
GC_2_95 b_2 NI_2 NS_95 0 1.6124339558981966e-02
GC_2_96 b_2 NI_2 NS_96 0 1.6774830659395820e-02
GC_2_97 b_2 NI_2 NS_97 0 1.2055181074532427e-02
GC_2_98 b_2 NI_2 NS_98 0 -2.4727523415190031e-03
GC_2_99 b_2 NI_2 NS_99 0 -8.3469690050764090e-03
GC_2_100 b_2 NI_2 NS_100 0 8.5428143282707689e-05
GC_2_101 b_2 NI_2 NS_101 0 1.1349985622472167e-02
GC_2_102 b_2 NI_2 NS_102 0 7.3343135439746642e-03
GC_2_103 b_2 NI_2 NS_103 0 -4.6479119448414883e-03
GC_2_104 b_2 NI_2 NS_104 0 7.3636028614354754e-03
GC_2_105 b_2 NI_2 NS_105 0 -8.0750687174886496e-03
GC_2_106 b_2 NI_2 NS_106 0 -3.7254203551445827e-03
GC_2_107 b_2 NI_2 NS_107 0 1.5991406060769514e-02
GC_2_108 b_2 NI_2 NS_108 0 -7.7330131665281666e-03
GC_2_109 b_2 NI_2 NS_109 0 -1.5530868320839141e-02
GC_2_110 b_2 NI_2 NS_110 0 6.4872575665567750e-09
GC_2_111 b_2 NI_2 NS_111 0 -1.0780988234711171e-06
GC_2_112 b_2 NI_2 NS_112 0 -2.3175274109547320e-05
GC_2_113 b_2 NI_2 NS_113 0 3.3380760479896800e-04
GC_2_114 b_2 NI_2 NS_114 0 -2.0548502423849409e-04
GC_2_115 b_2 NI_2 NS_115 0 -1.5862582242396593e-03
GC_2_116 b_2 NI_2 NS_116 0 -2.3361772915297943e-03
GC_2_117 b_2 NI_2 NS_117 0 -6.3216355249788909e-05
GC_2_118 b_2 NI_2 NS_118 0 4.3863825431021044e-03
GC_2_119 b_2 NI_2 NS_119 0 1.5399048802873115e-03
GC_2_120 b_2 NI_2 NS_120 0 -5.9456443665762051e-03
GC_2_121 b_2 NI_2 NS_121 0 -4.9710137030513201e-03
GC_2_122 b_2 NI_2 NS_122 0 6.5658943387615068e-03
GC_2_123 b_2 NI_2 NS_123 0 1.1033049601677752e-03
GC_2_124 b_2 NI_2 NS_124 0 -4.8869713796917793e-04
GC_2_125 b_2 NI_2 NS_125 0 2.8351211271457504e-03
GC_2_126 b_2 NI_2 NS_126 0 2.3742295355823253e-03
GC_2_127 b_2 NI_2 NS_127 0 -4.4219508017685934e-03
GC_2_128 b_2 NI_2 NS_128 0 -1.3476668926753766e-02
GC_2_129 b_2 NI_2 NS_129 0 1.7485551924607125e-03
GC_2_130 b_2 NI_2 NS_130 0 1.7702185490222150e-02
GC_2_131 b_2 NI_2 NS_131 0 9.8282594327939853e-03
GC_2_132 b_2 NI_2 NS_132 0 -2.3328386621705405e-03
GC_2_133 b_2 NI_2 NS_133 0 -1.3062251318156800e-02
GC_2_134 b_2 NI_2 NS_134 0 2.3406843805528796e-03
GC_2_135 b_2 NI_2 NS_135 0 9.2233753890635980e-03
GC_2_136 b_2 NI_2 NS_136 0 1.9112827881353511e-03
GC_2_137 b_2 NI_2 NS_137 0 -1.7997095998237681e-02
GC_2_138 b_2 NI_2 NS_138 0 -6.3439019430812761e-03
GC_2_139 b_2 NI_2 NS_139 0 1.5754262105909599e-02
GC_2_140 b_2 NI_2 NS_140 0 6.4095337182158525e-03
GC_2_141 b_2 NI_2 NS_141 0 8.1027183200186072e-03
GC_2_142 b_2 NI_2 NS_142 0 -4.2190611020471230e-03
GC_2_143 b_2 NI_2 NS_143 0 -7.4948915553305828e-03
GC_2_144 b_2 NI_2 NS_144 0 2.0941339334176095e-03
GC_2_145 b_2 NI_2 NS_145 0 6.7044800415872975e-03
GC_2_146 b_2 NI_2 NS_146 0 -2.7628606905911817e-03
GC_2_147 b_2 NI_2 NS_147 0 -6.5432407834933350e-03
GC_2_148 b_2 NI_2 NS_148 0 2.9299446522589906e-03
GC_2_149 b_2 NI_2 NS_149 0 7.6773806179843695e-03
GC_2_150 b_2 NI_2 NS_150 0 4.6375265103131344e-04
GC_2_151 b_2 NI_2 NS_151 0 -9.3401575977012079e-03
GC_2_152 b_2 NI_2 NS_152 0 -5.1079553032413027e-03
GC_2_153 b_2 NI_2 NS_153 0 6.8551899767938370e-03
GC_2_154 b_2 NI_2 NS_154 0 4.0869854575191055e-03
GC_2_155 b_2 NI_2 NS_155 0 -3.8349360358270643e-04
GC_2_156 b_2 NI_2 NS_156 0 -9.2299662211743183e-04
GC_2_157 b_2 NI_2 NS_157 0 5.6963375693308872e-03
GC_2_158 b_2 NI_2 NS_158 0 -1.3852990128852335e-03
GC_2_159 b_2 NI_2 NS_159 0 -9.1011041743309894e-03
GC_2_160 b_2 NI_2 NS_160 0 -1.2296019020128397e-03
GC_2_161 b_2 NI_2 NS_161 0 6.0201772757163870e-03
GC_2_162 b_2 NI_2 NS_162 0 7.1817299147971787e-04
GC_2_163 b_2 NI_2 NS_163 0 -2.6199046907130611e-03
GC_2_164 b_2 NI_2 NS_164 0 2.4600285323152221e-04
GC_2_165 b_2 NI_2 NS_165 0 6.7218299050604410e-03
GC_2_166 b_2 NI_2 NS_166 0 -2.2667453976546949e-03
GC_2_167 b_2 NI_2 NS_167 0 -9.2254204622589167e-03
GC_2_168 b_2 NI_2 NS_168 0 1.5046090677215530e-03
GC_2_169 b_2 NI_2 NS_169 0 5.7525390025045114e-03
GC_2_170 b_2 NI_2 NS_170 0 -1.5177985015858199e-03
GC_2_171 b_2 NI_2 NS_171 0 -3.2852539079674583e-03
GC_2_172 b_2 NI_2 NS_172 0 2.3899132658383392e-03
GC_2_173 b_2 NI_2 NS_173 0 7.2874270495532929e-03
GC_2_174 b_2 NI_2 NS_174 0 -4.1034629640530123e-03
GC_2_175 b_2 NI_2 NS_175 0 -8.5232791386860574e-03
GC_2_176 b_2 NI_2 NS_176 0 4.1574394236146162e-03
GC_2_177 b_2 NI_2 NS_177 0 4.8370647226199876e-03
GC_2_178 b_2 NI_2 NS_178 0 -3.8866667833394011e-03
GC_2_179 b_2 NI_2 NS_179 0 -2.3786687275305809e-03
GC_2_180 b_2 NI_2 NS_180 0 4.7281088504794551e-03
GC_2_181 b_2 NI_2 NS_181 0 7.0803230103502219e-03
GC_2_182 b_2 NI_2 NS_182 0 -7.3558602091557965e-03
GC_2_183 b_2 NI_2 NS_183 0 -7.0931612742461932e-03
GC_2_184 b_2 NI_2 NS_184 0 6.8359962682753694e-03
GC_2_185 b_2 NI_2 NS_185 0 1.6811451238135423e-03
GC_2_186 b_2 NI_2 NS_186 0 -5.3216376516711569e-03
GC_2_187 b_2 NI_2 NS_187 0 5.9853529083184751e-04
GC_2_188 b_2 NI_2 NS_188 0 5.4496392043412601e-03
GC_2_189 b_2 NI_2 NS_189 0 -4.1282353587583988e-09
GC_2_190 b_2 NI_2 NS_190 0 -1.3976314252434924e-08
GC_2_191 b_2 NI_2 NS_191 0 2.7262643674318752e-03
GC_2_192 b_2 NI_2 NS_192 0 -8.5984900355557843e-03
GC_2_193 b_2 NI_2 NS_193 0 8.7601828765639935e-04
GC_2_194 b_2 NI_2 NS_194 0 -3.4431550566540793e-03
GC_2_195 b_2 NI_2 NS_195 0 6.3792143208039767e-04
GC_2_196 b_2 NI_2 NS_196 0 4.0228569547313651e-03
GC_2_197 b_2 NI_2 NS_197 0 2.1875522053167824e-03
GC_2_198 b_2 NI_2 NS_198 0 -8.1664821177312892e-03
GC_2_199 b_2 NI_2 NS_199 0 -3.4772864743812170e-03
GC_2_200 b_2 NI_2 NS_200 0 6.9937177099683992e-03
GC_2_201 b_2 NI_2 NS_201 0 -8.5503727188458092e-08
GC_2_202 b_2 NI_2 NS_202 0 -3.1420283073461758e-07
GC_2_203 b_2 NI_2 NS_203 0 -7.9941562802591515e-03
GC_2_204 b_2 NI_2 NS_204 0 5.3784297957891851e-03
GC_2_205 b_2 NI_2 NS_205 0 4.1818213559482245e-03
GC_2_206 b_2 NI_2 NS_206 0 -6.8548439330208127e-03
GC_2_207 b_2 NI_2 NS_207 0 5.3337133193830906e-03
GC_2_208 b_2 NI_2 NS_208 0 7.4258455792824279e-04
GC_2_209 b_2 NI_2 NS_209 0 -2.3535039763463070e-03
GC_2_210 b_2 NI_2 NS_210 0 6.8399075503824194e-03
GC_2_211 b_2 NI_2 NS_211 0 -1.4841908740740228e-03
GC_2_212 b_2 NI_2 NS_212 0 -4.2255112512419365e-03
GC_2_213 b_2 NI_2 NS_213 0 2.3638870734322553e-03
GC_2_214 b_2 NI_2 NS_214 0 5.0284973543176003e-03
GC_2_215 b_2 NI_2 NS_215 0 -1.9828423531963834e-03
GC_2_216 b_2 NI_2 NS_216 0 -8.9598437406871994e-03
GC_2_217 b_2 NI_2 NS_217 0 -3.3036297565861997e-03
GC_2_218 b_2 NI_2 NS_218 0 1.8493831346309659e-09
GC_2_219 b_2 NI_2 NS_219 0 5.6032190423226659e-08
GC_2_220 b_2 NI_2 NS_220 0 1.8929692337150968e-06
GC_2_221 b_2 NI_2 NS_221 0 -9.1167690568746707e-05
GC_2_222 b_2 NI_2 NS_222 0 -5.7737975891099830e-05
GC_2_223 b_2 NI_2 NS_223 0 -1.2657733206401850e-03
GC_2_224 b_2 NI_2 NS_224 0 -2.9559391462452973e-04
GC_2_225 b_2 NI_2 NS_225 0 -1.6792135372403661e-03
GC_2_226 b_2 NI_2 NS_226 0 2.6464976116021394e-03
GC_2_227 b_2 NI_2 NS_227 0 5.1121143896497648e-04
GC_2_228 b_2 NI_2 NS_228 0 5.4276088285740336e-03
GC_2_229 b_2 NI_2 NS_229 0 7.1034883331695543e-03
GC_2_230 b_2 NI_2 NS_230 0 6.3629271575771059e-04
GC_2_231 b_2 NI_2 NS_231 0 6.4432994603425518e-04
GC_2_232 b_2 NI_2 NS_232 0 -6.6091923874630511e-04
GC_2_233 b_2 NI_2 NS_233 0 1.0576980594074721e-03
GC_2_234 b_2 NI_2 NS_234 0 1.5711404866409924e-03
GC_2_235 b_2 NI_2 NS_235 0 1.2687514030059778e-02
GC_2_236 b_2 NI_2 NS_236 0 1.3123213085017986e-02
GC_2_237 b_2 NI_2 NS_237 0 8.7187976265509382e-03
GC_2_238 b_2 NI_2 NS_238 0 -2.0392080386768058e-02
GC_2_239 b_2 NI_2 NS_239 0 8.3891005356606096e-03
GC_2_240 b_2 NI_2 NS_240 0 -2.9045256325944779e-03
GC_2_241 b_2 NI_2 NS_241 0 -1.2701288428712775e-02
GC_2_242 b_2 NI_2 NS_242 0 -3.8806698120404284e-02
GC_2_243 b_2 NI_2 NS_243 0 -7.2523388521349161e-03
GC_2_244 b_2 NI_2 NS_244 0 -2.1332751224029684e-03
GC_2_245 b_2 NI_2 NS_245 0 -5.2307197827227481e-02
GC_2_246 b_2 NI_2 NS_246 0 -1.7936177184318678e-03
GC_2_247 b_2 NI_2 NS_247 0 1.4914414729235725e-02
GC_2_248 b_2 NI_2 NS_248 0 8.6735769550041093e-03
GC_2_249 b_2 NI_2 NS_249 0 -5.9233531366575005e-03
GC_2_250 b_2 NI_2 NS_250 0 5.0044969310335157e-03
GC_2_251 b_2 NI_2 NS_251 0 8.3724191979080969e-03
GC_2_252 b_2 NI_2 NS_252 0 1.1688363789504238e-02
GC_2_253 b_2 NI_2 NS_253 0 4.5592641881590287e-03
GC_2_254 b_2 NI_2 NS_254 0 -2.9327403911450695e-03
GC_2_255 b_2 NI_2 NS_255 0 -7.8986719502985060e-03
GC_2_256 b_2 NI_2 NS_256 0 -8.1490659263202744e-03
GC_2_257 b_2 NI_2 NS_257 0 -5.6808133994830532e-03
GC_2_258 b_2 NI_2 NS_258 0 -6.1281063168011054e-04
GC_2_259 b_2 NI_2 NS_259 0 -1.8070850020868806e-02
GC_2_260 b_2 NI_2 NS_260 0 1.3578962034020302e-02
GC_2_261 b_2 NI_2 NS_261 0 4.7069857005425228e-03
GC_2_262 b_2 NI_2 NS_262 0 4.3794388164699518e-03
GC_2_263 b_2 NI_2 NS_263 0 6.5015843406849021e-04
GC_2_264 b_2 NI_2 NS_264 0 -1.0995433234541353e-04
GC_2_265 b_2 NI_2 NS_265 0 -3.7963995382206696e-03
GC_2_266 b_2 NI_2 NS_266 0 8.8498815951218598e-04
GC_2_267 b_2 NI_2 NS_267 0 -1.1178289603676467e-03
GC_2_268 b_2 NI_2 NS_268 0 1.6699686387568056e-02
GC_2_269 b_2 NI_2 NS_269 0 4.4472800679289355e-03
GC_2_270 b_2 NI_2 NS_270 0 7.0796428713336597e-04
GC_2_271 b_2 NI_2 NS_271 0 -5.1995857862934360e-04
GC_2_272 b_2 NI_2 NS_272 0 -2.2477513394626226e-03
GC_2_273 b_2 NI_2 NS_273 0 -4.9864559359745365e-03
GC_2_274 b_2 NI_2 NS_274 0 2.1108873302017155e-03
GC_2_275 b_2 NI_2 NS_275 0 7.3425263600871314e-03
GC_2_276 b_2 NI_2 NS_276 0 1.4345854912224685e-02
GC_2_277 b_2 NI_2 NS_277 0 4.1872274196254212e-03
GC_2_278 b_2 NI_2 NS_278 0 -1.6838584350453612e-03
GC_2_279 b_2 NI_2 NS_279 0 -3.3981251384694773e-03
GC_2_280 b_2 NI_2 NS_280 0 -2.1006235094581864e-03
GC_2_281 b_2 NI_2 NS_281 0 -5.4204257484207936e-03
GC_2_282 b_2 NI_2 NS_282 0 4.3817240944628629e-03
GC_2_283 b_2 NI_2 NS_283 0 1.3196871299294649e-02
GC_2_284 b_2 NI_2 NS_284 0 8.4333073908177437e-03
GC_2_285 b_2 NI_2 NS_285 0 2.8324336116298094e-03
GC_2_286 b_2 NI_2 NS_286 0 -4.1306060181108386e-03
GC_2_287 b_2 NI_2 NS_287 0 -5.3207863179017710e-03
GC_2_288 b_2 NI_2 NS_288 0 1.1381587447007421e-03
GC_2_289 b_2 NI_2 NS_289 0 -4.4310206647043392e-03
GC_2_290 b_2 NI_2 NS_290 0 8.3104309118741237e-03
GC_2_291 b_2 NI_2 NS_291 0 1.4612785667001091e-02
GC_2_292 b_2 NI_2 NS_292 0 -4.6824709735628290e-04
GC_2_293 b_2 NI_2 NS_293 0 -1.1845320506053819e-03
GC_2_294 b_2 NI_2 NS_294 0 -4.5473899300001010e-03
GC_2_295 b_2 NI_2 NS_295 0 -2.2825678116614638e-03
GC_2_296 b_2 NI_2 NS_296 0 4.3832546986360549e-03
GC_2_297 b_2 NI_2 NS_297 0 1.3571272571424782e-10
GC_2_298 b_2 NI_2 NS_298 0 -1.5466655106724164e-09
GC_2_299 b_2 NI_2 NS_299 0 1.4460257388538458e-03
GC_2_300 b_2 NI_2 NS_300 0 8.2165466843820093e-03
GC_2_301 b_2 NI_2 NS_301 0 -8.7895047316881368e-04
GC_2_302 b_2 NI_2 NS_302 0 -2.2072124535102121e-03
GC_2_303 b_2 NI_2 NS_303 0 -1.4679135477936311e-03
GC_2_304 b_2 NI_2 NS_304 0 2.7519861855207985e-03
GC_2_305 b_2 NI_2 NS_305 0 1.7320143439264737e-03
GC_2_306 b_2 NI_2 NS_306 0 7.6059325955026196e-03
GC_2_307 b_2 NI_2 NS_307 0 7.5874084276754657e-03
GC_2_308 b_2 NI_2 NS_308 0 -3.8276823066387120e-03
GC_2_309 b_2 NI_2 NS_309 0 -5.2101074820902505e-08
GC_2_310 b_2 NI_2 NS_310 0 -2.0817223764005466e-08
GC_2_311 b_2 NI_2 NS_311 0 1.1391243238784123e-02
GC_2_312 b_2 NI_2 NS_312 0 4.4700330704608368e-03
GC_2_313 b_2 NI_2 NS_313 0 -8.6185054262807707e-04
GC_2_314 b_2 NI_2 NS_314 0 6.4916224677959598e-03
GC_2_315 b_2 NI_2 NS_315 0 3.6263738295167626e-03
GC_2_316 b_2 NI_2 NS_316 0 4.0710468891073996e-04
GC_2_317 b_2 NI_2 NS_317 0 6.0525109540083121e-03
GC_2_318 b_2 NI_2 NS_318 0 -4.6635402185558851e-03
GC_2_319 b_2 NI_2 NS_319 0 -3.3929752213477057e-03
GC_2_320 b_2 NI_2 NS_320 0 -1.3533960294535986e-03
GC_2_321 b_2 NI_2 NS_321 0 1.1237962578393752e-04
GC_2_322 b_2 NI_2 NS_322 0 4.4958002644244774e-03
GC_2_323 b_2 NI_2 NS_323 0 7.2795568416792614e-03
GC_2_324 b_2 NI_2 NS_324 0 5.5305047722385365e-03
GC_2_325 b_2 NI_2 NS_325 0 1.1808946086173740e-03
GC_2_326 b_2 NI_2 NS_326 0 -3.5561529341731014e-09
GC_2_327 b_2 NI_2 NS_327 0 -4.8002191774797389e-08
GC_2_328 b_2 NI_2 NS_328 0 -3.4752340704546351e-06
GC_2_329 b_2 NI_2 NS_329 0 -3.6811901364778671e-04
GC_2_330 b_2 NI_2 NS_330 0 1.3598187543189329e-04
GC_2_331 b_2 NI_2 NS_331 0 1.1297146933370772e-03
GC_2_332 b_2 NI_2 NS_332 0 1.9432462846757804e-03
GC_2_333 b_2 NI_2 NS_333 0 -6.5024476552759974e-05
GC_2_334 b_2 NI_2 NS_334 0 -3.4937331271818937e-03
GC_2_335 b_2 NI_2 NS_335 0 -1.5644021981815197e-03
GC_2_336 b_2 NI_2 NS_336 0 5.0905624229486725e-03
GC_2_337 b_2 NI_2 NS_337 0 4.2534128653169447e-03
GC_2_338 b_2 NI_2 NS_338 0 -4.9937799992362886e-03
GC_2_339 b_2 NI_2 NS_339 0 -1.0085407529908234e-03
GC_2_340 b_2 NI_2 NS_340 0 5.6396386094322969e-04
GC_2_341 b_2 NI_2 NS_341 0 -2.0807406583216526e-03
GC_2_342 b_2 NI_2 NS_342 0 -1.8633318893576997e-03
GC_2_343 b_2 NI_2 NS_343 0 3.6453771295847080e-03
GC_2_344 b_2 NI_2 NS_344 0 1.1647296882442272e-02
GC_2_345 b_2 NI_2 NS_345 0 -8.9809614803268889e-04
GC_2_346 b_2 NI_2 NS_346 0 -1.4854265632828947e-02
GC_2_347 b_2 NI_2 NS_347 0 -8.1235076431967462e-03
GC_2_348 b_2 NI_2 NS_348 0 1.9195537939136612e-03
GC_2_349 b_2 NI_2 NS_349 0 1.1262993530090932e-02
GC_2_350 b_2 NI_2 NS_350 0 -1.8122069155800170e-03
GC_2_351 b_2 NI_2 NS_351 0 -7.5672398442390900e-03
GC_2_352 b_2 NI_2 NS_352 0 -1.6812116993683054e-03
GC_2_353 b_2 NI_2 NS_353 0 1.5281604976723692e-02
GC_2_354 b_2 NI_2 NS_354 0 5.3008405645795431e-03
GC_2_355 b_2 NI_2 NS_355 0 -1.3082790953757063e-02
GC_2_356 b_2 NI_2 NS_356 0 -5.4613178963360621e-03
GC_2_357 b_2 NI_2 NS_357 0 -6.6370644564244397e-03
GC_2_358 b_2 NI_2 NS_358 0 3.4566475701970811e-03
GC_2_359 b_2 NI_2 NS_359 0 6.3615644356748314e-03
GC_2_360 b_2 NI_2 NS_360 0 -1.8793118019296005e-03
GC_2_361 b_2 NI_2 NS_361 0 -5.4737186445375187e-03
GC_2_362 b_2 NI_2 NS_362 0 2.1829946686461677e-03
GC_2_363 b_2 NI_2 NS_363 0 5.3937393709662246e-03
GC_2_364 b_2 NI_2 NS_364 0 -2.6324117744461837e-03
GC_2_365 b_2 NI_2 NS_365 0 -6.3064431411678926e-03
GC_2_366 b_2 NI_2 NS_366 0 -4.8383735656623344e-04
GC_2_367 b_2 NI_2 NS_367 0 7.6452220984870754e-03
GC_2_368 b_2 NI_2 NS_368 0 3.6298705718534534e-03
GC_2_369 b_2 NI_2 NS_369 0 -5.8336093149022675e-03
GC_2_370 b_2 NI_2 NS_370 0 -3.4646024563500504e-03
GC_2_371 b_2 NI_2 NS_371 0 2.9619348919140569e-04
GC_2_372 b_2 NI_2 NS_372 0 5.5809941025784196e-04
GC_2_373 b_2 NI_2 NS_373 0 -4.9270657872239184e-03
GC_2_374 b_2 NI_2 NS_374 0 8.9217852429801937e-04
GC_2_375 b_2 NI_2 NS_375 0 6.2062929702045794e-03
GC_2_376 b_2 NI_2 NS_376 0 6.8828400938346313e-04
GC_2_377 b_2 NI_2 NS_377 0 -5.3209611644941439e-03
GC_2_378 b_2 NI_2 NS_378 0 -4.8420318236978767e-04
GC_2_379 b_2 NI_2 NS_379 0 1.5503149071470397e-03
GC_2_380 b_2 NI_2 NS_380 0 -4.3204677706377475e-05
GC_2_381 b_2 NI_2 NS_381 0 -6.0223419042159353e-03
GC_2_382 b_2 NI_2 NS_382 0 1.9232193706755134e-03
GC_2_383 b_2 NI_2 NS_383 0 6.2616196388788356e-03
GC_2_384 b_2 NI_2 NS_384 0 2.1739983894834415e-04
GC_2_385 b_2 NI_2 NS_385 0 -5.0592028594619387e-03
GC_2_386 b_2 NI_2 NS_386 0 1.7016087774868469e-03
GC_2_387 b_2 NI_2 NS_387 0 2.4884687136955738e-03
GC_2_388 b_2 NI_2 NS_388 0 -9.5763254243005002e-04
GC_2_389 b_2 NI_2 NS_389 0 -6.5329693358750556e-03
GC_2_390 b_2 NI_2 NS_390 0 3.8846207766478919e-03
GC_2_391 b_2 NI_2 NS_391 0 7.4932573120102507e-03
GC_2_392 b_2 NI_2 NS_392 0 -1.0959984792704128e-03
GC_2_393 b_2 NI_2 NS_393 0 -3.9851238840564202e-03
GC_2_394 b_2 NI_2 NS_394 0 4.0409678506999188e-03
GC_2_395 b_2 NI_2 NS_395 0 2.8633256063447339e-03
GC_2_396 b_2 NI_2 NS_396 0 -3.0534816325069694e-03
GC_2_397 b_2 NI_2 NS_397 0 -6.0227369844528872e-03
GC_2_398 b_2 NI_2 NS_398 0 7.2373641985871758e-03
GC_2_399 b_2 NI_2 NS_399 0 7.9896920165465641e-03
GC_2_400 b_2 NI_2 NS_400 0 -4.8114430249764605e-03
GC_2_401 b_2 NI_2 NS_401 0 -5.3743583256991737e-04
GC_2_402 b_2 NI_2 NS_402 0 5.0204619083621810e-03
GC_2_403 b_2 NI_2 NS_403 0 2.4825093756646038e-04
GC_2_404 b_2 NI_2 NS_404 0 -4.7581881502030531e-03
GC_2_405 b_2 NI_2 NS_405 0 1.8107800231229806e-09
GC_2_406 b_2 NI_2 NS_406 0 3.2741335365231206e-09
GC_2_407 b_2 NI_2 NS_407 0 -1.4272202680225157e-03
GC_2_408 b_2 NI_2 NS_408 0 7.8707216177804282e-03
GC_2_409 b_2 NI_2 NS_409 0 -1.7999315117172193e-04
GC_2_410 b_2 NI_2 NS_410 0 3.0272430884242330e-03
GC_2_411 b_2 NI_2 NS_411 0 -1.3039334253086570e-04
GC_2_412 b_2 NI_2 NS_412 0 -3.3752918432831962e-03
GC_2_413 b_2 NI_2 NS_413 0 -8.7633853397992803e-04
GC_2_414 b_2 NI_2 NS_414 0 7.5304799097414919e-03
GC_2_415 b_2 NI_2 NS_415 0 3.7887927327915566e-03
GC_2_416 b_2 NI_2 NS_416 0 -6.1573976215615906e-03
GC_2_417 b_2 NI_2 NS_417 0 8.6224686718229576e-08
GC_2_418 b_2 NI_2 NS_418 0 -3.5295555329358196e-07
GC_2_419 b_2 NI_2 NS_419 0 6.7186820305058341e-03
GC_2_420 b_2 NI_2 NS_420 0 -5.3194053991502989e-03
GC_2_421 b_2 NI_2 NS_421 0 -2.6111752847584736e-03
GC_2_422 b_2 NI_2 NS_422 0 6.0542436034969026e-03
GC_2_423 b_2 NI_2 NS_423 0 -4.2922721356863985e-03
GC_2_424 b_2 NI_2 NS_424 0 1.4428603149853243e-05
GC_2_425 b_2 NI_2 NS_425 0 2.7173857208233404e-03
GC_2_426 b_2 NI_2 NS_426 0 -6.2039921813178698e-03
GC_2_427 b_2 NI_2 NS_427 0 2.0957199164176000e-03
GC_2_428 b_2 NI_2 NS_428 0 3.2562861580773994e-03
GC_2_429 b_2 NI_2 NS_429 0 -1.9700288835581160e-03
GC_2_430 b_2 NI_2 NS_430 0 -4.4205333652797864e-03
GC_2_431 b_2 NI_2 NS_431 0 2.8640817371894025e-03
GC_2_432 b_2 NI_2 NS_432 0 8.0083593647128498e-03
GC_2_433 b_2 NI_2 NS_433 0 -1.5264059909676010e-04
GC_2_434 b_2 NI_2 NS_434 0 3.6649250947427022e-11
GC_2_435 b_2 NI_2 NS_435 0 1.8927352423826123e-11
GC_2_436 b_2 NI_2 NS_436 0 9.3057851778229996e-10
GC_2_437 b_2 NI_2 NS_437 0 -2.3228436259396465e-06
GC_2_438 b_2 NI_2 NS_438 0 -1.6428399936041074e-06
GC_2_439 b_2 NI_2 NS_439 0 1.4316455539952408e-06
GC_2_440 b_2 NI_2 NS_440 0 3.8987617022654576e-06
GC_2_441 b_2 NI_2 NS_441 0 3.0058882387408538e-06
GC_2_442 b_2 NI_2 NS_442 0 5.4029776935402072e-06
GC_2_443 b_2 NI_2 NS_443 0 5.4599134369355556e-06
GC_2_444 b_2 NI_2 NS_444 0 -8.4815362835491988e-06
GC_2_445 b_2 NI_2 NS_445 0 -2.3141895319938047e-06
GC_2_446 b_2 NI_2 NS_446 0 -1.2723709007438416e-05
GC_2_447 b_2 NI_2 NS_447 0 -3.7422369672879436e-06
GC_2_448 b_2 NI_2 NS_448 0 2.7238933259210947e-06
GC_2_449 b_2 NI_2 NS_449 0 4.5150284837565436e-06
GC_2_450 b_2 NI_2 NS_450 0 1.5307784709553071e-06
GC_2_451 b_2 NI_2 NS_451 0 8.7546471814393509e-06
GC_2_452 b_2 NI_2 NS_452 0 -3.8479441360790094e-05
GC_2_453 b_2 NI_2 NS_453 0 -4.3264345003444065e-05
GC_2_454 b_2 NI_2 NS_454 0 -1.4454245746019744e-06
GC_2_455 b_2 NI_2 NS_455 0 -1.4749708908304301e-05
GC_2_456 b_2 NI_2 NS_456 0 -8.4841759693453510e-06
GC_2_457 b_2 NI_2 NS_457 0 -7.0816021676349999e-05
GC_2_458 b_2 NI_2 NS_458 0 7.5581834242249385e-05
GC_2_459 b_2 NI_2 NS_459 0 4.8531178978863821e-06
GC_2_460 b_2 NI_2 NS_460 0 1.3247714630832833e-05
GC_2_461 b_2 NI_2 NS_461 0 6.5373791785026472e-05
GC_2_462 b_2 NI_2 NS_462 0 1.2307919584281818e-04
GC_2_463 b_2 NI_2 NS_463 0 -1.3647831700912228e-07
GC_2_464 b_2 NI_2 NS_464 0 -3.7823400640714276e-05
GC_2_465 b_2 NI_2 NS_465 0 1.6963538378843118e-05
GC_2_466 b_2 NI_2 NS_466 0 4.3618135286846765e-06
GC_2_467 b_2 NI_2 NS_467 0 2.5306405973596128e-05
GC_2_468 b_2 NI_2 NS_468 0 -3.1223662848819990e-05
GC_2_469 b_2 NI_2 NS_469 0 -8.6240524053637949e-06
GC_2_470 b_2 NI_2 NS_470 0 -2.7321969061800880e-06
GC_2_471 b_2 NI_2 NS_471 0 -8.1952294324779061e-06
GC_2_472 b_2 NI_2 NS_472 0 2.4464290128826777e-05
GC_2_473 b_2 NI_2 NS_473 0 6.0408727036470373e-06
GC_2_474 b_2 NI_2 NS_474 0 8.5944397194718999e-06
GC_2_475 b_2 NI_2 NS_475 0 5.7640092850800437e-05
GC_2_476 b_2 NI_2 NS_476 0 2.4091332394611368e-05
GC_2_477 b_2 NI_2 NS_477 0 3.6448050105617273e-06
GC_2_478 b_2 NI_2 NS_478 0 -1.2427225761286242e-05
GC_2_479 b_2 NI_2 NS_479 0 -7.2857785254247174e-08
GC_2_480 b_2 NI_2 NS_480 0 -1.3777536301121229e-06
GC_2_481 b_2 NI_2 NS_481 0 7.2151358017104518e-06
GC_2_482 b_2 NI_2 NS_482 0 2.9209036423094103e-06
GC_2_483 b_2 NI_2 NS_483 0 4.2719686590668904e-05
GC_2_484 b_2 NI_2 NS_484 0 -1.9006737334600494e-05
GC_2_485 b_2 NI_2 NS_485 0 -2.4853121532619056e-06
GC_2_486 b_2 NI_2 NS_486 0 -7.7712935209613263e-06
GC_2_487 b_2 NI_2 NS_487 0 -2.8170038562572319e-06
GC_2_488 b_2 NI_2 NS_488 0 1.1098437794990879e-06
GC_2_489 b_2 NI_2 NS_489 0 9.8836157050574172e-06
GC_2_490 b_2 NI_2 NS_490 0 2.6879024280177039e-06
GC_2_491 b_2 NI_2 NS_491 0 2.2660359756362080e-05
GC_2_492 b_2 NI_2 NS_492 0 -3.3266180569539460e-05
GC_2_493 b_2 NI_2 NS_493 0 -5.7340471794034670e-06
GC_2_494 b_2 NI_2 NS_494 0 -4.2992020704315137e-06
GC_2_495 b_2 NI_2 NS_495 0 -8.7798796691319815e-07
GC_2_496 b_2 NI_2 NS_496 0 4.2823121323874668e-06
GC_2_497 b_2 NI_2 NS_497 0 1.2543409560615316e-05
GC_2_498 b_2 NI_2 NS_498 0 -1.7550097091284672e-07
GC_2_499 b_2 NI_2 NS_499 0 6.1353681763887499e-07
GC_2_500 b_2 NI_2 NS_500 0 -3.3003914400517607e-05
GC_2_501 b_2 NI_2 NS_501 0 -6.9295699343804712e-06
GC_2_502 b_2 NI_2 NS_502 0 3.5370250123400997e-07
GC_2_503 b_2 NI_2 NS_503 0 3.8626384805772639e-06
GC_2_504 b_2 NI_2 NS_504 0 3.5637504740584866e-06
GC_2_505 b_2 NI_2 NS_505 0 1.4168026167722718e-05
GC_2_506 b_2 NI_2 NS_506 0 -6.6370209643289753e-06
GC_2_507 b_2 NI_2 NS_507 0 -1.5560847131577804e-05
GC_2_508 b_2 NI_2 NS_508 0 -1.9131787682402759e-05
GC_2_509 b_2 NI_2 NS_509 0 -2.9829616559151911e-06
GC_2_510 b_2 NI_2 NS_510 0 5.0701953962194832e-06
GC_2_511 b_2 NI_2 NS_511 0 4.2041743023603063e-06
GC_2_512 b_2 NI_2 NS_512 0 -1.9025773224664296e-06
GC_2_513 b_2 NI_2 NS_513 0 -2.7722055034348729e-11
GC_2_514 b_2 NI_2 NS_514 0 5.4087853819111099e-12
GC_2_515 b_2 NI_2 NS_515 0 4.8942906611717730e-06
GC_2_516 b_2 NI_2 NS_516 0 -1.1671147140389076e-05
GC_2_517 b_2 NI_2 NS_517 0 -5.0227426463347653e-07
GC_2_518 b_2 NI_2 NS_518 0 2.7925967650250114e-06
GC_2_519 b_2 NI_2 NS_519 0 2.3625581383825972e-06
GC_2_520 b_2 NI_2 NS_520 0 -1.5932302746864846e-06
GC_2_521 b_2 NI_2 NS_521 0 2.1702322545798011e-06
GC_2_522 b_2 NI_2 NS_522 0 -9.8796052160840254e-06
GC_2_523 b_2 NI_2 NS_523 0 -1.0601719710009091e-05
GC_2_524 b_2 NI_2 NS_524 0 -3.5478351847340119e-06
GC_2_525 b_2 NI_2 NS_525 0 -2.2615902101428535e-10
GC_2_526 b_2 NI_2 NS_526 0 4.2340234659478055e-10
GC_2_527 b_2 NI_2 NS_527 0 -9.1524874679389915e-06
GC_2_528 b_2 NI_2 NS_528 0 -5.6556584272127806e-06
GC_2_529 b_2 NI_2 NS_529 0 2.0112931055641023e-06
GC_2_530 b_2 NI_2 NS_530 0 -6.6968698929928597e-06
GC_2_531 b_2 NI_2 NS_531 0 -3.3581515191916081e-06
GC_2_532 b_2 NI_2 NS_532 0 -1.8350317146664258e-07
GC_2_533 b_2 NI_2 NS_533 0 -8.5821414196137109e-06
GC_2_534 b_2 NI_2 NS_534 0 5.9057852029230802e-07
GC_2_535 b_2 NI_2 NS_535 0 2.6252866822582102e-06
GC_2_536 b_2 NI_2 NS_536 0 2.8291308586512676e-06
GC_2_537 b_2 NI_2 NS_537 0 1.0192572746453698e-06
GC_2_538 b_2 NI_2 NS_538 0 -3.7248594031091969e-06
GC_2_539 b_2 NI_2 NS_539 0 -5.3998924909666910e-06
GC_2_540 b_2 NI_2 NS_540 0 -4.2209438624270128e-06
GC_2_541 b_2 NI_2 NS_541 0 -5.3680148918507863e-05
GC_2_542 b_2 NI_2 NS_542 0 -6.9833890984395251e-12
GC_2_543 b_2 NI_2 NS_543 0 -2.0805242394142046e-10
GC_2_544 b_2 NI_2 NS_544 0 9.8195269689431029e-09
GC_2_545 b_2 NI_2 NS_545 0 5.4711420020554162e-07
GC_2_546 b_2 NI_2 NS_546 0 4.2979641221810599e-08
GC_2_547 b_2 NI_2 NS_547 0 2.9239402662686304e-06
GC_2_548 b_2 NI_2 NS_548 0 -1.5091403382315435e-06
GC_2_549 b_2 NI_2 NS_549 0 -3.2045440946769001e-06
GC_2_550 b_2 NI_2 NS_550 0 -2.6196626459764562e-06
GC_2_551 b_2 NI_2 NS_551 0 4.6037977989660501e-06
GC_2_552 b_2 NI_2 NS_552 0 -4.0622268036109197e-07
GC_2_553 b_2 NI_2 NS_553 0 -7.4630335363038579e-06
GC_2_554 b_2 NI_2 NS_554 0 -7.5110658663679312e-06
GC_2_555 b_2 NI_2 NS_555 0 -2.6104614285469585e-07
GC_2_556 b_2 NI_2 NS_556 0 -1.3674921167180174e-06
GC_2_557 b_2 NI_2 NS_557 0 -5.9022051450393476e-06
GC_2_558 b_2 NI_2 NS_558 0 2.4898542504364121e-06
GC_2_559 b_2 NI_2 NS_559 0 5.2248128844570150e-06
GC_2_560 b_2 NI_2 NS_560 0 -5.0757007729459463e-06
GC_2_561 b_2 NI_2 NS_561 0 -1.6698149014293829e-05
GC_2_562 b_2 NI_2 NS_562 0 5.0787233794060739e-06
GC_2_563 b_2 NI_2 NS_563 0 -1.1561006176557503e-06
GC_2_564 b_2 NI_2 NS_564 0 7.5339646385570131e-06
GC_2_565 b_2 NI_2 NS_565 0 -6.6315684809492327e-06
GC_2_566 b_2 NI_2 NS_566 0 -4.0455605144711167e-06
GC_2_567 b_2 NI_2 NS_567 0 -3.2762113619772893e-06
GC_2_568 b_2 NI_2 NS_568 0 8.3571835885538507e-06
GC_2_569 b_2 NI_2 NS_569 0 -1.2997326394665963e-06
GC_2_570 b_2 NI_2 NS_570 0 -4.1162266943387727e-06
GC_2_571 b_2 NI_2 NS_571 0 -4.0024793514721365e-06
GC_2_572 b_2 NI_2 NS_572 0 1.1510740089973521e-05
GC_2_573 b_2 NI_2 NS_573 0 -2.4919204434659386e-08
GC_2_574 b_2 NI_2 NS_574 0 7.6861978937888198e-06
GC_2_575 b_2 NI_2 NS_575 0 -3.6434499159561939e-06
GC_2_576 b_2 NI_2 NS_576 0 1.4544315758291052e-06
GC_2_577 b_2 NI_2 NS_577 0 -3.5977796240554267e-07
GC_2_578 b_2 NI_2 NS_578 0 8.4286792415002643e-06
GC_2_579 b_2 NI_2 NS_579 0 -5.7518764427415522e-07
GC_2_580 b_2 NI_2 NS_580 0 2.1383300461926783e-06
GC_2_581 b_2 NI_2 NS_581 0 -2.3055743211593522e-06
GC_2_582 b_2 NI_2 NS_582 0 8.5102689283654486e-06
GC_2_583 b_2 NI_2 NS_583 0 7.1416288937222019e-07
GC_2_584 b_2 NI_2 NS_584 0 9.9220600975978281e-06
GC_2_585 b_2 NI_2 NS_585 0 -7.2144955486400724e-07
GC_2_586 b_2 NI_2 NS_586 0 8.9744372920914628e-06
GC_2_587 b_2 NI_2 NS_587 0 -1.2319737328660207e-06
GC_2_588 b_2 NI_2 NS_588 0 4.0766588757546660e-06
GC_2_589 b_2 NI_2 NS_589 0 1.2869279991661903e-06
GC_2_590 b_2 NI_2 NS_590 0 1.2351987669226296e-05
GC_2_591 b_2 NI_2 NS_591 0 1.8775556970997107e-05
GC_2_592 b_2 NI_2 NS_592 0 1.7032811245905632e-05
GC_2_593 b_2 NI_2 NS_593 0 5.0360269554456945e-06
GC_2_594 b_2 NI_2 NS_594 0 7.9043932987977459e-06
GC_2_595 b_2 NI_2 NS_595 0 1.0383334512299281e-05
GC_2_596 b_2 NI_2 NS_596 0 3.9003797609757263e-06
GC_2_597 b_2 NI_2 NS_597 0 6.8650996833830896e-06
GC_2_598 b_2 NI_2 NS_598 0 1.1089491431996154e-05
GC_2_599 b_2 NI_2 NS_599 0 3.3649743751093911e-05
GC_2_600 b_2 NI_2 NS_600 0 -6.1820207246496883e-06
GC_2_601 b_2 NI_2 NS_601 0 8.2297386927206094e-06
GC_2_602 b_2 NI_2 NS_602 0 3.4992007200141556e-06
GC_2_603 b_2 NI_2 NS_603 0 1.2051430309704073e-05
GC_2_604 b_2 NI_2 NS_604 0 -1.0349766247841768e-05
GC_2_605 b_2 NI_2 NS_605 0 1.0852241982769824e-05
GC_2_606 b_2 NI_2 NS_606 0 6.5921150383941055e-06
GC_2_607 b_2 NI_2 NS_607 0 1.7121437770927938e-05
GC_2_608 b_2 NI_2 NS_608 0 -3.0976643221370809e-05
GC_2_609 b_2 NI_2 NS_609 0 8.1822977592515548e-06
GC_2_610 b_2 NI_2 NS_610 0 -2.9067682591994178e-06
GC_2_611 b_2 NI_2 NS_611 0 -3.1851360745655842e-06
GC_2_612 b_2 NI_2 NS_612 0 -1.6366048732522685e-05
GC_2_613 b_2 NI_2 NS_613 0 1.1873639163725063e-05
GC_2_614 b_2 NI_2 NS_614 0 -1.5391800324437953e-06
GC_2_615 b_2 NI_2 NS_615 0 -1.2633532187013224e-05
GC_2_616 b_2 NI_2 NS_616 0 -2.5267040209687112e-05
GC_2_617 b_2 NI_2 NS_617 0 -1.0375362211167122e-07
GC_2_618 b_2 NI_2 NS_618 0 -6.6315508796360722e-06
GC_2_619 b_2 NI_2 NS_619 0 -9.5776935861330427e-06
GC_2_620 b_2 NI_2 NS_620 0 -2.6846437585399511e-06
GC_2_621 b_2 NI_2 NS_621 0 1.0229010229634231e-10
GC_2_622 b_2 NI_2 NS_622 0 4.5737895256498577e-11
GC_2_623 b_2 NI_2 NS_623 0 1.5527387690105963e-06
GC_2_624 b_2 NI_2 NS_624 0 -4.6900203821407739e-06
GC_2_625 b_2 NI_2 NS_625 0 -1.3369744123422507e-06
GC_2_626 b_2 NI_2 NS_626 0 -1.3619262346034412e-06
GC_2_627 b_2 NI_2 NS_627 0 -4.8411289832191756e-06
GC_2_628 b_2 NI_2 NS_628 0 -1.0239410457651672e-06
GC_2_629 b_2 NI_2 NS_629 0 -1.0645238548729452e-06
GC_2_630 b_2 NI_2 NS_630 0 -2.7299682350110506e-06
GC_2_631 b_2 NI_2 NS_631 0 -9.9885535081012305e-06
GC_2_632 b_2 NI_2 NS_632 0 -4.1154654211191204e-06
GC_2_633 b_2 NI_2 NS_633 0 6.6961071601763567e-09
GC_2_634 b_2 NI_2 NS_634 0 5.4062567297803794e-09
GC_2_635 b_2 NI_2 NS_635 0 1.7786610493453163e-06
GC_2_636 b_2 NI_2 NS_636 0 4.4250622698061336e-07
GC_2_637 b_2 NI_2 NS_637 0 -1.5845644611654238e-06
GC_2_638 b_2 NI_2 NS_638 0 3.2301030030196001e-06
GC_2_639 b_2 NI_2 NS_639 0 -8.2746728581535882e-07
GC_2_640 b_2 NI_2 NS_640 0 6.9450322144797785e-07
GC_2_641 b_2 NI_2 NS_641 0 -7.6658750747788203e-06
GC_2_642 b_2 NI_2 NS_642 0 4.7706462351983550e-07
GC_2_643 b_2 NI_2 NS_643 0 -2.2026811037295904e-06
GC_2_644 b_2 NI_2 NS_644 0 1.9565058125547174e-06
GC_2_645 b_2 NI_2 NS_645 0 -2.0865320114532855e-06
GC_2_646 b_2 NI_2 NS_646 0 1.9644979924126693e-06
GC_2_647 b_2 NI_2 NS_647 0 1.2958344248134552e-06
GC_2_648 b_2 NI_2 NS_648 0 2.8412087143176768e-06
GC_2_649 b_2 NI_2 NS_649 0 -8.9827468083850589e-05
GC_2_650 b_2 NI_2 NS_650 0 3.3242388762782999e-12
GC_2_651 b_2 NI_2 NS_651 0 -4.3152816916174019e-11
GC_2_652 b_2 NI_2 NS_652 0 3.0280991730753974e-10
GC_2_653 b_2 NI_2 NS_653 0 -1.5652910975210236e-06
GC_2_654 b_2 NI_2 NS_654 0 -1.5563383539810244e-06
GC_2_655 b_2 NI_2 NS_655 0 9.4716896351500681e-07
GC_2_656 b_2 NI_2 NS_656 0 7.1437281944483234e-07
GC_2_657 b_2 NI_2 NS_657 0 -2.7263877785632212e-06
GC_2_658 b_2 NI_2 NS_658 0 3.0058182166188174e-06
GC_2_659 b_2 NI_2 NS_659 0 -3.0650219949577188e-06
GC_2_660 b_2 NI_2 NS_660 0 -2.5788312482720560e-06
GC_2_661 b_2 NI_2 NS_661 0 1.4936480411254476e-06
GC_2_662 b_2 NI_2 NS_662 0 1.1480593084388789e-07
GC_2_663 b_2 NI_2 NS_663 0 -1.6611499224799247e-06
GC_2_664 b_2 NI_2 NS_664 0 1.7822125321512191e-06
GC_2_665 b_2 NI_2 NS_665 0 8.5990102132008360e-07
GC_2_666 b_2 NI_2 NS_666 0 4.1352244838465338e-06
GC_2_667 b_2 NI_2 NS_667 0 -4.3810577929588096e-06
GC_2_668 b_2 NI_2 NS_668 0 -1.9846182233964798e-06
GC_2_669 b_2 NI_2 NS_669 0 2.4929774276254572e-06
GC_2_670 b_2 NI_2 NS_670 0 -1.8455304248686424e-06
GC_2_671 b_2 NI_2 NS_671 0 -1.1634626127984459e-06
GC_2_672 b_2 NI_2 NS_672 0 3.2977038671005872e-06
GC_2_673 b_2 NI_2 NS_673 0 -8.1358031374312896e-06
GC_2_674 b_2 NI_2 NS_674 0 1.1093584760801024e-05
GC_2_675 b_2 NI_2 NS_675 0 1.2697843626668844e-06
GC_2_676 b_2 NI_2 NS_676 0 -1.6862485305155529e-06
GC_2_677 b_2 NI_2 NS_677 0 9.8771713689990207e-06
GC_2_678 b_2 NI_2 NS_678 0 1.6972999014487681e-05
GC_2_679 b_2 NI_2 NS_679 0 -7.1199368189717621e-07
GC_2_680 b_2 NI_2 NS_680 0 -4.4201291242784158e-07
GC_2_681 b_2 NI_2 NS_681 0 4.0869143639958436e-07
GC_2_682 b_2 NI_2 NS_682 0 -1.4042434840785583e-06
GC_2_683 b_2 NI_2 NS_683 0 6.8711702234450113e-06
GC_2_684 b_2 NI_2 NS_684 0 -1.2534677617471113e-07
GC_2_685 b_2 NI_2 NS_685 0 7.0588007212297565e-07
GC_2_686 b_2 NI_2 NS_686 0 3.0247964121506604e-06
GC_2_687 b_2 NI_2 NS_687 0 5.1851343432709852e-07
GC_2_688 b_2 NI_2 NS_688 0 2.8703473613948622e-06
GC_2_689 b_2 NI_2 NS_689 0 1.1686964565936318e-06
GC_2_690 b_2 NI_2 NS_690 0 -1.4312841411903238e-06
GC_2_691 b_2 NI_2 NS_691 0 9.2306188248958126e-06
GC_2_692 b_2 NI_2 NS_692 0 5.0868136459615429e-06
GC_2_693 b_2 NI_2 NS_693 0 5.3876456987471382e-07
GC_2_694 b_2 NI_2 NS_694 0 1.1688118005202273e-06
GC_2_695 b_2 NI_2 NS_695 0 4.7181770037985700e-08
GC_2_696 b_2 NI_2 NS_696 0 4.6163535883103090e-07
GC_2_697 b_2 NI_2 NS_697 0 1.2781453000993395e-06
GC_2_698 b_2 NI_2 NS_698 0 -8.5245090866915243e-07
GC_2_699 b_2 NI_2 NS_699 0 9.0033515432507473e-06
GC_2_700 b_2 NI_2 NS_700 0 7.1340603177595024e-07
GC_2_701 b_2 NI_2 NS_701 0 8.3038762750384371e-07
GC_2_702 b_2 NI_2 NS_702 0 1.4741772378198283e-06
GC_2_703 b_2 NI_2 NS_703 0 1.0390721096933457e-06
GC_2_704 b_2 NI_2 NS_704 0 6.2172567302981309e-07
GC_2_705 b_2 NI_2 NS_705 0 1.3551387413034891e-06
GC_2_706 b_2 NI_2 NS_706 0 -9.5010633379826864e-07
GC_2_707 b_2 NI_2 NS_707 0 7.9167086642955705e-06
GC_2_708 b_2 NI_2 NS_708 0 -2.0394105896414073e-06
GC_2_709 b_2 NI_2 NS_709 0 1.1753922149180199e-06
GC_2_710 b_2 NI_2 NS_710 0 1.5633839077602338e-06
GC_2_711 b_2 NI_2 NS_711 0 1.6188827790092419e-06
GC_2_712 b_2 NI_2 NS_712 0 -2.2250201100245137e-07
GC_2_713 b_2 NI_2 NS_713 0 1.3149917611376081e-06
GC_2_714 b_2 NI_2 NS_714 0 -9.9060498971953319e-07
GC_2_715 b_2 NI_2 NS_715 0 5.7974609435553820e-06
GC_2_716 b_2 NI_2 NS_716 0 -3.8075746014400229e-06
GC_2_717 b_2 NI_2 NS_717 0 1.8131060124394818e-06
GC_2_718 b_2 NI_2 NS_718 0 1.4425458892991014e-06
GC_2_719 b_2 NI_2 NS_719 0 1.1283349717535107e-06
GC_2_720 b_2 NI_2 NS_720 0 -1.3977641256769866e-06
GC_2_721 b_2 NI_2 NS_721 0 1.4102958481908516e-06
GC_2_722 b_2 NI_2 NS_722 0 -1.1060929479851104e-06
GC_2_723 b_2 NI_2 NS_723 0 2.9944053187759162e-06
GC_2_724 b_2 NI_2 NS_724 0 -4.1483178427597037e-06
GC_2_725 b_2 NI_2 NS_725 0 2.2296565583187967e-06
GC_2_726 b_2 NI_2 NS_726 0 3.1298529299200520e-07
GC_2_727 b_2 NI_2 NS_727 0 -3.1154060950536583e-07
GC_2_728 b_2 NI_2 NS_728 0 -1.1926002544107613e-06
GC_2_729 b_2 NI_2 NS_729 0 2.5423235012407930e-11
GC_2_730 b_2 NI_2 NS_730 0 -4.1101372456919574e-11
GC_2_731 b_2 NI_2 NS_731 0 8.0347366981199437e-07
GC_2_732 b_2 NI_2 NS_732 0 -1.5695283080541707e-06
GC_2_733 b_2 NI_2 NS_733 0 1.2661376925616862e-06
GC_2_734 b_2 NI_2 NS_734 0 2.2070185928085424e-07
GC_2_735 b_2 NI_2 NS_735 0 1.6021715491726533e-07
GC_2_736 b_2 NI_2 NS_736 0 -5.5094559320927357e-07
GC_2_737 b_2 NI_2 NS_737 0 5.5034160022115000e-07
GC_2_738 b_2 NI_2 NS_738 0 -8.6165088569733382e-07
GC_2_739 b_2 NI_2 NS_739 0 1.3129429368564499e-06
GC_2_740 b_2 NI_2 NS_740 0 -2.0695656031951000e-06
GC_2_741 b_2 NI_2 NS_741 0 4.8974761356722538e-10
GC_2_742 b_2 NI_2 NS_742 0 -1.2287954004229491e-09
GC_2_743 b_2 NI_2 NS_743 0 5.5017531752595661e-07
GC_2_744 b_2 NI_2 NS_744 0 -8.6030227580424755e-07
GC_2_745 b_2 NI_2 NS_745 0 7.1448111508134015e-07
GC_2_746 b_2 NI_2 NS_746 0 -9.5257238884992228e-07
GC_2_747 b_2 NI_2 NS_747 0 9.1157448155551550e-08
GC_2_748 b_2 NI_2 NS_748 0 4.9897344545016035e-08
GC_2_749 b_2 NI_2 NS_749 0 1.3758223121093978e-06
GC_2_750 b_2 NI_2 NS_750 0 -1.2408293087170797e-06
GC_2_751 b_2 NI_2 NS_751 0 1.6631100862632038e-06
GC_2_752 b_2 NI_2 NS_752 0 -3.1895778366467009e-07
GC_2_753 b_2 NI_2 NS_753 0 -2.4124534813619705e-07
GC_2_754 b_2 NI_2 NS_754 0 -7.4502411307049133e-07
GC_2_755 b_2 NI_2 NS_755 0 7.3810203011955735e-07
GC_2_756 b_2 NI_2 NS_756 0 2.9282314616645471e-07
GC_2_757 b_2 NI_2 NS_757 0 4.7631967211169404e-05
GC_2_758 b_2 NI_2 NS_758 0 7.4845184748417771e-12
GC_2_759 b_2 NI_2 NS_759 0 -1.8841428462713639e-11
GC_2_760 b_2 NI_2 NS_760 0 9.9252948208562532e-10
GC_2_761 b_2 NI_2 NS_761 0 -6.5468917747166326e-08
GC_2_762 b_2 NI_2 NS_762 0 2.4788335269587764e-07
GC_2_763 b_2 NI_2 NS_763 0 2.2310538344480537e-07
GC_2_764 b_2 NI_2 NS_764 0 4.0419327282969437e-07
GC_2_765 b_2 NI_2 NS_765 0 -1.7538224384143338e-07
GC_2_766 b_2 NI_2 NS_766 0 2.7605816883567987e-07
GC_2_767 b_2 NI_2 NS_767 0 7.2646981302421024e-07
GC_2_768 b_2 NI_2 NS_768 0 1.4718717419413265e-06
GC_2_769 b_2 NI_2 NS_769 0 1.0323109138538557e-06
GC_2_770 b_2 NI_2 NS_770 0 -4.2531107468690361e-07
GC_2_771 b_2 NI_2 NS_771 0 3.0287118778673699e-07
GC_2_772 b_2 NI_2 NS_772 0 9.1872025476586388e-07
GC_2_773 b_2 NI_2 NS_773 0 7.8010433398637654e-07
GC_2_774 b_2 NI_2 NS_774 0 -3.1455707642790671e-07
GC_2_775 b_2 NI_2 NS_775 0 4.3375164702701631e-06
GC_2_776 b_2 NI_2 NS_776 0 1.5052412022989740e-06
GC_2_777 b_2 NI_2 NS_777 0 -1.5165560267163152e-06
GC_2_778 b_2 NI_2 NS_778 0 -3.5706885586724622e-06
GC_2_779 b_2 NI_2 NS_779 0 2.4327997497182536e-07
GC_2_780 b_2 NI_2 NS_780 0 1.5795052183834780e-06
GC_2_781 b_2 NI_2 NS_781 0 3.1040271575717472e-06
GC_2_782 b_2 NI_2 NS_782 0 -4.6709510655039919e-06
GC_2_783 b_2 NI_2 NS_783 0 -7.4669661283175022e-07
GC_2_784 b_2 NI_2 NS_784 0 5.6972901705695263e-07
GC_2_785 b_2 NI_2 NS_785 0 5.7308732371598993e-06
GC_2_786 b_2 NI_2 NS_786 0 -5.7318871579747926e-06
GC_2_787 b_2 NI_2 NS_787 0 -3.3217238130045424e-06
GC_2_788 b_2 NI_2 NS_788 0 1.7569737519535379e-06
GC_2_789 b_2 NI_2 NS_789 0 8.8313631327707197e-07
GC_2_790 b_2 NI_2 NS_790 0 1.2588766235932832e-06
GC_2_791 b_2 NI_2 NS_791 0 1.6940415339634784e-06
GC_2_792 b_2 NI_2 NS_792 0 -4.0841763153681260e-06
GC_2_793 b_2 NI_2 NS_793 0 6.1060205423306521e-07
GC_2_794 b_2 NI_2 NS_794 0 2.1519043228951638e-07
GC_2_795 b_2 NI_2 NS_795 0 2.5345194552140135e-07
GC_2_796 b_2 NI_2 NS_796 0 -4.0636606842269682e-06
GC_2_797 b_2 NI_2 NS_797 0 -1.5617933837542172e-07
GC_2_798 b_2 NI_2 NS_798 0 1.7811619097919468e-07
GC_2_799 b_2 NI_2 NS_799 0 4.7913304011945142e-06
GC_2_800 b_2 NI_2 NS_800 0 -6.3202229303396484e-06
GC_2_801 b_2 NI_2 NS_801 0 -1.7962215285876295e-06
GC_2_802 b_2 NI_2 NS_802 0 -1.3136346625103587e-06
GC_2_803 b_2 NI_2 NS_803 0 1.4000600174780987e-06
GC_2_804 b_2 NI_2 NS_804 0 -1.1889559188322494e-06
GC_2_805 b_2 NI_2 NS_805 0 4.3422459042924698e-07
GC_2_806 b_2 NI_2 NS_806 0 -2.1045341564048078e-06
GC_2_807 b_2 NI_2 NS_807 0 -1.3395086610239982e-06
GC_2_808 b_2 NI_2 NS_808 0 -1.1872484907843843e-05
GC_2_809 b_2 NI_2 NS_809 0 -2.2432650101201733e-06
GC_2_810 b_2 NI_2 NS_810 0 -1.7314843809664899e-06
GC_2_811 b_2 NI_2 NS_811 0 -2.3524777991959496e-06
GC_2_812 b_2 NI_2 NS_812 0 -4.0390076862698562e-06
GC_2_813 b_2 NI_2 NS_813 0 -1.4499765319380358e-06
GC_2_814 b_2 NI_2 NS_814 0 -2.4370093373296220e-06
GC_2_815 b_2 NI_2 NS_815 0 -1.0683069914011476e-05
GC_2_816 b_2 NI_2 NS_816 0 -7.2200570971946704e-06
GC_2_817 b_2 NI_2 NS_817 0 -3.1781717162869398e-06
GC_2_818 b_2 NI_2 NS_818 0 -8.7729185586018519e-07
GC_2_819 b_2 NI_2 NS_819 0 -5.7541059756425336e-06
GC_2_820 b_2 NI_2 NS_820 0 -4.1607477118385378e-07
GC_2_821 b_2 NI_2 NS_821 0 -3.0997358080529845e-06
GC_2_822 b_2 NI_2 NS_822 0 -1.7555841183882858e-06
GC_2_823 b_2 NI_2 NS_823 0 -1.0627585456873123e-05
GC_2_824 b_2 NI_2 NS_824 0 3.2953775393521609e-06
GC_2_825 b_2 NI_2 NS_825 0 -3.6183714574175445e-06
GC_2_826 b_2 NI_2 NS_826 0 8.1870300191568695e-07
GC_2_827 b_2 NI_2 NS_827 0 -2.8814468519269859e-06
GC_2_828 b_2 NI_2 NS_828 0 3.9140068782209620e-06
GC_2_829 b_2 NI_2 NS_829 0 -4.3309340116361066e-06
GC_2_830 b_2 NI_2 NS_830 0 1.7127372693529064e-07
GC_2_831 b_2 NI_2 NS_831 0 -1.8671475711621386e-06
GC_2_832 b_2 NI_2 NS_832 0 7.2126083373818885e-06
GC_2_833 b_2 NI_2 NS_833 0 -1.5633431934076137e-06
GC_2_834 b_2 NI_2 NS_834 0 2.7935670736713233e-06
GC_2_835 b_2 NI_2 NS_835 0 9.2396525160328970e-07
GC_2_836 b_2 NI_2 NS_836 0 1.8140040965059768e-06
GC_2_837 b_2 NI_2 NS_837 0 -3.0213683703323362e-11
GC_2_838 b_2 NI_2 NS_838 0 -3.9931407287309175e-12
GC_2_839 b_2 NI_2 NS_839 0 -1.7134382661104784e-06
GC_2_840 b_2 NI_2 NS_840 0 2.1404406734212688e-06
GC_2_841 b_2 NI_2 NS_841 0 -3.2436348444069431e-07
GC_2_842 b_2 NI_2 NS_842 0 1.0487455156694508e-06
GC_2_843 b_2 NI_2 NS_843 0 1.4400269415284230e-07
GC_2_844 b_2 NI_2 NS_844 0 6.2111555074067658e-07
GC_2_845 b_2 NI_2 NS_845 0 -1.0462325207281919e-06
GC_2_846 b_2 NI_2 NS_846 0 1.2710924290666532e-06
GC_2_847 b_2 NI_2 NS_847 0 9.7965226657001122e-07
GC_2_848 b_2 NI_2 NS_848 0 1.8189637173085212e-06
GC_2_849 b_2 NI_2 NS_849 0 -1.5165329109324390e-09
GC_2_850 b_2 NI_2 NS_850 0 -7.8078247529220138e-10
GC_2_851 b_2 NI_2 NS_851 0 -4.8470485227436257e-07
GC_2_852 b_2 NI_2 NS_852 0 -2.7510956096647908e-08
GC_2_853 b_2 NI_2 NS_853 0 -3.1050717334027580e-07
GC_2_854 b_2 NI_2 NS_854 0 1.7476044163326472e-07
GC_2_855 b_2 NI_2 NS_855 0 -5.5079980901020085e-07
GC_2_856 b_2 NI_2 NS_856 0 1.5190552017230558e-07
GC_2_857 b_2 NI_2 NS_857 0 6.6424982604752738e-07
GC_2_858 b_2 NI_2 NS_858 0 8.1076613420865270e-07
GC_2_859 b_2 NI_2 NS_859 0 2.1776812687208374e-07
GC_2_860 b_2 NI_2 NS_860 0 6.9571018535766756e-07
GC_2_861 b_2 NI_2 NS_861 0 1.0940401563117955e-08
GC_2_862 b_2 NI_2 NS_862 0 -1.3810931503120307e-07
GC_2_863 b_2 NI_2 NS_863 0 -3.4771225928816090e-07
GC_2_864 b_2 NI_2 NS_864 0 2.9453656932721368e-07
GC_2_865 b_2 NI_2 NS_865 0 -6.4269092628253203e-05
GC_2_866 b_2 NI_2 NS_866 0 3.5608406934374015e-12
GC_2_867 b_2 NI_2 NS_867 0 5.0181514078696002e-11
GC_2_868 b_2 NI_2 NS_868 0 -1.5818276212038676e-09
GC_2_869 b_2 NI_2 NS_869 0 -1.0723782699604021e-06
GC_2_870 b_2 NI_2 NS_870 0 -1.0588571026391746e-06
GC_2_871 b_2 NI_2 NS_871 0 4.0966366695342191e-07
GC_2_872 b_2 NI_2 NS_872 0 3.5700932894109992e-07
GC_2_873 b_2 NI_2 NS_873 0 -2.2606362745160545e-06
GC_2_874 b_2 NI_2 NS_874 0 2.1080746227810320e-06
GC_2_875 b_2 NI_2 NS_875 0 -2.5321214514125417e-06
GC_2_876 b_2 NI_2 NS_876 0 -1.2387521298054199e-06
GC_2_877 b_2 NI_2 NS_877 0 1.3985158302281725e-06
GC_2_878 b_2 NI_2 NS_878 0 9.9856745625617237e-07
GC_2_879 b_2 NI_2 NS_879 0 -1.1234359115194083e-06
GC_2_880 b_2 NI_2 NS_880 0 1.3407147876607138e-06
GC_2_881 b_2 NI_2 NS_881 0 7.2716643962069052e-07
GC_2_882 b_2 NI_2 NS_882 0 3.0410821181981169e-06
GC_2_883 b_2 NI_2 NS_883 0 -2.8465638675320721e-06
GC_2_884 b_2 NI_2 NS_884 0 4.7261201386732017e-07
GC_2_885 b_2 NI_2 NS_885 0 3.6885489202302895e-06
GC_2_886 b_2 NI_2 NS_886 0 -2.0179826469499808e-06
GC_2_887 b_2 NI_2 NS_887 0 -1.8785557096617489e-07
GC_2_888 b_2 NI_2 NS_888 0 2.5632246650593485e-06
GC_2_889 b_2 NI_2 NS_889 0 -4.0642264071974584e-06
GC_2_890 b_2 NI_2 NS_890 0 4.8362694060220626e-06
GC_2_891 b_2 NI_2 NS_891 0 6.4243496159519318e-07
GC_2_892 b_2 NI_2 NS_892 0 -1.5864767827387881e-06
GC_2_893 b_2 NI_2 NS_893 0 4.6099971557655398e-06
GC_2_894 b_2 NI_2 NS_894 0 9.9431092317207427e-06
GC_2_895 b_2 NI_2 NS_895 0 -1.1100938602049560e-07
GC_2_896 b_2 NI_2 NS_896 0 5.2381783863710291e-07
GC_2_897 b_2 NI_2 NS_897 0 -6.3538796392971496e-09
GC_2_898 b_2 NI_2 NS_898 0 -7.8555928612125367e-07
GC_2_899 b_2 NI_2 NS_899 0 5.3519103420519223e-06
GC_2_900 b_2 NI_2 NS_900 0 4.9535139138572908e-07
GC_2_901 b_2 NI_2 NS_901 0 8.4640881472673305e-07
GC_2_902 b_2 NI_2 NS_902 0 1.9176171516763559e-06
GC_2_903 b_2 NI_2 NS_903 0 3.0833320891232296e-08
GC_2_904 b_2 NI_2 NS_904 0 1.1331864978723540e-06
GC_2_905 b_2 NI_2 NS_905 0 5.8507601778278788e-07
GC_2_906 b_2 NI_2 NS_906 0 -1.1108574297628668e-06
GC_2_907 b_2 NI_2 NS_907 0 5.8253822749684695e-06
GC_2_908 b_2 NI_2 NS_908 0 4.0748118360952951e-06
GC_2_909 b_2 NI_2 NS_909 0 6.0627970101075105e-07
GC_2_910 b_2 NI_2 NS_910 0 8.5953121070053967e-07
GC_2_911 b_2 NI_2 NS_911 0 1.9692893426054382e-07
GC_2_912 b_2 NI_2 NS_912 0 2.4097972380520093e-07
GC_2_913 b_2 NI_2 NS_913 0 8.4525729703706317e-07
GC_2_914 b_2 NI_2 NS_914 0 -6.7218108376738187e-07
GC_2_915 b_2 NI_2 NS_915 0 6.6650749215095394e-06
GC_2_916 b_2 NI_2 NS_916 0 7.5449015724542241e-07
GC_2_917 b_2 NI_2 NS_917 0 7.7455796337469608e-07
GC_2_918 b_2 NI_2 NS_918 0 7.4913720248292653e-07
GC_2_919 b_2 NI_2 NS_919 0 6.6483736001556071e-07
GC_2_920 b_2 NI_2 NS_920 0 -6.6211269594495361e-08
GC_2_921 b_2 NI_2 NS_921 0 8.7154192574259609e-07
GC_2_922 b_2 NI_2 NS_922 0 -6.4040101410243955e-07
GC_2_923 b_2 NI_2 NS_923 0 5.7751839948254314e-06
GC_2_924 b_2 NI_2 NS_924 0 -1.5909509344961629e-06
GC_2_925 b_2 NI_2 NS_925 0 8.2383155437985982e-07
GC_2_926 b_2 NI_2 NS_926 0 5.6703933565284397e-07
GC_2_927 b_2 NI_2 NS_927 0 6.2584013262323562e-07
GC_2_928 b_2 NI_2 NS_928 0 -5.5330933463191563e-07
GC_2_929 b_2 NI_2 NS_929 0 9.3776460874447493e-07
GC_2_930 b_2 NI_2 NS_930 0 -4.4580251940547866e-07
GC_2_931 b_2 NI_2 NS_931 0 3.9036758157894758e-06
GC_2_932 b_2 NI_2 NS_932 0 -2.9906819507770748e-06
GC_2_933 b_2 NI_2 NS_933 0 8.9572281240235294e-07
GC_2_934 b_2 NI_2 NS_934 0 3.2737878629660738e-07
GC_2_935 b_2 NI_2 NS_935 0 2.1610615748314066e-07
GC_2_936 b_2 NI_2 NS_936 0 -7.9557897123551339e-07
GC_2_937 b_2 NI_2 NS_937 0 1.1598899640331187e-06
GC_2_938 b_2 NI_2 NS_938 0 -3.2475253085540276e-07
GC_2_939 b_2 NI_2 NS_939 0 1.6774751361372448e-06
GC_2_940 b_2 NI_2 NS_940 0 -3.0902015968516628e-06
GC_2_941 b_2 NI_2 NS_941 0 7.9113685686455224e-07
GC_2_942 b_2 NI_2 NS_942 0 -1.0639338682710535e-07
GC_2_943 b_2 NI_2 NS_943 0 -1.9702242485336103e-07
GC_2_944 b_2 NI_2 NS_944 0 -4.0861369463894068e-07
GC_2_945 b_2 NI_2 NS_945 0 8.5879931557846641e-12
GC_2_946 b_2 NI_2 NS_946 0 -1.5730252519887665e-11
GC_2_947 b_2 NI_2 NS_947 0 8.3871903948815762e-07
GC_2_948 b_2 NI_2 NS_948 0 -5.9378051126155802e-07
GC_2_949 b_2 NI_2 NS_949 0 4.9464458870302777e-07
GC_2_950 b_2 NI_2 NS_950 0 -3.5993947725900411e-08
GC_2_951 b_2 NI_2 NS_951 0 1.7009729198001391e-08
GC_2_952 b_2 NI_2 NS_952 0 -8.9112184055742712e-08
GC_2_953 b_2 NI_2 NS_953 0 5.2142197188677951e-07
GC_2_954 b_2 NI_2 NS_954 0 -1.7667516491162101e-08
GC_2_955 b_2 NI_2 NS_955 0 7.0518044516258357e-07
GC_2_956 b_2 NI_2 NS_956 0 -1.5614003193223022e-06
GC_2_957 b_2 NI_2 NS_957 0 4.0969060627040163e-10
GC_2_958 b_2 NI_2 NS_958 0 -5.8070619298653978e-10
GC_2_959 b_2 NI_2 NS_959 0 1.0099567738810058e-06
GC_2_960 b_2 NI_2 NS_960 0 -2.7386378669318229e-07
GC_2_961 b_2 NI_2 NS_961 0 3.5400718244926328e-07
GC_2_962 b_2 NI_2 NS_962 0 -1.7369760227443887e-07
GC_2_963 b_2 NI_2 NS_963 0 2.5492754540144677e-07
GC_2_964 b_2 NI_2 NS_964 0 2.6554722141477669e-08
GC_2_965 b_2 NI_2 NS_965 0 1.0857942061550350e-06
GC_2_966 b_2 NI_2 NS_966 0 -1.1750267745720936e-06
GC_2_967 b_2 NI_2 NS_967 0 6.5375615807763627e-07
GC_2_968 b_2 NI_2 NS_968 0 -3.3455315114027505e-07
GC_2_969 b_2 NI_2 NS_969 0 -2.1221673335596836e-07
GC_2_970 b_2 NI_2 NS_970 0 -9.8558054621562662e-08
GC_2_971 b_2 NI_2 NS_971 0 7.5732176357716613e-07
GC_2_972 b_2 NI_2 NS_972 0 3.2283786323913744e-07
GC_2_973 b_2 NI_2 NS_973 0 8.6319239668171558e-06
GC_2_974 b_2 NI_2 NS_974 0 3.7625738811611550e-12
GC_2_975 b_2 NI_2 NS_975 0 -7.8512210792112541e-11
GC_2_976 b_2 NI_2 NS_976 0 2.5462456855673132e-09
GC_2_977 b_2 NI_2 NS_977 0 1.6079122184073875e-08
GC_2_978 b_2 NI_2 NS_978 0 -8.4902434808340893e-08
GC_2_979 b_2 NI_2 NS_979 0 -2.4705995134384564e-07
GC_2_980 b_2 NI_2 NS_980 0 2.7069003967134670e-07
GC_2_981 b_2 NI_2 NS_981 0 7.4260412219869012e-07
GC_2_982 b_2 NI_2 NS_982 0 -2.8637944563746641e-07
GC_2_983 b_2 NI_2 NS_983 0 -9.6682268060897678e-07
GC_2_984 b_2 NI_2 NS_984 0 -2.3726250224732226e-07
GC_2_985 b_2 NI_2 NS_985 0 1.0246327538233228e-06
GC_2_986 b_2 NI_2 NS_986 0 3.9650951922694945e-07
GC_2_987 b_2 NI_2 NS_987 0 -1.1998889647043288e-07
GC_2_988 b_2 NI_2 NS_988 0 -2.7403626654674282e-07
GC_2_989 b_2 NI_2 NS_989 0 1.0759529442381578e-07
GC_2_990 b_2 NI_2 NS_990 0 -5.1241292923312745e-07
GC_2_991 b_2 NI_2 NS_991 0 -2.0819735050443634e-06
GC_2_992 b_2 NI_2 NS_992 0 8.5957045050781611e-07
GC_2_993 b_2 NI_2 NS_993 0 2.4262767128568447e-06
GC_2_994 b_2 NI_2 NS_994 0 -6.0722251583277222e-07
GC_2_995 b_2 NI_2 NS_995 0 -6.6432106432316933e-07
GC_2_996 b_2 NI_2 NS_996 0 -1.3962518540964886e-06
GC_2_997 b_2 NI_2 NS_997 0 4.2621836416800958e-07
GC_2_998 b_2 NI_2 NS_998 0 1.8418704456912199e-06
GC_2_999 b_2 NI_2 NS_999 0 -3.2462193796712085e-08
GC_2_1000 b_2 NI_2 NS_1000 0 -1.3222089130024778e-06
GC_2_1001 b_2 NI_2 NS_1001 0 -6.3303673300800601e-07
GC_2_1002 b_2 NI_2 NS_1002 0 2.5875889208784986e-06
GC_2_1003 b_2 NI_2 NS_1003 0 4.5137924751336441e-07
GC_2_1004 b_2 NI_2 NS_1004 0 -2.2404791696986206e-06
GC_2_1005 b_2 NI_2 NS_1005 0 -7.9996206319866257e-07
GC_2_1006 b_2 NI_2 NS_1006 0 -9.3018042260180963e-07
GC_2_1007 b_2 NI_2 NS_1007 0 3.5769664718248218e-07
GC_2_1008 b_2 NI_2 NS_1008 0 9.1028105253903247e-07
GC_2_1009 b_2 NI_2 NS_1009 0 -5.5738521278485627e-07
GC_2_1010 b_2 NI_2 NS_1010 0 -7.2412991612391158e-07
GC_2_1011 b_2 NI_2 NS_1011 0 4.7554902722723841e-07
GC_2_1012 b_2 NI_2 NS_1012 0 7.3859787623895480e-07
GC_2_1013 b_2 NI_2 NS_1013 0 -1.7484843260658391e-07
GC_2_1014 b_2 NI_2 NS_1014 0 -8.7651974915068891e-07
GC_2_1015 b_2 NI_2 NS_1015 0 -3.3814247393909940e-07
GC_2_1016 b_2 NI_2 NS_1016 0 1.1560695489137161e-06
GC_2_1017 b_2 NI_2 NS_1017 0 2.5205990216550691e-07
GC_2_1018 b_2 NI_2 NS_1018 0 -8.4271732187995356e-07
GC_2_1019 b_2 NI_2 NS_1019 0 -6.4710312475756564e-08
GC_2_1020 b_2 NI_2 NS_1020 0 6.6992795528361729e-08
GC_2_1021 b_2 NI_2 NS_1021 0 -2.6027266487143805e-07
GC_2_1022 b_2 NI_2 NS_1022 0 -5.4871439342483016e-07
GC_2_1023 b_2 NI_2 NS_1023 0 1.8495503957512165e-07
GC_2_1024 b_2 NI_2 NS_1024 0 7.1500832625097783e-07
GC_2_1025 b_2 NI_2 NS_1025 0 -8.1315650366532080e-08
GC_2_1026 b_2 NI_2 NS_1026 0 -6.3403653700625403e-07
GC_2_1027 b_2 NI_2 NS_1027 0 1.0163446187314390e-07
GC_2_1028 b_2 NI_2 NS_1028 0 1.0359706185105970e-07
GC_2_1029 b_2 NI_2 NS_1029 0 -2.9116962363753871e-07
GC_2_1030 b_2 NI_2 NS_1030 0 -5.9231303199042808e-07
GC_2_1031 b_2 NI_2 NS_1031 0 1.5984706379636336e-07
GC_2_1032 b_2 NI_2 NS_1032 0 2.2926874095312133e-07
GC_2_1033 b_2 NI_2 NS_1033 0 -2.5752755371262594e-07
GC_2_1034 b_2 NI_2 NS_1034 0 -5.0661427038115576e-07
GC_2_1035 b_2 NI_2 NS_1035 0 4.7616359965993490e-08
GC_2_1036 b_2 NI_2 NS_1036 0 -4.9953552374349561e-08
GC_2_1037 b_2 NI_2 NS_1037 0 -3.6863259072414881e-07
GC_2_1038 b_2 NI_2 NS_1038 0 -5.5617336543789011e-07
GC_2_1039 b_2 NI_2 NS_1039 0 -2.3513370721663774e-07
GC_2_1040 b_2 NI_2 NS_1040 0 2.1281484805818312e-08
GC_2_1041 b_2 NI_2 NS_1041 0 -4.3378983351412353e-07
GC_2_1042 b_2 NI_2 NS_1042 0 -3.3905174856867897e-07
GC_2_1043 b_2 NI_2 NS_1043 0 -1.2438512688947321e-07
GC_2_1044 b_2 NI_2 NS_1044 0 1.6436495466990805e-08
GC_2_1045 b_2 NI_2 NS_1045 0 -5.6302285171167278e-07
GC_2_1046 b_2 NI_2 NS_1046 0 -4.3710301771149704e-07
GC_2_1047 b_2 NI_2 NS_1047 0 -3.1810682541383807e-07
GC_2_1048 b_2 NI_2 NS_1048 0 3.1491338738510486e-07
GC_2_1049 b_2 NI_2 NS_1049 0 -4.9916041756513076e-07
GC_2_1050 b_2 NI_2 NS_1050 0 3.8171750508580279e-08
GC_2_1051 b_2 NI_2 NS_1051 0 -1.1417308030734969e-08
GC_2_1052 b_2 NI_2 NS_1052 0 6.1722029437335553e-08
GC_2_1053 b_2 NI_2 NS_1053 0 -3.2599618526275623e-12
GC_2_1054 b_2 NI_2 NS_1054 0 3.2063195259332840e-12
GC_2_1055 b_2 NI_2 NS_1055 0 -5.7550681637799765e-07
GC_2_1056 b_2 NI_2 NS_1056 0 4.7702822098232909e-08
GC_2_1057 b_2 NI_2 NS_1057 0 -2.8964044819166363e-07
GC_2_1058 b_2 NI_2 NS_1058 0 1.1817129868178611e-07
GC_2_1059 b_2 NI_2 NS_1059 0 -6.6619936328457415e-09
GC_2_1060 b_2 NI_2 NS_1060 0 -6.8741047558722803e-08
GC_2_1061 b_2 NI_2 NS_1061 0 -6.6032069327273894e-07
GC_2_1062 b_2 NI_2 NS_1062 0 1.4099350408295729e-07
GC_2_1063 b_2 NI_2 NS_1063 0 2.8402088883853708e-08
GC_2_1064 b_2 NI_2 NS_1064 0 1.2370025882417019e-07
GC_2_1065 b_2 NI_2 NS_1065 0 -6.1319778457243189e-11
GC_2_1066 b_2 NI_2 NS_1066 0 1.2860108091953063e-10
GC_2_1067 b_2 NI_2 NS_1067 0 -3.4592603838805253e-08
GC_2_1068 b_2 NI_2 NS_1068 0 1.9617178166767861e-07
GC_2_1069 b_2 NI_2 NS_1069 0 -3.6672498889331957e-07
GC_2_1070 b_2 NI_2 NS_1070 0 -4.3542182269177626e-08
GC_2_1071 b_2 NI_2 NS_1071 0 -1.8660687519087212e-07
GC_2_1072 b_2 NI_2 NS_1072 0 -2.4842575704888162e-09
GC_2_1073 b_2 NI_2 NS_1073 0 1.9220361337150877e-07
GC_2_1074 b_2 NI_2 NS_1074 0 8.1573257487476201e-08
GC_2_1075 b_2 NI_2 NS_1075 0 -2.6531311879155728e-07
GC_2_1076 b_2 NI_2 NS_1076 0 3.1380216125374722e-07
GC_2_1077 b_2 NI_2 NS_1077 0 1.2493604919903394e-07
GC_2_1078 b_2 NI_2 NS_1078 0 -1.4405378303049769e-07
GC_2_1079 b_2 NI_2 NS_1079 0 -5.7943637891672715e-08
GC_2_1080 b_2 NI_2 NS_1080 0 2.3859210183219623e-07
GC_2_1081 b_2 NI_2 NS_1081 0 -2.9908322173509678e-05
GC_2_1082 b_2 NI_2 NS_1082 0 1.1048079077931725e-11
GC_2_1083 b_2 NI_2 NS_1083 0 -3.3938026252157550e-11
GC_2_1084 b_2 NI_2 NS_1084 0 2.1486272689790518e-10
GC_2_1085 b_2 NI_2 NS_1085 0 -4.0816353789364114e-07
GC_2_1086 b_2 NI_2 NS_1086 0 -2.7824134145082082e-07
GC_2_1087 b_2 NI_2 NS_1087 0 -1.0588618034171463e-07
GC_2_1088 b_2 NI_2 NS_1088 0 5.6550176910298998e-07
GC_2_1089 b_2 NI_2 NS_1089 0 2.3813388588375208e-07
GC_2_1090 b_2 NI_2 NS_1090 0 1.4039358153473941e-06
GC_2_1091 b_2 NI_2 NS_1091 0 1.1109697996188631e-06
GC_2_1092 b_2 NI_2 NS_1092 0 -3.7454545637452611e-07
GC_2_1093 b_2 NI_2 NS_1093 0 6.7784042260002690e-07
GC_2_1094 b_2 NI_2 NS_1094 0 -2.0281319495739519e-06
GC_2_1095 b_2 NI_2 NS_1095 0 -6.4680863842927353e-07
GC_2_1096 b_2 NI_2 NS_1096 0 2.8098202343888970e-07
GC_2_1097 b_2 NI_2 NS_1097 0 9.9940330132008075e-07
GC_2_1098 b_2 NI_2 NS_1098 0 6.6416447314337982e-07
GC_2_1099 b_2 NI_2 NS_1099 0 3.8974620475536669e-06
GC_2_1100 b_2 NI_2 NS_1100 0 -3.7311349483032212e-06
GC_2_1101 b_2 NI_2 NS_1101 0 -5.5969153812496244e-06
GC_2_1102 b_2 NI_2 NS_1102 0 -3.8629264829764545e-06
GC_2_1103 b_2 NI_2 NS_1103 0 -9.2017134413358040e-07
GC_2_1104 b_2 NI_2 NS_1104 0 -2.0450965298398121e-06
GC_2_1105 b_2 NI_2 NS_1105 0 -1.3600398180363280e-05
GC_2_1106 b_2 NI_2 NS_1106 0 5.3801239297614193e-06
GC_2_1107 b_2 NI_2 NS_1107 0 -5.3844155589257947e-07
GC_2_1108 b_2 NI_2 NS_1108 0 1.8937674490603650e-06
GC_2_1109 b_2 NI_2 NS_1109 0 7.8172915364680246e-07
GC_2_1110 b_2 NI_2 NS_1110 0 1.9309075104469618e-05
GC_2_1111 b_2 NI_2 NS_1111 0 2.7666959355892811e-06
GC_2_1112 b_2 NI_2 NS_1112 0 -4.5945382077923062e-06
GC_2_1113 b_2 NI_2 NS_1113 0 1.4653345467342847e-06
GC_2_1114 b_2 NI_2 NS_1114 0 1.7112797626894646e-06
GC_2_1115 b_2 NI_2 NS_1115 0 5.3166453433960013e-06
GC_2_1116 b_2 NI_2 NS_1116 0 -2.2410313097344438e-06
GC_2_1117 b_2 NI_2 NS_1117 0 -4.1276255128942088e-07
GC_2_1118 b_2 NI_2 NS_1118 0 -8.1224333706608351e-07
GC_2_1119 b_2 NI_2 NS_1119 0 -2.0565664958506803e-06
GC_2_1120 b_2 NI_2 NS_1120 0 2.3251987796950080e-06
GC_2_1121 b_2 NI_2 NS_1121 0 -3.0284606030003597e-08
GC_2_1122 b_2 NI_2 NS_1122 0 1.2397142346099484e-06
GC_2_1123 b_2 NI_2 NS_1123 0 5.2803288489021499e-06
GC_2_1124 b_2 NI_2 NS_1124 0 5.9467815075317083e-06
GC_2_1125 b_2 NI_2 NS_1125 0 1.4516667812858841e-06
GC_2_1126 b_2 NI_2 NS_1126 0 -1.0225308412720461e-06
GC_2_1127 b_2 NI_2 NS_1127 0 1.1386249758805848e-07
GC_2_1128 b_2 NI_2 NS_1128 0 -4.7252921723568218e-08
GC_2_1129 b_2 NI_2 NS_1129 0 5.0776014492051103e-07
GC_2_1130 b_2 NI_2 NS_1130 0 7.4654450907593413e-07
GC_2_1131 b_2 NI_2 NS_1131 0 6.0590694621455445e-06
GC_2_1132 b_2 NI_2 NS_1132 0 4.9646363864062875e-07
GC_2_1133 b_2 NI_2 NS_1133 0 5.5787787662670389e-07
GC_2_1134 b_2 NI_2 NS_1134 0 -8.6741809359676037e-07
GC_2_1135 b_2 NI_2 NS_1135 0 -1.2579149204150366e-07
GC_2_1136 b_2 NI_2 NS_1136 0 -3.6410547378789043e-08
GC_2_1137 b_2 NI_2 NS_1137 0 6.7967556675370402e-07
GC_2_1138 b_2 NI_2 NS_1138 0 8.5001315458588886e-07
GC_2_1139 b_2 NI_2 NS_1139 0 4.7885039996556304e-06
GC_2_1140 b_2 NI_2 NS_1140 0 -1.9381605613468887e-06
GC_2_1141 b_2 NI_2 NS_1141 0 1.3610400555033126e-07
GC_2_1142 b_2 NI_2 NS_1142 0 -7.2191626562384194e-07
GC_2_1143 b_2 NI_2 NS_1143 0 -1.2100627669030458e-07
GC_2_1144 b_2 NI_2 NS_1144 0 1.4828056816996923e-07
GC_2_1145 b_2 NI_2 NS_1145 0 9.4361677591473579e-07
GC_2_1146 b_2 NI_2 NS_1146 0 7.7731628098622940e-07
GC_2_1147 b_2 NI_2 NS_1147 0 2.7625444003342120e-06
GC_2_1148 b_2 NI_2 NS_1148 0 -3.0182470804862878e-06
GC_2_1149 b_2 NI_2 NS_1149 0 -1.0350572748502878e-07
GC_2_1150 b_2 NI_2 NS_1150 0 -4.8431821613935087e-07
GC_2_1151 b_2 NI_2 NS_1151 0 8.8979733004626948e-08
GC_2_1152 b_2 NI_2 NS_1152 0 2.0122321141347971e-07
GC_2_1153 b_2 NI_2 NS_1153 0 1.3138892514620009e-06
GC_2_1154 b_2 NI_2 NS_1154 0 5.1136391387892178e-07
GC_2_1155 b_2 NI_2 NS_1155 0 6.6547015123361122e-07
GC_2_1156 b_2 NI_2 NS_1156 0 -2.7705953734868426e-06
GC_2_1157 b_2 NI_2 NS_1157 0 -1.6498847987596784e-07
GC_2_1158 b_2 NI_2 NS_1158 0 -1.3966200621689580e-07
GC_2_1159 b_2 NI_2 NS_1159 0 2.2753878427132159e-07
GC_2_1160 b_2 NI_2 NS_1160 0 2.2626917737803636e-08
GC_2_1161 b_2 NI_2 NS_1161 0 1.6154000795154830e-12
GC_2_1162 b_2 NI_2 NS_1162 0 -6.1877302402298734e-12
GC_2_1163 b_2 NI_2 NS_1163 0 9.8103601235537330e-07
GC_2_1164 b_2 NI_2 NS_1164 0 -2.6426789463219528e-07
GC_2_1165 b_2 NI_2 NS_1165 0 -2.6851718558245062e-08
GC_2_1166 b_2 NI_2 NS_1166 0 4.9057065588672041e-08
GC_2_1167 b_2 NI_2 NS_1167 0 2.6314501913932904e-07
GC_2_1168 b_2 NI_2 NS_1168 0 1.1130651523524751e-08
GC_2_1169 b_2 NI_2 NS_1169 0 8.3328275951927573e-07
GC_2_1170 b_2 NI_2 NS_1170 0 -1.5920615920179657e-07
GC_2_1171 b_2 NI_2 NS_1171 0 -6.3069986628787706e-08
GC_2_1172 b_2 NI_2 NS_1172 0 -1.0947720472250063e-06
GC_2_1173 b_2 NI_2 NS_1173 0 7.6562681223389180e-11
GC_2_1174 b_2 NI_2 NS_1174 0 -1.9340927072710480e-10
GC_2_1175 b_2 NI_2 NS_1175 0 6.8042313436485811e-07
GC_2_1176 b_2 NI_2 NS_1176 0 -4.3030881336575155e-07
GC_2_1177 b_2 NI_2 NS_1177 0 4.2741733489893168e-07
GC_2_1178 b_2 NI_2 NS_1178 0 1.6120708409827470e-07
GC_2_1179 b_2 NI_2 NS_1179 0 1.4000296594107019e-07
GC_2_1180 b_2 NI_2 NS_1180 0 -8.2544163703832244e-08
GC_2_1181 b_2 NI_2 NS_1181 0 -1.4336568375280853e-07
GC_2_1182 b_2 NI_2 NS_1182 0 -6.7656556214547719e-07
GC_2_1183 b_2 NI_2 NS_1183 0 2.4257999185698915e-08
GC_2_1184 b_2 NI_2 NS_1184 0 2.3623466406401552e-07
GC_2_1185 b_2 NI_2 NS_1185 0 3.3298105659080921e-07
GC_2_1186 b_2 NI_2 NS_1186 0 -5.5339150723010937e-08
GC_2_1187 b_2 NI_2 NS_1187 0 4.0223383360991688e-07
GC_2_1188 b_2 NI_2 NS_1188 0 2.2651200227343684e-07
GC_2_1189 b_2 NI_2 NS_1189 0 1.0244824934496132e-05
GC_2_1190 b_2 NI_2 NS_1190 0 -4.7957565763202459e-12
GC_2_1191 b_2 NI_2 NS_1191 0 1.0352148763988975e-11
GC_2_1192 b_2 NI_2 NS_1192 0 3.7845711167222202e-10
GC_2_1193 b_2 NI_2 NS_1193 0 1.3512321934705165e-07
GC_2_1194 b_2 NI_2 NS_1194 0 1.0761650325971493e-07
GC_2_1195 b_2 NI_2 NS_1195 0 7.2007404806331167e-07
GC_2_1196 b_2 NI_2 NS_1196 0 -1.8726838075764485e-07
GC_2_1197 b_2 NI_2 NS_1197 0 -5.9814066807743202e-07
GC_2_1198 b_2 NI_2 NS_1198 0 -3.6306370048057923e-07
GC_2_1199 b_2 NI_2 NS_1199 0 1.3989866212219598e-06
GC_2_1200 b_2 NI_2 NS_1200 0 3.2532209312422334e-07
GC_2_1201 b_2 NI_2 NS_1201 0 -9.9970706584993768e-07
GC_2_1202 b_2 NI_2 NS_1202 0 -1.7789575773254586e-06
GC_2_1203 b_2 NI_2 NS_1203 0 2.5545141588688196e-07
GC_2_1204 b_2 NI_2 NS_1204 0 -5.4832305061169047e-09
GC_2_1205 b_2 NI_2 NS_1205 0 -8.7354451166881868e-07
GC_2_1206 b_2 NI_2 NS_1206 0 9.7910779282313118e-08
GC_2_1207 b_2 NI_2 NS_1207 0 2.5713350827444533e-06
GC_2_1208 b_2 NI_2 NS_1208 0 -1.1143659200583766e-06
GC_2_1209 b_2 NI_2 NS_1209 0 -3.9892769091067626e-06
GC_2_1210 b_2 NI_2 NS_1210 0 -2.3994112659313797e-07
GC_2_1211 b_2 NI_2 NS_1211 0 1.2120432369672162e-08
GC_2_1212 b_2 NI_2 NS_1212 0 1.6053768143519848e-06
GC_2_1213 b_2 NI_2 NS_1213 0 -8.3045130368967740e-07
GC_2_1214 b_2 NI_2 NS_1214 0 -2.6088612769950412e-06
GC_2_1215 b_2 NI_2 NS_1215 0 -7.8261801526069435e-07
GC_2_1216 b_2 NI_2 NS_1216 0 1.4932821202601290e-06
GC_2_1217 b_2 NI_2 NS_1217 0 5.8174643423570085e-07
GC_2_1218 b_2 NI_2 NS_1218 0 -3.0275227691380212e-06
GC_2_1219 b_2 NI_2 NS_1219 0 -1.4471015755140149e-06
GC_2_1220 b_2 NI_2 NS_1220 0 2.5661999337405026e-06
GC_2_1221 b_2 NI_2 NS_1221 0 2.3925623353524561e-07
GC_2_1222 b_2 NI_2 NS_1222 0 1.2705126103062140e-06
GC_2_1223 b_2 NI_2 NS_1223 0 -6.9731504057197362e-07
GC_2_1224 b_2 NI_2 NS_1224 0 -1.1693000850529994e-06
GC_2_1225 b_2 NI_2 NS_1225 0 -5.8078006464813672e-08
GC_2_1226 b_2 NI_2 NS_1226 0 1.0861776755153817e-06
GC_2_1227 b_2 NI_2 NS_1227 0 -6.5276871785912375e-07
GC_2_1228 b_2 NI_2 NS_1228 0 -7.6713787148156828e-07
GC_2_1229 b_2 NI_2 NS_1229 0 -5.1252571434248895e-07
GC_2_1230 b_2 NI_2 NS_1230 0 1.1060714675576454e-06
GC_2_1231 b_2 NI_2 NS_1231 0 4.5034093264547863e-08
GC_2_1232 b_2 NI_2 NS_1232 0 -8.8826783616456403e-07
GC_2_1233 b_2 NI_2 NS_1233 0 -9.1170823675592514e-07
GC_2_1234 b_2 NI_2 NS_1234 0 1.0678781809196017e-06
GC_2_1235 b_2 NI_2 NS_1235 0 -1.1157811836972003e-07
GC_2_1236 b_2 NI_2 NS_1236 0 7.9119377002730953e-09
GC_2_1237 b_2 NI_2 NS_1237 0 -3.3924077476787524e-07
GC_2_1238 b_2 NI_2 NS_1238 0 1.0187665714722790e-06
GC_2_1239 b_2 NI_2 NS_1239 0 -9.8122861495842536e-08
GC_2_1240 b_2 NI_2 NS_1240 0 1.1222945452419873e-07
GC_2_1241 b_2 NI_2 NS_1241 0 -3.0038754229376790e-07
GC_2_1242 b_2 NI_2 NS_1242 0 1.0059083970110860e-06
GC_2_1243 b_2 NI_2 NS_1243 0 8.0898666509573745e-08
GC_2_1244 b_2 NI_2 NS_1244 0 1.6439233762079382e-07
GC_2_1245 b_2 NI_2 NS_1245 0 -7.9032862418838515e-08
GC_2_1246 b_2 NI_2 NS_1246 0 1.1304511617387262e-06
GC_2_1247 b_2 NI_2 NS_1247 0 7.8465136125993836e-07
GC_2_1248 b_2 NI_2 NS_1248 0 -9.7832270792976779e-09
GC_2_1249 b_2 NI_2 NS_1249 0 8.4849804829692911e-08
GC_2_1250 b_2 NI_2 NS_1250 0 8.2101088913914990e-07
GC_2_1251 b_2 NI_2 NS_1251 0 3.1725535918735979e-07
GC_2_1252 b_2 NI_2 NS_1252 0 -1.9311026931794494e-07
GC_2_1253 b_2 NI_2 NS_1253 0 1.9073686926552513e-07
GC_2_1254 b_2 NI_2 NS_1254 0 1.0069325065051334e-06
GC_2_1255 b_2 NI_2 NS_1255 0 7.9531953128704692e-07
GC_2_1256 b_2 NI_2 NS_1256 0 -8.1781933285187677e-07
GC_2_1257 b_2 NI_2 NS_1257 0 3.2999046153352693e-07
GC_2_1258 b_2 NI_2 NS_1258 0 5.3261459660956006e-07
GC_2_1259 b_2 NI_2 NS_1259 0 -5.5979513397727754e-09
GC_2_1260 b_2 NI_2 NS_1260 0 -5.5297846681131321e-07
GC_2_1261 b_2 NI_2 NS_1261 0 4.5646394560483840e-07
GC_2_1262 b_2 NI_2 NS_1262 0 7.5300337674904394e-07
GC_2_1263 b_2 NI_2 NS_1263 0 -9.7913843885014036e-09
GC_2_1264 b_2 NI_2 NS_1264 0 -1.1014051210591523e-06
GC_2_1265 b_2 NI_2 NS_1265 0 3.1840338285168282e-07
GC_2_1266 b_2 NI_2 NS_1266 0 1.0304772551896797e-07
GC_2_1267 b_2 NI_2 NS_1267 0 -3.9308701979062608e-07
GC_2_1268 b_2 NI_2 NS_1268 0 -2.5353725938864523e-07
GC_2_1269 b_2 NI_2 NS_1269 0 1.4515475232757400e-12
GC_2_1270 b_2 NI_2 NS_1270 0 3.4001924355163612e-12
GC_2_1271 b_2 NI_2 NS_1271 0 3.9032022788949963e-07
GC_2_1272 b_2 NI_2 NS_1272 0 2.2951820705211356e-07
GC_2_1273 b_2 NI_2 NS_1273 0 1.1980276775096197e-07
GC_2_1274 b_2 NI_2 NS_1274 0 3.5450076689256875e-08
GC_2_1275 b_2 NI_2 NS_1275 0 -2.7884556592683239e-07
GC_2_1276 b_2 NI_2 NS_1276 0 -1.0897736393118806e-07
GC_2_1277 b_2 NI_2 NS_1277 0 3.2156250776848966e-07
GC_2_1278 b_2 NI_2 NS_1278 0 6.8215122957652735e-08
GC_2_1279 b_2 NI_2 NS_1279 0 -3.5585251451820418e-07
GC_2_1280 b_2 NI_2 NS_1280 0 -4.5136761047083471e-07
GC_2_1281 b_2 NI_2 NS_1281 0 -1.0584885327622276e-11
GC_2_1282 b_2 NI_2 NS_1282 0 3.2224318836283975e-10
GC_2_1283 b_2 NI_2 NS_1283 0 1.8885838195295883e-07
GC_2_1284 b_2 NI_2 NS_1284 0 -1.9034133280025442e-07
GC_2_1285 b_2 NI_2 NS_1285 0 -7.7178688033747115e-08
GC_2_1286 b_2 NI_2 NS_1286 0 3.9129202774792946e-07
GC_2_1287 b_2 NI_2 NS_1287 0 -1.7579598023333728e-07
GC_2_1288 b_2 NI_2 NS_1288 0 6.2408050580644958e-08
GC_2_1289 b_2 NI_2 NS_1289 0 -5.3348898414776999e-07
GC_2_1290 b_2 NI_2 NS_1290 0 -2.6042883839867589e-07
GC_2_1291 b_2 NI_2 NS_1291 0 5.9193997305081484e-08
GC_2_1292 b_2 NI_2 NS_1292 0 2.3071477802606987e-08
GC_2_1293 b_2 NI_2 NS_1293 0 -3.6617573323885000e-07
GC_2_1294 b_2 NI_2 NS_1294 0 6.6093771623615222e-08
GC_2_1295 b_2 NI_2 NS_1295 0 1.0697458194248928e-07
GC_2_1296 b_2 NI_2 NS_1296 0 3.2656960588728474e-07
GD_2_1 b_2 NI_2 NA_1 0 -4.9159171881793104e-03
GD_2_2 b_2 NI_2 NA_2 0 -1.0697627826309042e-02
GD_2_3 b_2 NI_2 NA_3 0 -1.1524177943753036e-03
GD_2_4 b_2 NI_2 NA_4 0 1.0616349053176282e-02
GD_2_5 b_2 NI_2 NA_5 0 1.9211933082206064e-05
GD_2_6 b_2 NI_2 NA_6 0 3.1568060439406801e-06
GD_2_7 b_2 NI_2 NA_7 0 1.1360090622450836e-05
GD_2_8 b_2 NI_2 NA_8 0 -2.6035568648901429e-06
GD_2_9 b_2 NI_2 NA_9 0 8.8077176040343653e-06
GD_2_10 b_2 NI_2 NA_10 0 -1.1809799684390413e-06
GD_2_11 b_2 NI_2 NA_11 0 3.3591010288444652e-06
GD_2_12 b_2 NI_2 NA_12 0 -2.2825072134952614e-06
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 1.1808946086155321e-03
GC_3_2 b_3 NI_3 NS_2 0 -3.5561529341965672e-09
GC_3_3 b_3 NI_3 NS_3 0 -4.8002191774701852e-08
GC_3_4 b_3 NI_3 NS_4 0 -3.4752340704549879e-06
GC_3_5 b_3 NI_3 NS_5 0 -3.6811901364780004e-04
GC_3_6 b_3 NI_3 NS_6 0 1.3598187543188193e-04
GC_3_7 b_3 NI_3 NS_7 0 1.1297146933370728e-03
GC_3_8 b_3 NI_3 NS_8 0 1.9432462846757893e-03
GC_3_9 b_3 NI_3 NS_9 0 -6.5024476552742058e-05
GC_3_10 b_3 NI_3 NS_10 0 -3.4937331271818863e-03
GC_3_11 b_3 NI_3 NS_11 0 -1.5644021981814785e-03
GC_3_12 b_3 NI_3 NS_12 0 5.0905624229486447e-03
GC_3_13 b_3 NI_3 NS_13 0 4.2534128653169048e-03
GC_3_14 b_3 NI_3 NS_14 0 -4.9937799992363406e-03
GC_3_15 b_3 NI_3 NS_15 0 -1.0085407529908136e-03
GC_3_16 b_3 NI_3 NS_16 0 5.6396386094321722e-04
GC_3_17 b_3 NI_3 NS_17 0 -2.0807406583217081e-03
GC_3_18 b_3 NI_3 NS_18 0 -1.8633318893576912e-03
GC_3_19 b_3 NI_3 NS_19 0 3.6453771295848012e-03
GC_3_20 b_3 NI_3 NS_20 0 1.1647296882442261e-02
GC_3_21 b_3 NI_3 NS_21 0 -8.9809614803279699e-04
GC_3_22 b_3 NI_3 NS_22 0 -1.4854265632828951e-02
GC_3_23 b_3 NI_3 NS_23 0 -8.1235076431966733e-03
GC_3_24 b_3 NI_3 NS_24 0 1.9195537939136588e-03
GC_3_25 b_3 NI_3 NS_25 0 1.1262993530090817e-02
GC_3_26 b_3 NI_3 NS_26 0 -1.8122069155800812e-03
GC_3_27 b_3 NI_3 NS_27 0 -7.5672398442390380e-03
GC_3_28 b_3 NI_3 NS_28 0 -1.6812116993683219e-03
GC_3_29 b_3 NI_3 NS_29 0 1.5281604976723493e-02
GC_3_30 b_3 NI_3 NS_30 0 5.3008405645793124e-03
GC_3_31 b_3 NI_3 NS_31 0 -1.3082790953757006e-02
GC_3_32 b_3 NI_3 NS_32 0 -5.4613178963359979e-03
GC_3_33 b_3 NI_3 NS_33 0 -6.6370644564244250e-03
GC_3_34 b_3 NI_3 NS_34 0 3.4566475701970282e-03
GC_3_35 b_3 NI_3 NS_35 0 6.3615644356746727e-03
GC_3_36 b_3 NI_3 NS_36 0 -1.8793118019297607e-03
GC_3_37 b_3 NI_3 NS_37 0 -5.4737186445375967e-03
GC_3_38 b_3 NI_3 NS_38 0 2.1829946686460931e-03
GC_3_39 b_3 NI_3 NS_39 0 5.3937393709659678e-03
GC_3_40 b_3 NI_3 NS_40 0 -2.6324117744461828e-03
GC_3_41 b_3 NI_3 NS_41 0 -6.3064431411680019e-03
GC_3_42 b_3 NI_3 NS_42 0 -4.8383735656624700e-04
GC_3_43 b_3 NI_3 NS_43 0 7.6452220984865853e-03
GC_3_44 b_3 NI_3 NS_44 0 3.6298705718534338e-03
GC_3_45 b_3 NI_3 NS_45 0 -5.8336093149023447e-03
GC_3_46 b_3 NI_3 NS_46 0 -3.4646024563499194e-03
GC_3_47 b_3 NI_3 NS_47 0 2.9619348919130833e-04
GC_3_48 b_3 NI_3 NS_48 0 5.5809941025782397e-04
GC_3_49 b_3 NI_3 NS_49 0 -4.9270657872240815e-03
GC_3_50 b_3 NI_3 NS_50 0 8.9217852429806111e-04
GC_3_51 b_3 NI_3 NS_51 0 6.2062929702040252e-03
GC_3_52 b_3 NI_3 NS_52 0 6.8828400938386754e-04
GC_3_53 b_3 NI_3 NS_53 0 -5.3209611644942463e-03
GC_3_54 b_3 NI_3 NS_54 0 -4.8420318236961778e-04
GC_3_55 b_3 NI_3 NS_55 0 1.5503149071468792e-03
GC_3_56 b_3 NI_3 NS_56 0 -4.3204677706099045e-05
GC_3_57 b_3 NI_3 NS_57 0 -6.0223419042160498e-03
GC_3_58 b_3 NI_3 NS_58 0 1.9232193706757007e-03
GC_3_59 b_3 NI_3 NS_59 0 6.2616196388788651e-03
GC_3_60 b_3 NI_3 NS_60 0 2.1739983894910730e-04
GC_3_61 b_3 NI_3 NS_61 0 -5.0592028594619205e-03
GC_3_62 b_3 NI_3 NS_62 0 1.7016087774869965e-03
GC_3_63 b_3 NI_3 NS_63 0 2.4884687136956488e-03
GC_3_64 b_3 NI_3 NS_64 0 -9.5763254242980402e-04
GC_3_65 b_3 NI_3 NS_65 0 -6.5329693358752014e-03
GC_3_66 b_3 NI_3 NS_66 0 3.8846207766480272e-03
GC_3_67 b_3 NI_3 NS_67 0 7.4932573120104866e-03
GC_3_68 b_3 NI_3 NS_68 0 -1.0959984792696749e-03
GC_3_69 b_3 NI_3 NS_69 0 -3.9851238840564549e-03
GC_3_70 b_3 NI_3 NS_70 0 4.0409678507002085e-03
GC_3_71 b_3 NI_3 NS_71 0 2.8633256063451220e-03
GC_3_72 b_3 NI_3 NS_72 0 -3.0534816325066467e-03
GC_3_73 b_3 NI_3 NS_73 0 -6.0227369844529791e-03
GC_3_74 b_3 NI_3 NS_74 0 7.2373641985876416e-03
GC_3_75 b_3 NI_3 NS_75 0 7.9896920165475442e-03
GC_3_76 b_3 NI_3 NS_76 0 -4.8114430249762054e-03
GC_3_77 b_3 NI_3 NS_77 0 -5.3743583256955492e-04
GC_3_78 b_3 NI_3 NS_78 0 5.0204619083623909e-03
GC_3_79 b_3 NI_3 NS_79 0 2.4825093756679020e-04
GC_3_80 b_3 NI_3 NS_80 0 -4.7581881502032578e-03
GC_3_81 b_3 NI_3 NS_81 0 1.8107800231420959e-09
GC_3_82 b_3 NI_3 NS_82 0 3.2741335365165904e-09
GC_3_83 b_3 NI_3 NS_83 0 -1.4272202680221762e-03
GC_3_84 b_3 NI_3 NS_84 0 7.8707216177806346e-03
GC_3_85 b_3 NI_3 NS_85 0 -1.7999315117155415e-04
GC_3_86 b_3 NI_3 NS_86 0 3.0272430884242282e-03
GC_3_87 b_3 NI_3 NS_87 0 -1.3039334253071925e-04
GC_3_88 b_3 NI_3 NS_88 0 -3.3752918432832890e-03
GC_3_89 b_3 NI_3 NS_89 0 -8.7633853397964809e-04
GC_3_90 b_3 NI_3 NS_90 0 7.5304799097416532e-03
GC_3_91 b_3 NI_3 NS_91 0 3.7887927327919127e-03
GC_3_92 b_3 NI_3 NS_92 0 -6.1573976215618647e-03
GC_3_93 b_3 NI_3 NS_93 0 8.6224686718153012e-08
GC_3_94 b_3 NI_3 NS_94 0 -3.5295555329375523e-07
GC_3_95 b_3 NI_3 NS_95 0 6.7186820305059434e-03
GC_3_96 b_3 NI_3 NS_96 0 -5.3194053991504568e-03
GC_3_97 b_3 NI_3 NS_97 0 -2.6111752847583652e-03
GC_3_98 b_3 NI_3 NS_98 0 6.0542436034968930e-03
GC_3_99 b_3 NI_3 NS_99 0 -4.2922721356863733e-03
GC_3_100 b_3 NI_3 NS_100 0 1.4428603149831981e-05
GC_3_101 b_3 NI_3 NS_101 0 2.7173857208235988e-03
GC_3_102 b_3 NI_3 NS_102 0 -6.2039921813181508e-03
GC_3_103 b_3 NI_3 NS_103 0 2.0957199164177666e-03
GC_3_104 b_3 NI_3 NS_104 0 3.2562861580772711e-03
GC_3_105 b_3 NI_3 NS_105 0 -1.9700288835581008e-03
GC_3_106 b_3 NI_3 NS_106 0 -4.4205333652799191e-03
GC_3_107 b_3 NI_3 NS_107 0 2.8640817371894936e-03
GC_3_108 b_3 NI_3 NS_108 0 8.0083593647129053e-03
GC_3_109 b_3 NI_3 NS_109 0 -3.3036181833295221e-03
GC_3_110 b_3 NI_3 NS_110 0 1.8493832879736667e-09
GC_3_111 b_3 NI_3 NS_111 0 5.6032189439071558e-08
GC_3_112 b_3 NI_3 NS_112 0 1.8929692746408944e-06
GC_3_113 b_3 NI_3 NS_113 0 -9.1167736727195163e-05
GC_3_114 b_3 NI_3 NS_114 0 -5.7737685973767697e-05
GC_3_115 b_3 NI_3 NS_115 0 -1.2657732146135821e-03
GC_3_116 b_3 NI_3 NS_116 0 -2.9559335286384196e-04
GC_3_117 b_3 NI_3 NS_117 0 -1.6792127358340608e-03
GC_3_118 b_3 NI_3 NS_118 0 2.6464980981649299e-03
GC_3_119 b_3 NI_3 NS_119 0 5.1121264671097376e-04
GC_3_120 b_3 NI_3 NS_120 0 5.4276095793636559e-03
GC_3_121 b_3 NI_3 NS_121 0 7.1034902484533547e-03
GC_3_122 b_3 NI_3 NS_122 0 6.3629124964924104e-04
GC_3_123 b_3 NI_3 NS_123 0 6.4433103928248010e-04
GC_3_124 b_3 NI_3 NS_124 0 -6.6091960612429219e-04
GC_3_125 b_3 NI_3 NS_125 0 1.0576976554500499e-03
GC_3_126 b_3 NI_3 NS_126 0 1.5711389928360555e-03
GC_3_127 b_3 NI_3 NS_127 0 1.2687515819068761e-02
GC_3_128 b_3 NI_3 NS_128 0 1.3123211167354478e-02
GC_3_129 b_3 NI_3 NS_129 0 8.7187952734211881e-03
GC_3_130 b_3 NI_3 NS_130 0 -2.0392082084500836e-02
GC_3_131 b_3 NI_3 NS_131 0 8.3891008488131656e-03
GC_3_132 b_3 NI_3 NS_132 0 -2.9045265252446023e-03
GC_3_133 b_3 NI_3 NS_133 0 -1.2701292160154020e-02
GC_3_134 b_3 NI_3 NS_134 0 -3.8806700449034136e-02
GC_3_135 b_3 NI_3 NS_135 0 -7.2523394845434280e-03
GC_3_136 b_3 NI_3 NS_136 0 -2.1332749811690133e-03
GC_3_137 b_3 NI_3 NS_137 0 -5.2307202174282016e-02
GC_3_138 b_3 NI_3 NS_138 0 -1.7936179654169594e-03
GC_3_139 b_3 NI_3 NS_139 0 1.4914415696362647e-02
GC_3_140 b_3 NI_3 NS_140 0 8.6735776585703528e-03
GC_3_141 b_3 NI_3 NS_141 0 -5.9233536280776386e-03
GC_3_142 b_3 NI_3 NS_142 0 5.0044967064219520e-03
GC_3_143 b_3 NI_3 NS_143 0 8.3724176249584861e-03
GC_3_144 b_3 NI_3 NS_144 0 1.1688364630635445e-02
GC_3_145 b_3 NI_3 NS_145 0 4.5592636074217579e-03
GC_3_146 b_3 NI_3 NS_146 0 -2.9327401707393550e-03
GC_3_147 b_3 NI_3 NS_147 0 -7.8986726013831141e-03
GC_3_148 b_3 NI_3 NS_148 0 -8.1490644502030963e-03
GC_3_149 b_3 NI_3 NS_149 0 -5.6808136154436620e-03
GC_3_150 b_3 NI_3 NS_150 0 -6.1281013974292837e-04
GC_3_151 b_3 NI_3 NS_151 0 -1.8070849982267680e-02
GC_3_152 b_3 NI_3 NS_152 0 1.3578963963608619e-02
GC_3_153 b_3 NI_3 NS_153 0 4.7069861997291644e-03
GC_3_154 b_3 NI_3 NS_154 0 4.3794387167996555e-03
GC_3_155 b_3 NI_3 NS_155 0 6.5015854709090228e-04
GC_3_156 b_3 NI_3 NS_156 0 -1.0995439796376788e-04
GC_3_157 b_3 NI_3 NS_157 0 -3.7963997125100798e-03
GC_3_158 b_3 NI_3 NS_158 0 8.8498808546380885e-04
GC_3_159 b_3 NI_3 NS_159 0 -1.1178294413854567e-03
GC_3_160 b_3 NI_3 NS_160 0 1.6699687323271033e-02
GC_3_161 b_3 NI_3 NS_161 0 4.4472802773569782e-03
GC_3_162 b_3 NI_3 NS_162 0 7.0796477313533727e-04
GC_3_163 b_3 NI_3 NS_163 0 -5.1995788897902064e-04
GC_3_164 b_3 NI_3 NS_164 0 -2.2477510487971630e-03
GC_3_165 b_3 NI_3 NS_165 0 -4.9864555048166528e-03
GC_3_166 b_3 NI_3 NS_166 0 2.1108871260369223e-03
GC_3_167 b_3 NI_3 NS_167 0 7.3425260205902190e-03
GC_3_168 b_3 NI_3 NS_168 0 1.4345854451170230e-02
GC_3_169 b_3 NI_3 NS_169 0 4.1872272120768352e-03
GC_3_170 b_3 NI_3 NS_170 0 -1.6838581543015731e-03
GC_3_171 b_3 NI_3 NS_171 0 -3.3981246404814779e-03
GC_3_172 b_3 NI_3 NS_172 0 -2.1006230650192324e-03
GC_3_173 b_3 NI_3 NS_173 0 -5.4204251570271695e-03
GC_3_174 b_3 NI_3 NS_174 0 4.3817243815421998e-03
GC_3_175 b_3 NI_3 NS_175 0 1.3196871855987086e-02
GC_3_176 b_3 NI_3 NS_176 0 8.4333056400068898e-03
GC_3_177 b_3 NI_3 NS_177 0 2.8324335654533821e-03
GC_3_178 b_3 NI_3 NS_178 0 -4.1306068390157460e-03
GC_3_179 b_3 NI_3 NS_179 0 -5.3207874827182330e-03
GC_3_180 b_3 NI_3 NS_180 0 1.1381584245146693e-03
GC_3_181 b_3 NI_3 NS_181 0 -4.4310212078039705e-03
GC_3_182 b_3 NI_3 NS_182 0 8.3104301820648829e-03
GC_3_183 b_3 NI_3 NS_183 0 1.4612784280878520e-02
GC_3_184 b_3 NI_3 NS_184 0 -4.6824611923794820e-04
GC_3_185 b_3 NI_3 NS_185 0 -1.1845326088367103e-03
GC_3_186 b_3 NI_3 NS_186 0 -4.5473896408065465e-03
GC_3_187 b_3 NI_3 NS_187 0 -2.2825677842982042e-03
GC_3_188 b_3 NI_3 NS_188 0 4.3832552601853671e-03
GC_3_189 b_3 NI_3 NS_189 0 1.3569687558105462e-10
GC_3_190 b_3 NI_3 NS_190 0 -1.5466153752760475e-09
GC_3_191 b_3 NI_3 NS_191 0 1.4460253089716940e-03
GC_3_192 b_3 NI_3 NS_192 0 8.2165469699566462e-03
GC_3_193 b_3 NI_3 NS_193 0 -8.7895048513280912e-04
GC_3_194 b_3 NI_3 NS_194 0 -2.2072123262807941e-03
GC_3_195 b_3 NI_3 NS_195 0 -1.4679135645063882e-03
GC_3_196 b_3 NI_3 NS_196 0 2.7519863036413899e-03
GC_3_197 b_3 NI_3 NS_197 0 1.7320140142980558e-03
GC_3_198 b_3 NI_3 NS_198 0 7.6059327070770273e-03
GC_3_199 b_3 NI_3 NS_199 0 7.5874085960345389e-03
GC_3_200 b_3 NI_3 NS_200 0 -3.8276817810715849e-03
GC_3_201 b_3 NI_3 NS_201 0 -5.2100999515094752e-08
GC_3_202 b_3 NI_3 NS_202 0 -2.0817381263197200e-08
GC_3_203 b_3 NI_3 NS_203 0 1.1391243329703342e-02
GC_3_204 b_3 NI_3 NS_204 0 4.4700330877502394e-03
GC_3_205 b_3 NI_3 NS_205 0 -8.6185050719419728e-04
GC_3_206 b_3 NI_3 NS_206 0 6.4916225462376582e-03
GC_3_207 b_3 NI_3 NS_207 0 3.6263738391833660e-03
GC_3_208 b_3 NI_3 NS_208 0 4.0710469134965757e-04
GC_3_209 b_3 NI_3 NS_209 0 6.0525110494710210e-03
GC_3_210 b_3 NI_3 NS_210 0 -4.6635397706706275e-03
GC_3_211 b_3 NI_3 NS_211 0 -3.3929751249081128e-03
GC_3_212 b_3 NI_3 NS_212 0 -1.3533957840833777e-03
GC_3_213 b_3 NI_3 NS_213 0 1.1237978020494131e-04
GC_3_214 b_3 NI_3 NS_214 0 4.4958002916889034e-03
GC_3_215 b_3 NI_3 NS_215 0 7.2795568499957209e-03
GC_3_216 b_3 NI_3 NS_216 0 5.5305047826560714e-03
GC_3_217 b_3 NI_3 NS_217 0 -1.4246404788190137e-02
GC_3_218 b_3 NI_3 NS_218 0 6.2292709467693438e-09
GC_3_219 b_3 NI_3 NS_219 0 -1.0771398389488892e-06
GC_3_220 b_3 NI_3 NS_220 0 -2.3238216360955719e-05
GC_3_221 b_3 NI_3 NS_221 0 3.4199237682638851e-04
GC_3_222 b_3 NI_3 NS_222 0 -1.9835152991894148e-04
GC_3_223 b_3 NI_3 NS_223 0 -1.5573879029213886e-03
GC_3_224 b_3 NI_3 NS_224 0 -2.3367654356295561e-03
GC_3_225 b_3 NI_3 NS_225 0 -6.7659612820981498e-05
GC_3_226 b_3 NI_3 NS_226 0 4.3764657852802952e-03
GC_3_227 b_3 NI_3 NS_227 0 1.6012883084795251e-03
GC_3_228 b_3 NI_3 NS_228 0 -5.9363758342384065e-03
GC_3_229 b_3 NI_3 NS_229 0 -4.9862911833464555e-03
GC_3_230 b_3 NI_3 NS_230 0 6.4938614129152108e-03
GC_3_231 b_3 NI_3 NS_231 0 1.1242578186705604e-03
GC_3_232 b_3 NI_3 NS_232 0 -4.9042040139159854e-04
GC_3_233 b_3 NI_3 NS_233 0 2.8092111687197160e-03
GC_3_234 b_3 NI_3 NS_234 0 2.3585345818559742e-03
GC_3_235 b_3 NI_3 NS_235 0 -4.3182654913180765e-03
GC_3_236 b_3 NI_3 NS_236 0 -1.3539568144360713e-02
GC_3_237 b_3 NI_3 NS_237 0 1.6031664291940662e-03
GC_3_238 b_3 NI_3 NS_238 0 1.7677771464974880e-02
GC_3_239 b_3 NI_3 NS_239 0 9.8386848386797544e-03
GC_3_240 b_3 NI_3 NS_240 0 -2.2919450913237000e-03
GC_3_241 b_3 NI_3 NS_241 0 -1.3104488469257020e-02
GC_3_242 b_3 NI_3 NS_242 0 2.2186341526220857e-03
GC_3_243 b_3 NI_3 NS_243 0 9.2001452439411102e-03
GC_3_244 b_3 NI_3 NS_244 0 1.9506157451927521e-03
GC_3_245 b_3 NI_3 NS_245 0 -1.7998042638951106e-02
GC_3_246 b_3 NI_3 NS_246 0 -6.4920168015484758e-03
GC_3_247 b_3 NI_3 NS_247 0 1.5711165321299542e-02
GC_3_248 b_3 NI_3 NS_248 0 6.4981562116889586e-03
GC_3_249 b_3 NI_3 NS_249 0 8.1166009630611689e-03
GC_3_250 b_3 NI_3 NS_250 0 -4.1938588857842359e-03
GC_3_251 b_3 NI_3 NS_251 0 -7.5320606970618329e-03
GC_3_252 b_3 NI_3 NS_252 0 2.0324568159714802e-03
GC_3_253 b_3 NI_3 NS_253 0 6.7023910841256277e-03
GC_3_254 b_3 NI_3 NS_254 0 -2.7451381598351788e-03
GC_3_255 b_3 NI_3 NS_255 0 -6.5840253691331124e-03
GC_3_256 b_3 NI_3 NS_256 0 2.8920130832389610e-03
GC_3_257 b_3 NI_3 NS_257 0 7.6634840947172652e-03
GC_3_258 b_3 NI_3 NS_258 0 4.8601872493886480e-04
GC_3_259 b_3 NI_3 NS_259 0 -9.3542511629111005e-03
GC_3_260 b_3 NI_3 NS_260 0 -5.1821771855507679e-03
GC_3_261 b_3 NI_3 NS_261 0 6.8205103837088556e-03
GC_3_262 b_3 NI_3 NS_262 0 4.1105940199482119e-03
GC_3_263 b_3 NI_3 NS_263 0 -3.8505207999989211e-04
GC_3_264 b_3 NI_3 NS_264 0 -9.3423363189745724e-04
GC_3_265 b_3 NI_3 NS_265 0 5.6830631042289175e-03
GC_3_266 b_3 NI_3 NS_266 0 -1.3773228603985617e-03
GC_3_267 b_3 NI_3 NS_267 0 -9.1525454294963966e-03
GC_3_268 b_3 NI_3 NS_268 0 -1.2845789187939623e-03
GC_3_269 b_3 NI_3 NS_269 0 5.9995882824452201e-03
GC_3_270 b_3 NI_3 NS_270 0 7.3474304397222598e-04
GC_3_271 b_3 NI_3 NS_271 0 -2.6407567579049590e-03
GC_3_272 b_3 NI_3 NS_272 0 2.3245280178851732e-04
GC_3_273 b_3 NI_3 NS_273 0 6.7119805317866930e-03
GC_3_274 b_3 NI_3 NS_274 0 -2.2566103582136125e-03
GC_3_275 b_3 NI_3 NS_275 0 -9.2876884338962788e-03
GC_3_276 b_3 NI_3 NS_276 0 1.4716553638636878e-03
GC_3_277 b_3 NI_3 NS_277 0 5.7396080224354105e-03
GC_3_278 b_3 NI_3 NS_278 0 -1.5055505373886822e-03
GC_3_279 b_3 NI_3 NS_279 0 -3.3169949944616165e-03
GC_3_280 b_3 NI_3 NS_280 0 2.3821032594906612e-03
GC_3_281 b_3 NI_3 NS_281 0 7.2818918524707368e-03
GC_3_282 b_3 NI_3 NS_282 0 -4.0976815561999938e-03
GC_3_283 b_3 NI_3 NS_283 0 -8.5931435656783003e-03
GC_3_284 b_3 NI_3 NS_284 0 4.1427791364409168e-03
GC_3_285 b_3 NI_3 NS_285 0 4.8244372078949547e-03
GC_3_286 b_3 NI_3 NS_286 0 -3.8807298253234995e-03
GC_3_287 b_3 NI_3 NS_287 0 -2.4175657565250206e-03
GC_3_288 b_3 NI_3 NS_288 0 4.7355224271885951e-03
GC_3_289 b_3 NI_3 NS_289 0 7.0698650818165083e-03
GC_3_290 b_3 NI_3 NS_290 0 -7.3594023641601692e-03
GC_3_291 b_3 NI_3 NS_291 0 -7.1573594779305210e-03
GC_3_292 b_3 NI_3 NS_292 0 6.8575806727567273e-03
GC_3_293 b_3 NI_3 NS_293 0 1.6629093812802708e-03
GC_3_294 b_3 NI_3 NS_294 0 -5.3099129266202588e-03
GC_3_295 b_3 NI_3 NS_295 0 5.8005275187170515e-04
GC_3_296 b_3 NI_3 NS_296 0 5.4707651829512972e-03
GC_3_297 b_3 NI_3 NS_297 0 -4.5823953993093211e-09
GC_3_298 b_3 NI_3 NS_298 0 -1.3467243226169073e-08
GC_3_299 b_3 NI_3 NS_299 0 2.7089353287053312e-03
GC_3_300 b_3 NI_3 NS_300 0 -8.5910076750722805e-03
GC_3_301 b_3 NI_3 NS_301 0 8.6608621310463459e-04
GC_3_302 b_3 NI_3 NS_302 0 -3.4347601326466400e-03
GC_3_303 b_3 NI_3 NS_303 0 6.2756504024883265e-04
GC_3_304 b_3 NI_3 NS_304 0 4.0313421846025887e-03
GC_3_305 b_3 NI_3 NS_305 0 2.1670469590617755e-03
GC_3_306 b_3 NI_3 NS_306 0 -8.1665277303215999e-03
GC_3_307 b_3 NI_3 NS_307 0 -3.4991650927440393e-03
GC_3_308 b_3 NI_3 NS_308 0 7.0126800881225729e-03
GC_3_309 b_3 NI_3 NS_309 0 -1.0829953942196049e-07
GC_3_310 b_3 NI_3 NS_310 0 -3.0048136554613643e-07
GC_3_311 b_3 NI_3 NS_311 0 -8.0240637224034510e-03
GC_3_312 b_3 NI_3 NS_312 0 5.3776064418065367e-03
GC_3_313 b_3 NI_3 NS_313 0 4.1768099630321185e-03
GC_3_314 b_3 NI_3 NS_314 0 -6.8620735186216029e-03
GC_3_315 b_3 NI_3 NS_315 0 5.3214176226709818e-03
GC_3_316 b_3 NI_3 NS_316 0 7.4369290354656201e-04
GC_3_317 b_3 NI_3 NS_317 0 -2.3651598819094924e-03
GC_3_318 b_3 NI_3 NS_318 0 6.8561912681334479e-03
GC_3_319 b_3 NI_3 NS_319 0 -1.4960018488860982e-03
GC_3_320 b_3 NI_3 NS_320 0 -4.2193419650894022e-03
GC_3_321 b_3 NI_3 NS_321 0 2.3601154435927822e-03
GC_3_322 b_3 NI_3 NS_322 0 5.0361471043600383e-03
GC_3_323 b_3 NI_3 NS_323 0 -2.0068775958371663e-03
GC_3_324 b_3 NI_3 NS_324 0 -8.9761633823016284e-03
GC_3_325 b_3 NI_3 NS_325 0 -1.0575519490685487e-02
GC_3_326 b_3 NI_3 NS_326 0 9.5500174528559330e-09
GC_3_327 b_3 NI_3 NS_327 0 9.8517531287614878e-07
GC_3_328 b_3 NI_3 NS_328 0 3.6184004029527964e-05
GC_3_329 b_3 NI_3 NS_329 0 4.3796852742098375e-03
GC_3_330 b_3 NI_3 NS_330 0 -3.4738125656410329e-03
GC_3_331 b_3 NI_3 NS_331 0 -3.7302977077457514e-03
GC_3_332 b_3 NI_3 NS_332 0 6.2452121993507477e-03
GC_3_333 b_3 NI_3 NS_333 0 -8.7505764070591480e-03
GC_3_334 b_3 NI_3 NS_334 0 -5.9709435532982200e-03
GC_3_335 b_3 NI_3 NS_335 0 9.2221610592950146e-03
GC_3_336 b_3 NI_3 NS_336 0 -5.9539729889409787e-03
GC_3_337 b_3 NI_3 NS_337 0 7.1416129620862825e-03
GC_3_338 b_3 NI_3 NS_338 0 1.1891219389718237e-02
GC_3_339 b_3 NI_3 NS_339 0 -4.2237329887351875e-03
GC_3_340 b_3 NI_3 NS_340 0 -1.1434264180499299e-03
GC_3_341 b_3 NI_3 NS_341 0 -8.8759584327553955e-03
GC_3_342 b_3 NI_3 NS_342 0 -4.8952956482121372e-04
GC_3_343 b_3 NI_3 NS_343 0 1.4613686258044616e-02
GC_3_344 b_3 NI_3 NS_344 0 -1.0366838854078960e-02
GC_3_345 b_3 NI_3 NS_345 0 1.6418018674665510e-02
GC_3_346 b_3 NI_3 NS_346 0 4.0448172865586891e-03
GC_3_347 b_3 NI_3 NS_347 0 -1.1484854341614854e-02
GC_3_348 b_3 NI_3 NS_348 0 -2.5534353699577705e-04
GC_3_349 b_3 NI_3 NS_349 0 -1.6636009386018336e-02
GC_3_350 b_3 NI_3 NS_350 0 -4.4594539468441413e-02
GC_3_351 b_3 NI_3 NS_351 0 1.0649430532553393e-02
GC_3_352 b_3 NI_3 NS_352 0 1.1312881341626984e-03
GC_3_353 b_3 NI_3 NS_353 0 -4.8338803818630101e-02
GC_3_354 b_3 NI_3 NS_354 0 1.1008215930981165e-02
GC_3_355 b_3 NI_3 NS_355 0 -1.0431912427998033e-02
GC_3_356 b_3 NI_3 NS_356 0 4.9178883291357291e-04
GC_3_357 b_3 NI_3 NS_357 0 9.7750246819467389e-03
GC_3_358 b_3 NI_3 NS_358 0 -5.7662818420000316e-04
GC_3_359 b_3 NI_3 NS_359 0 4.5630430109836716e-03
GC_3_360 b_3 NI_3 NS_360 0 2.4175266327969170e-02
GC_3_361 b_3 NI_3 NS_361 0 -1.0747445242586886e-02
GC_3_362 b_3 NI_3 NS_362 0 1.9593637663349200e-03
GC_3_363 b_3 NI_3 NS_363 0 -8.4818331395541211e-03
GC_3_364 b_3 NI_3 NS_364 0 -1.3531518511156521e-02
GC_3_365 b_3 NI_3 NS_365 0 1.0144353937138121e-02
GC_3_366 b_3 NI_3 NS_366 0 9.9163601991735786e-04
GC_3_367 b_3 NI_3 NS_367 0 -1.9215707611688757e-02
GC_3_368 b_3 NI_3 NS_368 0 2.8664621017311140e-02
GC_3_369 b_3 NI_3 NS_369 0 -9.6176097883424461e-03
GC_3_370 b_3 NI_3 NS_370 0 -9.6669099453875428e-04
GC_3_371 b_3 NI_3 NS_371 0 1.8850151805706343e-03
GC_3_372 b_3 NI_3 NS_372 0 -1.3790908817360261e-03
GC_3_373 b_3 NI_3 NS_373 0 9.4567889505828718e-03
GC_3_374 b_3 NI_3 NS_374 0 -2.3684573212387041e-04
GC_3_375 b_3 NI_3 NS_375 0 -2.0771813499441036e-04
GC_3_376 b_3 NI_3 NS_376 0 3.0287235260256323e-02
GC_3_377 b_3 NI_3 NS_377 0 -8.5365101452413768e-03
GC_3_378 b_3 NI_3 NS_378 0 1.5565781410542261e-04
GC_3_379 b_3 NI_3 NS_379 0 2.0684736114498078e-04
GC_3_380 b_3 NI_3 NS_380 0 -5.4692179914387507e-03
GC_3_381 b_3 NI_3 NS_381 0 1.0024589320747970e-02
GC_3_382 b_3 NI_3 NS_382 0 -3.2644304845964259e-04
GC_3_383 b_3 NI_3 NS_383 0 8.8940718003618340e-03
GC_3_384 b_3 NI_3 NS_384 0 2.6408657373320269e-02
GC_3_385 b_3 NI_3 NS_385 0 -8.3634747997869009e-03
GC_3_386 b_3 NI_3 NS_386 0 1.3809555879928470e-03
GC_3_387 b_3 NI_3 NS_387 0 -2.5880188543615473e-03
GC_3_388 b_3 NI_3 NS_388 0 -7.3315810760288223e-03
GC_3_389 b_3 NI_3 NS_389 0 1.0540515336797666e-02
GC_3_390 b_3 NI_3 NS_390 0 -8.1040481809333518e-04
GC_3_391 b_3 NI_3 NS_391 0 1.4431101689994390e-02
GC_3_392 b_3 NI_3 NS_392 0 2.0002744912694111e-02
GC_3_393 b_3 NI_3 NS_393 0 -8.2822253361821713e-03
GC_3_394 b_3 NI_3 NS_394 0 2.9406940584838477e-03
GC_3_395 b_3 NI_3 NS_395 0 -5.5808215669255444e-03
GC_3_396 b_3 NI_3 NS_396 0 -6.8969143321972607e-03
GC_3_397 b_3 NI_3 NS_397 0 1.1228129967359635e-02
GC_3_398 b_3 NI_3 NS_398 0 -1.3571857960940519e-03
GC_3_399 b_3 NI_3 NS_399 0 1.5726428598145797e-02
GC_3_400 b_3 NI_3 NS_400 0 1.2982469555517450e-02
GC_3_401 b_3 NI_3 NS_401 0 -7.1842587552582117e-03
GC_3_402 b_3 NI_3 NS_402 0 5.1249277034737355e-03
GC_3_403 b_3 NI_3 NS_403 0 -6.8612317657539322e-03
GC_3_404 b_3 NI_3 NS_404 0 -4.8303542718685869e-03
GC_3_405 b_3 NI_3 NS_405 0 5.1299879581948227e-09
GC_3_406 b_3 NI_3 NS_406 0 4.4376477008264907e-08
GC_3_407 b_3 NI_3 NS_407 0 1.2002066367289146e-02
GC_3_408 b_3 NI_3 NS_408 0 -2.5554094200757925e-03
GC_3_409 b_3 NI_3 NS_409 0 -5.2431655551256357e-03
GC_3_410 b_3 NI_3 NS_410 0 4.7077253049496535e-03
GC_3_411 b_3 NI_3 NS_411 0 -6.1541411405470385e-03
GC_3_412 b_3 NI_3 NS_412 0 -4.3159764406445356e-03
GC_3_413 b_3 NI_3 NS_413 0 1.1759646160199927e-02
GC_3_414 b_3 NI_3 NS_414 0 -3.7148872059305773e-03
GC_3_415 b_3 NI_3 NS_415 0 1.3000704175392007e-02
GC_3_416 b_3 NI_3 NS_416 0 9.4708329982350365e-03
GC_3_417 b_3 NI_3 NS_417 0 3.9444945149576896e-06
GC_3_418 b_3 NI_3 NS_418 0 -9.3341531512143170e-07
GC_3_419 b_3 NI_3 NS_419 0 1.6111754337009596e-02
GC_3_420 b_3 NI_3 NS_420 0 1.6784786344276582e-02
GC_3_421 b_3 NI_3 NS_421 0 1.2052343780144359e-02
GC_3_422 b_3 NI_3 NS_422 0 -2.4747684933194899e-03
GC_3_423 b_3 NI_3 NS_423 0 -8.3473638986931668e-03
GC_3_424 b_3 NI_3 NS_424 0 8.3965897925197575e-05
GC_3_425 b_3 NI_3 NS_425 0 1.1340540049644776e-02
GC_3_426 b_3 NI_3 NS_426 0 7.3400048894673442e-03
GC_3_427 b_3 NI_3 NS_427 0 -4.6549307283898890e-03
GC_3_428 b_3 NI_3 NS_428 0 7.3654587140112035e-03
GC_3_429 b_3 NI_3 NS_429 0 -8.0793093651674776e-03
GC_3_430 b_3 NI_3 NS_430 0 -3.7190000439631414e-03
GC_3_431 b_3 NI_3 NS_431 0 1.5982957914344887e-02
GC_3_432 b_3 NI_3 NS_432 0 -7.7385034283743628e-03
GC_3_433 b_3 NI_3 NS_433 0 7.9288748341783754e-05
GC_3_434 b_3 NI_3 NS_434 0 -1.2174290498918229e-10
GC_3_435 b_3 NI_3 NS_435 0 -2.0288821135085861e-09
GC_3_436 b_3 NI_3 NS_436 0 3.4022340611109259e-08
GC_3_437 b_3 NI_3 NS_437 0 -3.3983706540759051e-07
GC_3_438 b_3 NI_3 NS_438 0 -3.3574280506251254e-07
GC_3_439 b_3 NI_3 NS_439 0 -5.7584237066819604e-07
GC_3_440 b_3 NI_3 NS_440 0 9.6675316399059596e-06
GC_3_441 b_3 NI_3 NS_441 0 1.3105676203469716e-05
GC_3_442 b_3 NI_3 NS_442 0 -1.2342181898532230e-05
GC_3_443 b_3 NI_3 NS_443 0 -1.7112606669997782e-05
GC_3_444 b_3 NI_3 NS_444 0 8.5764475609902259e-06
GC_3_445 b_3 NI_3 NS_445 0 2.8663170574135972e-05
GC_3_446 b_3 NI_3 NS_446 0 -7.4194705102769838e-06
GC_3_447 b_3 NI_3 NS_447 0 -2.8956659037482216e-06
GC_3_448 b_3 NI_3 NS_448 0 -3.4130743251428452e-06
GC_3_449 b_3 NI_3 NS_449 0 -3.2449805614179802e-06
GC_3_450 b_3 NI_3 NS_450 0 -1.5090311680546233e-05
GC_3_451 b_3 NI_3 NS_451 0 -2.4828337522431015e-05
GC_3_452 b_3 NI_3 NS_452 0 3.9221720996960387e-05
GC_3_453 b_3 NI_3 NS_453 0 3.6987644135395511e-05
GC_3_454 b_3 NI_3 NS_454 0 -4.7225340727116541e-05
GC_3_455 b_3 NI_3 NS_455 0 -3.0518339486996669e-05
GC_3_456 b_3 NI_3 NS_456 0 -2.1425302238833142e-05
GC_3_457 b_3 NI_3 NS_457 0 3.2014657783478431e-05
GC_3_458 b_3 NI_3 NS_458 0 2.6387854880322412e-05
GC_3_459 b_3 NI_3 NS_459 0 -1.8545633870928283e-05
GC_3_460 b_3 NI_3 NS_460 0 -2.9076395091484659e-05
GC_3_461 b_3 NI_3 NS_461 0 2.0026492549390195e-05
GC_3_462 b_3 NI_3 NS_462 0 5.9804794277143845e-05
GC_3_463 b_3 NI_3 NS_463 0 -2.0977330446605740e-05
GC_3_464 b_3 NI_3 NS_464 0 -5.5613753317647659e-05
GC_3_465 b_3 NI_3 NS_465 0 -3.1646152877825364e-05
GC_3_466 b_3 NI_3 NS_466 0 -1.2116541129766774e-05
GC_3_467 b_3 NI_3 NS_467 0 1.9561870604874970e-05
GC_3_468 b_3 NI_3 NS_468 0 1.3806626372669835e-05
GC_3_469 b_3 NI_3 NS_469 0 -2.4957198229610124e-05
GC_3_470 b_3 NI_3 NS_470 0 -1.1262318003650680e-05
GC_3_471 b_3 NI_3 NS_471 0 2.0179937061848243e-05
GC_3_472 b_3 NI_3 NS_472 0 1.0341638971073189e-05
GC_3_473 b_3 NI_3 NS_473 0 -1.8434218520807260e-05
GC_3_474 b_3 NI_3 NS_474 0 -2.1152540806707857e-05
GC_3_475 b_3 NI_3 NS_475 0 4.2957734764276978e-06
GC_3_476 b_3 NI_3 NS_476 0 3.1958081815041139e-05
GC_3_477 b_3 NI_3 NS_477 0 -8.4065274554809462e-06
GC_3_478 b_3 NI_3 NS_478 0 -2.6582396550238322e-05
GC_3_479 b_3 NI_3 NS_479 0 -2.0402889636585728e-06
GC_3_480 b_3 NI_3 NS_480 0 1.5416007903730722e-06
GC_3_481 b_3 NI_3 NS_481 0 -1.9679904543878262e-05
GC_3_482 b_3 NI_3 NS_482 0 -1.2198708946806058e-05
GC_3_483 b_3 NI_3 NS_483 0 5.5390013850228335e-06
GC_3_484 b_3 NI_3 NS_484 0 2.1304114163880079e-05
GC_3_485 b_3 NI_3 NS_485 0 -1.6263704465232622e-05
GC_3_486 b_3 NI_3 NS_486 0 -1.4842861466753822e-05
GC_3_487 b_3 NI_3 NS_487 0 9.0210293868592366e-07
GC_3_488 b_3 NI_3 NS_488 0 5.5179733349875214e-06
GC_3_489 b_3 NI_3 NS_489 0 -2.5230906486445864e-05
GC_3_490 b_3 NI_3 NS_490 0 -1.0007044019372768e-05
GC_3_491 b_3 NI_3 NS_491 0 7.5032639170213123e-06
GC_3_492 b_3 NI_3 NS_492 0 2.3878271962760899e-05
GC_3_493 b_3 NI_3 NS_493 0 -2.0944112847441730e-05
GC_3_494 b_3 NI_3 NS_494 0 -5.6385636149592013e-06
GC_3_495 b_3 NI_3 NS_495 0 5.9392842791228235e-06
GC_3_496 b_3 NI_3 NS_496 0 7.9059437617353887e-06
GC_3_497 b_3 NI_3 NS_497 0 -3.0918933331932639e-05
GC_3_498 b_3 NI_3 NS_498 0 -2.7455168685233037e-06
GC_3_499 b_3 NI_3 NS_499 0 1.8051694416579107e-05
GC_3_500 b_3 NI_3 NS_500 0 2.6172444898805574e-05
GC_3_501 b_3 NI_3 NS_501 0 -2.2120772574608656e-05
GC_3_502 b_3 NI_3 NS_502 0 6.9971038447442136e-06
GC_3_503 b_3 NI_3 NS_503 0 1.5076743764700976e-05
GC_3_504 b_3 NI_3 NS_504 0 4.4857559945435255e-06
GC_3_505 b_3 NI_3 NS_505 0 -3.5006192574239558e-05
GC_3_506 b_3 NI_3 NS_506 0 1.3594831215997829e-05
GC_3_507 b_3 NI_3 NS_507 0 3.7185054377027495e-05
GC_3_508 b_3 NI_3 NS_508 0 1.3344808135759734e-05
GC_3_509 b_3 NI_3 NS_509 0 -7.9971580078133745e-06
GC_3_510 b_3 NI_3 NS_510 0 1.9077538238115875e-05
GC_3_511 b_3 NI_3 NS_511 0 1.2877243884352367e-05
GC_3_512 b_3 NI_3 NS_512 0 -1.0947055945521094e-05
GC_3_513 b_3 NI_3 NS_513 0 1.1098886880365967e-10
GC_3_514 b_3 NI_3 NS_514 0 4.4127842986745474e-11
GC_3_515 b_3 NI_3 NS_515 0 -1.3992975810812636e-05
GC_3_516 b_3 NI_3 NS_516 0 2.6116738052306620e-05
GC_3_517 b_3 NI_3 NS_517 0 -2.1466200625312570e-06
GC_3_518 b_3 NI_3 NS_518 0 1.0636847987244859e-05
GC_3_519 b_3 NI_3 NS_519 0 6.1623437997495518e-06
GC_3_520 b_3 NI_3 NS_520 0 -8.3666721060721817e-06
GC_3_521 b_3 NI_3 NS_521 0 -8.3609173283029481e-06
GC_3_522 b_3 NI_3 NS_522 0 2.5491814870143550e-05
GC_3_523 b_3 NI_3 NS_523 0 2.5015772430524796e-05
GC_3_524 b_3 NI_3 NS_524 0 -9.9981297101173857e-06
GC_3_525 b_3 NI_3 NS_525 0 4.8733518400475768e-09
GC_3_526 b_3 NI_3 NS_526 0 -1.1063144989205645e-09
GC_3_527 b_3 NI_3 NS_527 0 2.6321680400281924e-05
GC_3_528 b_3 NI_3 NS_528 0 -1.2477251716174242e-05
GC_3_529 b_3 NI_3 NS_529 0 -8.3190505039735985e-06
GC_3_530 b_3 NI_3 NS_530 0 1.8150061678833330e-05
GC_3_531 b_3 NI_3 NS_531 0 -1.0398845371621847e-05
GC_3_532 b_3 NI_3 NS_532 0 -2.8340376542205747e-07
GC_3_533 b_3 NI_3 NS_533 0 1.9410929087432574e-05
GC_3_534 b_3 NI_3 NS_534 0 -1.4077513684575097e-05
GC_3_535 b_3 NI_3 NS_535 0 7.1590830116475085e-06
GC_3_536 b_3 NI_3 NS_536 0 1.1754924633469265e-05
GC_3_537 b_3 NI_3 NS_537 0 -1.8100728828436785e-07
GC_3_538 b_3 NI_3 NS_538 0 -1.4547290501063122e-05
GC_3_539 b_3 NI_3 NS_539 0 1.3082934467548369e-05
GC_3_540 b_3 NI_3 NS_540 0 2.7942030080176412e-05
GC_3_541 b_3 NI_3 NS_541 0 -6.4096519279402203e-04
GC_3_542 b_3 NI_3 NS_542 0 -9.7194678094467582e-11
GC_3_543 b_3 NI_3 NS_543 0 3.8858048973612838e-09
GC_3_544 b_3 NI_3 NS_544 0 -6.7398839160299627e-08
GC_3_545 b_3 NI_3 NS_545 0 -1.1319905633218811e-05
GC_3_546 b_3 NI_3 NS_546 0 -9.3647684152654186e-06
GC_3_547 b_3 NI_3 NS_547 0 -2.2431735877849280e-06
GC_3_548 b_3 NI_3 NS_548 0 2.0358449381248975e-07
GC_3_549 b_3 NI_3 NS_549 0 -3.0429847449436261e-05
GC_3_550 b_3 NI_3 NS_550 0 2.7128787601797520e-05
GC_3_551 b_3 NI_3 NS_551 0 -3.3446191161219447e-05
GC_3_552 b_3 NI_3 NS_552 0 8.1023558296294296e-06
GC_3_553 b_3 NI_3 NS_553 0 3.1775639518541672e-05
GC_3_554 b_3 NI_3 NS_554 0 2.7493584539289286e-05
GC_3_555 b_3 NI_3 NS_555 0 -9.1079431664587748e-06
GC_3_556 b_3 NI_3 NS_556 0 1.4797969144889177e-05
GC_3_557 b_3 NI_3 NS_557 0 1.2654200668661801e-05
GC_3_558 b_3 NI_3 NS_558 0 3.7136155294312760e-05
GC_3_559 b_3 NI_3 NS_559 0 -1.1049973462363621e-05
GC_3_560 b_3 NI_3 NS_560 0 6.8460617275802066e-05
GC_3_561 b_3 NI_3 NS_561 0 9.6052096916483432e-05
GC_3_562 b_3 NI_3 NS_562 0 -6.6220028657107001e-05
GC_3_563 b_3 NI_3 NS_563 0 2.7188453061815506e-05
GC_3_564 b_3 NI_3 NS_564 0 3.2025518863967084e-05
GC_3_565 b_3 NI_3 NS_565 0 -6.9721051049947644e-06
GC_3_566 b_3 NI_3 NS_566 0 -7.2660798313216936e-05
GC_3_567 b_3 NI_3 NS_567 0 -9.8238618683368669e-06
GC_3_568 b_3 NI_3 NS_568 0 -3.4299021975996833e-05
GC_3_569 b_3 NI_3 NS_569 0 -7.6898749304986813e-05
GC_3_570 b_3 NI_3 NS_570 0 1.8642126554274563e-05
GC_3_571 b_3 NI_3 NS_571 0 2.4833373731533620e-05
GC_3_572 b_3 NI_3 NS_572 0 5.1420164959051402e-05
GC_3_573 b_3 NI_3 NS_573 0 -2.3340307786250049e-05
GC_3_574 b_3 NI_3 NS_574 0 -3.7721117528948561e-06
GC_3_575 b_3 NI_3 NS_575 0 7.0064431078953023e-05
GC_3_576 b_3 NI_3 NS_576 0 4.4958994735634309e-05
GC_3_577 b_3 NI_3 NS_577 0 2.9394323101390281e-05
GC_3_578 b_3 NI_3 NS_578 0 1.9999802850201240e-05
GC_3_579 b_3 NI_3 NS_579 0 -7.2203598085392578e-06
GC_3_580 b_3 NI_3 NS_580 0 -2.5839480579585212e-05
GC_3_581 b_3 NI_3 NS_581 0 -7.5634334036366812e-06
GC_3_582 b_3 NI_3 NS_582 0 -2.5468696398961454e-05
GC_3_583 b_3 NI_3 NS_583 0 6.9064332007064558e-06
GC_3_584 b_3 NI_3 NS_584 0 4.9199292095002321e-05
GC_3_585 b_3 NI_3 NS_585 0 1.2870888594969830e-05
GC_3_586 b_3 NI_3 NS_586 0 2.7631523311755763e-05
GC_3_587 b_3 NI_3 NS_587 0 5.8803260015810867e-06
GC_3_588 b_3 NI_3 NS_588 0 2.1449596447860135e-06
GC_3_589 b_3 NI_3 NS_589 0 -6.1110748726733272e-07
GC_3_590 b_3 NI_3 NS_590 0 -1.5594150858490844e-05
GC_3_591 b_3 NI_3 NS_591 0 5.6392040310862021e-05
GC_3_592 b_3 NI_3 NS_592 0 3.8210555801440701e-05
GC_3_593 b_3 NI_3 NS_593 0 1.9988519947754532e-05
GC_3_594 b_3 NI_3 NS_594 0 1.5010231953626078e-05
GC_3_595 b_3 NI_3 NS_595 0 8.4379867511083121e-06
GC_3_596 b_3 NI_3 NS_596 0 -1.2896798787930660e-05
GC_3_597 b_3 NI_3 NS_597 0 -5.6459236552622443e-06
GC_3_598 b_3 NI_3 NS_598 0 -1.4204662005227251e-05
GC_3_599 b_3 NI_3 NS_599 0 6.6278849803423341e-05
GC_3_600 b_3 NI_3 NS_600 0 1.2995847847199136e-05
GC_3_601 b_3 NI_3 NS_601 0 2.2839924688685369e-05
GC_3_602 b_3 NI_3 NS_602 0 5.0561044121262851e-06
GC_3_603 b_3 NI_3 NS_603 0 -5.5482128057890352e-06
GC_3_604 b_3 NI_3 NS_604 0 -2.2088160755117591e-05
GC_3_605 b_3 NI_3 NS_605 0 -9.1406501875523818e-06
GC_3_606 b_3 NI_3 NS_606 0 -7.2230791469077473e-06
GC_3_607 b_3 NI_3 NS_607 0 6.0751022676375617e-05
GC_3_608 b_3 NI_3 NS_608 0 -9.5212285484179220e-06
GC_3_609 b_3 NI_3 NS_609 0 2.1480532300696621e-05
GC_3_610 b_3 NI_3 NS_610 0 -7.3371799289233979e-06
GC_3_611 b_3 NI_3 NS_611 0 -2.3109770418999255e-05
GC_3_612 b_3 NI_3 NS_612 0 -1.3195890149297649e-05
GC_3_613 b_3 NI_3 NS_613 0 -8.6441676931997166e-06
GC_3_614 b_3 NI_3 NS_614 0 4.3874538123759307e-06
GC_3_615 b_3 NI_3 NS_615 0 4.5483159545880018e-05
GC_3_616 b_3 NI_3 NS_616 0 -2.5698442967621768e-05
GC_3_617 b_3 NI_3 NS_617 0 6.0412477482498822e-06
GC_3_618 b_3 NI_3 NS_618 0 -1.6494038841537749e-05
GC_3_619 b_3 NI_3 NS_619 0 -1.8742827362044494e-05
GC_3_620 b_3 NI_3 NS_620 0 8.5986466268740750e-06
GC_3_621 b_3 NI_3 NS_621 0 -4.6792761378612171e-11
GC_3_622 b_3 NI_3 NS_622 0 -1.7807240794879957e-10
GC_3_623 b_3 NI_3 NS_623 0 1.7713032240626713e-06
GC_3_624 b_3 NI_3 NS_624 0 8.7581319339666863e-06
GC_3_625 b_3 NI_3 NS_625 0 2.2084503476230542e-06
GC_3_626 b_3 NI_3 NS_626 0 -7.0117486289654574e-06
GC_3_627 b_3 NI_3 NS_627 0 -9.0106068019312138e-06
GC_3_628 b_3 NI_3 NS_628 0 5.7573252376648386e-06
GC_3_629 b_3 NI_3 NS_629 0 4.7874443214052022e-06
GC_3_630 b_3 NI_3 NS_630 0 1.1558466898826803e-05
GC_3_631 b_3 NI_3 NS_631 0 2.4565262871639701e-05
GC_3_632 b_3 NI_3 NS_632 0 -2.1165220938800276e-05
GC_3_633 b_3 NI_3 NS_633 0 -5.7150012037119728e-09
GC_3_634 b_3 NI_3 NS_634 0 -5.6483319108174473e-09
GC_3_635 b_3 NI_3 NS_635 0 3.0655890404757572e-05
GC_3_636 b_3 NI_3 NS_636 0 7.4872133548011052e-06
GC_3_637 b_3 NI_3 NS_637 0 -2.6797308961936641e-06
GC_3_638 b_3 NI_3 NS_638 0 1.1045237531599606e-05
GC_3_639 b_3 NI_3 NS_639 0 8.0410643541720206e-06
GC_3_640 b_3 NI_3 NS_640 0 1.1946460101207240e-06
GC_3_641 b_3 NI_3 NS_641 0 1.9120714183249608e-05
GC_3_642 b_3 NI_3 NS_642 0 -2.1559499832323254e-05
GC_3_643 b_3 NI_3 NS_643 0 -6.5502994872348925e-06
GC_3_644 b_3 NI_3 NS_644 0 -7.4615405536929573e-06
GC_3_645 b_3 NI_3 NS_645 0 -5.3942508467503822e-06
GC_3_646 b_3 NI_3 NS_646 0 1.2484971087039410e-05
GC_3_647 b_3 NI_3 NS_647 0 1.6111580163334561e-05
GC_3_648 b_3 NI_3 NS_648 0 7.3766059220711541e-06
GC_3_649 b_3 NI_3 NS_649 0 -2.7355542573336887e-05
GC_3_650 b_3 NI_3 NS_650 0 -9.2005620290625430e-13
GC_3_651 b_3 NI_3 NS_651 0 -2.3520837613857581e-10
GC_3_652 b_3 NI_3 NS_652 0 1.0469206461162468e-08
GC_3_653 b_3 NI_3 NS_653 0 7.2942592001678264e-07
GC_3_654 b_3 NI_3 NS_654 0 1.1057573129455704e-07
GC_3_655 b_3 NI_3 NS_655 0 3.2329357560442220e-06
GC_3_656 b_3 NI_3 NS_656 0 -1.3955668005341952e-06
GC_3_657 b_3 NI_3 NS_657 0 -2.7334272216021501e-06
GC_3_658 b_3 NI_3 NS_658 0 -2.8887391788089376e-06
GC_3_659 b_3 NI_3 NS_659 0 5.0379778952158204e-06
GC_3_660 b_3 NI_3 NS_660 0 -5.9339261020989814e-07
GC_3_661 b_3 NI_3 NS_661 0 -7.0890001648592670e-06
GC_3_662 b_3 NI_3 NS_662 0 -8.3126031260027058e-06
GC_3_663 b_3 NI_3 NS_663 0 8.1233576627629320e-08
GC_3_664 b_3 NI_3 NS_664 0 -1.6105145685008275e-06
GC_3_665 b_3 NI_3 NS_665 0 -6.1810004255555138e-06
GC_3_666 b_3 NI_3 NS_666 0 1.8479511773914306e-06
GC_3_667 b_3 NI_3 NS_667 0 5.4033093663502904e-06
GC_3_668 b_3 NI_3 NS_668 0 -6.0039261741008855e-06
GC_3_669 b_3 NI_3 NS_669 0 -1.7425745696427919e-05
GC_3_670 b_3 NI_3 NS_670 0 4.6515785310191588e-06
GC_3_671 b_3 NI_3 NS_671 0 -1.1775863834592140e-06
GC_3_672 b_3 NI_3 NS_672 0 7.0644007074382843e-06
GC_3_673 b_3 NI_3 NS_673 0 -7.5195205679586350e-06
GC_3_674 b_3 NI_3 NS_674 0 -4.7823989772047162e-06
GC_3_675 b_3 NI_3 NS_675 0 -3.4396136734242288e-06
GC_3_676 b_3 NI_3 NS_676 0 8.0393796503332119e-06
GC_3_677 b_3 NI_3 NS_677 0 -2.5304451111156507e-06
GC_3_678 b_3 NI_3 NS_678 0 -4.9642139260598833e-06
GC_3_679 b_3 NI_3 NS_679 0 -3.8886555572790891e-06
GC_3_680 b_3 NI_3 NS_680 0 1.1491298838636697e-05
GC_3_681 b_3 NI_3 NS_681 0 -1.9009350759163734e-07
GC_3_682 b_3 NI_3 NS_682 0 7.1731153291547707e-06
GC_3_683 b_3 NI_3 NS_683 0 -4.3615428945145289e-06
GC_3_684 b_3 NI_3 NS_684 0 1.1394832480417147e-06
GC_3_685 b_3 NI_3 NS_685 0 -6.9161343786112695e-07
GC_3_686 b_3 NI_3 NS_686 0 7.9938192472556748e-06
GC_3_687 b_3 NI_3 NS_687 0 -1.2344330937587836e-06
GC_3_688 b_3 NI_3 NS_688 0 2.1996720984501816e-06
GC_3_689 b_3 NI_3 NS_689 0 -2.4841809849453658e-06
GC_3_690 b_3 NI_3 NS_690 0 8.1284198547710831e-06
GC_3_691 b_3 NI_3 NS_691 0 -4.1621104739951376e-07
GC_3_692 b_3 NI_3 NS_692 0 9.3187005230972797e-06
GC_3_693 b_3 NI_3 NS_693 0 -9.6408205333558304e-07
GC_3_694 b_3 NI_3 NS_694 0 8.8146488298289406e-06
GC_3_695 b_3 NI_3 NS_695 0 -1.3883421605481633e-06
GC_3_696 b_3 NI_3 NS_696 0 3.8439571781940877e-06
GC_3_697 b_3 NI_3 NS_697 0 8.6419624895523205e-07
GC_3_698 b_3 NI_3 NS_698 0 1.1901958874041500e-05
GC_3_699 b_3 NI_3 NS_699 0 1.7097639557248967e-05
GC_3_700 b_3 NI_3 NS_700 0 1.6762494103210088e-05
GC_3_701 b_3 NI_3 NS_701 0 4.6416751531732292e-06
GC_3_702 b_3 NI_3 NS_702 0 7.7284891826678090e-06
GC_3_703 b_3 NI_3 NS_703 0 9.7558221382078173e-06
GC_3_704 b_3 NI_3 NS_704 0 3.9053282543285631e-06
GC_3_705 b_3 NI_3 NS_705 0 6.3770740827166772e-06
GC_3_706 b_3 NI_3 NS_706 0 1.0690285666587357e-05
GC_3_707 b_3 NI_3 NS_707 0 3.1851231961764098e-05
GC_3_708 b_3 NI_3 NS_708 0 -5.6094616373767788e-06
GC_3_709 b_3 NI_3 NS_709 0 7.7676140594365746e-06
GC_3_710 b_3 NI_3 NS_710 0 3.4156071244945016e-06
GC_3_711 b_3 NI_3 NS_711 0 1.1409487215695193e-05
GC_3_712 b_3 NI_3 NS_712 0 -9.8749569507264013e-06
GC_3_713 b_3 NI_3 NS_713 0 1.0301967532235236e-05
GC_3_714 b_3 NI_3 NS_714 0 6.2888523140750239e-06
GC_3_715 b_3 NI_3 NS_715 0 1.5924361430783647e-05
GC_3_716 b_3 NI_3 NS_716 0 -2.9747673328769177e-05
GC_3_717 b_3 NI_3 NS_717 0 7.6974769090524504e-06
GC_3_718 b_3 NI_3 NS_718 0 -2.8352585871025316e-06
GC_3_719 b_3 NI_3 NS_719 0 -3.4077947491967134e-06
GC_3_720 b_3 NI_3 NS_720 0 -1.5676420398830460e-05
GC_3_721 b_3 NI_3 NS_721 0 1.1261363855137156e-05
GC_3_722 b_3 NI_3 NS_722 0 -1.6843785186933320e-06
GC_3_723 b_3 NI_3 NS_723 0 -1.2932102918271445e-05
GC_3_724 b_3 NI_3 NS_724 0 -2.4084153779413579e-05
GC_3_725 b_3 NI_3 NS_725 0 -4.1147783057531965e-07
GC_3_726 b_3 NI_3 NS_726 0 -6.3604259976744664e-06
GC_3_727 b_3 NI_3 NS_727 0 -9.4858826249718311e-06
GC_3_728 b_3 NI_3 NS_728 0 -2.3359061317560598e-06
GC_3_729 b_3 NI_3 NS_729 0 9.8167963223250750e-11
GC_3_730 b_3 NI_3 NS_730 0 5.4215162430425681e-11
GC_3_731 b_3 NI_3 NS_731 0 1.1810241566230886e-06
GC_3_732 b_3 NI_3 NS_732 0 -4.5943645360185014e-06
GC_3_733 b_3 NI_3 NS_733 0 -1.4778925100888582e-06
GC_3_734 b_3 NI_3 NS_734 0 -1.2797106260282140e-06
GC_3_735 b_3 NI_3 NS_735 0 -4.9247464723251121e-06
GC_3_736 b_3 NI_3 NS_736 0 -8.6882657284496607e-07
GC_3_737 b_3 NI_3 NS_737 0 -1.3801285827474389e-06
GC_3_738 b_3 NI_3 NS_738 0 -2.8355643244125362e-06
GC_3_739 b_3 NI_3 NS_739 0 -1.0039741583070359e-05
GC_3_740 b_3 NI_3 NS_740 0 -3.6814540166324874e-06
GC_3_741 b_3 NI_3 NS_741 0 6.6579466416904979e-09
GC_3_742 b_3 NI_3 NS_742 0 5.7676980937849128e-09
GC_3_743 b_3 NI_3 NS_743 0 1.3984242907929010e-06
GC_3_744 b_3 NI_3 NS_744 0 6.7801360111326123e-07
GC_3_745 b_3 NI_3 NS_745 0 -1.7284101334476144e-06
GC_3_746 b_3 NI_3 NS_746 0 3.1540252409498978e-06
GC_3_747 b_3 NI_3 NS_747 0 -9.2400628204016724e-07
GC_3_748 b_3 NI_3 NS_748 0 7.7572763025873638e-07
GC_3_749 b_3 NI_3 NS_749 0 -7.9033350197252917e-06
GC_3_750 b_3 NI_3 NS_750 0 8.3212762913432852e-07
GC_3_751 b_3 NI_3 NS_751 0 -2.4107255645528072e-06
GC_3_752 b_3 NI_3 NS_752 0 2.0829180595171174e-06
GC_3_753 b_3 NI_3 NS_753 0 -2.1271854147244160e-06
GC_3_754 b_3 NI_3 NS_754 0 2.1516734688725426e-06
GC_3_755 b_3 NI_3 NS_755 0 1.1284198633010088e-06
GC_3_756 b_3 NI_3 NS_756 0 2.8125734757496343e-06
GC_3_757 b_3 NI_3 NS_757 0 -1.4436375625828516e-04
GC_3_758 b_3 NI_3 NS_758 0 3.3291262807282880e-11
GC_3_759 b_3 NI_3 NS_759 0 3.9882304085378514e-11
GC_3_760 b_3 NI_3 NS_760 0 9.0903451459516971e-10
GC_3_761 b_3 NI_3 NS_761 0 -2.1100781772492012e-06
GC_3_762 b_3 NI_3 NS_762 0 -1.6555673626595899e-06
GC_3_763 b_3 NI_3 NS_763 0 1.8947206183832116e-06
GC_3_764 b_3 NI_3 NS_764 0 3.8512917548461082e-06
GC_3_765 b_3 NI_3 NS_765 0 3.3113004589310871e-06
GC_3_766 b_3 NI_3 NS_766 0 4.9314150725341936e-06
GC_3_767 b_3 NI_3 NS_767 0 5.8708133977770993e-06
GC_3_768 b_3 NI_3 NS_768 0 -9.1115743321420913e-06
GC_3_769 b_3 NI_3 NS_769 0 -2.5609911787096947e-06
GC_3_770 b_3 NI_3 NS_770 0 -1.3919625232812814e-05
GC_3_771 b_3 NI_3 NS_771 0 -3.5429291322449613e-06
GC_3_772 b_3 NI_3 NS_772 0 2.1898060105718448e-06
GC_3_773 b_3 NI_3 NS_773 0 3.6501944544711360e-06
GC_3_774 b_3 NI_3 NS_774 0 1.2869477834530357e-06
GC_3_775 b_3 NI_3 NS_775 0 8.0000509509074179e-06
GC_3_776 b_3 NI_3 NS_776 0 -3.9897559213308073e-05
GC_3_777 b_3 NI_3 NS_777 0 -4.4313712016731078e-05
GC_3_778 b_3 NI_3 NS_778 0 -9.3697261704138949e-07
GC_3_779 b_3 NI_3 NS_779 0 -1.4827741223220499e-05
GC_3_780 b_3 NI_3 NS_780 0 -8.5761185394940832e-06
GC_3_781 b_3 NI_3 NS_781 0 -7.2939514907894413e-05
GC_3_782 b_3 NI_3 NS_782 0 7.5520236112830468e-05
GC_3_783 b_3 NI_3 NS_783 0 4.6289615426040011e-06
GC_3_784 b_3 NI_3 NS_784 0 1.3120054088590003e-05
GC_3_785 b_3 NI_3 NS_785 0 6.2840278321967362e-05
GC_3_786 b_3 NI_3 NS_786 0 1.2319963836453509e-04
GC_3_787 b_3 NI_3 NS_787 0 3.6326948481249521e-07
GC_3_788 b_3 NI_3 NS_788 0 -3.7019877498736819e-05
GC_3_789 b_3 NI_3 NS_789 0 1.6508678116810902e-05
GC_3_790 b_3 NI_3 NS_790 0 3.9672161038711577e-06
GC_3_791 b_3 NI_3 NS_791 0 2.4447787489406659e-05
GC_3_792 b_3 NI_3 NS_792 0 -3.0457961836901388e-05
GC_3_793 b_3 NI_3 NS_793 0 -8.8967728077273195e-06
GC_3_794 b_3 NI_3 NS_794 0 -2.3402119593525554e-06
GC_3_795 b_3 NI_3 NS_795 0 -8.8832896256785692e-06
GC_3_796 b_3 NI_3 NS_796 0 2.5237309406570649e-05
GC_3_797 b_3 NI_3 NS_797 0 5.8267206950776330e-06
GC_3_798 b_3 NI_3 NS_798 0 8.4670732341507218e-06
GC_3_799 b_3 NI_3 NS_799 0 5.6328289039083256e-05
GC_3_800 b_3 NI_3 NS_800 0 2.4970028923784872e-05
GC_3_801 b_3 NI_3 NS_801 0 3.5271326637809141e-06
GC_3_802 b_3 NI_3 NS_802 0 -1.1687101824654425e-05
GC_3_803 b_3 NI_3 NS_803 0 -4.0893823518938578e-07
GC_3_804 b_3 NI_3 NS_804 0 -1.3155542605580849e-06
GC_3_805 b_3 NI_3 NS_805 0 6.8059479317462960e-06
GC_3_806 b_3 NI_3 NS_806 0 3.0643166767038212e-06
GC_3_807 b_3 NI_3 NS_807 0 4.1947328182121476e-05
GC_3_808 b_3 NI_3 NS_808 0 -1.7198850686061673e-05
GC_3_809 b_3 NI_3 NS_809 0 -2.5587381648522656e-06
GC_3_810 b_3 NI_3 NS_810 0 -7.0969089496108462e-06
GC_3_811 b_3 NI_3 NS_811 0 -3.0311305667412328e-06
GC_3_812 b_3 NI_3 NS_812 0 1.7555145239758741e-06
GC_3_813 b_3 NI_3 NS_813 0 9.5694183774174486e-06
GC_3_814 b_3 NI_3 NS_814 0 2.9161061638379040e-06
GC_3_815 b_3 NI_3 NS_815 0 2.2975734843631131e-05
GC_3_816 b_3 NI_3 NS_816 0 -3.1187525516132392e-05
GC_3_817 b_3 NI_3 NS_817 0 -5.6937387719374329e-06
GC_3_818 b_3 NI_3 NS_818 0 -3.6756787372355002e-06
GC_3_819 b_3 NI_3 NS_819 0 -5.6139609185501988e-07
GC_3_820 b_3 NI_3 NS_820 0 5.0284658224451405e-06
GC_3_821 b_3 NI_3 NS_821 0 1.2292599868045946e-05
GC_3_822 b_3 NI_3 NS_822 0 2.0421157533764655e-07
GC_3_823 b_3 NI_3 NS_823 0 1.9184489557658854e-06
GC_3_824 b_3 NI_3 NS_824 0 -3.1503446941607862e-05
GC_3_825 b_3 NI_3 NS_825 0 -6.7231145433544231e-06
GC_3_826 b_3 NI_3 NS_826 0 9.4627912001846438e-07
GC_3_827 b_3 NI_3 NS_827 0 4.5912669843495469e-06
GC_3_828 b_3 NI_3 NS_828 0 3.8667933862349351e-06
GC_3_829 b_3 NI_3 NS_829 0 1.4096552359487495e-05
GC_3_830 b_3 NI_3 NS_830 0 -6.0051965043248030e-06
GC_3_831 b_3 NI_3 NS_831 0 -1.3991398843112036e-05
GC_3_832 b_3 NI_3 NS_832 0 -1.8834214408005415e-05
GC_3_833 b_3 NI_3 NS_833 0 -2.5005337400052953e-06
GC_3_834 b_3 NI_3 NS_834 0 5.3959384179046051e-06
GC_3_835 b_3 NI_3 NS_835 0 4.6402364167576557e-06
GC_3_836 b_3 NI_3 NS_836 0 -2.0953558108470921e-06
GC_3_837 b_3 NI_3 NS_837 0 -1.4466664248636737e-11
GC_3_838 b_3 NI_3 NS_838 0 3.9862275905169703e-12
GC_3_839 b_3 NI_3 NS_839 0 5.2050488123223110e-06
GC_3_840 b_3 NI_3 NS_840 0 -1.1255636414838616e-05
GC_3_841 b_3 NI_3 NS_841 0 -2.6207638208057526e-07
GC_3_842 b_3 NI_3 NS_842 0 2.9240728178134803e-06
GC_3_843 b_3 NI_3 NS_843 0 2.6491372006687385e-06
GC_3_844 b_3 NI_3 NS_844 0 -1.6106173652973849e-06
GC_3_845 b_3 NI_3 NS_845 0 2.4311226641432671e-06
GC_3_846 b_3 NI_3 NS_846 0 -9.4257142084186216e-06
GC_3_847 b_3 NI_3 NS_847 0 -9.9190992713045025e-06
GC_3_848 b_3 NI_3 NS_848 0 -3.6952579499555889e-06
GC_3_849 b_3 NI_3 NS_849 0 3.1959411841289133e-10
GC_3_850 b_3 NI_3 NS_850 0 2.6405667791978424e-10
GC_3_851 b_3 NI_3 NS_851 0 -8.5810808148530714e-06
GC_3_852 b_3 NI_3 NS_852 0 -5.7196684179012733e-06
GC_3_853 b_3 NI_3 NS_853 0 2.2759099727273564e-06
GC_3_854 b_3 NI_3 NS_854 0 -6.4442878822626431e-06
GC_3_855 b_3 NI_3 NS_855 0 -3.0692757627501459e-06
GC_3_856 b_3 NI_3 NS_856 0 -1.3767164209917423e-07
GC_3_857 b_3 NI_3 NS_857 0 -7.9175932172841623e-06
GC_3_858 b_3 NI_3 NS_858 0 4.8805172798943057e-07
GC_3_859 b_3 NI_3 NS_859 0 3.0157393054437787e-06
GC_3_860 b_3 NI_3 NS_860 0 2.8670353497504996e-06
GC_3_861 b_3 NI_3 NS_861 0 1.2342978936950965e-06
GC_3_862 b_3 NI_3 NS_862 0 -3.9109824204664124e-06
GC_3_863 b_3 NI_3 NS_863 0 -4.8692441102399873e-06
GC_3_864 b_3 NI_3 NS_864 0 -3.9053549780454923e-06
GC_3_865 b_3 NI_3 NS_865 0 3.7776222790710724e-05
GC_3_866 b_3 NI_3 NS_866 0 1.2388280370055701e-12
GC_3_867 b_3 NI_3 NS_867 0 -8.1190354709640468e-12
GC_3_868 b_3 NI_3 NS_868 0 3.0025196652102926e-09
GC_3_869 b_3 NI_3 NS_869 0 3.6863547882124271e-07
GC_3_870 b_3 NI_3 NS_870 0 9.8381726677865538e-08
GC_3_871 b_3 NI_3 NS_871 0 6.5833304502979685e-07
GC_3_872 b_3 NI_3 NS_872 0 3.5826080842055159e-07
GC_3_873 b_3 NI_3 NS_873 0 1.2346308091382786e-06
GC_3_874 b_3 NI_3 NS_874 0 -8.6742346445105313e-07
GC_3_875 b_3 NI_3 NS_875 0 7.8269096416576094e-07
GC_3_876 b_3 NI_3 NS_876 0 -5.3019532045051225e-07
GC_3_877 b_3 NI_3 NS_877 0 8.2387689112440912e-07
GC_3_878 b_3 NI_3 NS_878 0 -2.1815866444211061e-06
GC_3_879 b_3 NI_3 NS_879 0 6.7226784670630556e-07
GC_3_880 b_3 NI_3 NS_880 0 -8.4320817793078804e-07
GC_3_881 b_3 NI_3 NS_881 0 -1.1291288293265790e-06
GC_3_882 b_3 NI_3 NS_882 0 -1.5078760062049339e-06
GC_3_883 b_3 NI_3 NS_883 0 -4.8952415384633402e-07
GC_3_884 b_3 NI_3 NS_884 0 -2.1009697921562839e-06
GC_3_885 b_3 NI_3 NS_885 0 -1.7840493830481467e-06
GC_3_886 b_3 NI_3 NS_886 0 -6.5665285373097617e-07
GC_3_887 b_3 NI_3 NS_887 0 -5.8884953617470710e-07
GC_3_888 b_3 NI_3 NS_888 0 -1.1663418110810802e-06
GC_3_889 b_3 NI_3 NS_889 0 -2.5817961377111298e-06
GC_3_890 b_3 NI_3 NS_890 0 -7.0824187744159758e-07
GC_3_891 b_3 NI_3 NS_891 0 -7.1488745881563720e-07
GC_3_892 b_3 NI_3 NS_892 0 -6.2488999257849105e-07
GC_3_893 b_3 NI_3 NS_893 0 -3.5724825167704720e-06
GC_3_894 b_3 NI_3 NS_894 0 -4.6955722117234718e-07
GC_3_895 b_3 NI_3 NS_895 0 2.3206426217299902e-07
GC_3_896 b_3 NI_3 NS_896 0 -2.1172238407580988e-07
GC_3_897 b_3 NI_3 NS_897 0 -9.1741046374630796e-07
GC_3_898 b_3 NI_3 NS_898 0 -9.0467139706927681e-07
GC_3_899 b_3 NI_3 NS_899 0 -1.9019403968467026e-06
GC_3_900 b_3 NI_3 NS_900 0 1.9080868144942685e-07
GC_3_901 b_3 NI_3 NS_901 0 -1.1727181468160984e-06
GC_3_902 b_3 NI_3 NS_902 0 -4.8227513482540420e-07
GC_3_903 b_3 NI_3 NS_903 0 -1.3189682515202162e-06
GC_3_904 b_3 NI_3 NS_904 0 9.6812054033274870e-07
GC_3_905 b_3 NI_3 NS_905 0 -7.9967177663019193e-07
GC_3_906 b_3 NI_3 NS_906 0 -4.7982923320930618e-07
GC_3_907 b_3 NI_3 NS_907 0 -3.1176527339319567e-06
GC_3_908 b_3 NI_3 NS_908 0 3.9717198822221583e-07
GC_3_909 b_3 NI_3 NS_909 0 -6.0260904189941901e-07
GC_3_910 b_3 NI_3 NS_910 0 1.6123368550211962e-07
GC_3_911 b_3 NI_3 NS_911 0 -6.6727495681390236e-07
GC_3_912 b_3 NI_3 NS_912 0 -1.5680990842856341e-07
GC_3_913 b_3 NI_3 NS_913 0 -1.3447840090612345e-06
GC_3_914 b_3 NI_3 NS_914 0 -7.5287365575698812e-08
GC_3_915 b_3 NI_3 NS_915 0 -3.0786966619551189e-06
GC_3_916 b_3 NI_3 NS_916 0 2.3443908374620578e-06
GC_3_917 b_3 NI_3 NS_917 0 -7.5437662909605286e-07
GC_3_918 b_3 NI_3 NS_918 0 3.5807607488619968e-07
GC_3_919 b_3 NI_3 NS_919 0 -7.9998423574099369e-07
GC_3_920 b_3 NI_3 NS_920 0 1.0728522241788252e-06
GC_3_921 b_3 NI_3 NS_921 0 -1.2382061479513159e-06
GC_3_922 b_3 NI_3 NS_922 0 1.6928415056705649e-07
GC_3_923 b_3 NI_3 NS_923 0 -1.0794847344650845e-06
GC_3_924 b_3 NI_3 NS_924 0 3.5772854438353349e-06
GC_3_925 b_3 NI_3 NS_925 0 -6.8449389517398655e-07
GC_3_926 b_3 NI_3 NS_926 0 4.6095713084164014e-07
GC_3_927 b_3 NI_3 NS_927 0 1.7789024250573081e-07
GC_3_928 b_3 NI_3 NS_928 0 1.4971619466248406e-06
GC_3_929 b_3 NI_3 NS_929 0 -1.1956477713831067e-06
GC_3_930 b_3 NI_3 NS_930 0 3.1705883244986402e-07
GC_3_931 b_3 NI_3 NS_931 0 9.5835726607784762e-07
GC_3_932 b_3 NI_3 NS_932 0 3.0172743890091853e-06
GC_3_933 b_3 NI_3 NS_933 0 -5.5639024543631065e-07
GC_3_934 b_3 NI_3 NS_934 0 6.1270807965315119e-07
GC_3_935 b_3 NI_3 NS_935 0 1.0073479982968640e-06
GC_3_936 b_3 NI_3 NS_936 0 8.4907982015368514e-07
GC_3_937 b_3 NI_3 NS_937 0 -1.1354555495305376e-06
GC_3_938 b_3 NI_3 NS_938 0 5.7364218300795430e-07
GC_3_939 b_3 NI_3 NS_939 0 1.7677940433646317e-06
GC_3_940 b_3 NI_3 NS_940 0 1.3974054775249589e-06
GC_3_941 b_3 NI_3 NS_941 0 -1.4090127388564067e-07
GC_3_942 b_3 NI_3 NS_942 0 6.5188720854770371e-07
GC_3_943 b_3 NI_3 NS_943 0 6.9857260745744239e-07
GC_3_944 b_3 NI_3 NS_944 0 -1.8049690655976513e-08
GC_3_945 b_3 NI_3 NS_945 0 2.1846611416864390e-11
GC_3_946 b_3 NI_3 NS_946 0 1.4146787456525498e-11
GC_3_947 b_3 NI_3 NS_947 0 -5.3444760789157378e-07
GC_3_948 b_3 NI_3 NS_948 0 6.6480172208968075e-07
GC_3_949 b_3 NI_3 NS_949 0 -1.6743782653948774e-08
GC_3_950 b_3 NI_3 NS_950 0 3.0212233598687809e-07
GC_3_951 b_3 NI_3 NS_951 0 2.1121849120581602e-07
GC_3_952 b_3 NI_3 NS_952 0 1.5832456301732411e-07
GC_3_953 b_3 NI_3 NS_953 0 -1.8419257652695752e-07
GC_3_954 b_3 NI_3 NS_954 0 5.6372796205443902e-07
GC_3_955 b_3 NI_3 NS_955 0 8.6157895329540425e-07
GC_3_956 b_3 NI_3 NS_956 0 4.0476723482266600e-07
GC_3_957 b_3 NI_3 NS_957 0 7.9125353242157232e-10
GC_3_958 b_3 NI_3 NS_958 0 5.1026245196820690e-10
GC_3_959 b_3 NI_3 NS_959 0 1.2590914088367804e-06
GC_3_960 b_3 NI_3 NS_960 0 1.3277196209865256e-07
GC_3_961 b_3 NI_3 NS_961 0 -1.4104096100947847e-07
GC_3_962 b_3 NI_3 NS_962 0 8.3427622792184973e-07
GC_3_963 b_3 NI_3 NS_963 0 8.2109873274970467e-08
GC_3_964 b_3 NI_3 NS_964 0 4.1437007751141209e-08
GC_3_965 b_3 NI_3 NS_965 0 3.4449300199387227e-07
GC_3_966 b_3 NI_3 NS_966 0 3.3673157679931018e-07
GC_3_967 b_3 NI_3 NS_967 0 3.0905491444128004e-07
GC_3_968 b_3 NI_3 NS_968 0 4.0929893610800702e-07
GC_3_969 b_3 NI_3 NS_969 0 6.5355092528818810e-08
GC_3_970 b_3 NI_3 NS_970 0 5.9257322080320180e-08
GC_3_971 b_3 NI_3 NS_971 0 7.1106668021220484e-07
GC_3_972 b_3 NI_3 NS_972 0 8.9929617045272205e-07
GC_3_973 b_3 NI_3 NS_973 0 -7.7897460602936231e-06
GC_3_974 b_3 NI_3 NS_974 0 -1.0504404246097737e-11
GC_3_975 b_3 NI_3 NS_975 0 7.2834329729233129e-11
GC_3_976 b_3 NI_3 NS_976 0 -4.8050176450523578e-09
GC_3_977 b_3 NI_3 NS_977 0 -9.4013963263522155e-07
GC_3_978 b_3 NI_3 NS_978 0 -7.1654544445758566e-07
GC_3_979 b_3 NI_3 NS_979 0 6.8854927603549055e-07
GC_3_980 b_3 NI_3 NS_980 0 1.1986218366004547e-06
GC_3_981 b_3 NI_3 NS_981 0 -6.6100523350219126e-07
GC_3_982 b_3 NI_3 NS_982 0 2.7641655265257155e-06
GC_3_983 b_3 NI_3 NS_983 0 -1.7497783360340520e-07
GC_3_984 b_3 NI_3 NS_984 0 -8.3646173559544305e-07
GC_3_985 b_3 NI_3 NS_985 0 3.2529131648917475e-06
GC_3_986 b_3 NI_3 NS_986 0 -1.7247887960412427e-06
GC_3_987 b_3 NI_3 NS_987 0 -2.9874485528217751e-07
GC_3_988 b_3 NI_3 NS_988 0 1.3039975296795281e-06
GC_3_989 b_3 NI_3 NS_989 0 1.3767976956268477e-06
GC_3_990 b_3 NI_3 NS_990 0 1.3767912930843363e-06
GC_3_991 b_3 NI_3 NS_991 0 2.3876662560583894e-06
GC_3_992 b_3 NI_3 NS_992 0 -3.3964994200775705e-06
GC_3_993 b_3 NI_3 NS_993 0 -2.0837789902873759e-06
GC_3_994 b_3 NI_3 NS_994 0 -6.2972652196937665e-06
GC_3_995 b_3 NI_3 NS_995 0 -1.0479874754594366e-07
GC_3_996 b_3 NI_3 NS_996 0 5.0287943102723625e-07
GC_3_997 b_3 NI_3 NS_997 0 -1.2562660211608749e-05
GC_3_998 b_3 NI_3 NS_998 0 3.3121634140489698e-06
GC_3_999 b_3 NI_3 NS_999 0 -1.5084748753430245e-07
GC_3_1000 b_3 NI_3 NS_1000 0 -6.4681545986168911e-07
GC_3_1001 b_3 NI_3 NS_1001 0 3.1495019498380424e-06
GC_3_1002 b_3 NI_3 NS_1002 0 1.5214615784353130e-05
GC_3_1003 b_3 NI_3 NS_1003 0 1.0368157573845136e-06
GC_3_1004 b_3 NI_3 NS_1004 0 -1.0548128391773940e-06
GC_3_1005 b_3 NI_3 NS_1005 0 1.1266686940483934e-06
GC_3_1006 b_3 NI_3 NS_1006 0 -3.1888276530659319e-07
GC_3_1007 b_3 NI_3 NS_1007 0 6.6856521282576532e-06
GC_3_1008 b_3 NI_3 NS_1008 0 -3.1044316446760741e-06
GC_3_1009 b_3 NI_3 NS_1009 0 3.3082679062150847e-07
GC_3_1010 b_3 NI_3 NS_1010 0 3.9509228777037399e-07
GC_3_1011 b_3 NI_3 NS_1011 0 -2.9432347110329884e-06
GC_3_1012 b_3 NI_3 NS_1012 0 8.3276129263639849e-07
GC_3_1013 b_3 NI_3 NS_1013 0 1.7555365923548180e-07
GC_3_1014 b_3 NI_3 NS_1014 0 -8.8267390770487047e-07
GC_3_1015 b_3 NI_3 NS_1015 0 6.7910523980651372e-06
GC_3_1016 b_3 NI_3 NS_1016 0 3.5401113980618714e-06
GC_3_1017 b_3 NI_3 NS_1017 0 3.3550365840873807e-07
GC_3_1018 b_3 NI_3 NS_1018 0 8.9056883457498513e-09
GC_3_1019 b_3 NI_3 NS_1019 0 2.4547458644948968e-07
GC_3_1020 b_3 NI_3 NS_1020 0 -6.0588414723250036e-07
GC_3_1021 b_3 NI_3 NS_1021 0 4.0057090471419302e-07
GC_3_1022 b_3 NI_3 NS_1022 0 -1.3949646898614506e-06
GC_3_1023 b_3 NI_3 NS_1023 0 6.0103699139181961e-06
GC_3_1024 b_3 NI_3 NS_1024 0 -2.3488802021605365e-06
GC_3_1025 b_3 NI_3 NS_1025 0 2.3332715056637053e-08
GC_3_1026 b_3 NI_3 NS_1026 0 -2.5588152599198745e-07
GC_3_1027 b_3 NI_3 NS_1027 0 -9.3826675512032715e-07
GC_3_1028 b_3 NI_3 NS_1028 0 -1.1597830283820277e-06
GC_3_1029 b_3 NI_3 NS_1029 0 3.0914660580504447e-07
GC_3_1030 b_3 NI_3 NS_1030 0 -1.3347744735062569e-06
GC_3_1031 b_3 NI_3 NS_1031 0 3.0251058319142003e-06
GC_3_1032 b_3 NI_3 NS_1032 0 -4.1459941916636855e-06
GC_3_1033 b_3 NI_3 NS_1033 0 -1.7543349986346702e-07
GC_3_1034 b_3 NI_3 NS_1034 0 -3.4365969410298041e-07
GC_3_1035 b_3 NI_3 NS_1035 0 -1.9736550400930781e-06
GC_3_1036 b_3 NI_3 NS_1036 0 -6.6869864132916716e-07
GC_3_1037 b_3 NI_3 NS_1037 0 2.0799747702129498e-07
GC_3_1038 b_3 NI_3 NS_1038 0 -1.4276250279220612e-06
GC_3_1039 b_3 NI_3 NS_1039 0 9.0918056111690689e-08
GC_3_1040 b_3 NI_3 NS_1040 0 -3.5637761455539293e-06
GC_3_1041 b_3 NI_3 NS_1041 0 -4.5635407912012426e-07
GC_3_1042 b_3 NI_3 NS_1042 0 -3.7736056133564476e-07
GC_3_1043 b_3 NI_3 NS_1043 0 -2.1515974290425873e-06
GC_3_1044 b_3 NI_3 NS_1044 0 5.3436192736069731e-07
GC_3_1045 b_3 NI_3 NS_1045 0 -6.9689773924364562e-08
GC_3_1046 b_3 NI_3 NS_1046 0 -1.6164299370035435e-06
GC_3_1047 b_3 NI_3 NS_1047 0 -1.2654804703885673e-06
GC_3_1048 b_3 NI_3 NS_1048 0 -1.4050915596212297e-06
GC_3_1049 b_3 NI_3 NS_1049 0 -8.0777193497780135e-07
GC_3_1050 b_3 NI_3 NS_1050 0 9.5484822515542580e-08
GC_3_1051 b_3 NI_3 NS_1051 0 -9.4861252523542362e-07
GC_3_1052 b_3 NI_3 NS_1052 0 1.0889515400129353e-06
GC_3_1053 b_3 NI_3 NS_1053 0 -1.7801506037942984e-11
GC_3_1054 b_3 NI_3 NS_1054 0 1.0630295236820815e-11
GC_3_1055 b_3 NI_3 NS_1055 0 -5.7532605447189263e-07
GC_3_1056 b_3 NI_3 NS_1056 0 -1.1642954789164241e-06
GC_3_1057 b_3 NI_3 NS_1057 0 -3.7975234194194798e-07
GC_3_1058 b_3 NI_3 NS_1058 0 2.2310889389967782e-07
GC_3_1059 b_3 NI_3 NS_1059 0 -5.0948369190502705e-07
GC_3_1060 b_3 NI_3 NS_1060 0 3.9880801697257150e-07
GC_3_1061 b_3 NI_3 NS_1061 0 -1.9110900316247429e-07
GC_3_1062 b_3 NI_3 NS_1062 0 -1.0234485524849850e-06
GC_3_1063 b_3 NI_3 NS_1063 0 -4.4605829437820637e-07
GC_3_1064 b_3 NI_3 NS_1064 0 -2.0182507942765925e-07
GC_3_1065 b_3 NI_3 NS_1065 0 -9.1683270903032988e-10
GC_3_1066 b_3 NI_3 NS_1066 0 1.5474504414939049e-10
GC_3_1067 b_3 NI_3 NS_1067 0 -2.2824735863381844e-07
GC_3_1068 b_3 NI_3 NS_1068 0 -1.9835481794455212e-07
GC_3_1069 b_3 NI_3 NS_1069 0 -1.7951620406705508e-07
GC_3_1070 b_3 NI_3 NS_1070 0 -3.4653915566061284e-07
GC_3_1071 b_3 NI_3 NS_1071 0 -3.9555957925644710e-07
GC_3_1072 b_3 NI_3 NS_1072 0 -1.3726968473554629e-07
GC_3_1073 b_3 NI_3 NS_1073 0 -9.9082674201513068e-07
GC_3_1074 b_3 NI_3 NS_1074 0 5.0308194601258428e-08
GC_3_1075 b_3 NI_3 NS_1075 0 -5.8387941439370568e-07
GC_3_1076 b_3 NI_3 NS_1076 0 4.7571089200241364e-07
GC_3_1077 b_3 NI_3 NS_1077 0 -1.3188422079152970e-08
GC_3_1078 b_3 NI_3 NS_1078 0 4.1222560361601918e-07
GC_3_1079 b_3 NI_3 NS_1079 0 -8.6504628654947213e-07
GC_3_1080 b_3 NI_3 NS_1080 0 -9.7526961363991539e-07
GC_3_1081 b_3 NI_3 NS_1081 0 8.6499760697279228e-06
GC_3_1082 b_3 NI_3 NS_1082 0 3.7611075939792824e-12
GC_3_1083 b_3 NI_3 NS_1083 0 -7.8508192241374158e-11
GC_3_1084 b_3 NI_3 NS_1084 0 2.5460399000505486e-09
GC_3_1085 b_3 NI_3 NS_1085 0 1.6514174522185145e-08
GC_3_1086 b_3 NI_3 NS_1086 0 -8.5494770527429905e-08
GC_3_1087 b_3 NI_3 NS_1087 0 -2.4857697333612501e-07
GC_3_1088 b_3 NI_3 NS_1088 0 2.6957994950094591e-07
GC_3_1089 b_3 NI_3 NS_1089 0 7.4441982656586475e-07
GC_3_1090 b_3 NI_3 NS_1090 0 -2.8507177006602925e-07
GC_3_1091 b_3 NI_3 NS_1091 0 -9.6886905768051224e-07
GC_3_1092 b_3 NI_3 NS_1092 0 -2.4196041195101523e-07
GC_3_1093 b_3 NI_3 NS_1093 0 1.0238384473795697e-06
GC_3_1094 b_3 NI_3 NS_1094 0 4.0092170339491546e-07
GC_3_1095 b_3 NI_3 NS_1095 0 -1.2005343089181322e-07
GC_3_1096 b_3 NI_3 NS_1096 0 -2.7540994466566224e-07
GC_3_1097 b_3 NI_3 NS_1097 0 1.0875932140459285e-07
GC_3_1098 b_3 NI_3 NS_1098 0 -5.1234262679653527e-07
GC_3_1099 b_3 NI_3 NS_1099 0 -2.0908861925245252e-06
GC_3_1100 b_3 NI_3 NS_1100 0 8.5580367426962479e-07
GC_3_1101 b_3 NI_3 NS_1101 0 2.4337654523400269e-06
GC_3_1102 b_3 NI_3 NS_1102 0 -6.0045388771755636e-07
GC_3_1103 b_3 NI_3 NS_1103 0 -6.6288729138483703e-07
GC_3_1104 b_3 NI_3 NS_1104 0 -1.4012567872296981e-06
GC_3_1105 b_3 NI_3 NS_1105 0 4.2235826892230442e-07
GC_3_1106 b_3 NI_3 NS_1106 0 1.8489190228542526e-06
GC_3_1107 b_3 NI_3 NS_1107 0 -2.9760464947141977e-08
GC_3_1108 b_3 NI_3 NS_1108 0 -1.3254973002998511e-06
GC_3_1109 b_3 NI_3 NS_1109 0 -6.4020208284293644e-07
GC_3_1110 b_3 NI_3 NS_1110 0 2.5950866923641724e-06
GC_3_1111 b_3 NI_3 NS_1111 0 4.5705235832528088e-07
GC_3_1112 b_3 NI_3 NS_1112 0 -2.2460566847200263e-06
GC_3_1113 b_3 NI_3 NS_1113 0 -8.0117683248625152e-07
GC_3_1114 b_3 NI_3 NS_1114 0 -9.3397538516266902e-07
GC_3_1115 b_3 NI_3 NS_1115 0 3.5739864232911778e-07
GC_3_1116 b_3 NI_3 NS_1116 0 9.1444694454686937e-07
GC_3_1117 b_3 NI_3 NS_1117 0 -5.5834208011740468e-07
GC_3_1118 b_3 NI_3 NS_1118 0 -7.2678594532431835e-07
GC_3_1119 b_3 NI_3 NS_1119 0 4.7648087055231108e-07
GC_3_1120 b_3 NI_3 NS_1120 0 7.4219333533512872e-07
GC_3_1121 b_3 NI_3 NS_1121 0 -1.7459567228683978e-07
GC_3_1122 b_3 NI_3 NS_1122 0 -8.7943212307325200e-07
GC_3_1123 b_3 NI_3 NS_1123 0 -3.4060715996318504e-07
GC_3_1124 b_3 NI_3 NS_1124 0 1.1609613803212248e-06
GC_3_1125 b_3 NI_3 NS_1125 0 2.5385913164736568e-07
GC_3_1126 b_3 NI_3 NS_1126 0 -8.4525455204049069e-07
GC_3_1127 b_3 NI_3 NS_1127 0 -6.5148072035354393e-08
GC_3_1128 b_3 NI_3 NS_1128 0 6.7372794732604432e-08
GC_3_1129 b_3 NI_3 NS_1129 0 -2.6093310149635805e-07
GC_3_1130 b_3 NI_3 NS_1130 0 -5.5061992592262972e-07
GC_3_1131 b_3 NI_3 NS_1131 0 1.8491349427419658e-07
GC_3_1132 b_3 NI_3 NS_1132 0 7.1949277637286105e-07
GC_3_1133 b_3 NI_3 NS_1133 0 -8.1165289169303187e-08
GC_3_1134 b_3 NI_3 NS_1134 0 -6.3616031756413865e-07
GC_3_1135 b_3 NI_3 NS_1135 0 1.0184234117242053e-07
GC_3_1136 b_3 NI_3 NS_1136 0 1.0497370014197878e-07
GC_3_1137 b_3 NI_3 NS_1137 0 -2.9217446022889237e-07
GC_3_1138 b_3 NI_3 NS_1138 0 -5.9433384667843912e-07
GC_3_1139 b_3 NI_3 NS_1139 0 1.6155144070273117e-07
GC_3_1140 b_3 NI_3 NS_1140 0 2.3346996145255165e-07
GC_3_1141 b_3 NI_3 NS_1141 0 -2.5774766101751143e-07
GC_3_1142 b_3 NI_3 NS_1142 0 -5.0844982427349114e-07
GC_3_1143 b_3 NI_3 NS_1143 0 4.9022073733313104e-08
GC_3_1144 b_3 NI_3 NS_1144 0 -4.9060768080724659e-08
GC_3_1145 b_3 NI_3 NS_1145 0 -3.6949396826847419e-07
GC_3_1146 b_3 NI_3 NS_1146 0 -5.5863800674157284e-07
GC_3_1147 b_3 NI_3 NS_1147 0 -2.3397484042252079e-07
GC_3_1148 b_3 NI_3 NS_1148 0 2.3113987072223356e-08
GC_3_1149 b_3 NI_3 NS_1149 0 -4.3492502539818341e-07
GC_3_1150 b_3 NI_3 NS_1150 0 -3.4101525093031211e-07
GC_3_1151 b_3 NI_3 NS_1151 0 -1.2370426653621801e-07
GC_3_1152 b_3 NI_3 NS_1152 0 1.7270977904652627e-08
GC_3_1153 b_3 NI_3 NS_1153 0 -5.6511183252999882e-07
GC_3_1154 b_3 NI_3 NS_1154 0 -4.3986483555540997e-07
GC_3_1155 b_3 NI_3 NS_1155 0 -3.1751839557889779e-07
GC_3_1156 b_3 NI_3 NS_1156 0 3.1817909095396322e-07
GC_3_1157 b_3 NI_3 NS_1157 0 -5.0074805465218262e-07
GC_3_1158 b_3 NI_3 NS_1158 0 3.7787320355561914e-08
GC_3_1159 b_3 NI_3 NS_1159 0 -9.9072878410843799e-09
GC_3_1160 b_3 NI_3 NS_1160 0 6.2428894188219412e-08
GC_3_1161 b_3 NI_3 NS_1161 0 -3.2503510851902601e-12
GC_3_1162 b_3 NI_3 NS_1162 0 3.2070864704850453e-12
GC_3_1163 b_3 NI_3 NS_1163 0 -5.7741465318644939e-07
GC_3_1164 b_3 NI_3 NS_1164 0 4.6881106833645316e-08
GC_3_1165 b_3 NI_3 NS_1165 0 -2.9017231532812806e-07
GC_3_1166 b_3 NI_3 NS_1166 0 1.1797445271751377e-07
GC_3_1167 b_3 NI_3 NS_1167 0 -5.7762666152895780e-09
GC_3_1168 b_3 NI_3 NS_1168 0 -6.8374774520683980e-08
GC_3_1169 b_3 NI_3 NS_1169 0 -6.6136365822173070e-07
GC_3_1170 b_3 NI_3 NS_1170 0 1.4039123820852317e-07
GC_3_1171 b_3 NI_3 NS_1171 0 2.9868708380503248e-08
GC_3_1172 b_3 NI_3 NS_1172 0 1.2538985853118363e-07
GC_3_1173 b_3 NI_3 NS_1173 0 -6.1347532197929273e-11
GC_3_1174 b_3 NI_3 NS_1174 0 1.2844605143310803e-10
GC_3_1175 b_3 NI_3 NS_1175 0 -3.4935699546006341e-08
GC_3_1176 b_3 NI_3 NS_1176 0 1.9709080761443364e-07
GC_3_1177 b_3 NI_3 NS_1177 0 -3.6685714270277736e-07
GC_3_1178 b_3 NI_3 NS_1178 0 -4.4445749137693096e-08
GC_3_1179 b_3 NI_3 NS_1179 0 -1.8614734309373757e-07
GC_3_1180 b_3 NI_3 NS_1180 0 -2.6651584315545898e-09
GC_3_1181 b_3 NI_3 NS_1181 0 1.9333586809877323e-07
GC_3_1182 b_3 NI_3 NS_1182 0 8.2525006304740327e-08
GC_3_1183 b_3 NI_3 NS_1183 0 -2.6572625664130416e-07
GC_3_1184 b_3 NI_3 NS_1184 0 3.1365990297398866e-07
GC_3_1185 b_3 NI_3 NS_1185 0 1.2571479188084991e-07
GC_3_1186 b_3 NI_3 NS_1186 0 -1.4398641671776392e-07
GC_3_1187 b_3 NI_3 NS_1187 0 -5.8257020153597384e-08
GC_3_1188 b_3 NI_3 NS_1188 0 2.3778827371725476e-07
GC_3_1189 b_3 NI_3 NS_1189 0 -6.4297412272203272e-05
GC_3_1190 b_3 NI_3 NS_1190 0 3.5514235869631269e-12
GC_3_1191 b_3 NI_3 NS_1191 0 5.0206486791833467e-11
GC_3_1192 b_3 NI_3 NS_1192 0 -1.5827698920948701e-09
GC_3_1193 b_3 NI_3 NS_1193 0 -1.0722828933200687e-06
GC_3_1194 b_3 NI_3 NS_1194 0 -1.0608507475561062e-06
GC_3_1195 b_3 NI_3 NS_1195 0 4.1036076311628142e-07
GC_3_1196 b_3 NI_3 NS_1196 0 3.5893571377090403e-07
GC_3_1197 b_3 NI_3 NS_1197 0 -2.2645833124840754e-06
GC_3_1198 b_3 NI_3 NS_1198 0 2.1075513920262079e-06
GC_3_1199 b_3 NI_3 NS_1199 0 -2.5340137861648331e-06
GC_3_1200 b_3 NI_3 NS_1200 0 -1.2433708025262304e-06
GC_3_1201 b_3 NI_3 NS_1201 0 1.3995740030758579e-06
GC_3_1202 b_3 NI_3 NS_1202 0 1.0022088387151152e-06
GC_3_1203 b_3 NI_3 NS_1203 0 -1.1248412643989546e-06
GC_3_1204 b_3 NI_3 NS_1204 0 1.3421231783428241e-06
GC_3_1205 b_3 NI_3 NS_1205 0 7.2528849444911206e-07
GC_3_1206 b_3 NI_3 NS_1206 0 3.0434862611068877e-06
GC_3_1207 b_3 NI_3 NS_1207 0 -2.8542769913363534e-06
GC_3_1208 b_3 NI_3 NS_1208 0 4.6950197875806584e-07
GC_3_1209 b_3 NI_3 NS_1209 0 3.6961210083111703e-06
GC_3_1210 b_3 NI_3 NS_1210 0 -2.0128609171382267e-06
GC_3_1211 b_3 NI_3 NS_1211 0 -1.9025399234708104e-07
GC_3_1212 b_3 NI_3 NS_1212 0 2.5688277011651937e-06
GC_3_1213 b_3 NI_3 NS_1213 0 -4.0608190676609042e-06
GC_3_1214 b_3 NI_3 NS_1214 0 4.8420445497625661e-06
GC_3_1215 b_3 NI_3 NS_1215 0 6.4548938524185092e-07
GC_3_1216 b_3 NI_3 NS_1216 0 -1.5900718915782203e-06
GC_3_1217 b_3 NI_3 NS_1217 0 4.6200332807073634e-06
GC_3_1218 b_3 NI_3 NS_1218 0 9.9425470176513199e-06
GC_3_1219 b_3 NI_3 NS_1219 0 -1.1566708036379689e-07
GC_3_1220 b_3 NI_3 NS_1220 0 5.2797010234067277e-07
GC_3_1221 b_3 NI_3 NS_1221 0 -6.9202510556828457e-09
GC_3_1222 b_3 NI_3 NS_1222 0 -7.8936878282899767e-07
GC_3_1223 b_3 NI_3 NS_1223 0 5.3542038007278873e-06
GC_3_1224 b_3 NI_3 NS_1224 0 4.9601575613463205e-07
GC_3_1225 b_3 NI_3 NS_1225 0 8.4752708507068303e-07
GC_3_1226 b_3 NI_3 NS_1226 0 1.9215332741914785e-06
GC_3_1227 b_3 NI_3 NS_1227 0 3.1631761985099379e-08
GC_3_1228 b_3 NI_3 NS_1228 0 1.1340872726601043e-06
GC_3_1229 b_3 NI_3 NS_1229 0 5.8569848670761818e-07
GC_3_1230 b_3 NI_3 NS_1230 0 -1.1142344034648720e-06
GC_3_1231 b_3 NI_3 NS_1231 0 5.8308848426238781e-06
GC_3_1232 b_3 NI_3 NS_1232 0 4.0738777187664284e-06
GC_3_1233 b_3 NI_3 NS_1233 0 6.0565117509307706e-07
GC_3_1234 b_3 NI_3 NS_1234 0 8.6240374159637696e-07
GC_3_1235 b_3 NI_3 NS_1235 0 1.9671298752514494e-07
GC_3_1236 b_3 NI_3 NS_1236 0 2.4104642474440342e-07
GC_3_1237 b_3 NI_3 NS_1237 0 8.4506760537914294e-07
GC_3_1238 b_3 NI_3 NS_1238 0 -6.7479264361511128e-07
GC_3_1239 b_3 NI_3 NS_1239 0 6.6692115150788596e-06
GC_3_1240 b_3 NI_3 NS_1240 0 7.5282429197950534e-07
GC_3_1241 b_3 NI_3 NS_1241 0 7.7512228865918122e-07
GC_3_1242 b_3 NI_3 NS_1242 0 7.5176083678239308e-07
GC_3_1243 b_3 NI_3 NS_1243 0 6.6485040734087620e-07
GC_3_1244 b_3 NI_3 NS_1244 0 -6.6043563420037758e-08
GC_3_1245 b_3 NI_3 NS_1245 0 8.7117258289697854e-07
GC_3_1246 b_3 NI_3 NS_1246 0 -6.4327579308889517e-07
GC_3_1247 b_3 NI_3 NS_1247 0 5.7782949123236246e-06
GC_3_1248 b_3 NI_3 NS_1248 0 -1.5930752002140226e-06
GC_3_1249 b_3 NI_3 NS_1249 0 8.2495328550066645e-07
GC_3_1250 b_3 NI_3 NS_1250 0 5.6932086635125915e-07
GC_3_1251 b_3 NI_3 NS_1251 0 6.2573263056524826e-07
GC_3_1252 b_3 NI_3 NS_1252 0 -5.5367383576110764e-07
GC_3_1253 b_3 NI_3 NS_1253 0 9.3726572126018233e-07
GC_3_1254 b_3 NI_3 NS_1254 0 -4.4873224448415382e-07
GC_3_1255 b_3 NI_3 NS_1255 0 3.9054793162363959e-06
GC_3_1256 b_3 NI_3 NS_1256 0 -2.9926331407550171e-06
GC_3_1257 b_3 NI_3 NS_1257 0 8.9723679786252013e-07
GC_3_1258 b_3 NI_3 NS_1258 0 3.2914489375119446e-07
GC_3_1259 b_3 NI_3 NS_1259 0 2.1534206229511193e-07
GC_3_1260 b_3 NI_3 NS_1260 0 -7.9633593698850240e-07
GC_3_1261 b_3 NI_3 NS_1261 0 1.1591902992846267e-06
GC_3_1262 b_3 NI_3 NS_1262 0 -3.2770578886019402e-07
GC_3_1263 b_3 NI_3 NS_1263 0 1.6782711498448465e-06
GC_3_1264 b_3 NI_3 NS_1264 0 -3.0911768582879330e-06
GC_3_1265 b_3 NI_3 NS_1265 0 7.9264307790817912e-07
GC_3_1266 b_3 NI_3 NS_1266 0 -1.0570197213793237e-07
GC_3_1267 b_3 NI_3 NS_1267 0 -1.9831575567156398e-07
GC_3_1268 b_3 NI_3 NS_1268 0 -4.0881219681125173e-07
GC_3_1269 b_3 NI_3 NS_1269 0 8.5890829174839454e-12
GC_3_1270 b_3 NI_3 NS_1270 0 -1.5739957282276767e-11
GC_3_1271 b_3 NI_3 NS_1271 0 8.3767062242451204e-07
GC_3_1272 b_3 NI_3 NS_1272 0 -5.9585114205071387e-07
GC_3_1273 b_3 NI_3 NS_1273 0 4.9537093177233497e-07
GC_3_1274 b_3 NI_3 NS_1274 0 -3.5565908055820252e-08
GC_3_1275 b_3 NI_3 NS_1275 0 1.6374041304240207e-08
GC_3_1276 b_3 NI_3 NS_1276 0 -8.9212636100079678e-08
GC_3_1277 b_3 NI_3 NS_1277 0 5.2071353167670246e-07
GC_3_1278 b_3 NI_3 NS_1278 0 -1.9287637196135125e-08
GC_3_1279 b_3 NI_3 NS_1279 0 7.0590608121788305e-07
GC_3_1280 b_3 NI_3 NS_1280 0 -1.5618062318983539e-06
GC_3_1281 b_3 NI_3 NS_1281 0 4.0958055597296431e-10
GC_3_1282 b_3 NI_3 NS_1282 0 -5.8094691120126357e-10
GC_3_1283 b_3 NI_3 NS_1283 0 1.0094261923604203e-06
GC_3_1284 b_3 NI_3 NS_1284 0 -2.7418423606128643e-07
GC_3_1285 b_3 NI_3 NS_1285 0 3.5391568538188004e-07
GC_3_1286 b_3 NI_3 NS_1286 0 -1.7487869350401040e-07
GC_3_1287 b_3 NI_3 NS_1287 0 2.5449981903220582e-07
GC_3_1288 b_3 NI_3 NS_1288 0 2.6674265458372448e-08
GC_3_1289 b_3 NI_3 NS_1289 0 1.0861096271302963e-06
GC_3_1290 b_3 NI_3 NS_1290 0 -1.1751132122605891e-06
GC_3_1291 b_3 NI_3 NS_1291 0 6.5444226169251881e-07
GC_3_1292 b_3 NI_3 NS_1292 0 -3.3449157854871962e-07
GC_3_1293 b_3 NI_3 NS_1293 0 -2.1289964648260744e-07
GC_3_1294 b_3 NI_3 NS_1294 0 -9.8626048028037387e-08
GC_3_1295 b_3 NI_3 NS_1295 0 7.5675679485447304e-07
GC_3_1296 b_3 NI_3 NS_1296 0 3.2207287586360221e-07
GD_3_1 b_3 NI_3 NA_1 0 1.0616349053176422e-02
GD_3_2 b_3 NI_3 NA_2 0 -1.1524190478452503e-03
GD_3_3 b_3 NI_3 NA_3 0 -1.0894627888821864e-02
GD_3_4 b_3 NI_3 NA_4 0 -5.0003252503784748e-03
GD_3_5 b_3 NI_3 NA_5 0 2.2219274415387805e-05
GD_3_6 b_3 NI_3 NA_6 0 1.0510730226758834e-04
GD_3_7 b_3 NI_3 NA_7 0 -1.0996159851898246e-06
GD_3_8 b_3 NI_3 NA_8 0 1.6002510073223825e-05
GD_3_9 b_3 NI_3 NA_9 0 -7.3787017813712797e-06
GD_3_10 b_3 NI_3 NA_10 0 2.0978230138391877e-06
GD_3_11 b_3 NI_3 NA_11 0 -1.1882831422966855e-06
GD_3_12 b_3 NI_3 NA_12 0 8.8115119568417009e-06
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 -3.3036299659495202e-03
GC_4_2 b_4 NI_4 NS_2 0 1.8493831333748727e-09
GC_4_3 b_4 NI_4 NS_3 0 5.6032190447337941e-08
GC_4_4 b_4 NI_4 NS_4 0 1.8929692330477028e-06
GC_4_5 b_4 NI_4 NS_5 0 -9.1167689772451752e-05
GC_4_6 b_4 NI_4 NS_6 0 -5.7737977656453684e-05
GC_4_7 b_4 NI_4 NS_7 0 -1.2657733195001227e-03
GC_4_8 b_4 NI_4 NS_8 0 -2.9559391758780817e-04
GC_4_9 b_4 NI_4 NS_9 0 -1.6792135386434644e-03
GC_4_10 b_4 NI_4 NS_10 0 2.6464976074095409e-03
GC_4_11 b_4 NI_4 NS_11 0 5.1121143940030262e-04
GC_4_12 b_4 NI_4 NS_12 0 5.4276088234639433e-03
GC_4_13 b_4 NI_4 NS_13 0 7.1034883281088619e-03
GC_4_14 b_4 NI_4 NS_14 0 6.3629270836289883e-04
GC_4_15 b_4 NI_4 NS_15 0 6.4432995071112399e-04
GC_4_16 b_4 NI_4 NS_16 0 -6.6091924438288756e-04
GC_4_17 b_4 NI_4 NS_17 0 1.0576980463265408e-03
GC_4_18 b_4 NI_4 NS_18 0 1.5711404780115884e-03
GC_4_19 b_4 NI_4 NS_19 0 1.2687514002831107e-02
GC_4_20 b_4 NI_4 NS_20 0 1.3123213057122857e-02
GC_4_21 b_4 NI_4 NS_21 0 8.7187976086676080e-03
GC_4_22 b_4 NI_4 NS_22 0 -2.0392080353350578e-02
GC_4_23 b_4 NI_4 NS_23 0 8.3891005278679300e-03
GC_4_24 b_4 NI_4 NS_24 0 -2.9045256335337236e-03
GC_4_25 b_4 NI_4 NS_25 0 -1.2701288451032579e-02
GC_4_26 b_4 NI_4 NS_26 0 -3.8806698093156539e-02
GC_4_27 b_4 NI_4 NS_27 0 -7.2523388538709909e-03
GC_4_28 b_4 NI_4 NS_28 0 -2.1332751200162136e-03
GC_4_29 b_4 NI_4 NS_29 0 -5.2307197882006391e-02
GC_4_30 b_4 NI_4 NS_30 0 -1.7936176889304968e-03
GC_4_31 b_4 NI_4 NS_31 0 1.4914414747264045e-02
GC_4_32 b_4 NI_4 NS_32 0 8.6735769599791158e-03
GC_4_33 b_4 NI_4 NS_33 0 -5.9233531499012495e-03
GC_4_34 b_4 NI_4 NS_34 0 5.0044969318290998e-03
GC_4_35 b_4 NI_4 NS_35 0 8.3724191777758035e-03
GC_4_36 b_4 NI_4 NS_36 0 1.1688363832600418e-02
GC_4_37 b_4 NI_4 NS_37 0 4.5592641793986838e-03
GC_4_38 b_4 NI_4 NS_38 0 -2.9327403765924500e-03
GC_4_39 b_4 NI_4 NS_39 0 -7.8986719439334430e-03
GC_4_40 b_4 NI_4 NS_40 0 -8.1490658831921709e-03
GC_4_41 b_4 NI_4 NS_41 0 -5.6808134019349418e-03
GC_4_42 b_4 NI_4 NS_42 0 -6.1281061858789758e-04
GC_4_43 b_4 NI_4 NS_43 0 -1.8070850038082717e-02
GC_4_44 b_4 NI_4 NS_44 0 1.3578962120178121e-02
GC_4_45 b_4 NI_4 NS_45 0 4.7069857203916304e-03
GC_4_46 b_4 NI_4 NS_46 0 4.3794388360163285e-03
GC_4_47 b_4 NI_4 NS_47 0 6.5015842441291092e-04
GC_4_48 b_4 NI_4 NS_48 0 -1.0995431105456216e-04
GC_4_49 b_4 NI_4 NS_49 0 -3.7963995323925122e-03
GC_4_50 b_4 NI_4 NS_50 0 8.8498820079000189e-04
GC_4_51 b_4 NI_4 NS_51 0 -1.1178288590647377e-03
GC_4_52 b_4 NI_4 NS_52 0 1.6699686524908212e-02
GC_4_53 b_4 NI_4 NS_53 0 4.4472801150505269e-03
GC_4_54 b_4 NI_4 NS_54 0 7.0796431371151450e-04
GC_4_55 b_4 NI_4 NS_55 0 -5.1995848568804832e-04
GC_4_56 b_4 NI_4 NS_56 0 -2.2477513013483062e-03
GC_4_57 b_4 NI_4 NS_57 0 -4.9864558426922822e-03
GC_4_58 b_4 NI_4 NS_58 0 2.1108873628474536e-03
GC_4_59 b_4 NI_4 NS_59 0 7.3425265677526915e-03
GC_4_60 b_4 NI_4 NS_60 0 1.4345854693753225e-02
GC_4_61 b_4 NI_4 NS_61 0 4.1872274284202255e-03
GC_4_62 b_4 NI_4 NS_62 0 -1.6838585093975735e-03
GC_4_63 b_4 NI_4 NS_63 0 -3.3981251905511904e-03
GC_4_64 b_4 NI_4 NS_64 0 -2.1006235889358240e-03
GC_4_65 b_4 NI_4 NS_65 0 -5.4204257559384806e-03
GC_4_66 b_4 NI_4 NS_66 0 4.3817240576716193e-03
GC_4_67 b_4 NI_4 NS_67 0 1.3196871230933565e-02
GC_4_68 b_4 NI_4 NS_68 0 8.4333073603318834e-03
GC_4_69 b_4 NI_4 NS_69 0 2.8324336032150752e-03
GC_4_70 b_4 NI_4 NS_70 0 -4.1306060240013185e-03
GC_4_71 b_4 NI_4 NS_71 0 -5.3207863284678459e-03
GC_4_72 b_4 NI_4 NS_72 0 1.1381587447445594e-03
GC_4_73 b_4 NI_4 NS_73 0 -4.4310206572533784e-03
GC_4_74 b_4 NI_4 NS_74 0 8.3104309072311762e-03
GC_4_75 b_4 NI_4 NS_75 0 1.4612785651422731e-02
GC_4_76 b_4 NI_4 NS_76 0 -4.6824711949203538e-04
GC_4_77 b_4 NI_4 NS_77 0 -1.1845320565709938e-03
GC_4_78 b_4 NI_4 NS_78 0 -4.5473899410772975e-03
GC_4_79 b_4 NI_4 NS_79 0 -2.2825678225249111e-03
GC_4_80 b_4 NI_4 NS_80 0 4.3832546992168030e-03
GC_4_81 b_4 NI_4 NS_81 0 1.3571252026534121e-10
GC_4_82 b_4 NI_4 NS_82 0 -1.5466654416853168e-09
GC_4_83 b_4 NI_4 NS_83 0 1.4460257346634263e-03
GC_4_84 b_4 NI_4 NS_84 0 8.2165466761966767e-03
GC_4_85 b_4 NI_4 NS_85 0 -8.7895047602657155e-04
GC_4_86 b_4 NI_4 NS_86 0 -2.2072124549669964e-03
GC_4_87 b_4 NI_4 NS_87 0 -1.4679135508807010e-03
GC_4_88 b_4 NI_4 NS_88 0 2.7519861857558908e-03
GC_4_89 b_4 NI_4 NS_89 0 1.7320143417073920e-03
GC_4_90 b_4 NI_4 NS_90 0 7.6059325919460010e-03
GC_4_91 b_4 NI_4 NS_91 0 7.5874084177808788e-03
GC_4_92 b_4 NI_4 NS_92 0 -3.8276823056536346e-03
GC_4_93 b_4 NI_4 NS_93 0 -5.2101075106709342e-08
GC_4_94 b_4 NI_4 NS_94 0 -2.0817222334933978e-08
GC_4_95 b_4 NI_4 NS_95 0 1.1391243237851206e-02
GC_4_96 b_4 NI_4 NS_96 0 4.4700330710704247e-03
GC_4_97 b_4 NI_4 NS_97 0 -8.6185054339452561e-04
GC_4_98 b_4 NI_4 NS_98 0 6.4916224675031975e-03
GC_4_99 b_4 NI_4 NS_99 0 3.6263738293742221e-03
GC_4_100 b_4 NI_4 NS_100 0 4.0710468898222672e-04
GC_4_101 b_4 NI_4 NS_101 0 6.0525109496231966e-03
GC_4_102 b_4 NI_4 NS_102 0 -4.6635402172840448e-03
GC_4_103 b_4 NI_4 NS_103 0 -3.3929752234436081e-03
GC_4_104 b_4 NI_4 NS_104 0 -1.3533960292098190e-03
GC_4_105 b_4 NI_4 NS_105 0 1.1237962504259089e-04
GC_4_106 b_4 NI_4 NS_106 0 4.4958002654125083e-03
GC_4_107 b_4 NI_4 NS_107 0 7.2795568413537189e-03
GC_4_108 b_4 NI_4 NS_108 0 5.5305047720051372e-03
GC_4_109 b_4 NI_4 NS_109 0 1.1804733938835439e-03
GC_4_110 b_4 NI_4 NS_110 0 -3.5559930493000567e-09
GC_4_111 b_4 NI_4 NS_111 0 -4.8002576630688173e-08
GC_4_112 b_4 NI_4 NS_112 0 -3.4752160401910813e-06
GC_4_113 b_4 NI_4 NS_113 0 -3.6812594745616302e-04
GC_4_114 b_4 NI_4 NS_114 0 1.3598225788758885e-04
GC_4_115 b_4 NI_4 NS_115 0 1.1297229763767268e-03
GC_4_116 b_4 NI_4 NS_116 0 1.9432473205368420e-03
GC_4_117 b_4 NI_4 NS_117 0 -6.5058844844250330e-05
GC_4_118 b_4 NI_4 NS_118 0 -3.4937471194254246e-03
GC_4_119 b_4 NI_4 NS_119 0 -1.5644007768149523e-03
GC_4_120 b_4 NI_4 NS_120 0 5.0906039852630040e-03
GC_4_121 b_4 NI_4 NS_121 0 4.2533992707037326e-03
GC_4_122 b_4 NI_4 NS_122 0 -4.9938033549717332e-03
GC_4_123 b_4 NI_4 NS_123 0 -1.0085547500383015e-03
GC_4_124 b_4 NI_4 NS_124 0 5.6397878414695963e-04
GC_4_125 b_4 NI_4 NS_125 0 -2.0807515128245346e-03
GC_4_126 b_4 NI_4 NS_126 0 -1.8633117462639945e-03
GC_4_127 b_4 NI_4 NS_127 0 3.6454397848812324e-03
GC_4_128 b_4 NI_4 NS_128 0 1.1647366929189523e-02
GC_4_129 b_4 NI_4 NS_129 0 -8.9814148433892973e-04
GC_4_130 b_4 NI_4 NS_130 0 -1.4854322544909182e-02
GC_4_131 b_4 NI_4 NS_131 0 -8.1235361409249581e-03
GC_4_132 b_4 NI_4 NS_132 0 1.9196061448188558e-03
GC_4_133 b_4 NI_4 NS_133 0 1.1263056429845044e-02
GC_4_134 b_4 NI_4 NS_134 0 -1.8122318494942112e-03
GC_4_135 b_4 NI_4 NS_135 0 -7.5672718811669332e-03
GC_4_136 b_4 NI_4 NS_136 0 -1.6811818303357035e-03
GC_4_137 b_4 NI_4 NS_137 0 1.5281711114416554e-02
GC_4_138 b_4 NI_4 NS_138 0 5.3008448871395908e-03
GC_4_139 b_4 NI_4 NS_139 0 -1.3082856901286993e-02
GC_4_140 b_4 NI_4 NS_140 0 -5.4612973807671994e-03
GC_4_141 b_4 NI_4 NS_141 0 -6.6370717898199226e-03
GC_4_142 b_4 NI_4 NS_142 0 3.4566938999519591e-03
GC_4_143 b_4 NI_4 NS_143 0 6.3616039737471155e-03
GC_4_144 b_4 NI_4 NS_144 0 -1.8793243531983461e-03
GC_4_145 b_4 NI_4 NS_145 0 -5.4737176496378664e-03
GC_4_146 b_4 NI_4 NS_146 0 2.1830271440324328e-03
GC_4_147 b_4 NI_4 NS_147 0 5.3937683808071499e-03
GC_4_148 b_4 NI_4 NS_148 0 -2.6324374322198932e-03
GC_4_149 b_4 NI_4 NS_149 0 -6.3064546626286156e-03
GC_4_150 b_4 NI_4 NS_150 0 -4.8381472979925044e-04
GC_4_151 b_4 NI_4 NS_151 0 7.6452800868578369e-03
GC_4_152 b_4 NI_4 NS_152 0 3.6298731644361453e-03
GC_4_153 b_4 NI_4 NS_153 0 -5.8336241546881346e-03
GC_4_154 b_4 NI_4 NS_154 0 -3.4645948161465506e-03
GC_4_155 b_4 NI_4 NS_155 0 2.9620035999771311e-04
GC_4_156 b_4 NI_4 NS_156 0 5.5810466131066857e-04
GC_4_157 b_4 NI_4 NS_157 0 -4.9270628232564451e-03
GC_4_158 b_4 NI_4 NS_158 0 8.9219828285828483e-04
GC_4_159 b_4 NI_4 NS_159 0 6.2063416449247514e-03
GC_4_160 b_4 NI_4 NS_160 0 6.8827498974224747e-04
GC_4_161 b_4 NI_4 NS_161 0 -5.3209621302306052e-03
GC_4_162 b_4 NI_4 NS_162 0 -4.8418936157540796e-04
GC_4_163 b_4 NI_4 NS_163 0 1.5503327183282488e-03
GC_4_164 b_4 NI_4 NS_164 0 -4.3207881715928786e-05
GC_4_165 b_4 NI_4 NS_165 0 -6.0223328282395273e-03
GC_4_166 b_4 NI_4 NS_166 0 1.9232412388156532e-03
GC_4_167 b_4 NI_4 NS_167 0 6.2616666845880763e-03
GC_4_168 b_4 NI_4 NS_168 0 2.1736210808271910e-04
GC_4_169 b_4 NI_4 NS_169 0 -5.0591984910259803e-03
GC_4_170 b_4 NI_4 NS_170 0 1.7016163938301965e-03
GC_4_171 b_4 NI_4 NS_171 0 2.4884732755286248e-03
GC_4_172 b_4 NI_4 NS_172 0 -9.5765139659464288e-04
GC_4_173 b_4 NI_4 NS_173 0 -6.5329629517140875e-03
GC_4_174 b_4 NI_4 NS_174 0 3.8846376440248341e-03
GC_4_175 b_4 NI_4 NS_175 0 7.4932677112668307e-03
GC_4_176 b_4 NI_4 NS_176 0 -1.0960274168074187e-03
GC_4_177 b_4 NI_4 NS_177 0 -3.9851190206327764e-03
GC_4_178 b_4 NI_4 NS_178 0 4.0409800030220180e-03
GC_4_179 b_4 NI_4 NS_179 0 2.8633260159070047e-03
GC_4_180 b_4 NI_4 NS_180 0 -3.0534889780626405e-03
GC_4_181 b_4 NI_4 NS_181 0 -6.0227292283394698e-03
GC_4_182 b_4 NI_4 NS_182 0 7.2373892458611937e-03
GC_4_183 b_4 NI_4 NS_183 0 7.9897111884946852e-03
GC_4_184 b_4 NI_4 NS_184 0 -4.8114595179570294e-03
GC_4_185 b_4 NI_4 NS_185 0 -5.3741900587964044e-04
GC_4_186 b_4 NI_4 NS_186 0 5.0204728214654380e-03
GC_4_187 b_4 NI_4 NS_187 0 2.4825551867528546e-04
GC_4_188 b_4 NI_4 NS_188 0 -4.7581976238974862e-03
GC_4_189 b_4 NI_4 NS_189 0 1.8109240222801872e-09
GC_4_190 b_4 NI_4 NS_190 0 3.2744954075368164e-09
GC_4_191 b_4 NI_4 NS_191 0 -1.4271962552611062e-03
GC_4_192 b_4 NI_4 NS_192 0 7.8707399683173810e-03
GC_4_193 b_4 NI_4 NS_193 0 -1.7997930789362258e-04
GC_4_194 b_4 NI_4 NS_194 0 3.0272441092164255e-03
GC_4_195 b_4 NI_4 NS_195 0 -1.3038553844318902e-04
GC_4_196 b_4 NI_4 NS_196 0 -3.3753037109675575e-03
GC_4_197 b_4 NI_4 NS_197 0 -8.7631252272640835e-04
GC_4_198 b_4 NI_4 NS_198 0 7.5304828375111028e-03
GC_4_199 b_4 NI_4 NS_199 0 3.7888078333956901e-03
GC_4_200 b_4 NI_4 NS_200 0 -6.1574210765510187e-03
GC_4_201 b_4 NI_4 NS_201 0 8.6236229003774553e-08
GC_4_202 b_4 NI_4 NS_202 0 -3.5294047713599015e-07
GC_4_203 b_4 NI_4 NS_203 0 6.7186801410480043e-03
GC_4_204 b_4 NI_4 NS_204 0 -5.3194116319874403e-03
GC_4_205 b_4 NI_4 NS_205 0 -2.6111716282871795e-03
GC_4_206 b_4 NI_4 NS_206 0 6.0542407327173423e-03
GC_4_207 b_4 NI_4 NS_207 0 -4.2922714918981345e-03
GC_4_208 b_4 NI_4 NS_208 0 1.4429424531418159e-05
GC_4_209 b_4 NI_4 NS_209 0 2.7173890707041519e-03
GC_4_210 b_4 NI_4 NS_210 0 -6.2040229558799308e-03
GC_4_211 b_4 NI_4 NS_211 0 2.0957200635848047e-03
GC_4_212 b_4 NI_4 NS_212 0 3.2562725001881294e-03
GC_4_213 b_4 NI_4 NS_213 0 -1.9700344228987723e-03
GC_4_214 b_4 NI_4 NS_214 0 -4.4205369355976437e-03
GC_4_215 b_4 NI_4 NS_215 0 2.8640861853323207e-03
GC_4_216 b_4 NI_4 NS_216 0 8.0083630617668201e-03
GC_4_217 b_4 NI_4 NS_217 0 -1.0575543390287998e-02
GC_4_218 b_4 NI_4 NS_218 0 9.5500570048345293e-09
GC_4_219 b_4 NI_4 NS_219 0 9.8517511441656238e-07
GC_4_220 b_4 NI_4 NS_220 0 3.6184007362585494e-05
GC_4_221 b_4 NI_4 NS_221 0 4.3796968247234265e-03
GC_4_222 b_4 NI_4 NS_222 0 -3.4738253478814106e-03
GC_4_223 b_4 NI_4 NS_223 0 -3.7303117957833399e-03
GC_4_224 b_4 NI_4 NS_224 0 6.2452214585123735e-03
GC_4_225 b_4 NI_4 NS_225 0 -8.7506176751483717e-03
GC_4_226 b_4 NI_4 NS_226 0 -5.9709679155804714e-03
GC_4_227 b_4 NI_4 NS_227 0 9.2221539742008678e-03
GC_4_228 b_4 NI_4 NS_228 0 -5.9539856734248118e-03
GC_4_229 b_4 NI_4 NS_229 0 7.1416220231734547e-03
GC_4_230 b_4 NI_4 NS_230 0 1.1891292787261018e-02
GC_4_231 b_4 NI_4 NS_231 0 -4.2237377927143568e-03
GC_4_232 b_4 NI_4 NS_232 0 -1.1434228656134978e-03
GC_4_233 b_4 NI_4 NS_233 0 -8.8759855077183095e-03
GC_4_234 b_4 NI_4 NS_234 0 -4.8953453755559890e-04
GC_4_235 b_4 NI_4 NS_235 0 1.4613642594067168e-02
GC_4_236 b_4 NI_4 NS_236 0 -1.0366838583162360e-02
GC_4_237 b_4 NI_4 NS_237 0 1.6418112296657260e-02
GC_4_238 b_4 NI_4 NS_238 0 4.0449085810566419e-03
GC_4_239 b_4 NI_4 NS_239 0 -1.1484885842428880e-02
GC_4_240 b_4 NI_4 NS_240 0 -2.5530968993815934e-04
GC_4_241 b_4 NI_4 NS_241 0 -1.6635876461258185e-02
GC_4_242 b_4 NI_4 NS_242 0 -4.4594577683613426e-02
GC_4_243 b_4 NI_4 NS_243 0 1.0649468919889587e-02
GC_4_244 b_4 NI_4 NS_244 0 1.1312753596659174e-03
GC_4_245 b_4 NI_4 NS_245 0 -4.8338782796399311e-02
GC_4_246 b_4 NI_4 NS_246 0 1.1008133577368530e-02
GC_4_247 b_4 NI_4 NS_247 0 -1.0431967215636684e-02
GC_4_248 b_4 NI_4 NS_248 0 4.9180137810140938e-04
GC_4_249 b_4 NI_4 NS_249 0 9.7750322510752208e-03
GC_4_250 b_4 NI_4 NS_250 0 -5.7663577021140229e-04
GC_4_251 b_4 NI_4 NS_251 0 4.5630558426753608e-03
GC_4_252 b_4 NI_4 NS_252 0 2.4175329263178238e-02
GC_4_253 b_4 NI_4 NS_253 0 -1.0747433455818047e-02
GC_4_254 b_4 NI_4 NS_254 0 1.9593868633228091e-03
GC_4_255 b_4 NI_4 NS_255 0 -8.4817663253616837e-03
GC_4_256 b_4 NI_4 NS_256 0 -1.3531579896405481e-02
GC_4_257 b_4 NI_4 NS_257 0 1.0144386457718632e-02
GC_4_258 b_4 NI_4 NS_258 0 9.9161527106657581e-04
GC_4_259 b_4 NI_4 NS_259 0 -1.9215689083992179e-02
GC_4_260 b_4 NI_4 NS_260 0 2.8664526916828432e-02
GC_4_261 b_4 NI_4 NS_261 0 -9.6176497180131375e-03
GC_4_262 b_4 NI_4 NS_262 0 -9.6670704864721009e-04
GC_4_263 b_4 NI_4 NS_263 0 1.8850184091243186e-03
GC_4_264 b_4 NI_4 NS_264 0 -1.3791037344946439e-03
GC_4_265 b_4 NI_4 NS_265 0 9.4567927089606423e-03
GC_4_266 b_4 NI_4 NS_266 0 -2.3686791589521466e-04
GC_4_267 b_4 NI_4 NS_267 0 -2.0777099666938171e-04
GC_4_268 b_4 NI_4 NS_268 0 3.0287198920892912e-02
GC_4_269 b_4 NI_4 NS_269 0 -8.5365287638884801e-03
GC_4_270 b_4 NI_4 NS_270 0 1.5565498022713421e-04
GC_4_271 b_4 NI_4 NS_271 0 2.0683702788054732e-04
GC_4_272 b_4 NI_4 NS_272 0 -5.4692371141128789e-03
GC_4_273 b_4 NI_4 NS_273 0 1.0024582664773558e-02
GC_4_274 b_4 NI_4 NS_274 0 -3.2646570941148101e-04
GC_4_275 b_4 NI_4 NS_275 0 8.8939963060280930e-03
GC_4_276 b_4 NI_4 NS_276 0 2.6408684340642318e-02
GC_4_277 b_4 NI_4 NS_277 0 -8.3634846280485099e-03
GC_4_278 b_4 NI_4 NS_278 0 1.3809707151292219e-03
GC_4_279 b_4 NI_4 NS_279 0 -2.5880174875845593e-03
GC_4_280 b_4 NI_4 NS_280 0 -7.3315849346175417e-03
GC_4_281 b_4 NI_4 NS_281 0 1.0540510272077497e-02
GC_4_282 b_4 NI_4 NS_282 0 -8.1042019463104594e-04
GC_4_283 b_4 NI_4 NS_283 0 1.4431068337973474e-02
GC_4_284 b_4 NI_4 NS_284 0 2.0002785824478633e-02
GC_4_285 b_4 NI_4 NS_285 0 -8.2822297589726247e-03
GC_4_286 b_4 NI_4 NS_286 0 2.9407040205225447e-03
GC_4_287 b_4 NI_4 NS_287 0 -5.5808241983728562e-03
GC_4_288 b_4 NI_4 NS_288 0 -6.8969132264541586e-03
GC_4_289 b_4 NI_4 NS_289 0 1.1228113575450170e-02
GC_4_290 b_4 NI_4 NS_290 0 -1.3571866112998129e-03
GC_4_291 b_4 NI_4 NS_291 0 1.5726445902255297e-02
GC_4_292 b_4 NI_4 NS_292 0 1.2982511064230930e-02
GC_4_293 b_4 NI_4 NS_293 0 -7.1842451639626366e-03
GC_4_294 b_4 NI_4 NS_294 0 5.1249333809084540e-03
GC_4_295 b_4 NI_4 NS_295 0 -6.8612321581334561e-03
GC_4_296 b_4 NI_4 NS_296 0 -4.8303664787581113e-03
GC_4_297 b_4 NI_4 NS_297 0 5.1317157772654806e-09
GC_4_298 b_4 NI_4 NS_298 0 4.4376330546090372e-08
GC_4_299 b_4 NI_4 NS_299 0 1.2002064975706925e-02
GC_4_300 b_4 NI_4 NS_300 0 -2.5554093666726395e-03
GC_4_301 b_4 NI_4 NS_301 0 -5.2431620135277544e-03
GC_4_302 b_4 NI_4 NS_302 0 4.7077205115174780e-03
GC_4_303 b_4 NI_4 NS_303 0 -6.1541469583877651e-03
GC_4_304 b_4 NI_4 NS_304 0 -4.3159830596897044e-03
GC_4_305 b_4 NI_4 NS_305 0 1.1759634246399640e-02
GC_4_306 b_4 NI_4 NS_306 0 -3.7148948887488638e-03
GC_4_307 b_4 NI_4 NS_307 0 1.3000710298869456e-02
GC_4_308 b_4 NI_4 NS_308 0 9.4708365789193741e-03
GC_4_309 b_4 NI_4 NS_309 0 3.9444932660188372e-06
GC_4_310 b_4 NI_4 NS_310 0 -9.3342785565435420e-07
GC_4_311 b_4 NI_4 NS_311 0 1.6111756422071469e-02
GC_4_312 b_4 NI_4 NS_312 0 1.6784785992348825e-02
GC_4_313 b_4 NI_4 NS_313 0 1.2052345778950813e-02
GC_4_314 b_4 NI_4 NS_314 0 -2.4747668173413320e-03
GC_4_315 b_4 NI_4 NS_315 0 -8.3473636716150362e-03
GC_4_316 b_4 NI_4 NS_316 0 8.3965830747979455e-05
GC_4_317 b_4 NI_4 NS_317 0 1.1340533638883226e-02
GC_4_318 b_4 NI_4 NS_318 0 7.3400203287226429e-03
GC_4_319 b_4 NI_4 NS_319 0 -4.6549299349229320e-03
GC_4_320 b_4 NI_4 NS_320 0 7.3654668652397681e-03
GC_4_321 b_4 NI_4 NS_321 0 -8.0793046197459150e-03
GC_4_322 b_4 NI_4 NS_322 0 -3.7189982954207623e-03
GC_4_323 b_4 NI_4 NS_323 0 1.5982958496217253e-02
GC_4_324 b_4 NI_4 NS_324 0 -7.7385028191496825e-03
GC_4_325 b_4 NI_4 NS_325 0 -1.4246404788187667e-02
GC_4_326 b_4 NI_4 NS_326 0 6.2292709467999834e-09
GC_4_327 b_4 NI_4 NS_327 0 -1.0771398389490103e-06
GC_4_328 b_4 NI_4 NS_328 0 -2.3238216360955485e-05
GC_4_329 b_4 NI_4 NS_329 0 3.4199237682637295e-04
GC_4_330 b_4 NI_4 NS_330 0 -1.9835152991893974e-04
GC_4_331 b_4 NI_4 NS_331 0 -1.5573879029213494e-03
GC_4_332 b_4 NI_4 NS_332 0 -2.3367654356295526e-03
GC_4_333 b_4 NI_4 NS_333 0 -6.7659612820999238e-05
GC_4_334 b_4 NI_4 NS_334 0 4.3764657852802796e-03
GC_4_335 b_4 NI_4 NS_335 0 1.6012883084795394e-03
GC_4_336 b_4 NI_4 NS_336 0 -5.9363758342384264e-03
GC_4_337 b_4 NI_4 NS_337 0 -4.9862911833464937e-03
GC_4_338 b_4 NI_4 NS_338 0 6.4938614129151978e-03
GC_4_339 b_4 NI_4 NS_339 0 1.1242578186705355e-03
GC_4_340 b_4 NI_4 NS_340 0 -4.9042040139161286e-04
GC_4_341 b_4 NI_4 NS_341 0 2.8092111687196991e-03
GC_4_342 b_4 NI_4 NS_342 0 2.3585345818560068e-03
GC_4_343 b_4 NI_4 NS_343 0 -4.3182654913181510e-03
GC_4_344 b_4 NI_4 NS_344 0 -1.3539568144360628e-02
GC_4_345 b_4 NI_4 NS_345 0 1.6031664291941690e-03
GC_4_346 b_4 NI_4 NS_346 0 1.7677771464974915e-02
GC_4_347 b_4 NI_4 NS_347 0 9.8386848386797544e-03
GC_4_348 b_4 NI_4 NS_348 0 -2.2919450913236757e-03
GC_4_349 b_4 NI_4 NS_349 0 -1.3104488469256876e-02
GC_4_350 b_4 NI_4 NS_350 0 2.2186341526221525e-03
GC_4_351 b_4 NI_4 NS_351 0 9.2001452439411501e-03
GC_4_352 b_4 NI_4 NS_352 0 1.9506157451927473e-03
GC_4_353 b_4 NI_4 NS_353 0 -1.7998042638950867e-02
GC_4_354 b_4 NI_4 NS_354 0 -6.4920168015484619e-03
GC_4_355 b_4 NI_4 NS_355 0 1.5711165321299507e-02
GC_4_356 b_4 NI_4 NS_356 0 6.4981562116889040e-03
GC_4_357 b_4 NI_4 NS_357 0 8.1166009630612157e-03
GC_4_358 b_4 NI_4 NS_358 0 -4.1938588857842107e-03
GC_4_359 b_4 NI_4 NS_359 0 -7.5320606970616889e-03
GC_4_360 b_4 NI_4 NS_360 0 2.0324568159713814e-03
GC_4_361 b_4 NI_4 NS_361 0 6.7023910841256858e-03
GC_4_362 b_4 NI_4 NS_362 0 -2.7451381598352174e-03
GC_4_363 b_4 NI_4 NS_363 0 -6.5840253691330829e-03
GC_4_364 b_4 NI_4 NS_364 0 2.8920130832388014e-03
GC_4_365 b_4 NI_4 NS_365 0 7.6634840947172617e-03
GC_4_366 b_4 NI_4 NS_366 0 4.8601872493882306e-04
GC_4_367 b_4 NI_4 NS_367 0 -9.3542511629111005e-03
GC_4_368 b_4 NI_4 NS_368 0 -5.1821771855508677e-03
GC_4_369 b_4 NI_4 NS_369 0 6.8205103837088556e-03
GC_4_370 b_4 NI_4 NS_370 0 4.1105940199482162e-03
GC_4_371 b_4 NI_4 NS_371 0 -3.8505207999990567e-04
GC_4_372 b_4 NI_4 NS_372 0 -9.3423363189744173e-04
GC_4_373 b_4 NI_4 NS_373 0 5.6830631042289600e-03
GC_4_374 b_4 NI_4 NS_374 0 -1.3773228603985231e-03
GC_4_375 b_4 NI_4 NS_375 0 -9.1525454294961502e-03
GC_4_376 b_4 NI_4 NS_376 0 -1.2845789187938914e-03
GC_4_377 b_4 NI_4 NS_377 0 5.9995882824453407e-03
GC_4_378 b_4 NI_4 NS_378 0 7.3474304397221839e-04
GC_4_379 b_4 NI_4 NS_379 0 -2.6407567579047634e-03
GC_4_380 b_4 NI_4 NS_380 0 2.3245280178849426e-04
GC_4_381 b_4 NI_4 NS_381 0 6.7119805317869098e-03
GC_4_382 b_4 NI_4 NS_382 0 -2.2566103582135947e-03
GC_4_383 b_4 NI_4 NS_383 0 -9.2876884338957064e-03
GC_4_384 b_4 NI_4 NS_384 0 1.4716553638630440e-03
GC_4_385 b_4 NI_4 NS_385 0 5.7396080224355892e-03
GC_4_386 b_4 NI_4 NS_386 0 -1.5055505373888971e-03
GC_4_387 b_4 NI_4 NS_387 0 -3.3169949944615753e-03
GC_4_388 b_4 NI_4 NS_388 0 2.3821032594901143e-03
GC_4_389 b_4 NI_4 NS_389 0 7.2818918524709996e-03
GC_4_390 b_4 NI_4 NS_390 0 -4.0976815562003086e-03
GC_4_391 b_4 NI_4 NS_391 0 -8.5931435656789474e-03
GC_4_392 b_4 NI_4 NS_392 0 4.1427791364397988e-03
GC_4_393 b_4 NI_4 NS_393 0 4.8244372078948116e-03
GC_4_394 b_4 NI_4 NS_394 0 -3.8807298253238950e-03
GC_4_395 b_4 NI_4 NS_395 0 -2.4175657565256555e-03
GC_4_396 b_4 NI_4 NS_396 0 4.7355224271884381e-03
GC_4_397 b_4 NI_4 NS_397 0 7.0698650818163530e-03
GC_4_398 b_4 NI_4 NS_398 0 -7.3594023641606627e-03
GC_4_399 b_4 NI_4 NS_399 0 -7.1573594779315323e-03
GC_4_400 b_4 NI_4 NS_400 0 6.8575806727569433e-03
GC_4_401 b_4 NI_4 NS_401 0 1.6629093812799123e-03
GC_4_402 b_4 NI_4 NS_402 0 -5.3099129266202935e-03
GC_4_403 b_4 NI_4 NS_403 0 5.8005275187150045e-04
GC_4_404 b_4 NI_4 NS_404 0 5.4707651829515600e-03
GC_4_405 b_4 NI_4 NS_405 0 -4.5823953993476213e-09
GC_4_406 b_4 NI_4 NS_406 0 -1.3467243226158302e-08
GC_4_407 b_4 NI_4 NS_407 0 2.7089353287049868e-03
GC_4_408 b_4 NI_4 NS_408 0 -8.5910076750723742e-03
GC_4_409 b_4 NI_4 NS_409 0 8.6608621310450200e-04
GC_4_410 b_4 NI_4 NS_410 0 -3.4347601326465693e-03
GC_4_411 b_4 NI_4 NS_411 0 6.2756504024875069e-04
GC_4_412 b_4 NI_4 NS_412 0 4.0313421846027205e-03
GC_4_413 b_4 NI_4 NS_413 0 2.1670469590615825e-03
GC_4_414 b_4 NI_4 NS_414 0 -8.1665277303216172e-03
GC_4_415 b_4 NI_4 NS_415 0 -3.4991650927442843e-03
GC_4_416 b_4 NI_4 NS_416 0 7.0126800881229173e-03
GC_4_417 b_4 NI_4 NS_417 0 -1.0829953942224426e-07
GC_4_418 b_4 NI_4 NS_418 0 -3.0048136554598339e-07
GC_4_419 b_4 NI_4 NS_419 0 -8.0240637224035117e-03
GC_4_420 b_4 NI_4 NS_420 0 5.3776064418066642e-03
GC_4_421 b_4 NI_4 NS_421 0 4.1768099630320309e-03
GC_4_422 b_4 NI_4 NS_422 0 -6.8620735186215847e-03
GC_4_423 b_4 NI_4 NS_423 0 5.3214176226709601e-03
GC_4_424 b_4 NI_4 NS_424 0 7.4369290354658012e-04
GC_4_425 b_4 NI_4 NS_425 0 -2.3651598819096082e-03
GC_4_426 b_4 NI_4 NS_426 0 6.8561912681336483e-03
GC_4_427 b_4 NI_4 NS_427 0 -1.4960018488862027e-03
GC_4_428 b_4 NI_4 NS_428 0 -4.2193419650893085e-03
GC_4_429 b_4 NI_4 NS_429 0 2.3601154435927748e-03
GC_4_430 b_4 NI_4 NS_430 0 5.0361471043601381e-03
GC_4_431 b_4 NI_4 NS_431 0 -2.0068775958372222e-03
GC_4_432 b_4 NI_4 NS_432 0 -8.9761633823016562e-03
GC_4_433 b_4 NI_4 NS_433 0 -6.4105871955193823e-04
GC_4_434 b_4 NI_4 NS_434 0 -9.7197843542628142e-11
GC_4_435 b_4 NI_4 NS_435 0 3.8858267089041561e-09
GC_4_436 b_4 NI_4 NS_436 0 -6.7399752296316684e-08
GC_4_437 b_4 NI_4 NS_437 0 -1.1325348013250873e-05
GC_4_438 b_4 NI_4 NS_438 0 -9.3599518509370960e-06
GC_4_439 b_4 NI_4 NS_439 0 -2.2402039620116331e-06
GC_4_440 b_4 NI_4 NS_440 0 1.9787536243740949e-07
GC_4_441 b_4 NI_4 NS_441 0 -3.0414374000577836e-05
GC_4_442 b_4 NI_4 NS_442 0 2.7141385993251129e-05
GC_4_443 b_4 NI_4 NS_443 0 -3.3444223147780053e-05
GC_4_444 b_4 NI_4 NS_444 0 8.1131373725379616e-06
GC_4_445 b_4 NI_4 NS_445 0 3.1774136273666374e-05
GC_4_446 b_4 NI_4 NS_446 0 2.7463325592563718e-05
GC_4_447 b_4 NI_4 NS_447 0 -9.1036096296775066e-06
GC_4_448 b_4 NI_4 NS_448 0 1.4796420308263693e-05
GC_4_449 b_4 NI_4 NS_449 0 1.2667861992621178e-05
GC_4_450 b_4 NI_4 NS_450 0 3.7134953331918569e-05
GC_4_451 b_4 NI_4 NS_451 0 -1.1026758187655488e-05
GC_4_452 b_4 NI_4 NS_452 0 6.8453876774598430e-05
GC_4_453 b_4 NI_4 NS_453 0 9.5993846769765797e-05
GC_4_454 b_4 NI_4 NS_454 0 -6.6259875316651196e-05
GC_4_455 b_4 NI_4 NS_455 0 2.7201066028124882e-05
GC_4_456 b_4 NI_4 NS_456 0 3.2003861426467150e-05
GC_4_457 b_4 NI_4 NS_457 0 -7.0532285320554775e-06
GC_4_458 b_4 NI_4 NS_458 0 -7.2616526499663553e-05
GC_4_459 b_4 NI_4 NS_459 0 -9.8457000725717954e-06
GC_4_460 b_4 NI_4 NS_460 0 -3.4285198532702927e-05
GC_4_461 b_4 NI_4 NS_461 0 -7.6897184629675500e-05
GC_4_462 b_4 NI_4 NS_462 0 1.8745842335921118e-05
GC_4_463 b_4 NI_4 NS_463 0 2.4874738691381825e-05
GC_4_464 b_4 NI_4 NS_464 0 5.1393203366608012e-05
GC_4_465 b_4 NI_4 NS_465 0 -2.3342758699503438e-05
GC_4_466 b_4 NI_4 NS_466 0 -3.7551214972140018e-06
GC_4_467 b_4 NI_4 NS_467 0 7.0090133270947759e-05
GC_4_468 b_4 NI_4 NS_468 0 4.4926314733442104e-05
GC_4_469 b_4 NI_4 NS_469 0 2.9399642893565641e-05
GC_4_470 b_4 NI_4 NS_470 0 1.9985854366663746e-05
GC_4_471 b_4 NI_4 NS_471 0 -7.2378716798025511e-06
GC_4_472 b_4 NI_4 NS_472 0 -2.5815164602205658e-05
GC_4_473 b_4 NI_4 NS_473 0 -7.5769846525466491e-06
GC_4_474 b_4 NI_4 NS_474 0 -2.5457569325997269e-05
GC_4_475 b_4 NI_4 NS_475 0 6.9370997529349566e-06
GC_4_476 b_4 NI_4 NS_476 0 4.9224287066343327e-05
GC_4_477 b_4 NI_4 NS_477 0 1.2889462631622776e-05
GC_4_478 b_4 NI_4 NS_478 0 2.7625573325103871e-05
GC_4_479 b_4 NI_4 NS_479 0 5.8786694059064820e-06
GC_4_480 b_4 NI_4 NS_480 0 2.1442975906815052e-06
GC_4_481 b_4 NI_4 NS_481 0 -6.1843598330390246e-07
GC_4_482 b_4 NI_4 NS_482 0 -1.5585944012772863e-05
GC_4_483 b_4 NI_4 NS_483 0 5.6423068349288623e-05
GC_4_484 b_4 NI_4 NS_484 0 3.8203695310339558e-05
GC_4_485 b_4 NI_4 NS_485 0 1.9996590434712857e-05
GC_4_486 b_4 NI_4 NS_486 0 1.5002578511998205e-05
GC_4_487 b_4 NI_4 NS_487 0 8.4325782594416849e-06
GC_4_488 b_4 NI_4 NS_488 0 -1.2893607433814521e-05
GC_4_489 b_4 NI_4 NS_489 0 -5.6500498515618588e-06
GC_4_490 b_4 NI_4 NS_490 0 -1.4195057998907794e-05
GC_4_491 b_4 NI_4 NS_491 0 6.6301882329949501e-05
GC_4_492 b_4 NI_4 NS_492 0 1.2978523595337807e-05
GC_4_493 b_4 NI_4 NS_493 0 2.2841962253115839e-05
GC_4_494 b_4 NI_4 NS_494 0 5.0486960626144851e-06
GC_4_495 b_4 NI_4 NS_495 0 -5.5524339087341465e-06
GC_4_496 b_4 NI_4 NS_496 0 -2.2079814171582553e-05
GC_4_497 b_4 NI_4 NS_497 0 -9.1403007845713397e-06
GC_4_498 b_4 NI_4 NS_498 0 -7.2135381061985898e-06
GC_4_499 b_4 NI_4 NS_499 0 6.0763591083307558e-05
GC_4_500 b_4 NI_4 NS_500 0 -9.5421076452735131e-06
GC_4_501 b_4 NI_4 NS_501 0 2.1478231335777970e-05
GC_4_502 b_4 NI_4 NS_502 0 -7.3421663276382699e-06
GC_4_503 b_4 NI_4 NS_503 0 -2.3108207545479321e-05
GC_4_504 b_4 NI_4 NS_504 0 -1.3186417267361792e-05
GC_4_505 b_4 NI_4 NS_505 0 -8.6384518101472354e-06
GC_4_506 b_4 NI_4 NS_506 0 4.3948623318141781e-06
GC_4_507 b_4 NI_4 NS_507 0 4.5484326358845480e-05
GC_4_508 b_4 NI_4 NS_508 0 -2.5717099151481436e-05
GC_4_509 b_4 NI_4 NS_509 0 6.0380888824795451e-06
GC_4_510 b_4 NI_4 NS_510 0 -1.6494075837666420e-05
GC_4_511 b_4 NI_4 NS_511 0 -1.8737716665504468e-05
GC_4_512 b_4 NI_4 NS_512 0 8.6024230200458686e-06
GC_4_513 b_4 NI_4 NS_513 0 -4.6784672126388249e-11
GC_4_514 b_4 NI_4 NS_514 0 -1.7807452610673450e-10
GC_4_515 b_4 NI_4 NS_515 0 1.7771649176606838e-06
GC_4_516 b_4 NI_4 NS_516 0 8.7584987436129116e-06
GC_4_517 b_4 NI_4 NS_517 0 2.2074336392125781e-06
GC_4_518 b_4 NI_4 NS_518 0 -7.0114811359567639e-06
GC_4_519 b_4 NI_4 NS_519 0 -9.0081329858376935e-06
GC_4_520 b_4 NI_4 NS_520 0 5.7591250281312166e-06
GC_4_521 b_4 NI_4 NS_521 0 4.7915722883031584e-06
GC_4_522 b_4 NI_4 NS_522 0 1.1558576898963115e-05
GC_4_523 b_4 NI_4 NS_523 0 2.4562413509199697e-05
GC_4_524 b_4 NI_4 NS_524 0 -2.1173228386126995e-05
GC_4_525 b_4 NI_4 NS_525 0 -5.7146480984565196e-09
GC_4_526 b_4 NI_4 NS_526 0 -5.6481287784526978e-09
GC_4_527 b_4 NI_4 NS_527 0 3.0658429446850426e-05
GC_4_528 b_4 NI_4 NS_528 0 7.4840758206953014e-06
GC_4_529 b_4 NI_4 NS_529 0 -2.6776562550279763e-06
GC_4_530 b_4 NI_4 NS_530 0 1.1046089816291742e-05
GC_4_531 b_4 NI_4 NS_531 0 8.0413958588231210e-06
GC_4_532 b_4 NI_4 NS_532 0 1.1940898121836872e-06
GC_4_533 b_4 NI_4 NS_533 0 1.9118667208900317e-05
GC_4_534 b_4 NI_4 NS_534 0 -2.1563825631126743e-05
GC_4_535 b_4 NI_4 NS_535 0 -6.5506353172723640e-06
GC_4_536 b_4 NI_4 NS_536 0 -7.4600027307048289e-06
GC_4_537 b_4 NI_4 NS_537 0 -5.3917926200942202e-06
GC_4_538 b_4 NI_4 NS_538 0 1.2485350066167197e-05
GC_4_539 b_4 NI_4 NS_539 0 1.6112329650031604e-05
GC_4_540 b_4 NI_4 NS_540 0 7.3766605591956703e-06
GC_4_541 b_4 NI_4 NS_541 0 7.9312354140308633e-05
GC_4_542 b_4 NI_4 NS_542 0 -1.2174730800124704e-10
GC_4_543 b_4 NI_4 NS_543 0 -2.0288643689844102e-09
GC_4_544 b_4 NI_4 NS_544 0 3.4021536249681155e-08
GC_4_545 b_4 NI_4 NS_545 0 -3.3964217414573158e-07
GC_4_546 b_4 NI_4 NS_546 0 -3.3541268665674230e-07
GC_4_547 b_4 NI_4 NS_547 0 -5.7544868048069386e-07
GC_4_548 b_4 NI_4 NS_548 0 9.6680844876308566e-06
GC_4_549 b_4 NI_4 NS_549 0 1.3106737926963593e-05
GC_4_550 b_4 NI_4 NS_550 0 -1.2342131207504191e-05
GC_4_551 b_4 NI_4 NS_551 0 -1.7111534605521760e-05
GC_4_552 b_4 NI_4 NS_552 0 8.5766069078401313e-06
GC_4_553 b_4 NI_4 NS_553 0 2.8664513219108682e-05
GC_4_554 b_4 NI_4 NS_554 0 -7.4207270616274021e-06
GC_4_555 b_4 NI_4 NS_555 0 -2.8948009986762023e-06
GC_4_556 b_4 NI_4 NS_556 0 -3.4132500293480733e-06
GC_4_557 b_4 NI_4 NS_557 0 -3.2450867233653904e-06
GC_4_558 b_4 NI_4 NS_558 0 -1.5091692929919002e-05
GC_4_559 b_4 NI_4 NS_559 0 -2.4827137317764870e-05
GC_4_560 b_4 NI_4 NS_560 0 3.9219960424188521e-05
GC_4_561 b_4 NI_4 NS_561 0 3.6986155606637819e-05
GC_4_562 b_4 NI_4 NS_562 0 -4.7226452043939924e-05
GC_4_563 b_4 NI_4 NS_563 0 -3.0518033087277460e-05
GC_4_564 b_4 NI_4 NS_564 0 -2.1425944380860553e-05
GC_4_565 b_4 NI_4 NS_565 0 3.2013255772624888e-05
GC_4_566 b_4 NI_4 NS_566 0 2.6385821118264476e-05
GC_4_567 b_4 NI_4 NS_567 0 -1.8545782512122305e-05
GC_4_568 b_4 NI_4 NS_568 0 -2.9076767499538764e-05
GC_4_569 b_4 NI_4 NS_569 0 2.0024654870338550e-05
GC_4_570 b_4 NI_4 NS_570 0 5.9802323031988712e-05
GC_4_571 b_4 NI_4 NS_571 0 -2.0977171131556530e-05
GC_4_572 b_4 NI_4 NS_572 0 -5.5613239035211896e-05
GC_4_573 b_4 NI_4 NS_573 0 -3.1646088559443627e-05
GC_4_574 b_4 NI_4 NS_574 0 -1.2117270707260588e-05
GC_4_575 b_4 NI_4 NS_575 0 1.9560562117652856e-05
GC_4_576 b_4 NI_4 NS_576 0 1.3805678465381333e-05
GC_4_577 b_4 NI_4 NS_577 0 -2.4957519356724885e-05
GC_4_578 b_4 NI_4 NS_578 0 -1.1262954445134751e-05
GC_4_579 b_4 NI_4 NS_579 0 2.0178607426963257e-05
GC_4_580 b_4 NI_4 NS_580 0 1.0341431355727460e-05
GC_4_581 b_4 NI_4 NS_581 0 -1.8434399211936146e-05
GC_4_582 b_4 NI_4 NS_582 0 -2.1152962494996800e-05
GC_4_583 b_4 NI_4 NS_583 0 4.2938788822463120e-06
GC_4_584 b_4 NI_4 NS_584 0 3.1956498460129953e-05
GC_4_585 b_4 NI_4 NS_585 0 -8.4070372938940702e-06
GC_4_586 b_4 NI_4 NS_586 0 -2.6582372763677358e-05
GC_4_587 b_4 NI_4 NS_587 0 -2.0405921104077798e-06
GC_4_588 b_4 NI_4 NS_588 0 1.5411378349881855e-06
GC_4_589 b_4 NI_4 NS_589 0 -1.9680638295388679e-05
GC_4_590 b_4 NI_4 NS_590 0 -1.2199249561964079e-05
GC_4_591 b_4 NI_4 NS_591 0 5.5358510941108805e-06
GC_4_592 b_4 NI_4 NS_592 0 2.1303963920637647e-05
GC_4_593 b_4 NI_4 NS_593 0 -1.6264288581868473e-05
GC_4_594 b_4 NI_4 NS_594 0 -1.4842704419713367e-05
GC_4_595 b_4 NI_4 NS_595 0 9.0112775016787231e-07
GC_4_596 b_4 NI_4 NS_596 0 5.5183490818574919e-06
GC_4_597 b_4 NI_4 NS_597 0 -2.5231535237073046e-05
GC_4_598 b_4 NI_4 NS_598 0 -1.0007123607091233e-05
GC_4_599 b_4 NI_4 NS_599 0 7.5015448387752421e-06
GC_4_600 b_4 NI_4 NS_600 0 2.3879817458133976e-05
GC_4_601 b_4 NI_4 NS_601 0 -2.0944356704434570e-05
GC_4_602 b_4 NI_4 NS_602 0 -5.6383718377773360e-06
GC_4_603 b_4 NI_4 NS_603 0 5.9390405989491058e-06
GC_4_604 b_4 NI_4 NS_604 0 7.9065229387995411e-06
GC_4_605 b_4 NI_4 NS_605 0 -3.0919140146189074e-05
GC_4_606 b_4 NI_4 NS_606 0 -2.7456249925504910e-06
GC_4_607 b_4 NI_4 NS_607 0 1.8051019044687326e-05
GC_4_608 b_4 NI_4 NS_608 0 2.6173001484548499e-05
GC_4_609 b_4 NI_4 NS_609 0 -2.2120993396346091e-05
GC_4_610 b_4 NI_4 NS_610 0 6.9969215728855058e-06
GC_4_611 b_4 NI_4 NS_611 0 1.5076260638611982e-05
GC_4_612 b_4 NI_4 NS_612 0 4.4859632968719482e-06
GC_4_613 b_4 NI_4 NS_613 0 -3.5006554669752135e-05
GC_4_614 b_4 NI_4 NS_614 0 1.3594209053851188e-05
GC_4_615 b_4 NI_4 NS_615 0 3.7183707114711700e-05
GC_4_616 b_4 NI_4 NS_616 0 1.3345626770854664e-05
GC_4_617 b_4 NI_4 NS_617 0 -7.9978704203242382e-06
GC_4_618 b_4 NI_4 NS_618 0 1.9077609490381817e-05
GC_4_619 b_4 NI_4 NS_619 0 1.2877011139014643e-05
GC_4_620 b_4 NI_4 NS_620 0 -1.0946409545297071e-05
GC_4_621 b_4 NI_4 NS_621 0 1.1098384656710157e-10
GC_4_622 b_4 NI_4 NS_622 0 4.4145429538852414e-11
GC_4_623 b_4 NI_4 NS_623 0 -1.3993786649713629e-05
GC_4_624 b_4 NI_4 NS_624 0 2.6116714415893084e-05
GC_4_625 b_4 NI_4 NS_625 0 -2.1469383365712258e-06
GC_4_626 b_4 NI_4 NS_626 0 1.0637063121640112e-05
GC_4_627 b_4 NI_4 NS_627 0 6.1622217838455718e-06
GC_4_628 b_4 NI_4 NS_628 0 -8.3662943092668995e-06
GC_4_629 b_4 NI_4 NS_629 0 -8.3615490876427517e-06
GC_4_630 b_4 NI_4 NS_630 0 2.5491909469059216e-05
GC_4_631 b_4 NI_4 NS_631 0 2.5015462294645175e-05
GC_4_632 b_4 NI_4 NS_632 0 -9.9972203148208448e-06
GC_4_633 b_4 NI_4 NS_633 0 4.8733644028004104e-09
GC_4_634 b_4 NI_4 NS_634 0 -1.1064269176468085e-09
GC_4_635 b_4 NI_4 NS_635 0 2.6321438614123518e-05
GC_4_636 b_4 NI_4 NS_636 0 -1.2477166318948374e-05
GC_4_637 b_4 NI_4 NS_637 0 -8.3191199215644740e-06
GC_4_638 b_4 NI_4 NS_638 0 1.8150071152819179e-05
GC_4_639 b_4 NI_4 NS_639 0 -1.0398966348671650e-05
GC_4_640 b_4 NI_4 NS_640 0 -2.8340100322885316e-07
GC_4_641 b_4 NI_4 NS_641 0 1.9410890667805953e-05
GC_4_642 b_4 NI_4 NS_642 0 -1.4076803259079451e-05
GC_4_643 b_4 NI_4 NS_643 0 7.1589745469011103e-06
GC_4_644 b_4 NI_4 NS_644 0 1.1755238492955826e-05
GC_4_645 b_4 NI_4 NS_645 0 -1.8090536038880760e-07
GC_4_646 b_4 NI_4 NS_646 0 -1.4547113197340590e-05
GC_4_647 b_4 NI_4 NS_647 0 1.3082626884929554e-05
GC_4_648 b_4 NI_4 NS_648 0 2.7941805129107809e-05
GC_4_649 b_4 NI_4 NS_649 0 -1.4436789320089585e-04
GC_4_650 b_4 NI_4 NS_650 0 3.3291129847051269e-11
GC_4_651 b_4 NI_4 NS_651 0 3.9883491753353503e-11
GC_4_652 b_4 NI_4 NS_652 0 9.0899872849377275e-10
GC_4_653 b_4 NI_4 NS_653 0 -2.1101231866222947e-06
GC_4_654 b_4 NI_4 NS_654 0 -1.6555661739140185e-06
GC_4_655 b_4 NI_4 NS_655 0 1.8946759458589847e-06
GC_4_656 b_4 NI_4 NS_656 0 3.8512532527564929e-06
GC_4_657 b_4 NI_4 NS_657 0 3.3113087007890266e-06
GC_4_658 b_4 NI_4 NS_658 0 4.9314964068785536e-06
GC_4_659 b_4 NI_4 NS_659 0 5.8707440398216149e-06
GC_4_660 b_4 NI_4 NS_660 0 -9.1115054864706637e-06
GC_4_661 b_4 NI_4 NS_661 0 -2.5610780640025754e-06
GC_4_662 b_4 NI_4 NS_662 0 -1.3919644492729616e-05
GC_4_663 b_4 NI_4 NS_663 0 -3.5429760964838056e-06
GC_4_664 b_4 NI_4 NS_664 0 2.1898500155717740e-06
GC_4_665 b_4 NI_4 NS_665 0 3.6503630613476032e-06
GC_4_666 b_4 NI_4 NS_666 0 1.2870366146119357e-06
GC_4_667 b_4 NI_4 NS_667 0 8.0001994580517745e-06
GC_4_668 b_4 NI_4 NS_668 0 -3.9897463332545231e-05
GC_4_669 b_4 NI_4 NS_669 0 -4.4314027368061623e-05
GC_4_670 b_4 NI_4 NS_670 0 -9.3722982994154308e-07
GC_4_671 b_4 NI_4 NS_671 0 -1.4827665062907907e-05
GC_4_672 b_4 NI_4 NS_672 0 -8.5762707364395577e-06
GC_4_673 b_4 NI_4 NS_673 0 -7.2940073781811786e-05
GC_4_674 b_4 NI_4 NS_674 0 7.5520865743086441e-05
GC_4_675 b_4 NI_4 NS_675 0 4.6287952272922240e-06
GC_4_676 b_4 NI_4 NS_676 0 1.3120199142218354e-05
GC_4_677 b_4 NI_4 NS_677 0 6.2840585919585515e-05
GC_4_678 b_4 NI_4 NS_678 0 1.2320097405617202e-04
GC_4_679 b_4 NI_4 NS_679 0 3.6368075644057744e-07
GC_4_680 b_4 NI_4 NS_680 0 -3.7020256531051475e-05
GC_4_681 b_4 NI_4 NS_681 0 1.6508676413246590e-05
GC_4_682 b_4 NI_4 NS_682 0 3.9674577388750167e-06
GC_4_683 b_4 NI_4 NS_683 0 2.4448297276392644e-05
GC_4_684 b_4 NI_4 NS_684 0 -3.0458304662791298e-05
GC_4_685 b_4 NI_4 NS_685 0 -8.8966470072447820e-06
GC_4_686 b_4 NI_4 NS_686 0 -2.3403618709481641e-06
GC_4_687 b_4 NI_4 NS_687 0 -8.8833952611217703e-06
GC_4_688 b_4 NI_4 NS_688 0 2.5237533619490147e-05
GC_4_689 b_4 NI_4 NS_689 0 5.8265836605188677e-06
GC_4_690 b_4 NI_4 NS_690 0 8.4671999909409377e-06
GC_4_691 b_4 NI_4 NS_691 0 5.6328875453694550e-05
GC_4_692 b_4 NI_4 NS_692 0 2.4970423960460536e-05
GC_4_693 b_4 NI_4 NS_693 0 3.5274180692701278e-06
GC_4_694 b_4 NI_4 NS_694 0 -1.1687206742792962e-05
GC_4_695 b_4 NI_4 NS_695 0 -4.0890882826959990e-07
GC_4_696 b_4 NI_4 NS_696 0 -1.3155477319957977e-06
GC_4_697 b_4 NI_4 NS_697 0 6.8059239904187946e-06
GC_4_698 b_4 NI_4 NS_698 0 3.0643939017254706e-06
GC_4_699 b_4 NI_4 NS_699 0 4.1947964565774668e-05
GC_4_700 b_4 NI_4 NS_700 0 -1.7199000134301142e-05
GC_4_701 b_4 NI_4 NS_701 0 -2.5585878533281671e-06
GC_4_702 b_4 NI_4 NS_702 0 -7.0970298589025471e-06
GC_4_703 b_4 NI_4 NS_703 0 -3.0311256094387873e-06
GC_4_704 b_4 NI_4 NS_704 0 1.7554981243626457e-06
GC_4_705 b_4 NI_4 NS_705 0 9.5694277822978079e-06
GC_4_706 b_4 NI_4 NS_706 0 2.9162023207012282e-06
GC_4_707 b_4 NI_4 NS_707 0 2.2976236247144082e-05
GC_4_708 b_4 NI_4 NS_708 0 -3.1187894088032165e-05
GC_4_709 b_4 NI_4 NS_709 0 -5.6936511965148459e-06
GC_4_710 b_4 NI_4 NS_710 0 -3.6758095533814535e-06
GC_4_711 b_4 NI_4 NS_711 0 -5.6141489831843492e-07
GC_4_712 b_4 NI_4 NS_712 0 5.0284085631909380e-06
GC_4_713 b_4 NI_4 NS_713 0 1.2292663292051253e-05
GC_4_714 b_4 NI_4 NS_714 0 2.0426126159120290e-07
GC_4_715 b_4 NI_4 NS_715 0 1.9186165369991448e-06
GC_4_716 b_4 NI_4 NS_716 0 -3.1503873755539763e-05
GC_4_717 b_4 NI_4 NS_717 0 -6.7230962212731239e-06
GC_4_718 b_4 NI_4 NS_718 0 9.4617189644474709e-07
GC_4_719 b_4 NI_4 NS_719 0 4.5912196268598299e-06
GC_4_720 b_4 NI_4 NS_720 0 3.8667658402348100e-06
GC_4_721 b_4 NI_4 NS_721 0 1.4096640884216375e-05
GC_4_722 b_4 NI_4 NS_722 0 -6.0051917731777323e-06
GC_4_723 b_4 NI_4 NS_723 0 -1.3991434852604207e-05
GC_4_724 b_4 NI_4 NS_724 0 -1.8834469558181233e-05
GC_4_725 b_4 NI_4 NS_725 0 -2.5005431580136941e-06
GC_4_726 b_4 NI_4 NS_726 0 5.3958760513212211e-06
GC_4_727 b_4 NI_4 NS_727 0 4.6402114121465328e-06
GC_4_728 b_4 NI_4 NS_728 0 -2.0953703644950450e-06
GC_4_729 b_4 NI_4 NS_729 0 -1.4467290988382671e-11
GC_4_730 b_4 NI_4 NS_730 0 3.9854311259675119e-12
GC_4_731 b_4 NI_4 NS_731 0 5.2050945305161063e-06
GC_4_732 b_4 NI_4 NS_732 0 -1.1255676673576374e-05
GC_4_733 b_4 NI_4 NS_733 0 -2.6207647012538367e-07
GC_4_734 b_4 NI_4 NS_734 0 2.9240500451002252e-06
GC_4_735 b_4 NI_4 NS_735 0 2.6491334526366350e-06
GC_4_736 b_4 NI_4 NS_736 0 -1.6106315958801221e-06
GC_4_737 b_4 NI_4 NS_737 0 2.4311641080702080e-06
GC_4_738 b_4 NI_4 NS_738 0 -9.4257315615735216e-06
GC_4_739 b_4 NI_4 NS_739 0 -9.9191376567381823e-06
GC_4_740 b_4 NI_4 NS_740 0 -3.6953370973670289e-06
GC_4_741 b_4 NI_4 NS_741 0 3.1960030768076237e-10
GC_4_742 b_4 NI_4 NS_742 0 2.6398622099600089e-10
GC_4_743 b_4 NI_4 NS_743 0 -8.5810754083047748e-06
GC_4_744 b_4 NI_4 NS_744 0 -5.7196778758790075e-06
GC_4_745 b_4 NI_4 NS_745 0 2.2759195467606458e-06
GC_4_746 b_4 NI_4 NS_746 0 -6.4442955626889546e-06
GC_4_747 b_4 NI_4 NS_747 0 -3.0692683121084721e-06
GC_4_748 b_4 NI_4 NS_748 0 -1.3767743112562981e-07
GC_4_749 b_4 NI_4 NS_749 0 -7.9176040315324018e-06
GC_4_750 b_4 NI_4 NS_750 0 4.8798758098282946e-07
GC_4_751 b_4 NI_4 NS_751 0 3.0157302238879673e-06
GC_4_752 b_4 NI_4 NS_752 0 2.8670059690536483e-06
GC_4_753 b_4 NI_4 NS_753 0 1.2342825820782177e-06
GC_4_754 b_4 NI_4 NS_754 0 -3.9109850755549164e-06
GC_4_755 b_4 NI_4 NS_755 0 -4.8692367853999883e-06
GC_4_756 b_4 NI_4 NS_756 0 -3.9053572815086359e-06
GC_4_757 b_4 NI_4 NS_757 0 -2.8450100285876385e-05
GC_4_758 b_4 NI_4 NS_758 0 -9.0137948500863433e-13
GC_4_759 b_4 NI_4 NS_759 0 -2.3532348446608338e-10
GC_4_760 b_4 NI_4 NS_760 0 1.0469899375618505e-08
GC_4_761 b_4 NI_4 NS_761 0 7.2361380917118775e-07
GC_4_762 b_4 NI_4 NS_762 0 1.1682421364628972e-07
GC_4_763 b_4 NI_4 NS_763 0 3.2158789644032236e-06
GC_4_764 b_4 NI_4 NS_764 0 -1.3848969436930007e-06
GC_4_765 b_4 NI_4 NS_765 0 -2.7214325366975932e-06
GC_4_766 b_4 NI_4 NS_766 0 -2.8594433591596203e-06
GC_4_767 b_4 NI_4 NS_767 0 5.0260144190128289e-06
GC_4_768 b_4 NI_4 NS_768 0 -5.8504264162792141e-07
GC_4_769 b_4 NI_4 NS_769 0 -7.0572385605663288e-06
GC_4_770 b_4 NI_4 NS_770 0 -8.2657448865058530e-06
GC_4_771 b_4 NI_4 NS_771 0 8.4163828882739141e-08
GC_4_772 b_4 NI_4 NS_772 0 -1.5979811471661405e-06
GC_4_773 b_4 NI_4 NS_773 0 -6.1458564485398593e-06
GC_4_774 b_4 NI_4 NS_774 0 1.8452524484335932e-06
GC_4_775 b_4 NI_4 NS_775 0 5.3927006212414955e-06
GC_4_776 b_4 NI_4 NS_776 0 -5.9846568399380461e-06
GC_4_777 b_4 NI_4 NS_777 0 -1.7353900592704186e-05
GC_4_778 b_4 NI_4 NS_778 0 4.6493303203767928e-06
GC_4_779 b_4 NI_4 NS_779 0 -1.1603760686569871e-06
GC_4_780 b_4 NI_4 NS_780 0 7.0453709559157944e-06
GC_4_781 b_4 NI_4 NS_781 0 -7.4845946123030352e-06
GC_4_782 b_4 NI_4 NS_782 0 -4.7597386588678325e-06
GC_4_783 b_4 NI_4 NS_783 0 -3.4153041114888180e-06
GC_4_784 b_4 NI_4 NS_784 0 8.0176901642267886e-06
GC_4_785 b_4 NI_4 NS_785 0 -2.5103464003071635e-06
GC_4_786 b_4 NI_4 NS_786 0 -4.9392794617856809e-06
GC_4_787 b_4 NI_4 NS_787 0 -3.8632873102894556e-06
GC_4_788 b_4 NI_4 NS_788 0 1.1456367934286762e-05
GC_4_789 b_4 NI_4 NS_789 0 -1.7994801919577812e-07
GC_4_790 b_4 NI_4 NS_790 0 7.1537421787439271e-06
GC_4_791 b_4 NI_4 NS_791 0 -4.3372986742722093e-06
GC_4_792 b_4 NI_4 NS_792 0 1.1467062641791373e-06
GC_4_793 b_4 NI_4 NS_793 0 -6.7842090383139085e-07
GC_4_794 b_4 NI_4 NS_794 0 7.9730689376140297e-06
GC_4_795 b_4 NI_4 NS_795 0 -1.2189495232361543e-06
GC_4_796 b_4 NI_4 NS_796 0 2.1994248042174192e-06
GC_4_797 b_4 NI_4 NS_797 0 -2.4670331447698651e-06
GC_4_798 b_4 NI_4 NS_798 0 8.1096123793415715e-06
GC_4_799 b_4 NI_4 NS_799 0 -3.9818519746548869e-07
GC_4_800 b_4 NI_4 NS_800 0 9.3212475400813040e-06
GC_4_801 b_4 NI_4 NS_801 0 -9.4389266291860176e-07
GC_4_802 b_4 NI_4 NS_802 0 8.7939544443944619e-06
GC_4_803 b_4 NI_4 NS_803 0 -1.3825918476470598e-06
GC_4_804 b_4 NI_4 NS_804 0 3.8436284110541785e-06
GC_4_805 b_4 NI_4 NS_805 0 8.7890240013768223e-07
GC_4_806 b_4 NI_4 NS_806 0 1.1882941627578669e-05
GC_4_807 b_4 NI_4 NS_807 0 1.7118686912600169e-05
GC_4_808 b_4 NI_4 NS_808 0 1.6747351655185610e-05
GC_4_809 b_4 NI_4 NS_809 0 4.6531234863139869e-06
GC_4_810 b_4 NI_4 NS_810 0 7.7083937543199952e-06
GC_4_811 b_4 NI_4 NS_811 0 9.7617612481451089e-06
GC_4_812 b_4 NI_4 NS_812 0 3.8979694206781687e-06
GC_4_813 b_4 NI_4 NS_813 0 6.3871969782148112e-06
GC_4_814 b_4 NI_4 NS_814 0 1.0670550267386323e-05
GC_4_815 b_4 NI_4 NS_815 0 3.1859678013162793e-05
GC_4_816 b_4 NI_4 NS_816 0 -5.6285997110281860e-06
GC_4_817 b_4 NI_4 NS_817 0 7.7729849572903039e-06
GC_4_818 b_4 NI_4 NS_818 0 3.3978521782737480e-06
GC_4_819 b_4 NI_4 NS_819 0 1.1412306949832902e-05
GC_4_820 b_4 NI_4 NS_820 0 -9.8828255038134044e-06
GC_4_821 b_4 NI_4 NS_821 0 1.0308208664417088e-05
GC_4_822 b_4 NI_4 NS_822 0 6.2712890554383016e-06
GC_4_823 b_4 NI_4 NS_823 0 1.5926514861075614e-05
GC_4_824 b_4 NI_4 NS_824 0 -2.9763092166948447e-05
GC_4_825 b_4 NI_4 NS_825 0 7.6989671243662563e-06
GC_4_826 b_4 NI_4 NS_826 0 -2.8503569647558329e-06
GC_4_827 b_4 NI_4 NS_827 0 -3.4066362745780672e-06
GC_4_828 b_4 NI_4 NS_828 0 -1.5683575883372885e-05
GC_4_829 b_4 NI_4 NS_829 0 1.1265212126804300e-05
GC_4_830 b_4 NI_4 NS_830 0 -1.7001885885811120e-06
GC_4_831 b_4 NI_4 NS_831 0 -1.2934680419953016e-05
GC_4_832 b_4 NI_4 NS_832 0 -2.4095960773097591e-05
GC_4_833 b_4 NI_4 NS_833 0 -4.1482548544787354e-07
GC_4_834 b_4 NI_4 NS_834 0 -6.3721082533970489e-06
GC_4_835 b_4 NI_4 NS_835 0 -9.4862698340619314e-06
GC_4_836 b_4 NI_4 NS_836 0 -2.3404459049830899e-06
GC_4_837 b_4 NI_4 NS_837 0 9.7942947225488299e-11
GC_4_838 b_4 NI_4 NS_838 0 5.4145738050290924e-11
GC_4_839 b_4 NI_4 NS_839 0 1.1788420209417217e-06
GC_4_840 b_4 NI_4 NS_840 0 -4.6057061038761645e-06
GC_4_841 b_4 NI_4 NS_841 0 -1.4797998448848681e-06
GC_4_842 b_4 NI_4 NS_842 0 -1.2848524113343879e-06
GC_4_843 b_4 NI_4 NS_843 0 -4.9236172833793944e-06
GC_4_844 b_4 NI_4 NS_844 0 -8.7275546874503299e-07
GC_4_845 b_4 NI_4 NS_845 0 -1.3800578918317433e-06
GC_4_846 b_4 NI_4 NS_846 0 -2.8436546057436237e-06
GC_4_847 b_4 NI_4 NS_847 0 -1.0040390087403215e-05
GC_4_848 b_4 NI_4 NS_848 0 -3.6858166341084989e-06
GC_4_849 b_4 NI_4 NS_849 0 6.6581513573610846e-09
GC_4_850 b_4 NI_4 NS_850 0 5.7685223502924011e-09
GC_4_851 b_4 NI_4 NS_851 0 1.3973576184362228e-06
GC_4_852 b_4 NI_4 NS_852 0 6.7929610799409382e-07
GC_4_853 b_4 NI_4 NS_853 0 -1.7307673297152600e-06
GC_4_854 b_4 NI_4 NS_854 0 3.1503400468929027e-06
GC_4_855 b_4 NI_4 NS_855 0 -9.2380472965876257e-07
GC_4_856 b_4 NI_4 NS_856 0 7.7445357331619210e-07
GC_4_857 b_4 NI_4 NS_857 0 -7.9050290128140964e-06
GC_4_858 b_4 NI_4 NS_858 0 8.2698616757449617e-07
GC_4_859 b_4 NI_4 NS_859 0 -2.4152008553846792e-06
GC_4_860 b_4 NI_4 NS_860 0 2.0790177934044485e-06
GC_4_861 b_4 NI_4 NS_861 0 -2.1277773376149892e-06
GC_4_862 b_4 NI_4 NS_862 0 2.1503900431224540e-06
GC_4_863 b_4 NI_4 NS_863 0 1.1274193490781443e-06
GC_4_864 b_4 NI_4 NS_864 0 2.8111018105601150e-06
GC_4_865 b_4 NI_4 NS_865 0 -7.7926159179902931e-06
GC_4_866 b_4 NI_4 NS_866 0 -1.0504567516688305e-11
GC_4_867 b_4 NI_4 NS_867 0 7.2835225399892603e-11
GC_4_868 b_4 NI_4 NS_868 0 -4.8050674542472472e-09
GC_4_869 b_4 NI_4 NS_869 0 -9.4069098050652565e-07
GC_4_870 b_4 NI_4 NS_870 0 -7.1603741521707283e-07
GC_4_871 b_4 NI_4 NS_871 0 6.8892096163021496e-07
GC_4_872 b_4 NI_4 NS_872 0 1.1980952475655529e-06
GC_4_873 b_4 NI_4 NS_873 0 -6.5943742966164001e-07
GC_4_874 b_4 NI_4 NS_874 0 2.7654889816197687e-06
GC_4_875 b_4 NI_4 NS_875 0 -1.7473351717887798e-07
GC_4_876 b_4 NI_4 NS_876 0 -8.3537242995095756e-07
GC_4_877 b_4 NI_4 NS_877 0 3.2530571481039231e-06
GC_4_878 b_4 NI_4 NS_878 0 -1.7278309909604032e-06
GC_4_879 b_4 NI_4 NS_879 0 -2.9824533064594189e-07
GC_4_880 b_4 NI_4 NS_880 0 1.3038473833593245e-06
GC_4_881 b_4 NI_4 NS_881 0 1.3780595232154013e-06
GC_4_882 b_4 NI_4 NS_882 0 1.3766292405800571e-06
GC_4_883 b_4 NI_4 NS_883 0 2.3900013322690102e-06
GC_4_884 b_4 NI_4 NS_884 0 -3.3970769595674545e-06
GC_4_885 b_4 NI_4 NS_885 0 -2.0889412560141029e-06
GC_4_886 b_4 NI_4 NS_886 0 -6.3013833259020671e-06
GC_4_887 b_4 NI_4 NS_887 0 -1.0350513882184442e-07
GC_4_888 b_4 NI_4 NS_888 0 5.0098931152009965e-07
GC_4_889 b_4 NI_4 NS_889 0 -1.2570127043446414e-05
GC_4_890 b_4 NI_4 NS_890 0 3.3150842392318616e-06
GC_4_891 b_4 NI_4 NS_891 0 -1.5284518285673819e-07
GC_4_892 b_4 NI_4 NS_892 0 -6.4577854279343673e-07
GC_4_893 b_4 NI_4 NS_893 0 3.1485875008649454e-06
GC_4_894 b_4 NI_4 NS_894 0 1.5222932790048137e-05
GC_4_895 b_4 NI_4 NS_895 0 1.0404489520255369e-06
GC_4_896 b_4 NI_4 NS_896 0 -1.0566938643505030e-06
GC_4_897 b_4 NI_4 NS_897 0 1.1263378529574475e-06
GC_4_898 b_4 NI_4 NS_898 0 -3.1753763308410403e-07
GC_4_899 b_4 NI_4 NS_899 0 6.6877942117200017e-06
GC_4_900 b_4 NI_4 NS_900 0 -3.1068911899304123e-06
GC_4_901 b_4 NI_4 NS_901 0 3.3131614549104895e-07
GC_4_902 b_4 NI_4 NS_902 0 3.9398701535424651e-07
GC_4_903 b_4 NI_4 NS_903 0 -2.9448268398966087e-06
GC_4_904 b_4 NI_4 NS_904 0 8.3451713458542790e-07
GC_4_905 b_4 NI_4 NS_905 0 1.7440840746061067e-07
GC_4_906 b_4 NI_4 NS_906 0 -8.8189850390054780e-07
GC_4_907 b_4 NI_4 NS_907 0 6.7930744833962582e-06
GC_4_908 b_4 NI_4 NS_908 0 3.5420987152920701e-06
GC_4_909 b_4 NI_4 NS_909 0 3.3691999519314830e-07
GC_4_910 b_4 NI_4 NS_910 0 8.5660422284961213e-09
GC_4_911 b_4 NI_4 NS_911 0 2.4534062214753655e-07
GC_4_912 b_4 NI_4 NS_912 0 -6.0596859457518641e-07
GC_4_913 b_4 NI_4 NS_913 0 3.9992419372327795e-07
GC_4_914 b_4 NI_4 NS_914 0 -1.3944049527412173e-06
GC_4_915 b_4 NI_4 NS_915 0 6.0125071777102377e-06
GC_4_916 b_4 NI_4 NS_916 0 -2.3492494179680421e-06
GC_4_917 b_4 NI_4 NS_917 0 2.3930279562620700e-08
GC_4_918 b_4 NI_4 NS_918 0 -2.5641169875372038e-07
GC_4_919 b_4 NI_4 NS_919 0 -9.3874761233081881e-07
GC_4_920 b_4 NI_4 NS_920 0 -1.1595548975984106e-06
GC_4_921 b_4 NI_4 NS_921 0 3.0874894676903450e-07
GC_4_922 b_4 NI_4 NS_922 0 -1.3340634186771026e-06
GC_4_923 b_4 NI_4 NS_923 0 3.0267241771448605e-06
GC_4_924 b_4 NI_4 NS_924 0 -4.1471321445646400e-06
GC_4_925 b_4 NI_4 NS_925 0 -1.7529086922029641e-07
GC_4_926 b_4 NI_4 NS_926 0 -3.4421193734291835e-07
GC_4_927 b_4 NI_4 NS_927 0 -1.9740564028270501e-06
GC_4_928 b_4 NI_4 NS_928 0 -6.6802046630289222e-07
GC_4_929 b_4 NI_4 NS_929 0 2.0794817930956727e-07
GC_4_930 b_4 NI_4 NS_930 0 -1.4268869549192797e-06
GC_4_931 b_4 NI_4 NS_931 0 9.1798302375271167e-08
GC_4_932 b_4 NI_4 NS_932 0 -3.5652572604445051e-06
GC_4_933 b_4 NI_4 NS_933 0 -4.5658114072864160e-07
GC_4_934 b_4 NI_4 NS_934 0 -3.7774913773830578e-07
GC_4_935 b_4 NI_4 NS_935 0 -2.1515201890565538e-06
GC_4_936 b_4 NI_4 NS_936 0 5.3521040599585412e-07
GC_4_937 b_4 NI_4 NS_937 0 -6.9312958551068174e-08
GC_4_938 b_4 NI_4 NS_938 0 -1.6158294067057565e-06
GC_4_939 b_4 NI_4 NS_939 0 -1.2654290843152699e-06
GC_4_940 b_4 NI_4 NS_940 0 -1.4064575387577185e-06
GC_4_941 b_4 NI_4 NS_941 0 -8.0808689204840966e-07
GC_4_942 b_4 NI_4 NS_942 0 9.5516005577720104e-08
GC_4_943 b_4 NI_4 NS_943 0 -9.4819654658998634e-07
GC_4_944 b_4 NI_4 NS_944 0 1.0893415376849940e-06
GC_4_945 b_4 NI_4 NS_945 0 -1.7800769069321416e-11
GC_4_946 b_4 NI_4 NS_946 0 1.0630963777700579e-11
GC_4_947 b_4 NI_4 NS_947 0 -5.7491710357202749e-07
GC_4_948 b_4 NI_4 NS_948 0 -1.1642133951151643e-06
GC_4_949 b_4 NI_4 NS_949 0 -3.7984302256871036e-07
GC_4_950 b_4 NI_4 NS_950 0 2.2312123541984687e-07
GC_4_951 b_4 NI_4 NS_951 0 -5.0935820818637061e-07
GC_4_952 b_4 NI_4 NS_952 0 3.9895582617836314e-07
GC_4_953 b_4 NI_4 NS_953 0 -1.9090303874476833e-07
GC_4_954 b_4 NI_4 NS_954 0 -1.0234021327292337e-06
GC_4_955 b_4 NI_4 NS_955 0 -4.4623499589194629e-07
GC_4_956 b_4 NI_4 NS_956 0 -2.0241835529338344e-07
GC_4_957 b_4 NI_4 NS_957 0 -9.1682537174289672e-10
GC_4_958 b_4 NI_4 NS_958 0 1.5482592843341583e-10
GC_4_959 b_4 NI_4 NS_959 0 -2.2810780228117700e-07
GC_4_960 b_4 NI_4 NS_960 0 -1.9852514227026701e-07
GC_4_961 b_4 NI_4 NS_961 0 -1.7941683102278825e-07
GC_4_962 b_4 NI_4 NS_962 0 -3.4649133068211604e-07
GC_4_963 b_4 NI_4 NS_963 0 -3.9554549994668822e-07
GC_4_964 b_4 NI_4 NS_964 0 -1.3729803224296584e-07
GC_4_965 b_4 NI_4 NS_965 0 -9.9086737000275319e-07
GC_4_966 b_4 NI_4 NS_966 0 5.0092585810630463e-08
GC_4_967 b_4 NI_4 NS_967 0 -5.8386569656609457e-07
GC_4_968 b_4 NI_4 NS_968 0 4.7577268793018504e-07
GC_4_969 b_4 NI_4 NS_969 0 -1.3073904613417549e-08
GC_4_970 b_4 NI_4 NS_970 0 4.1221603217133393e-07
GC_4_971 b_4 NI_4 NS_971 0 -8.6500709046588344e-07
GC_4_972 b_4 NI_4 NS_972 0 -9.7526648351566145e-07
GC_4_973 b_4 NI_4 NS_973 0 3.7776795408648213e-05
GC_4_974 b_4 NI_4 NS_974 0 1.2387413188554956e-12
GC_4_975 b_4 NI_4 NS_975 0 -8.1186813964375236e-12
GC_4_976 b_4 NI_4 NS_976 0 3.0025136893961746e-09
GC_4_977 b_4 NI_4 NS_977 0 3.6864096194820298e-07
GC_4_978 b_4 NI_4 NS_978 0 9.8384374040999766e-08
GC_4_979 b_4 NI_4 NS_979 0 6.5834108499363600e-07
GC_4_980 b_4 NI_4 NS_980 0 3.5826322847139055e-07
GC_4_981 b_4 NI_4 NS_981 0 1.2346444758001889e-06
GC_4_982 b_4 NI_4 NS_982 0 -8.6742584579019163e-07
GC_4_983 b_4 NI_4 NS_983 0 7.8270820209508065e-07
GC_4_984 b_4 NI_4 NS_984 0 -5.3020286248025818e-07
GC_4_985 b_4 NI_4 NS_985 0 8.2388487014267913e-07
GC_4_986 b_4 NI_4 NS_986 0 -2.1816060537801400e-06
GC_4_987 b_4 NI_4 NS_987 0 6.7227947773523825e-07
GC_4_988 b_4 NI_4 NS_988 0 -8.4321341330774050e-07
GC_4_989 b_4 NI_4 NS_989 0 -1.1291327276327577e-06
GC_4_990 b_4 NI_4 NS_990 0 -1.5078928913904593e-06
GC_4_991 b_4 NI_4 NS_991 0 -4.8950885583937881e-07
GC_4_992 b_4 NI_4 NS_992 0 -2.1010055379788596e-06
GC_4_993 b_4 NI_4 NS_993 0 -1.7840769101827864e-06
GC_4_994 b_4 NI_4 NS_994 0 -6.5666044581262571e-07
GC_4_995 b_4 NI_4 NS_995 0 -5.8884157266514735e-07
GC_4_996 b_4 NI_4 NS_996 0 -1.1663525150801964e-06
GC_4_997 b_4 NI_4 NS_997 0 -2.5818290690411881e-06
GC_4_998 b_4 NI_4 NS_998 0 -7.0827742407870420e-07
GC_4_999 b_4 NI_4 NS_999 0 -7.1488913509691582e-07
GC_4_1000 b_4 NI_4 NS_1000 0 -6.2489467249722050e-07
GC_4_1001 b_4 NI_4 NS_1001 0 -3.5725261224585766e-06
GC_4_1002 b_4 NI_4 NS_1002 0 -4.6960428513226054e-07
GC_4_1003 b_4 NI_4 NS_1003 0 2.3207021216132403e-07
GC_4_1004 b_4 NI_4 NS_1004 0 -2.1170865853287728e-07
GC_4_1005 b_4 NI_4 NS_1005 0 -9.1740994821439016e-07
GC_4_1006 b_4 NI_4 NS_1006 0 -9.0468419265576172e-07
GC_4_1007 b_4 NI_4 NS_1007 0 -1.9019681522001721e-06
GC_4_1008 b_4 NI_4 NS_1008 0 1.9079371730842782e-07
GC_4_1009 b_4 NI_4 NS_1009 0 -1.1727248604565507e-06
GC_4_1010 b_4 NI_4 NS_1010 0 -4.8228536068642879e-07
GC_4_1011 b_4 NI_4 NS_1011 0 -1.3189943529962266e-06
GC_4_1012 b_4 NI_4 NS_1012 0 9.6811830772631986e-07
GC_4_1013 b_4 NI_4 NS_1013 0 -7.9967652913991844e-07
GC_4_1014 b_4 NI_4 NS_1014 0 -4.7983612628878510e-07
GC_4_1015 b_4 NI_4 NS_1015 0 -3.1176929082812009e-06
GC_4_1016 b_4 NI_4 NS_1016 0 3.9714418083652692e-07
GC_4_1017 b_4 NI_4 NS_1017 0 -6.0262008628194347e-07
GC_4_1018 b_4 NI_4 NS_1018 0 1.6123614284049951e-07
GC_4_1019 b_4 NI_4 NS_1019 0 -6.6728210798391818e-07
GC_4_1020 b_4 NI_4 NS_1020 0 -1.5681802658974241e-07
GC_4_1021 b_4 NI_4 NS_1021 0 -1.3447997254328266e-06
GC_4_1022 b_4 NI_4 NS_1022 0 -7.5295239971009302e-08
GC_4_1023 b_4 NI_4 NS_1023 0 -3.0787565670071368e-06
GC_4_1024 b_4 NI_4 NS_1024 0 2.3443931989140608e-06
GC_4_1025 b_4 NI_4 NS_1025 0 -7.5438804173783701e-07
GC_4_1026 b_4 NI_4 NS_1026 0 3.5807956977346084e-07
GC_4_1027 b_4 NI_4 NS_1027 0 -8.0000261720679889e-07
GC_4_1028 b_4 NI_4 NS_1028 0 1.0728587023832996e-06
GC_4_1029 b_4 NI_4 NS_1029 0 -1.2382199160539569e-06
GC_4_1030 b_4 NI_4 NS_1030 0 1.6928091058958507e-07
GC_4_1031 b_4 NI_4 NS_1031 0 -1.0795275182692306e-06
GC_4_1032 b_4 NI_4 NS_1032 0 3.5773154919472768e-06
GC_4_1033 b_4 NI_4 NS_1033 0 -6.8450357193569094e-07
GC_4_1034 b_4 NI_4 NS_1034 0 4.6096044356220265e-07
GC_4_1035 b_4 NI_4 NS_1035 0 1.7787768101544438e-07
GC_4_1036 b_4 NI_4 NS_1036 0 1.4971787380896512e-06
GC_4_1037 b_4 NI_4 NS_1037 0 -1.1956615028030994e-06
GC_4_1038 b_4 NI_4 NS_1038 0 3.1705683238850231e-07
GC_4_1039 b_4 NI_4 NS_1039 0 9.5833849873155620e-07
GC_4_1040 b_4 NI_4 NS_1040 0 3.0173138592281795e-06
GC_4_1041 b_4 NI_4 NS_1041 0 -5.5639889058937207e-07
GC_4_1042 b_4 NI_4 NS_1042 0 6.1271390672560921e-07
GC_4_1043 b_4 NI_4 NS_1043 0 1.0073492164972070e-06
GC_4_1044 b_4 NI_4 NS_1044 0 8.4909697209418866e-07
GC_4_1045 b_4 NI_4 NS_1045 0 -1.1354681295249996e-06
GC_4_1046 b_4 NI_4 NS_1046 0 5.7364268067109195e-07
GC_4_1047 b_4 NI_4 NS_1047 0 1.7677957675825010e-06
GC_4_1048 b_4 NI_4 NS_1048 0 1.3974325712397891e-06
GC_4_1049 b_4 NI_4 NS_1049 0 -1.4090601651171649e-07
GC_4_1050 b_4 NI_4 NS_1050 0 6.5189401693343375e-07
GC_4_1051 b_4 NI_4 NS_1051 0 6.9857706290626552e-07
GC_4_1052 b_4 NI_4 NS_1052 0 -1.8042587816957940e-08
GC_4_1053 b_4 NI_4 NS_1053 0 2.1846689154877313e-11
GC_4_1054 b_4 NI_4 NS_1054 0 1.4146800150368978e-11
GC_4_1055 b_4 NI_4 NS_1055 0 -5.3445544311549725e-07
GC_4_1056 b_4 NI_4 NS_1056 0 6.6480542462743993e-07
GC_4_1057 b_4 NI_4 NS_1057 0 -1.6746246023394304e-08
GC_4_1058 b_4 NI_4 NS_1058 0 3.0212497585392171e-07
GC_4_1059 b_4 NI_4 NS_1059 0 2.1121846483217156e-07
GC_4_1060 b_4 NI_4 NS_1060 0 1.5832849794867022e-07
GC_4_1061 b_4 NI_4 NS_1061 0 -1.8419988079997154e-07
GC_4_1062 b_4 NI_4 NS_1062 0 5.6372901500620484e-07
GC_4_1063 b_4 NI_4 NS_1063 0 8.6158139571867219e-07
GC_4_1064 b_4 NI_4 NS_1064 0 4.0477759692772932e-07
GC_4_1065 b_4 NI_4 NS_1065 0 7.9125234611031185e-10
GC_4_1066 b_4 NI_4 NS_1066 0 5.1026693973273417e-10
GC_4_1067 b_4 NI_4 NS_1067 0 1.2590892390583516e-06
GC_4_1068 b_4 NI_4 NS_1068 0 1.3277674221216033e-07
GC_4_1069 b_4 NI_4 NS_1069 0 -1.4104382023288224e-07
GC_4_1070 b_4 NI_4 NS_1070 0 8.3427633851329014e-07
GC_4_1071 b_4 NI_4 NS_1071 0 8.2109247535414205e-08
GC_4_1072 b_4 NI_4 NS_1072 0 4.1437502332551882e-08
GC_4_1073 b_4 NI_4 NS_1073 0 3.4449293024734000e-07
GC_4_1074 b_4 NI_4 NS_1074 0 3.3674005947123369e-07
GC_4_1075 b_4 NI_4 NS_1075 0 3.0905305969895095e-07
GC_4_1076 b_4 NI_4 NS_1076 0 4.0930284728893024e-07
GC_4_1077 b_4 NI_4 NS_1077 0 6.5356222967029092e-08
GC_4_1078 b_4 NI_4 NS_1078 0 5.9259710059430064e-08
GC_4_1079 b_4 NI_4 NS_1079 0 7.1106409178642460e-07
GC_4_1080 b_4 NI_4 NS_1080 0 8.9929453789909169e-07
GC_4_1081 b_4 NI_4 NS_1081 0 -6.4297371565516851e-05
GC_4_1082 b_4 NI_4 NS_1082 0 3.5514087114614693e-12
GC_4_1083 b_4 NI_4 NS_1083 0 5.0206447902918256e-11
GC_4_1084 b_4 NI_4 NS_1084 0 -1.5827700559032664e-09
GC_4_1085 b_4 NI_4 NS_1085 0 -1.0722887952863219e-06
GC_4_1086 b_4 NI_4 NS_1086 0 -1.0608550085816174e-06
GC_4_1087 b_4 NI_4 NS_1087 0 4.1036420206254637e-07
GC_4_1088 b_4 NI_4 NS_1088 0 3.5893460006623391e-07
GC_4_1089 b_4 NI_4 NS_1089 0 -2.2645998652798010e-06
GC_4_1090 b_4 NI_4 NS_1090 0 2.1075672924155170e-06
GC_4_1091 b_4 NI_4 NS_1091 0 -2.5340369455752492e-06
GC_4_1092 b_4 NI_4 NS_1092 0 -1.2433598111408819e-06
GC_4_1093 b_4 NI_4 NS_1093 0 1.3996047064213742e-06
GC_4_1094 b_4 NI_4 NS_1094 0 1.0022276631129546e-06
GC_4_1095 b_4 NI_4 NS_1095 0 -1.1248387970601809e-06
GC_4_1096 b_4 NI_4 NS_1096 0 1.3421363583486184e-06
GC_4_1097 b_4 NI_4 NS_1097 0 7.2530386736199405e-07
GC_4_1098 b_4 NI_4 NS_1098 0 3.0434992989625940e-06
GC_4_1099 b_4 NI_4 NS_1099 0 -2.8542607341886139e-06
GC_4_1100 b_4 NI_4 NS_1100 0 4.6955374882228885e-07
GC_4_1101 b_4 NI_4 NS_1101 0 3.6961799999206065e-06
GC_4_1102 b_4 NI_4 NS_1102 0 -2.0129312763040804e-06
GC_4_1103 b_4 NI_4 NS_1103 0 -1.9022277173228729e-07
GC_4_1104 b_4 NI_4 NS_1104 0 2.5688425481254821e-06
GC_4_1105 b_4 NI_4 NS_1105 0 -4.0608181929865969e-06
GC_4_1106 b_4 NI_4 NS_1106 0 4.8419384513215490e-06
GC_4_1107 b_4 NI_4 NS_1107 0 6.4547440780623923e-07
GC_4_1108 b_4 NI_4 NS_1108 0 -1.5900968484356856e-06
GC_4_1109 b_4 NI_4 NS_1109 0 4.6199468493712092e-06
GC_4_1110 b_4 NI_4 NS_1110 0 9.9424796524959636e-06
GC_4_1111 b_4 NI_4 NS_1111 0 -1.1565186269010674e-07
GC_4_1112 b_4 NI_4 NS_1112 0 5.2802063184841239e-07
GC_4_1113 b_4 NI_4 NS_1113 0 -6.9401161795082252e-09
GC_4_1114 b_4 NI_4 NS_1114 0 -7.8937763321376929e-07
GC_4_1115 b_4 NI_4 NS_1115 0 5.3542099454672398e-06
GC_4_1116 b_4 NI_4 NS_1116 0 4.9603705099770733e-07
GC_4_1117 b_4 NI_4 NS_1117 0 8.4754028904234389e-07
GC_4_1118 b_4 NI_4 NS_1118 0 1.9215377299852587e-06
GC_4_1119 b_4 NI_4 NS_1119 0 3.1612345903537793e-08
GC_4_1120 b_4 NI_4 NS_1120 0 1.1340680038340760e-06
GC_4_1121 b_4 NI_4 NS_1121 0 5.8568536317226121e-07
GC_4_1122 b_4 NI_4 NS_1122 0 -1.1142478322993033e-06
GC_4_1123 b_4 NI_4 NS_1123 0 5.8308429628669644e-06
GC_4_1124 b_4 NI_4 NS_1124 0 4.0738907110413064e-06
GC_4_1125 b_4 NI_4 NS_1125 0 6.0565470961144218e-07
GC_4_1126 b_4 NI_4 NS_1126 0 8.6242515345106142e-07
GC_4_1127 b_4 NI_4 NS_1127 0 1.9671091653058639e-07
GC_4_1128 b_4 NI_4 NS_1128 0 2.4105028168502230e-07
GC_4_1129 b_4 NI_4 NS_1129 0 8.4506367117109229e-07
GC_4_1130 b_4 NI_4 NS_1130 0 -6.7479248817862511e-07
GC_4_1131 b_4 NI_4 NS_1131 0 6.6692216197498819e-06
GC_4_1132 b_4 NI_4 NS_1132 0 7.5284376018501332e-07
GC_4_1133 b_4 NI_4 NS_1133 0 7.7512903406051550e-07
GC_4_1134 b_4 NI_4 NS_1134 0 7.5176299682890334e-07
GC_4_1135 b_4 NI_4 NS_1135 0 6.6484739796768046e-07
GC_4_1136 b_4 NI_4 NS_1136 0 -6.6049843280993862e-08
GC_4_1137 b_4 NI_4 NS_1137 0 8.7116464100625701e-07
GC_4_1138 b_4 NI_4 NS_1138 0 -6.4327917624388387e-07
GC_4_1139 b_4 NI_4 NS_1139 0 5.7782990046480806e-06
GC_4_1140 b_4 NI_4 NS_1140 0 -1.5930662829621499e-06
GC_4_1141 b_4 NI_4 NS_1141 0 8.2495579086625750e-07
GC_4_1142 b_4 NI_4 NS_1142 0 5.6931882879638832e-07
GC_4_1143 b_4 NI_4 NS_1143 0 6.2572122827219460e-07
GC_4_1144 b_4 NI_4 NS_1144 0 -5.5367418889514617e-07
GC_4_1145 b_4 NI_4 NS_1145 0 9.3725569699543907e-07
GC_4_1146 b_4 NI_4 NS_1146 0 -4.4873086326904109e-07
GC_4_1147 b_4 NI_4 NS_1147 0 3.9054872685110617e-06
GC_4_1148 b_4 NI_4 NS_1148 0 -2.9926171579729578e-06
GC_4_1149 b_4 NI_4 NS_1149 0 8.9723919541415289e-07
GC_4_1150 b_4 NI_4 NS_1150 0 3.2914617558044299e-07
GC_4_1151 b_4 NI_4 NS_1151 0 2.1534160440611062e-07
GC_4_1152 b_4 NI_4 NS_1152 0 -7.9633296115262362e-07
GC_4_1153 b_4 NI_4 NS_1153 0 1.1591892462855251e-06
GC_4_1154 b_4 NI_4 NS_1154 0 -3.2770153225568717e-07
GC_4_1155 b_4 NI_4 NS_1155 0 1.6782780586904946e-06
GC_4_1156 b_4 NI_4 NS_1156 0 -3.0911800886172362e-06
GC_4_1157 b_4 NI_4 NS_1157 0 7.9264100179165172e-07
GC_4_1158 b_4 NI_4 NS_1158 0 -1.0570297005218432e-07
GC_4_1159 b_4 NI_4 NS_1159 0 -1.9831591654114373e-07
GC_4_1160 b_4 NI_4 NS_1160 0 -4.0880811566481018e-07
GC_4_1161 b_4 NI_4 NS_1161 0 8.5889532986776189e-12
GC_4_1162 b_4 NI_4 NS_1162 0 -1.5739918258876974e-11
GC_4_1163 b_4 NI_4 NS_1163 0 8.3767146195560125e-07
GC_4_1164 b_4 NI_4 NS_1164 0 -5.9584797896411487e-07
GC_4_1165 b_4 NI_4 NS_1165 0 4.9537049655227477e-07
GC_4_1166 b_4 NI_4 NS_1166 0 -3.5566029171648482e-08
GC_4_1167 b_4 NI_4 NS_1167 0 1.6373891567663647e-08
GC_4_1168 b_4 NI_4 NS_1168 0 -8.9211328734574000e-08
GC_4_1169 b_4 NI_4 NS_1169 0 5.2071322385616317e-07
GC_4_1170 b_4 NI_4 NS_1170 0 -1.9285955239511106e-08
GC_4_1171 b_4 NI_4 NS_1171 0 7.0590856987879271e-07
GC_4_1172 b_4 NI_4 NS_1172 0 -1.5618081720456326e-06
GC_4_1173 b_4 NI_4 NS_1173 0 4.0957995068931890e-10
GC_4_1174 b_4 NI_4 NS_1174 0 -5.8094794254692826e-10
GC_4_1175 b_4 NI_4 NS_1175 0 1.0094269047470102e-06
GC_4_1176 b_4 NI_4 NS_1176 0 -2.7418463270180809e-07
GC_4_1177 b_4 NI_4 NS_1177 0 3.5391611156943077e-07
GC_4_1178 b_4 NI_4 NS_1178 0 -1.7487840651139988e-07
GC_4_1179 b_4 NI_4 NS_1179 0 2.5449991651368490e-07
GC_4_1180 b_4 NI_4 NS_1180 0 2.6674179513330830e-08
GC_4_1181 b_4 NI_4 NS_1181 0 1.0861112780627123e-06
GC_4_1182 b_4 NI_4 NS_1182 0 -1.1751131198194532e-06
GC_4_1183 b_4 NI_4 NS_1183 0 6.5444283849452822e-07
GC_4_1184 b_4 NI_4 NS_1184 0 -3.3449113832749875e-07
GC_4_1185 b_4 NI_4 NS_1185 0 -2.1289903082637366e-07
GC_4_1186 b_4 NI_4 NS_1186 0 -9.8626030054703732e-08
GC_4_1187 b_4 NI_4 NS_1187 0 7.5675695348973922e-07
GC_4_1188 b_4 NI_4 NS_1188 0 3.2207291425898510e-07
GC_4_1189 b_4 NI_4 NS_1189 0 8.5535251026678356e-06
GC_4_1190 b_4 NI_4 NS_1190 0 3.7642345460060006e-12
GC_4_1191 b_4 NI_4 NS_1191 0 -7.8551955575354626e-11
GC_4_1192 b_4 NI_4 NS_1192 0 2.5470430419923847e-09
GC_4_1193 b_4 NI_4 NS_1193 0 1.5926560601238302e-08
GC_4_1194 b_4 NI_4 NS_1194 0 -8.5340749401516645e-08
GC_4_1195 b_4 NI_4 NS_1195 0 -2.5044505624780498e-07
GC_4_1196 b_4 NI_4 NS_1196 0 2.6988969668559641e-07
GC_4_1197 b_4 NI_4 NS_1197 0 7.4472042717052957e-07
GC_4_1198 b_4 NI_4 NS_1198 0 -2.8257741925226350e-07
GC_4_1199 b_4 NI_4 NS_1199 0 -9.7076242329732492e-07
GC_4_1200 b_4 NI_4 NS_1200 0 -2.4180542177669113e-07
GC_4_1201 b_4 NI_4 NS_1201 0 1.0253000992931598e-06
GC_4_1202 b_4 NI_4 NS_1202 0 4.0598757009057696e-07
GC_4_1203 b_4 NI_4 NS_1203 0 -1.2043560723680874e-07
GC_4_1204 b_4 NI_4 NS_1204 0 -2.7435484755036492e-07
GC_4_1205 b_4 NI_4 NS_1205 0 1.1179344555102048e-07
GC_4_1206 b_4 NI_4 NS_1206 0 -5.1154211381903626e-07
GC_4_1207 b_4 NI_4 NS_1207 0 -2.0930621906035442e-06
GC_4_1208 b_4 NI_4 NS_1208 0 8.5810281787891552e-07
GC_4_1209 b_4 NI_4 NS_1209 0 2.4408886836524368e-06
GC_4_1210 b_4 NI_4 NS_1210 0 -5.9923555031653962e-07
GC_4_1211 b_4 NI_4 NS_1211 0 -6.6143704298275498e-07
GC_4_1212 b_4 NI_4 NS_1212 0 -1.4026137541655285e-06
GC_4_1213 b_4 NI_4 NS_1213 0 4.2548612107271359e-07
GC_4_1214 b_4 NI_4 NS_1214 0 1.8523053157468170e-06
GC_4_1215 b_4 NI_4 NS_1215 0 -2.7461843382734932e-08
GC_4_1216 b_4 NI_4 NS_1216 0 -1.3270320182956243e-06
GC_4_1217 b_4 NI_4 NS_1217 0 -6.3828670893419905e-07
GC_4_1218 b_4 NI_4 NS_1218 0 2.5986444830823258e-06
GC_4_1219 b_4 NI_4 NS_1219 0 4.5949660453535412e-07
GC_4_1220 b_4 NI_4 NS_1220 0 -2.2490727431925790e-06
GC_4_1221 b_4 NI_4 NS_1221 0 -8.0030287442929613e-07
GC_4_1222 b_4 NI_4 NS_1222 0 -9.3521755342913346e-07
GC_4_1223 b_4 NI_4 NS_1223 0 3.5980080130334052e-07
GC_4_1224 b_4 NI_4 NS_1224 0 9.1582450105394131e-07
GC_4_1225 b_4 NI_4 NS_1225 0 -5.5704122503349969e-07
GC_4_1226 b_4 NI_4 NS_1226 0 -7.2806113486252826e-07
GC_4_1227 b_4 NI_4 NS_1227 0 4.7834214323502626e-07
GC_4_1228 b_4 NI_4 NS_1228 0 7.4258410350247088e-07
GC_4_1229 b_4 NI_4 NS_1229 0 -1.7303766408728006e-07
GC_4_1230 b_4 NI_4 NS_1230 0 -8.8058541102887080e-07
GC_4_1231 b_4 NI_4 NS_1231 0 -3.3837653935993440e-07
GC_4_1232 b_4 NI_4 NS_1232 0 1.1624993516186430e-06
GC_4_1233 b_4 NI_4 NS_1233 0 2.5595331832502341e-07
GC_4_1234 b_4 NI_4 NS_1234 0 -8.4667910970690395e-07
GC_4_1235 b_4 NI_4 NS_1235 0 -6.4574651828145964e-08
GC_4_1236 b_4 NI_4 NS_1236 0 6.7761767230176621e-08
GC_4_1237 b_4 NI_4 NS_1237 0 -2.5919661646746070e-07
GC_4_1238 b_4 NI_4 NS_1238 0 -5.5152737422571217e-07
GC_4_1239 b_4 NI_4 NS_1239 0 1.8905503552331134e-07
GC_4_1240 b_4 NI_4 NS_1240 0 7.1901979693733687e-07
GC_4_1241 b_4 NI_4 NS_1241 0 -7.9602463118558724e-08
GC_4_1242 b_4 NI_4 NS_1242 0 -6.3772382306005291e-07
GC_4_1243 b_4 NI_4 NS_1243 0 1.0329815149581191e-07
GC_4_1244 b_4 NI_4 NS_1244 0 1.0426217753384269e-07
GC_4_1245 b_4 NI_4 NS_1245 0 -2.9062604459995502e-07
GC_4_1246 b_4 NI_4 NS_1246 0 -5.9569098033170643e-07
GC_4_1247 b_4 NI_4 NS_1247 0 1.6437698423303590e-07
GC_4_1248 b_4 NI_4 NS_1248 0 2.3048467726322929e-07
GC_4_1249 b_4 NI_4 NS_1249 0 -2.5683223043557350e-07
GC_4_1250 b_4 NI_4 NS_1250 0 -5.1013999720247193e-07
GC_4_1251 b_4 NI_4 NS_1251 0 4.9680099074328062e-08
GC_4_1252 b_4 NI_4 NS_1252 0 -5.0624163818209845e-08
GC_4_1253 b_4 NI_4 NS_1253 0 -3.6842305759398856e-07
GC_4_1254 b_4 NI_4 NS_1254 0 -5.6019338899945853e-07
GC_4_1255 b_4 NI_4 NS_1255 0 -2.3359372199038320e-07
GC_4_1256 b_4 NI_4 NS_1256 0 2.0119127649467396e-08
GC_4_1257 b_4 NI_4 NS_1257 0 -4.3463047173879170e-07
GC_4_1258 b_4 NI_4 NS_1258 0 -3.4260334924896520e-07
GC_4_1259 b_4 NI_4 NS_1259 0 -1.2394309247658259e-07
GC_4_1260 b_4 NI_4 NS_1260 0 1.6157692594390511e-08
GC_4_1261 b_4 NI_4 NS_1261 0 -5.6455863448733907e-07
GC_4_1262 b_4 NI_4 NS_1262 0 -4.4144307534123278e-07
GC_4_1263 b_4 NI_4 NS_1263 0 -3.1825758914346598e-07
GC_4_1264 b_4 NI_4 NS_1264 0 3.1675260939157244e-07
GC_4_1265 b_4 NI_4 NS_1265 0 -5.0108244255899548e-07
GC_4_1266 b_4 NI_4 NS_1266 0 3.6711580977003923e-08
GC_4_1267 b_4 NI_4 NS_1267 0 -1.0041276180611355e-08
GC_4_1268 b_4 NI_4 NS_1268 0 6.2080292532669981e-08
GC_4_1269 b_4 NI_4 NS_1269 0 -3.2608739409704240e-12
GC_4_1270 b_4 NI_4 NS_1270 0 3.1978332660848790e-12
GC_4_1271 b_4 NI_4 NS_1271 0 -5.7750182669162827e-07
GC_4_1272 b_4 NI_4 NS_1272 0 4.5921422231565011e-08
GC_4_1273 b_4 NI_4 NS_1273 0 -2.9018151337931570e-07
GC_4_1274 b_4 NI_4 NS_1274 0 1.1752550807071822e-07
GC_4_1275 b_4 NI_4 NS_1275 0 -5.6679600787596550e-09
GC_4_1276 b_4 NI_4 NS_1276 0 -6.8755103531708997e-08
GC_4_1277 b_4 NI_4 NS_1277 0 -6.6097126813590386e-07
GC_4_1278 b_4 NI_4 NS_1278 0 1.3969832672648536e-07
GC_4_1279 b_4 NI_4 NS_1279 0 2.9822753982354771e-08
GC_4_1280 b_4 NI_4 NS_1280 0 1.2499661750050685e-07
GC_4_1281 b_4 NI_4 NS_1281 0 -6.1662769042760649e-11
GC_4_1282 b_4 NI_4 NS_1282 0 1.2835945134397911e-10
GC_4_1283 b_4 NI_4 NS_1283 0 -3.4930435154169624e-08
GC_4_1284 b_4 NI_4 NS_1284 0 1.9717730284276584e-07
GC_4_1285 b_4 NI_4 NS_1285 0 -3.6700057485093794e-07
GC_4_1286 b_4 NI_4 NS_1286 0 -4.4689542768180213e-08
GC_4_1287 b_4 NI_4 NS_1287 0 -1.8607415866796081e-07
GC_4_1288 b_4 NI_4 NS_1288 0 -2.7291718937873618e-09
GC_4_1289 b_4 NI_4 NS_1289 0 1.9304457199515219e-07
GC_4_1290 b_4 NI_4 NS_1290 0 8.1847819164777949e-08
GC_4_1291 b_4 NI_4 NS_1291 0 -2.6597636016480522e-07
GC_4_1292 b_4 NI_4 NS_1292 0 3.1322701882741062e-07
GC_4_1293 b_4 NI_4 NS_1293 0 1.2554900436318668e-07
GC_4_1294 b_4 NI_4 NS_1294 0 -1.4412635641479203e-07
GC_4_1295 b_4 NI_4 NS_1295 0 -5.8147438627903279e-08
GC_4_1296 b_4 NI_4 NS_1296 0 2.3784873689179144e-07
GD_4_1 b_4 NI_4 NA_1 0 -1.1524177909361349e-03
GD_4_2 b_4 NI_4 NA_2 0 1.0616253484660441e-02
GD_4_3 b_4 NI_4 NA_3 0 -5.0003083239244838e-03
GD_4_4 b_4 NI_4 NA_4 0 -1.0894627888821886e-02
GD_4_5 b_4 NI_4 NA_5 0 1.0511509928807459e-04
GD_4_6 b_4 NI_4 NA_6 0 2.2219404053217939e-05
GD_4_7 b_4 NI_4 NA_7 0 1.6003148970072700e-05
GD_4_8 b_4 NI_4 NA_8 0 -6.7345471873276455e-07
GD_4_9 b_4 NI_4 NA_9 0 2.0977582185156723e-06
GD_4_10 b_4 NI_4 NA_10 0 -7.3787541409576805e-06
GD_4_11 b_4 NI_4 NA_11 0 8.8115123730307144e-06
GD_4_12 b_4 NI_4 NA_12 0 -1.1565256116698626e-06
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 -5.3680129526507305e-05
GC_5_2 b_5 NI_5 NS_2 0 -6.9833821954368458e-12
GC_5_3 b_5 NI_5 NS_3 0 -2.0805248769436771e-10
GC_5_4 b_5 NI_5 NS_4 0 9.8195269669862864e-09
GC_5_5 b_5 NI_5 NS_5 0 5.4711434452171201e-07
GC_5_6 b_5 NI_5 NS_6 0 4.2979795426208142e-08
GC_5_7 b_5 NI_5 NS_7 0 2.9239405765226281e-06
GC_5_8 b_5 NI_5 NS_8 0 -1.5091400525384371e-06
GC_5_9 b_5 NI_5 NS_9 0 -3.2045433958834257e-06
GC_5_10 b_5 NI_5 NS_10 0 -2.6196626924306725e-06
GC_5_11 b_5 NI_5 NS_11 0 4.6037988169203621e-06
GC_5_12 b_5 NI_5 NS_12 0 -4.0622264345346639e-07
GC_5_13 b_5 NI_5 NS_13 0 -7.4630326170180541e-06
GC_5_14 b_5 NI_5 NS_14 0 -7.5110674502945018e-06
GC_5_15 b_5 NI_5 NS_15 0 -2.6104519385237572e-07
GC_5_16 b_5 NI_5 NS_16 0 -1.3674927512381009e-06
GC_5_17 b_5 NI_5 NS_17 0 -5.9022061872817237e-06
GC_5_18 b_5 NI_5 NS_18 0 2.4898529331520114e-06
GC_5_19 b_5 NI_5 NS_19 0 5.2248128967619118e-06
GC_5_20 b_5 NI_5 NS_20 0 -5.0757034246097503e-06
GC_5_21 b_5 NI_5 NS_21 0 -1.6698151594636138e-05
GC_5_22 b_5 NI_5 NS_22 0 5.0787239778674043e-06
GC_5_23 b_5 NI_5 NS_23 0 -1.1561010181961655e-06
GC_5_24 b_5 NI_5 NS_24 0 7.5339642023526788e-06
GC_5_25 b_5 NI_5 NS_25 0 -6.6315705947812177e-06
GC_5_26 b_5 NI_5 NS_26 0 -4.0455597904254603e-06
GC_5_27 b_5 NI_5 NS_27 0 -3.2762114331238810e-06
GC_5_28 b_5 NI_5 NS_28 0 8.3571837732236706e-06
GC_5_29 b_5 NI_5 NS_29 0 -1.2997338688599877e-06
GC_5_30 b_5 NI_5 NS_30 0 -4.1162262108627993e-06
GC_5_31 b_5 NI_5 NS_31 0 -4.0024790282590336e-06
GC_5_32 b_5 NI_5 NS_32 0 1.1510740169044306e-05
GC_5_33 b_5 NI_5 NS_33 0 -2.4919345408249360e-08
GC_5_34 b_5 NI_5 NS_34 0 7.6861978975891924e-06
GC_5_35 b_5 NI_5 NS_35 0 -3.6434501054284942e-06
GC_5_36 b_5 NI_5 NS_36 0 1.4544318657644410e-06
GC_5_37 b_5 NI_5 NS_37 0 -3.5977796128677399e-07
GC_5_38 b_5 NI_5 NS_38 0 8.4286793072373902e-06
GC_5_39 b_5 NI_5 NS_39 0 -5.7518759418532002e-07
GC_5_40 b_5 NI_5 NS_40 0 2.1383299906348521e-06
GC_5_41 b_5 NI_5 NS_41 0 -2.3055742948009431e-06
GC_5_42 b_5 NI_5 NS_42 0 8.5102688271103796e-06
GC_5_43 b_5 NI_5 NS_43 0 7.1416267639705601e-07
GC_5_44 b_5 NI_5 NS_44 0 9.9220593592789660e-06
GC_5_45 b_5 NI_5 NS_45 0 -7.2144983203847427e-07
GC_5_46 b_5 NI_5 NS_46 0 8.9744372490638018e-06
GC_5_47 b_5 NI_5 NS_47 0 -1.2319738384149936e-06
GC_5_48 b_5 NI_5 NS_48 0 4.0766587113877439e-06
GC_5_49 b_5 NI_5 NS_49 0 1.2869277814799517e-06
GC_5_50 b_5 NI_5 NS_50 0 1.2351987567679139e-05
GC_5_51 b_5 NI_5 NS_51 0 1.8775556306236546e-05
GC_5_52 b_5 NI_5 NS_52 0 1.7032810916265126e-05
GC_5_53 b_5 NI_5 NS_53 0 5.0360268121533528e-06
GC_5_54 b_5 NI_5 NS_54 0 7.9043932325098961e-06
GC_5_55 b_5 NI_5 NS_55 0 1.0383334282888344e-05
GC_5_56 b_5 NI_5 NS_56 0 3.9003795528834498e-06
GC_5_57 b_5 NI_5 NS_57 0 6.8650995533498688e-06
GC_5_58 b_5 NI_5 NS_58 0 1.1089491143073741e-05
GC_5_59 b_5 NI_5 NS_59 0 3.3649742406185243e-05
GC_5_60 b_5 NI_5 NS_60 0 -6.1820210984330019e-06
GC_5_61 b_5 NI_5 NS_61 0 8.2297383182382039e-06
GC_5_62 b_5 NI_5 NS_62 0 3.4992006896258732e-06
GC_5_63 b_5 NI_5 NS_63 0 1.2051429772545331e-05
GC_5_64 b_5 NI_5 NS_64 0 -1.0349766034369781e-05
GC_5_65 b_5 NI_5 NS_65 0 1.0852241711164685e-05
GC_5_66 b_5 NI_5 NS_66 0 6.5921148528310469e-06
GC_5_67 b_5 NI_5 NS_67 0 1.7121436669823338e-05
GC_5_68 b_5 NI_5 NS_68 0 -3.0976642769810694e-05
GC_5_69 b_5 NI_5 NS_69 0 8.1822973300010053e-06
GC_5_70 b_5 NI_5 NS_70 0 -2.9067682434294393e-06
GC_5_71 b_5 NI_5 NS_71 0 -3.1851363784286997e-06
GC_5_72 b_5 NI_5 NS_72 0 -1.6366048166865836e-05
GC_5_73 b_5 NI_5 NS_73 0 1.1873638821207866e-05
GC_5_74 b_5 NI_5 NS_74 0 -1.5391800502810433e-06
GC_5_75 b_5 NI_5 NS_75 0 -1.2633532485136995e-05
GC_5_76 b_5 NI_5 NS_76 0 -2.5267039597519969e-05
GC_5_77 b_5 NI_5 NS_77 0 -1.0375386706889778e-07
GC_5_78 b_5 NI_5 NS_78 0 -6.6315508036872661e-06
GC_5_79 b_5 NI_5 NS_79 0 -9.5776936856794514e-06
GC_5_80 b_5 NI_5 NS_80 0 -2.6846435069995723e-06
GC_5_81 b_5 NI_5 NS_81 0 1.0229009790565136e-10
GC_5_82 b_5 NI_5 NS_82 0 4.5737902425820546e-11
GC_5_83 b_5 NI_5 NS_83 0 1.5527383944617813e-06
GC_5_84 b_5 NI_5 NS_84 0 -4.6900204114156573e-06
GC_5_85 b_5 NI_5 NS_85 0 -1.3369745545032063e-06
GC_5_86 b_5 NI_5 NS_86 0 -1.3619261726067078e-06
GC_5_87 b_5 NI_5 NS_87 0 -4.8411291129694053e-06
GC_5_88 b_5 NI_5 NS_88 0 -1.0239409184712528e-06
GC_5_89 b_5 NI_5 NS_89 0 -1.0645242413161073e-06
GC_5_90 b_5 NI_5 NS_90 0 -2.7299683602199877e-06
GC_5_91 b_5 NI_5 NS_91 0 -9.9885536925315942e-06
GC_5_92 b_5 NI_5 NS_92 0 -4.1154650085584920e-06
GC_5_93 b_5 NI_5 NS_93 0 6.6961072962745583e-09
GC_5_94 b_5 NI_5 NS_94 0 5.4062569618574502e-09
GC_5_95 b_5 NI_5 NS_95 0 1.7786609774380774e-06
GC_5_96 b_5 NI_5 NS_96 0 4.4250649018771524e-07
GC_5_97 b_5 NI_5 NS_97 0 -1.5845646268569676e-06
GC_5_98 b_5 NI_5 NS_98 0 3.2301030652529907e-06
GC_5_99 b_5 NI_5 NS_99 0 -8.2746730852375775e-07
GC_5_100 b_5 NI_5 NS_100 0 6.9450325756867244e-07
GC_5_101 b_5 NI_5 NS_101 0 -7.6658753291285927e-06
GC_5_102 b_5 NI_5 NS_102 0 4.7706505573280084e-07
GC_5_103 b_5 NI_5 NS_103 0 -2.2026813030470147e-06
GC_5_104 b_5 NI_5 NS_104 0 1.9565060225806608e-06
GC_5_105 b_5 NI_5 NS_105 0 -2.0865320009819402e-06
GC_5_106 b_5 NI_5 NS_106 0 1.9644981953767161e-06
GC_5_107 b_5 NI_5 NS_107 0 1.2958343286312508e-06
GC_5_108 b_5 NI_5 NS_108 0 2.8412086672532440e-06
GC_5_109 b_5 NI_5 NS_109 0 -1.5264422047903155e-04
GC_5_110 b_5 NI_5 NS_110 0 3.6649137353162220e-11
GC_5_111 b_5 NI_5 NS_111 0 1.8928535655547295e-11
GC_5_112 b_5 NI_5 NS_112 0 9.3054203097794671e-10
GC_5_113 b_5 NI_5 NS_113 0 -2.3228677220503136e-06
GC_5_114 b_5 NI_5 NS_114 0 -1.6428458717770513e-06
GC_5_115 b_5 NI_5 NS_115 0 1.4316064842889543e-06
GC_5_116 b_5 NI_5 NS_116 0 3.8987538068458981e-06
GC_5_117 b_5 NI_5 NS_117 0 3.0058959463940692e-06
GC_5_118 b_5 NI_5 NS_118 0 5.4030099742622810e-06
GC_5_119 b_5 NI_5 NS_119 0 5.4598831850726664e-06
GC_5_120 b_5 NI_5 NS_120 0 -8.4815313466336340e-06
GC_5_121 b_5 NI_5 NS_121 0 -2.3142976671272668e-06
GC_5_122 b_5 NI_5 NS_122 0 -1.2723712100652006e-05
GC_5_123 b_5 NI_5 NS_123 0 -3.7422796653128973e-06
GC_5_124 b_5 NI_5 NS_124 0 2.7239303112661160e-06
GC_5_125 b_5 NI_5 NS_125 0 4.5151411605317008e-06
GC_5_126 b_5 NI_5 NS_126 0 1.5308235720148332e-06
GC_5_127 b_5 NI_5 NS_127 0 8.7547077471954067e-06
GC_5_128 b_5 NI_5 NS_128 0 -3.8479491722355212e-05
GC_5_129 b_5 NI_5 NS_129 0 -4.3264676081735339e-05
GC_5_130 b_5 NI_5 NS_130 0 -1.4454839590956339e-06
GC_5_131 b_5 NI_5 NS_131 0 -1.4749716077453832e-05
GC_5_132 b_5 NI_5 NS_132 0 -8.4842962341677641e-06
GC_5_133 b_5 NI_5 NS_133 0 -7.0816465142272458e-05
GC_5_134 b_5 NI_5 NS_134 0 7.5582589814833227e-05
GC_5_135 b_5 NI_5 NS_135 0 4.8530268041117052e-06
GC_5_136 b_5 NI_5 NS_136 0 1.3247864620256898e-05
GC_5_137 b_5 NI_5 NS_137 0 6.5374364333054382e-05
GC_5_138 b_5 NI_5 NS_138 0 1.2308041375876515e-04
GC_5_139 b_5 NI_5 NS_139 0 -1.3621976358942521e-07
GC_5_140 b_5 NI_5 NS_140 0 -3.7823805209160376e-05
GC_5_141 b_5 NI_5 NS_141 0 1.6963590041203515e-05
GC_5_142 b_5 NI_5 NS_142 0 4.3619926062420418e-06
GC_5_143 b_5 NI_5 NS_143 0 2.5306791387095624e-05
GC_5_144 b_5 NI_5 NS_144 0 -3.1224056754734523e-05
GC_5_145 b_5 NI_5 NS_145 0 -8.6239867171775490e-06
GC_5_146 b_5 NI_5 NS_146 0 -2.7323224727029034e-06
GC_5_147 b_5 NI_5 NS_147 0 -8.1953080524118284e-06
GC_5_148 b_5 NI_5 NS_148 0 2.4464546783607928e-05
GC_5_149 b_5 NI_5 NS_149 0 6.0407833711090298e-06
GC_5_150 b_5 NI_5 NS_150 0 8.5945632963172084e-06
GC_5_151 b_5 NI_5 NS_151 0 5.7640723383354862e-05
GC_5_152 b_5 NI_5 NS_152 0 2.4091616569992172e-05
GC_5_153 b_5 NI_5 NS_153 0 3.6450300557564802e-06
GC_5_154 b_5 NI_5 NS_154 0 -1.2427359937450567e-05
GC_5_155 b_5 NI_5 NS_155 0 -7.2831135218646188e-08
GC_5_156 b_5 NI_5 NS_156 0 -1.3777686779702281e-06
GC_5_157 b_5 NI_5 NS_157 0 7.2151108210705061e-06
GC_5_158 b_5 NI_5 NS_158 0 2.9209455164854195e-06
GC_5_159 b_5 NI_5 NS_159 0 4.2720180349118585e-05
GC_5_160 b_5 NI_5 NS_160 0 -1.9006948890630886e-05
GC_5_161 b_5 NI_5 NS_161 0 -2.4852123198813042e-06
GC_5_162 b_5 NI_5 NS_162 0 -7.7713947895694157e-06
GC_5_163 b_5 NI_5 NS_163 0 -2.8170177173374440e-06
GC_5_164 b_5 NI_5 NS_164 0 1.1098437706058294e-06
GC_5_165 b_5 NI_5 NS_165 0 9.8836278162012447e-06
GC_5_166 b_5 NI_5 NS_166 0 2.6879779132640394e-06
GC_5_167 b_5 NI_5 NS_167 0 2.2660734701609785e-05
GC_5_168 b_5 NI_5 NS_168 0 -3.3266519774984321e-05
GC_5_169 b_5 NI_5 NS_169 0 -5.7339960180601794e-06
GC_5_170 b_5 NI_5 NS_170 0 -4.2993052421381814e-06
GC_5_171 b_5 NI_5 NS_171 0 -8.7801403861780995e-07
GC_5_172 b_5 NI_5 NS_172 0 4.2822873388479817e-06
GC_5_173 b_5 NI_5 NS_173 0 1.2543456932289933e-05
GC_5_174 b_5 NI_5 NS_174 0 -1.7546455034801471e-07
GC_5_175 b_5 NI_5 NS_175 0 6.1365437826763355e-07
GC_5_176 b_5 NI_5 NS_176 0 -3.3004235280196080e-05
GC_5_177 b_5 NI_5 NS_177 0 -6.9295586688150999e-06
GC_5_178 b_5 NI_5 NS_178 0 3.5363607827503736e-07
GC_5_179 b_5 NI_5 NS_179 0 3.8626225691404407e-06
GC_5_180 b_5 NI_5 NS_180 0 3.5637315396801641e-06
GC_5_181 b_5 NI_5 NS_181 0 1.4168104589277933e-05
GC_5_182 b_5 NI_5 NS_182 0 -6.6370225967526434e-06
GC_5_183 b_5 NI_5 NS_183 0 -1.5560877831113016e-05
GC_5_184 b_5 NI_5 NS_184 0 -1.9131984324151728e-05
GC_5_185 b_5 NI_5 NS_185 0 -2.9829633958296556e-06
GC_5_186 b_5 NI_5 NS_186 0 5.0701585869991597e-06
GC_5_187 b_5 NI_5 NS_187 0 4.2041653841236000e-06
GC_5_188 b_5 NI_5 NS_188 0 -1.9025970383808676e-06
GC_5_189 b_5 NI_5 NS_189 0 -2.7722208047355360e-11
GC_5_190 b_5 NI_5 NS_190 0 5.4080553477674832e-12
GC_5_191 b_5 NI_5 NS_191 0 4.8943359664259501e-06
GC_5_192 b_5 NI_5 NS_192 0 -1.1671179340103900e-05
GC_5_193 b_5 NI_5 NS_193 0 -5.0226823241890364e-07
GC_5_194 b_5 NI_5 NS_194 0 2.7925790778147635e-06
GC_5_195 b_5 NI_5 NS_195 0 2.3625602483794482e-06
GC_5_196 b_5 NI_5 NS_196 0 -1.5932471527649705e-06
GC_5_197 b_5 NI_5 NS_197 0 2.1702780011101765e-06
GC_5_198 b_5 NI_5 NS_198 0 -9.8796185581650037e-06
GC_5_199 b_5 NI_5 NS_199 0 -1.0601744018663884e-05
GC_5_200 b_5 NI_5 NS_200 0 -3.5479011364653381e-06
GC_5_201 b_5 NI_5 NS_201 0 -2.2615789175465848e-10
GC_5_202 b_5 NI_5 NS_202 0 4.2333637444384087e-10
GC_5_203 b_5 NI_5 NS_203 0 -9.1524845256411647e-06
GC_5_204 b_5 NI_5 NS_204 0 -5.6556645078108469e-06
GC_5_205 b_5 NI_5 NS_205 0 2.0113008664685177e-06
GC_5_206 b_5 NI_5 NS_206 0 -6.6968789551833710e-06
GC_5_207 b_5 NI_5 NS_207 0 -3.3581443855826444e-06
GC_5_208 b_5 NI_5 NS_208 0 -1.8350847420995814e-07
GC_5_209 b_5 NI_5 NS_209 0 -8.5821482181935273e-06
GC_5_210 b_5 NI_5 NS_210 0 5.9051085095420980e-07
GC_5_211 b_5 NI_5 NS_211 0 2.6252776974095459e-06
GC_5_212 b_5 NI_5 NS_212 0 2.8290990425750742e-06
GC_5_213 b_5 NI_5 NS_213 0 1.0192405083659929e-06
GC_5_214 b_5 NI_5 NS_214 0 -3.7248619913016149e-06
GC_5_215 b_5 NI_5 NS_215 0 -5.3998861522584640e-06
GC_5_216 b_5 NI_5 NS_216 0 -4.2209464232648554e-06
GC_5_217 b_5 NI_5 NS_217 0 7.9312340287385335e-05
GC_5_218 b_5 NI_5 NS_218 0 -1.2174728879028769e-10
GC_5_219 b_5 NI_5 NS_219 0 -2.0288642719533222e-09
GC_5_220 b_5 NI_5 NS_220 0 3.4021535716010720e-08
GC_5_221 b_5 NI_5 NS_221 0 -3.3964213887284576e-07
GC_5_222 b_5 NI_5 NS_222 0 -3.3541275618804137e-07
GC_5_223 b_5 NI_5 NS_223 0 -5.7544861153099127e-07
GC_5_224 b_5 NI_5 NS_224 0 9.6680843459861226e-06
GC_5_225 b_5 NI_5 NS_225 0 1.3106737842406999e-05
GC_5_226 b_5 NI_5 NS_226 0 -1.2342131449792206e-05
GC_5_227 b_5 NI_5 NS_227 0 -1.7111534650678110e-05
GC_5_228 b_5 NI_5 NS_228 0 8.5766065778295356e-06
GC_5_229 b_5 NI_5 NS_229 0 2.8664512720412465e-05
GC_5_230 b_5 NI_5 NS_230 0 -7.4207273445259304e-06
GC_5_231 b_5 NI_5 NS_231 0 -2.8948010736409704e-06
GC_5_232 b_5 NI_5 NS_232 0 -3.4132503440024330e-06
GC_5_233 b_5 NI_5 NS_233 0 -3.2450872673487185e-06
GC_5_234 b_5 NI_5 NS_234 0 -1.5091692824993239e-05
GC_5_235 b_5 NI_5 NS_235 0 -2.4827138350307669e-05
GC_5_236 b_5 NI_5 NS_236 0 3.9219959907066287e-05
GC_5_237 b_5 NI_5 NS_237 0 3.6986155281493279e-05
GC_5_238 b_5 NI_5 NS_238 0 -4.7226450976527001e-05
GC_5_239 b_5 NI_5 NS_239 0 -3.0518033319569036e-05
GC_5_240 b_5 NI_5 NS_240 0 -2.1425944494030440e-05
GC_5_241 b_5 NI_5 NS_241 0 3.2013254461636942e-05
GC_5_242 b_5 NI_5 NS_242 0 2.6385822254694680e-05
GC_5_243 b_5 NI_5 NS_243 0 -1.8545782640186131e-05
GC_5_244 b_5 NI_5 NS_244 0 -2.9076767252964962e-05
GC_5_245 b_5 NI_5 NS_245 0 2.0024652579897973e-05
GC_5_246 b_5 NI_5 NS_246 0 5.9802325505021992e-05
GC_5_247 b_5 NI_5 NS_247 0 -2.0977170143840720e-05
GC_5_248 b_5 NI_5 NS_248 0 -5.5613239106559751e-05
GC_5_249 b_5 NI_5 NS_249 0 -3.1646089244782871e-05
GC_5_250 b_5 NI_5 NS_250 0 -1.2117270378733763e-05
GC_5_251 b_5 NI_5 NS_251 0 1.9560562289148279e-05
GC_5_252 b_5 NI_5 NS_252 0 1.3805681165603732e-05
GC_5_253 b_5 NI_5 NS_253 0 -2.4957519127897135e-05
GC_5_254 b_5 NI_5 NS_254 0 -1.1262953470921864e-05
GC_5_255 b_5 NI_5 NS_255 0 2.0178609176623610e-05
GC_5_256 b_5 NI_5 NS_256 0 1.0341432468666392e-05
GC_5_257 b_5 NI_5 NS_257 0 -1.8434398821733068e-05
GC_5_258 b_5 NI_5 NS_258 0 -2.1152962142287066e-05
GC_5_259 b_5 NI_5 NS_259 0 4.2938807325511784e-06
GC_5_260 b_5 NI_5 NS_260 0 3.1956500207445692e-05
GC_5_261 b_5 NI_5 NS_261 0 -8.4070366811796401e-06
GC_5_262 b_5 NI_5 NS_262 0 -2.6582373016082145e-05
GC_5_263 b_5 NI_5 NS_263 0 -2.0405918550151595e-06
GC_5_264 b_5 NI_5 NS_264 0 1.5411381230737415e-06
GC_5_265 b_5 NI_5 NS_265 0 -1.9680637760611203e-05
GC_5_266 b_5 NI_5 NS_266 0 -1.2199249318004474e-05
GC_5_267 b_5 NI_5 NS_267 0 5.5358532311673602e-06
GC_5_268 b_5 NI_5 NS_268 0 2.1303964189302156e-05
GC_5_269 b_5 NI_5 NS_269 0 -1.6264288097054502e-05
GC_5_270 b_5 NI_5 NS_270 0 -1.4842704671931754e-05
GC_5_271 b_5 NI_5 NS_271 0 9.0112822626279403e-07
GC_5_272 b_5 NI_5 NS_272 0 5.5183487177882359e-06
GC_5_273 b_5 NI_5 NS_273 0 -2.5231535076039770e-05
GC_5_274 b_5 NI_5 NS_274 0 -1.0007123700603306e-05
GC_5_275 b_5 NI_5 NS_275 0 7.5015455301516696e-06
GC_5_276 b_5 NI_5 NS_276 0 2.3879817466643611e-05
GC_5_277 b_5 NI_5 NS_277 0 -2.0944356483758350e-05
GC_5_278 b_5 NI_5 NS_278 0 -5.6383716821824844e-06
GC_5_279 b_5 NI_5 NS_279 0 5.9390411813307787e-06
GC_5_280 b_5 NI_5 NS_280 0 7.9065229502285228e-06
GC_5_281 b_5 NI_5 NS_281 0 -3.0919139851502015e-05
GC_5_282 b_5 NI_5 NS_282 0 -2.7456247115619932e-06
GC_5_283 b_5 NI_5 NS_283 0 1.8051020262471785e-05
GC_5_284 b_5 NI_5 NS_284 0 2.6173001080867463e-05
GC_5_285 b_5 NI_5 NS_285 0 -2.2120993067776816e-05
GC_5_286 b_5 NI_5 NS_286 0 6.9969215974378713e-06
GC_5_287 b_5 NI_5 NS_287 0 1.5076261028388675e-05
GC_5_288 b_5 NI_5 NS_288 0 4.4859629687018865e-06
GC_5_289 b_5 NI_5 NS_289 0 -3.5006554378738130e-05
GC_5_290 b_5 NI_5 NS_290 0 1.3594209357041676e-05
GC_5_291 b_5 NI_5 NS_291 0 3.7183707988699120e-05
GC_5_292 b_5 NI_5 NS_292 0 1.3345626225646490e-05
GC_5_293 b_5 NI_5 NS_293 0 -7.9978699141781709e-06
GC_5_294 b_5 NI_5 NS_294 0 1.9077609464559750e-05
GC_5_295 b_5 NI_5 NS_295 0 1.2877011362647394e-05
GC_5_296 b_5 NI_5 NS_296 0 -1.0946410020861583e-05
GC_5_297 b_5 NI_5 NS_297 0 1.1098383904467769e-10
GC_5_298 b_5 NI_5 NS_298 0 4.4145416124398918e-11
GC_5_299 b_5 NI_5 NS_299 0 -1.3993786032243076e-05
GC_5_300 b_5 NI_5 NS_300 0 2.6116714369132735e-05
GC_5_301 b_5 NI_5 NS_301 0 -2.1469382270038087e-06
GC_5_302 b_5 NI_5 NS_302 0 1.0637062906842548e-05
GC_5_303 b_5 NI_5 NS_303 0 6.1622217285742884e-06
GC_5_304 b_5 NI_5 NS_304 0 -8.3662944813252374e-06
GC_5_305 b_5 NI_5 NS_305 0 -8.3615490223166079e-06
GC_5_306 b_5 NI_5 NS_306 0 2.5491909516699304e-05
GC_5_307 b_5 NI_5 NS_307 0 2.5015462421219589e-05
GC_5_308 b_5 NI_5 NS_308 0 -9.9972210299303892e-06
GC_5_309 b_5 NI_5 NS_309 0 4.8733647576968243e-09
GC_5_310 b_5 NI_5 NS_310 0 -1.1064268423560237e-09
GC_5_311 b_5 NI_5 NS_311 0 2.6321439058683769e-05
GC_5_312 b_5 NI_5 NS_312 0 -1.2477166441000342e-05
GC_5_313 b_5 NI_5 NS_313 0 -8.3191197590192563e-06
GC_5_314 b_5 NI_5 NS_314 0 1.8150071297753763e-05
GC_5_315 b_5 NI_5 NS_315 0 -1.0398966208042270e-05
GC_5_316 b_5 NI_5 NS_316 0 -2.8340099544356740e-07
GC_5_317 b_5 NI_5 NS_317 0 1.9410890875706547e-05
GC_5_318 b_5 NI_5 NS_318 0 -1.4076803304902632e-05
GC_5_319 b_5 NI_5 NS_319 0 7.1589747635440692e-06
GC_5_320 b_5 NI_5 NS_320 0 1.1755238511269529e-05
GC_5_321 b_5 NI_5 NS_321 0 -1.8090522501790801e-07
GC_5_322 b_5 NI_5 NS_322 0 -1.4547113308895627e-05
GC_5_323 b_5 NI_5 NS_323 0 1.3082627277679036e-05
GC_5_324 b_5 NI_5 NS_324 0 2.7941805431571423e-05
GC_5_325 b_5 NI_5 NS_325 0 -6.4096524188712964e-04
GC_5_326 b_5 NI_5 NS_326 0 -9.7194652103576596e-11
GC_5_327 b_5 NI_5 NS_327 0 3.8858046973773393e-09
GC_5_328 b_5 NI_5 NS_328 0 -6.7398838150045628e-08
GC_5_329 b_5 NI_5 NS_329 0 -1.1319906730508755e-05
GC_5_330 b_5 NI_5 NS_330 0 -9.3647686904640091e-06
GC_5_331 b_5 NI_5 NS_331 0 -2.2431758661141731e-06
GC_5_332 b_5 NI_5 NS_332 0 2.0358582925232762e-07
GC_5_333 b_5 NI_5 NS_333 0 -3.0429845588867101e-05
GC_5_334 b_5 NI_5 NS_334 0 2.7128791122381809e-05
GC_5_335 b_5 NI_5 NS_335 0 -3.3446187014487919e-05
GC_5_336 b_5 NI_5 NS_336 0 8.1023554136814512e-06
GC_5_337 b_5 NI_5 NS_337 0 3.1775636534477179e-05
GC_5_338 b_5 NI_5 NS_338 0 2.7493580026078690e-05
GC_5_339 b_5 NI_5 NS_339 0 -9.1079481586903514e-06
GC_5_340 b_5 NI_5 NS_340 0 1.4797967073144262e-05
GC_5_341 b_5 NI_5 NS_341 0 1.2654201149064630e-05
GC_5_342 b_5 NI_5 NS_342 0 3.7136163185928859e-05
GC_5_343 b_5 NI_5 NS_343 0 -1.1049969265257533e-05
GC_5_344 b_5 NI_5 NS_344 0 6.8460625983763772e-05
GC_5_345 b_5 NI_5 NS_345 0 9.6052101801470433e-05
GC_5_346 b_5 NI_5 NS_346 0 -6.6220034837778468e-05
GC_5_347 b_5 NI_5 NS_347 0 2.7188454434379573e-05
GC_5_348 b_5 NI_5 NS_348 0 3.2025518834109497e-05
GC_5_349 b_5 NI_5 NS_349 0 -6.9721036164181328e-06
GC_5_350 b_5 NI_5 NS_350 0 -7.2660803358987527e-05
GC_5_351 b_5 NI_5 NS_351 0 -9.8238622879540956e-06
GC_5_352 b_5 NI_5 NS_352 0 -3.4299022567157071e-05
GC_5_353 b_5 NI_5 NS_353 0 -7.6898752082057623e-05
GC_5_354 b_5 NI_5 NS_354 0 1.8642121849917050e-05
GC_5_355 b_5 NI_5 NS_355 0 2.4833373571420110e-05
GC_5_356 b_5 NI_5 NS_356 0 5.1420166605223892e-05
GC_5_357 b_5 NI_5 NS_357 0 -2.3340308167248569e-05
GC_5_358 b_5 NI_5 NS_358 0 -3.7721127675747912e-06
GC_5_359 b_5 NI_5 NS_359 0 7.0064427220874737e-05
GC_5_360 b_5 NI_5 NS_360 0 4.4958994560725184e-05
GC_5_361 b_5 NI_5 NS_361 0 2.9394321559782050e-05
GC_5_362 b_5 NI_5 NS_362 0 1.9999802746396495e-05
GC_5_363 b_5 NI_5 NS_363 0 -7.2203628846963043e-06
GC_5_364 b_5 NI_5 NS_364 0 -2.5839477841251672e-05
GC_5_365 b_5 NI_5 NS_365 0 -7.5634346949473650e-06
GC_5_366 b_5 NI_5 NS_366 0 -2.5468695720511736e-05
GC_5_367 b_5 NI_5 NS_367 0 6.9064251988408714e-06
GC_5_368 b_5 NI_5 NS_368 0 4.9199298330854250e-05
GC_5_369 b_5 NI_5 NS_369 0 1.2870889028669816e-05
GC_5_370 b_5 NI_5 NS_370 0 2.7631526925720403e-05
GC_5_371 b_5 NI_5 NS_371 0 5.8803230541565413e-06
GC_5_372 b_5 NI_5 NS_372 0 2.1449616235898124e-06
GC_5_373 b_5 NI_5 NS_373 0 -6.1110934648000879e-07
GC_5_374 b_5 NI_5 NS_374 0 -1.5594144304049277e-05
GC_5_375 b_5 NI_5 NS_375 0 5.6392053631215779e-05
GC_5_376 b_5 NI_5 NS_376 0 3.8210578508976788e-05
GC_5_377 b_5 NI_5 NS_377 0 1.9988529622808133e-05
GC_5_378 b_5 NI_5 NS_378 0 1.5010233907489081e-05
GC_5_379 b_5 NI_5 NS_379 0 8.4379987541403134e-06
GC_5_380 b_5 NI_5 NS_380 0 -1.2896802811186457e-05
GC_5_381 b_5 NI_5 NS_381 0 -5.6459176403866037e-06
GC_5_382 b_5 NI_5 NS_382 0 -1.4204665875109669e-05
GC_5_383 b_5 NI_5 NS_383 0 6.6278851865041673e-05
GC_5_384 b_5 NI_5 NS_384 0 1.2995832380157651e-05
GC_5_385 b_5 NI_5 NS_385 0 2.2839922936942664e-05
GC_5_386 b_5 NI_5 NS_386 0 5.0561016903861697e-06
GC_5_387 b_5 NI_5 NS_387 0 -5.5482171369921653e-06
GC_5_388 b_5 NI_5 NS_388 0 -2.2088161004867522e-05
GC_5_389 b_5 NI_5 NS_389 0 -9.1406537728618196e-06
GC_5_390 b_5 NI_5 NS_390 0 -7.2230786479206559e-06
GC_5_391 b_5 NI_5 NS_391 0 6.0751027178145810e-05
GC_5_392 b_5 NI_5 NS_392 0 -9.5212181549709886e-06
GC_5_393 b_5 NI_5 NS_393 0 2.1480537553740708e-05
GC_5_394 b_5 NI_5 NS_394 0 -7.3371752582271807e-06
GC_5_395 b_5 NI_5 NS_395 0 -2.3109762471187094e-05
GC_5_396 b_5 NI_5 NS_396 0 -1.3195896352784168e-05
GC_5_397 b_5 NI_5 NS_397 0 -8.6441610886410418e-06
GC_5_398 b_5 NI_5 NS_398 0 4.3874530325957994e-06
GC_5_399 b_5 NI_5 NS_399 0 4.5483158253399227e-05
GC_5_400 b_5 NI_5 NS_400 0 -2.5698454241879601e-05
GC_5_401 b_5 NI_5 NS_401 0 6.0412474105379190e-06
GC_5_402 b_5 NI_5 NS_402 0 -1.6494042023223898e-05
GC_5_403 b_5 NI_5 NS_403 0 -1.8742829615567515e-05
GC_5_404 b_5 NI_5 NS_404 0 8.5986458384940614e-06
GC_5_405 b_5 NI_5 NS_405 0 -4.6792901998604387e-11
GC_5_406 b_5 NI_5 NS_406 0 -1.7807207643411924e-10
GC_5_407 b_5 NI_5 NS_407 0 1.7713030730704860e-06
GC_5_408 b_5 NI_5 NS_408 0 8.7581308107499136e-06
GC_5_409 b_5 NI_5 NS_409 0 2.2084514150115554e-06
GC_5_410 b_5 NI_5 NS_410 0 -7.0117489405335226e-06
GC_5_411 b_5 NI_5 NS_411 0 -9.0106065282487055e-06
GC_5_412 b_5 NI_5 NS_412 0 5.7573236107450229e-06
GC_5_413 b_5 NI_5 NS_413 0 4.7874459814928740e-06
GC_5_414 b_5 NI_5 NS_414 0 1.1558464822946979e-05
GC_5_415 b_5 NI_5 NS_415 0 2.4565262552523318e-05
GC_5_416 b_5 NI_5 NS_416 0 -2.1165221313736700e-05
GC_5_417 b_5 NI_5 NS_417 0 -5.7149999727927585e-09
GC_5_418 b_5 NI_5 NS_418 0 -5.6483219370892215e-09
GC_5_419 b_5 NI_5 NS_419 0 3.0655889741418790e-05
GC_5_420 b_5 NI_5 NS_420 0 7.4872140595220056e-06
GC_5_421 b_5 NI_5 NS_421 0 -2.6797317153853448e-06
GC_5_422 b_5 NI_5 NS_422 0 1.1045236987708439e-05
GC_5_423 b_5 NI_5 NS_423 0 8.0410643091225191e-06
GC_5_424 b_5 NI_5 NS_424 0 1.1946460638839478e-06
GC_5_425 b_5 NI_5 NS_425 0 1.9120712051456026e-05
GC_5_426 b_5 NI_5 NS_426 0 -2.1559501970631235e-05
GC_5_427 b_5 NI_5 NS_427 0 -6.5503006494838480e-06
GC_5_428 b_5 NI_5 NS_428 0 -7.4615416082513339e-06
GC_5_429 b_5 NI_5 NS_429 0 -5.3942518305392882e-06
GC_5_430 b_5 NI_5 NS_430 0 1.2484971255732885e-05
GC_5_431 b_5 NI_5 NS_431 0 1.6111580009673562e-05
GC_5_432 b_5 NI_5 NS_432 0 7.3766058346903001e-06
GC_5_433 b_5 NI_5 NS_433 0 -1.3590038758593249e-02
GC_5_434 b_5 NI_5 NS_434 0 5.7574113574367023e-09
GC_5_435 b_5 NI_5 NS_435 0 -1.0755251955003008e-06
GC_5_436 b_5 NI_5 NS_436 0 -2.3265200914776547e-05
GC_5_437 b_5 NI_5 NS_437 0 3.4981851747783630e-04
GC_5_438 b_5 NI_5 NS_438 0 -1.9740598410815851e-04
GC_5_439 b_5 NI_5 NS_439 0 -1.5437483444288782e-03
GC_5_440 b_5 NI_5 NS_440 0 -2.3356983122441431e-03
GC_5_441 b_5 NI_5 NS_441 0 -5.1340364113444250e-05
GC_5_442 b_5 NI_5 NS_442 0 4.3605120496332042e-03
GC_5_443 b_5 NI_5 NS_443 0 1.6175824927349835e-03
GC_5_444 b_5 NI_5 NS_444 0 -5.9520405602870117e-03
GC_5_445 b_5 NI_5 NS_445 0 -4.9853593163292865e-03
GC_5_446 b_5 NI_5 NS_446 0 6.4563571009632866e-03
GC_5_447 b_5 NI_5 NS_447 0 1.1341380715634882e-03
GC_5_448 b_5 NI_5 NS_448 0 -5.0675425946490019e-04
GC_5_449 b_5 NI_5 NS_449 0 2.7871014128826818e-03
GC_5_450 b_5 NI_5 NS_450 0 2.3388044429882081e-03
GC_5_451 b_5 NI_5 NS_451 0 -4.3321682726310774e-03
GC_5_452 b_5 NI_5 NS_452 0 -1.3583565618000164e-02
GC_5_453 b_5 NI_5 NS_453 0 1.5695038276344019e-03
GC_5_454 b_5 NI_5 NS_454 0 1.7683041197579442e-02
GC_5_455 b_5 NI_5 NS_455 0 9.8323126131528420e-03
GC_5_456 b_5 NI_5 NS_456 0 -2.3109432708629794e-03
GC_5_457 b_5 NI_5 NS_457 0 -1.3157073609238330e-02
GC_5_458 b_5 NI_5 NS_458 0 2.2142408000816963e-03
GC_5_459 b_5 NI_5 NS_459 0 9.1925784034046949e-03
GC_5_460 b_5 NI_5 NS_460 0 1.9425112077200361e-03
GC_5_461 b_5 NI_5 NS_461 0 -1.8069422469017122e-02
GC_5_462 b_5 NI_5 NS_462 0 -6.4922283942858783e-03
GC_5_463 b_5 NI_5 NS_463 0 1.5725028675783109e-02
GC_5_464 b_5 NI_5 NS_464 0 6.4951447484251686e-03
GC_5_465 b_5 NI_5 NS_465 0 8.1032003105176095e-03
GC_5_466 b_5 NI_5 NS_466 0 -4.2110876475472802e-03
GC_5_467 b_5 NI_5 NS_467 0 -7.5660795372926573e-03
GC_5_468 b_5 NI_5 NS_468 0 2.0432100992714675e-03
GC_5_469 b_5 NI_5 NS_469 0 6.6854379760949885e-03
GC_5_470 b_5 NI_5 NS_470 0 -2.7541177502804033e-03
GC_5_471 b_5 NI_5 NS_471 0 -6.6055144911246078e-03
GC_5_472 b_5 NI_5 NS_472 0 2.9142121005506848e-03
GC_5_473 b_5 NI_5 NS_473 0 7.6544557708656900e-03
GC_5_474 b_5 NI_5 NS_474 0 4.7732052876346117e-04
GC_5_475 b_5 NI_5 NS_475 0 -9.4088268642744249e-03
GC_5_476 b_5 NI_5 NS_476 0 -5.1695959250252135e-03
GC_5_477 b_5 NI_5 NS_477 0 6.8169842482272642e-03
GC_5_478 b_5 NI_5 NS_478 0 4.1131794029750429e-03
GC_5_479 b_5 NI_5 NS_479 0 -3.9574846280538876e-04
GC_5_480 b_5 NI_5 NS_480 0 -9.3604180763591407e-04
GC_5_481 b_5 NI_5 NS_481 0 5.6653317207762338e-03
GC_5_482 b_5 NI_5 NS_482 0 -1.3801820683057744e-03
GC_5_483 b_5 NI_5 NS_483 0 -9.2023184182152221e-03
GC_5_484 b_5 NI_5 NS_484 0 -1.2456050726628426e-03
GC_5_485 b_5 NI_5 NS_485 0 5.9915313907571858e-03
GC_5_486 b_5 NI_5 NS_486 0 7.3808348578682185e-04
GC_5_487 b_5 NI_5 NS_487 0 -2.6544549900193856e-03
GC_5_488 b_5 NI_5 NS_488 0 2.4842222125145063e-04
GC_5_489 b_5 NI_5 NS_489 0 6.6958828091666237e-03
GC_5_490 b_5 NI_5 NS_490 0 -2.2582329946152272e-03
GC_5_491 b_5 NI_5 NS_491 0 -9.3158089924149767e-03
GC_5_492 b_5 NI_5 NS_492 0 1.5268648283366004e-03
GC_5_493 b_5 NI_5 NS_493 0 5.7300536260805291e-03
GC_5_494 b_5 NI_5 NS_494 0 -1.5007448373696784e-03
GC_5_495 b_5 NI_5 NS_495 0 -3.3211781925187741e-03
GC_5_496 b_5 NI_5 NS_496 0 2.4082389398275782e-03
GC_5_497 b_5 NI_5 NS_497 0 7.2643742621706269e-03
GC_5_498 b_5 NI_5 NS_498 0 -4.0966037542834134e-03
GC_5_499 b_5 NI_5 NS_499 0 -8.5936681109166930e-03
GC_5_500 b_5 NI_5 NS_500 0 4.2025452154415581e-03
GC_5_501 b_5 NI_5 NS_501 0 4.8158705784495260e-03
GC_5_502 b_5 NI_5 NS_502 0 -3.8696540515473087e-03
GC_5_503 b_5 NI_5 NS_503 0 -2.4037860168784767e-03
GC_5_504 b_5 NI_5 NS_504 0 4.7598874104292626e-03
GC_5_505 b_5 NI_5 NS_505 0 7.0540631349609731e-03
GC_5_506 b_5 NI_5 NS_506 0 -7.3479437791381073e-03
GC_5_507 b_5 NI_5 NS_507 0 -7.1271032067403610e-03
GC_5_508 b_5 NI_5 NS_508 0 6.8936503102674821e-03
GC_5_509 b_5 NI_5 NS_509 0 1.6683514128538954e-03
GC_5_510 b_5 NI_5 NS_510 0 -5.2972255960430170e-03
GC_5_511 b_5 NI_5 NS_511 0 5.9423078355015592e-04
GC_5_512 b_5 NI_5 NS_512 0 5.4734770636633212e-03
GC_5_513 b_5 NI_5 NS_513 0 -4.1996224590810328e-09
GC_5_514 b_5 NI_5 NS_514 0 -1.3215473074973935e-08
GC_5_515 b_5 NI_5 NS_515 0 2.7118324802203695e-03
GC_5_516 b_5 NI_5 NS_516 0 -8.5806166158300858e-03
GC_5_517 b_5 NI_5 NS_517 0 8.7189105151590663e-04
GC_5_518 b_5 NI_5 NS_518 0 -3.4318678539232007e-03
GC_5_519 b_5 NI_5 NS_519 0 6.2897431415977765e-04
GC_5_520 b_5 NI_5 NS_520 0 4.0346894477520413e-03
GC_5_521 b_5 NI_5 NS_521 0 2.1766535629687989e-03
GC_5_522 b_5 NI_5 NS_522 0 -8.1586516493607278e-03
GC_5_523 b_5 NI_5 NS_523 0 -3.4870480262388921e-03
GC_5_524 b_5 NI_5 NS_524 0 7.0184773261586387e-03
GC_5_525 b_5 NI_5 NS_525 0 -9.0338470133171919e-08
GC_5_526 b_5 NI_5 NS_526 0 -3.0340980818064251e-07
GC_5_527 b_5 NI_5 NS_527 0 -8.0011233891473764e-03
GC_5_528 b_5 NI_5 NS_528 0 5.3809331600617122e-03
GC_5_529 b_5 NI_5 NS_529 0 4.1753794557669987e-03
GC_5_530 b_5 NI_5 NS_530 0 -6.8471564425540178e-03
GC_5_531 b_5 NI_5 NS_531 0 5.3267679624766015e-03
GC_5_532 b_5 NI_5 NS_532 0 7.4221568060225062e-04
GC_5_533 b_5 NI_5 NS_533 0 -2.3672765884590399e-03
GC_5_534 b_5 NI_5 NS_534 0 6.8575175439453268e-03
GC_5_535 b_5 NI_5 NS_535 0 -1.4866281827222091e-03
GC_5_536 b_5 NI_5 NS_536 0 -4.2154555137040133e-03
GC_5_537 b_5 NI_5 NS_537 0 2.3568558413644310e-03
GC_5_538 b_5 NI_5 NS_538 0 5.0372669558086591e-03
GC_5_539 b_5 NI_5 NS_539 0 -1.9997035533975130e-03
GC_5_540 b_5 NI_5 NS_540 0 -8.9736637719760350e-03
GC_5_541 b_5 NI_5 NS_541 0 -1.0963064049019198e-02
GC_5_542 b_5 NI_5 NS_542 0 8.3276040449876566e-09
GC_5_543 b_5 NI_5 NS_543 0 9.8608103426122305e-07
GC_5_544 b_5 NI_5 NS_544 0 3.6177580226032927e-05
GC_5_545 b_5 NI_5 NS_545 0 4.3739109611715052e-03
GC_5_546 b_5 NI_5 NS_546 0 -3.4750186020288576e-03
GC_5_547 b_5 NI_5 NS_547 0 -3.7382698156534977e-03
GC_5_548 b_5 NI_5 NS_548 0 6.2463760221297786e-03
GC_5_549 b_5 NI_5 NS_549 0 -8.7586388741214237e-03
GC_5_550 b_5 NI_5 NS_550 0 -5.9567829542500539e-03
GC_5_551 b_5 NI_5 NS_551 0 9.2115253055727649e-03
GC_5_552 b_5 NI_5 NS_552 0 -5.9461326426276826e-03
GC_5_553 b_5 NI_5 NS_553 0 7.1478898347439521e-03
GC_5_554 b_5 NI_5 NS_554 0 1.1907375056175749e-02
GC_5_555 b_5 NI_5 NS_555 0 -4.2314190352109420e-03
GC_5_556 b_5 NI_5 NS_556 0 -1.1324176399823728e-03
GC_5_557 b_5 NI_5 NS_557 0 -8.8598375246884218e-03
GC_5_558 b_5 NI_5 NS_558 0 -4.7420113826033547e-04
GC_5_559 b_5 NI_5 NS_559 0 1.4618469427396467e-02
GC_5_560 b_5 NI_5 NS_560 0 -1.0343832302290327e-02
GC_5_561 b_5 NI_5 NS_561 0 1.6441807885684410e-02
GC_5_562 b_5 NI_5 NS_562 0 4.0224873813991579e-03
GC_5_563 b_5 NI_5 NS_563 0 -1.1482355556039063e-02
GC_5_564 b_5 NI_5 NS_564 0 -2.4511486411351929e-04
GC_5_565 b_5 NI_5 NS_565 0 -1.6636891788926068e-02
GC_5_566 b_5 NI_5 NS_566 0 -4.4573868505651218e-02
GC_5_567 b_5 NI_5 NS_567 0 1.0652631230489205e-02
GC_5_568 b_5 NI_5 NS_568 0 1.1245746841033893e-03
GC_5_569 b_5 NI_5 NS_569 0 -4.8294106848337529e-02
GC_5_570 b_5 NI_5 NS_570 0 1.1061711810642527e-02
GC_5_571 b_5 NI_5 NS_571 0 -1.0433752537752548e-02
GC_5_572 b_5 NI_5 NS_572 0 4.8882942819980047e-04
GC_5_573 b_5 NI_5 NS_573 0 9.7769907743760678e-03
GC_5_574 b_5 NI_5 NS_574 0 -5.7680205299312645e-04
GC_5_575 b_5 NI_5 NS_575 0 4.6095772202893433e-03
GC_5_576 b_5 NI_5 NS_576 0 2.4174004313286972e-02
GC_5_577 b_5 NI_5 NS_577 0 -1.0735354440562044e-02
GC_5_578 b_5 NI_5 NS_578 0 1.9692006570899779e-03
GC_5_579 b_5 NI_5 NS_579 0 -8.4727383217558967e-03
GC_5_580 b_5 NI_5 NS_580 0 -1.3537885007543816e-02
GC_5_581 b_5 NI_5 NS_581 0 1.0150130521780005e-02
GC_5_582 b_5 NI_5 NS_582 0 9.8140712602090042e-04
GC_5_583 b_5 NI_5 NS_583 0 -1.9163144483401562e-02
GC_5_584 b_5 NI_5 NS_584 0 2.8679170724212825e-02
GC_5_585 b_5 NI_5 NS_585 0 -9.6128548515520534e-03
GC_5_586 b_5 NI_5 NS_586 0 -9.6554385072997108e-04
GC_5_587 b_5 NI_5 NS_587 0 1.8914200218990637e-03
GC_5_588 b_5 NI_5 NS_588 0 -1.3780552719562279e-03
GC_5_589 b_5 NI_5 NS_589 0 9.4682970903075345e-03
GC_5_590 b_5 NI_5 NS_590 0 -2.4741583795876636e-04
GC_5_591 b_5 NI_5 NS_591 0 -1.4945957045042364e-04
GC_5_592 b_5 NI_5 NS_592 0 3.0270105339883772e-02
GC_5_593 b_5 NI_5 NS_593 0 -8.5288659060314461e-03
GC_5_594 b_5 NI_5 NS_594 0 1.5478659070894863e-04
GC_5_595 b_5 NI_5 NS_595 0 2.1681753052877524e-04
GC_5_596 b_5 NI_5 NS_596 0 -5.4812542014245364e-03
GC_5_597 b_5 NI_5 NS_597 0 1.0036166626380514e-02
GC_5_598 b_5 NI_5 NS_598 0 -3.3857521486935042e-04
GC_5_599 b_5 NI_5 NS_599 0 8.9341677935640459e-03
GC_5_600 b_5 NI_5 NS_600 0 2.6365823192744001e-02
GC_5_601 b_5 NI_5 NS_601 0 -8.3555383637252435e-03
GC_5_602 b_5 NI_5 NS_602 0 1.3766457737780589e-03
GC_5_603 b_5 NI_5 NS_603 0 -2.5869076875063598e-03
GC_5_604 b_5 NI_5 NS_604 0 -7.3539566536967573e-03
GC_5_605 b_5 NI_5 NS_605 0 1.0553563485746017e-02
GC_5_606 b_5 NI_5 NS_606 0 -8.2348944107654557e-04
GC_5_607 b_5 NI_5 NS_607 0 1.4439011550631426e-02
GC_5_608 b_5 NI_5 NS_608 0 1.9950607649539161e-02
GC_5_609 b_5 NI_5 NS_609 0 -8.2760873721814902e-03
GC_5_610 b_5 NI_5 NS_610 0 2.9305070575233690e-03
GC_5_611 b_5 NI_5 NS_611 0 -5.5941943284403958e-03
GC_5_612 b_5 NI_5 NS_612 0 -6.9177099727461859e-03
GC_5_613 b_5 NI_5 NS_613 0 1.1244063383513423e-02
GC_5_614 b_5 NI_5 NS_614 0 -1.3754142170368589e-03
GC_5_615 b_5 NI_5 NS_615 0 1.5700530413114439e-02
GC_5_616 b_5 NI_5 NS_616 0 1.2945594242576342e-02
GC_5_617 b_5 NI_5 NS_617 0 -7.1893619194723672e-03
GC_5_618 b_5 NI_5 NS_618 0 5.1106082376705074e-03
GC_5_619 b_5 NI_5 NS_619 0 -6.8765830029316648e-03
GC_5_620 b_5 NI_5 NS_620 0 -4.8360422681987128e-03
GC_5_621 b_5 NI_5 NS_621 0 4.7733278170655428e-09
GC_5_622 b_5 NI_5 NS_622 0 4.4199354920259731e-08
GC_5_623 b_5 NI_5 NS_623 0 1.2004105577491788e-02
GC_5_624 b_5 NI_5 NS_624 0 -2.5766622965509496e-03
GC_5_625 b_5 NI_5 NS_625 0 -5.2510754139268919e-03
GC_5_626 b_5 NI_5 NS_626 0 4.7015455809010015e-03
GC_5_627 b_5 NI_5 NS_627 0 -6.1588973822056829e-03
GC_5_628 b_5 NI_5 NS_628 0 -4.3232026021505420e-03
GC_5_629 b_5 NI_5 NS_629 0 1.1774219228665495e-02
GC_5_630 b_5 NI_5 NS_630 0 -3.7297226039134115e-03
GC_5_631 b_5 NI_5 NS_631 0 1.2978428438086245e-02
GC_5_632 b_5 NI_5 NS_632 0 9.4653971215730350e-03
GC_5_633 b_5 NI_5 NS_633 0 3.9180870575213841e-06
GC_5_634 b_5 NI_5 NS_634 0 -9.4184409370855057e-07
GC_5_635 b_5 NI_5 NS_635 0 1.6087880549333813e-02
GC_5_636 b_5 NI_5 NS_636 0 1.6769946127507041e-02
GC_5_637 b_5 NI_5 NS_637 0 1.2047068161880257e-02
GC_5_638 b_5 NI_5 NS_638 0 -2.4806927911000570e-03
GC_5_639 b_5 NI_5 NS_639 0 -8.3607714057994682e-03
GC_5_640 b_5 NI_5 NS_640 0 7.9691369514851043e-05
GC_5_641 b_5 NI_5 NS_641 0 1.1309400358354756e-02
GC_5_642 b_5 NI_5 NS_642 0 7.3306474354893920e-03
GC_5_643 b_5 NI_5 NS_643 0 -4.6732529370359282e-03
GC_5_644 b_5 NI_5 NS_644 0 7.3569230661379289e-03
GC_5_645 b_5 NI_5 NS_645 0 -8.0809726220005661e-03
GC_5_646 b_5 NI_5 NS_646 0 -3.7224016096122164e-03
GC_5_647 b_5 NI_5 NS_647 0 1.5958293471080159e-02
GC_5_648 b_5 NI_5 NS_648 0 -7.7554804179507282e-03
GC_5_649 b_5 NI_5 NS_649 0 1.4425743160263048e-03
GC_5_650 b_5 NI_5 NS_650 0 -3.5904351902060078e-09
GC_5_651 b_5 NI_5 NS_651 0 -4.7342043005218681e-08
GC_5_652 b_5 NI_5 NS_652 0 -3.5032371879168616e-06
GC_5_653 b_5 NI_5 NS_653 0 -3.6675402894641997e-04
GC_5_654 b_5 NI_5 NS_654 0 1.3531650072533770e-04
GC_5_655 b_5 NI_5 NS_655 0 1.1270906275200521e-03
GC_5_656 b_5 NI_5 NS_656 0 1.9466317895270150e-03
GC_5_657 b_5 NI_5 NS_657 0 -5.2133196348760781e-05
GC_5_658 b_5 NI_5 NS_658 0 -3.4959654221104592e-03
GC_5_659 b_5 NI_5 NS_659 0 -1.5728294468906720e-03
GC_5_660 b_5 NI_5 NS_660 0 5.0835061312654306e-03
GC_5_661 b_5 NI_5 NS_661 0 4.2660497518820471e-03
GC_5_662 b_5 NI_5 NS_662 0 -4.9897929468884199e-03
GC_5_663 b_5 NI_5 NS_663 0 -1.0071498220759407e-03
GC_5_664 b_5 NI_5 NS_664 0 5.5941855889055970e-04
GC_5_665 b_5 NI_5 NS_665 0 -2.0791294208185357e-03
GC_5_666 b_5 NI_5 NS_666 0 -1.8719561555056231e-03
GC_5_667 b_5 NI_5 NS_667 0 3.6235023872609852e-03
GC_5_668 b_5 NI_5 NS_668 0 1.1644121608893596e-02
GC_5_669 b_5 NI_5 NS_669 0 -8.7672707288597481e-04
GC_5_670 b_5 NI_5 NS_670 0 -1.4855229397094541e-02
GC_5_671 b_5 NI_5 NS_671 0 -8.1250075395500106e-03
GC_5_672 b_5 NI_5 NS_672 0 1.9028461769214050e-03
GC_5_673 b_5 NI_5 NS_673 0 1.1255574772855150e-02
GC_5_674 b_5 NI_5 NS_674 0 -1.8013331580535811e-03
GC_5_675 b_5 NI_5 NS_675 0 -7.5649379527732664e-03
GC_5_676 b_5 NI_5 NS_676 0 -1.6931181123028536e-03
GC_5_677 b_5 NI_5 NS_677 0 1.5263484583700327e-02
GC_5_678 b_5 NI_5 NS_678 0 5.3089269192999767e-03
GC_5_679 b_5 NI_5 NS_679 0 -1.3074208595461078e-02
GC_5_680 b_5 NI_5 NS_680 0 -5.4740973546442582e-03
GC_5_681 b_5 NI_5 NS_681 0 -6.6401728312199338e-03
GC_5_682 b_5 NI_5 NS_682 0 3.4469264611769962e-03
GC_5_683 b_5 NI_5 NS_683 0 6.3571561981593276e-03
GC_5_684 b_5 NI_5 NS_684 0 -1.8769364689314126e-03
GC_5_685 b_5 NI_5 NS_685 0 -5.4767784277633446e-03
GC_5_686 b_5 NI_5 NS_686 0 2.1761635009273222e-03
GC_5_687 b_5 NI_5 NS_687 0 5.3904709118370881e-03
GC_5_688 b_5 NI_5 NS_688 0 -2.6291409473562077e-03
GC_5_689 b_5 NI_5 NS_689 0 -6.3068613159885222e-03
GC_5_690 b_5 NI_5 NS_690 0 -4.8944545977235097e-04
GC_5_691 b_5 NI_5 NS_691 0 7.6383029679271538e-03
GC_5_692 b_5 NI_5 NS_692 0 3.6283278652218857e-03
GC_5_693 b_5 NI_5 NS_693 0 -5.8333234857385037e-03
GC_5_694 b_5 NI_5 NS_694 0 -3.4684301852644281e-03
GC_5_695 b_5 NI_5 NS_695 0 2.9592189498357574e-04
GC_5_696 b_5 NI_5 NS_696 0 5.5702925731862052e-04
GC_5_697 b_5 NI_5 NS_697 0 -4.9284028648938971e-03
GC_5_698 b_5 NI_5 NS_698 0 8.8733927749231483e-04
GC_5_699 b_5 NI_5 NS_699 0 6.2016451885352425e-03
GC_5_700 b_5 NI_5 NS_700 0 6.8248095452396503e-04
GC_5_701 b_5 NI_5 NS_701 0 -5.3226827125023987e-03
GC_5_702 b_5 NI_5 NS_702 0 -4.8918923172088262e-04
GC_5_703 b_5 NI_5 NS_703 0 1.5482736461424884e-03
GC_5_704 b_5 NI_5 NS_704 0 -4.6609139366061315e-05
GC_5_705 b_5 NI_5 NS_705 0 -6.0242735099147451e-03
GC_5_706 b_5 NI_5 NS_706 0 1.9161515657498500e-03
GC_5_707 b_5 NI_5 NS_707 0 6.2494033097373145e-03
GC_5_708 b_5 NI_5 NS_708 0 2.0850478901550696e-04
GC_5_709 b_5 NI_5 NS_709 0 -5.0636589797219888e-03
GC_5_710 b_5 NI_5 NS_710 0 1.6954532442548021e-03
GC_5_711 b_5 NI_5 NS_711 0 2.4806587508526558e-03
GC_5_712 b_5 NI_5 NS_712 0 -9.6015729719484729e-04
GC_5_713 b_5 NI_5 NS_713 0 -6.5381321213501629e-03
GC_5_714 b_5 NI_5 NS_714 0 3.8750074616022089e-03
GC_5_715 b_5 NI_5 NS_715 0 7.4722546541904928e-03
GC_5_716 b_5 NI_5 NS_716 0 -1.0944729819690833e-03
GC_5_717 b_5 NI_5 NS_717 0 -3.9943218736883607e-03
GC_5_718 b_5 NI_5 NS_718 0 4.0357752344017212e-03
GC_5_719 b_5 NI_5 NS_719 0 2.8552013767554744e-03
GC_5_720 b_5 NI_5 NS_720 0 -3.0472624895247729e-03
GC_5_721 b_5 NI_5 NS_721 0 -6.0351388958252575e-03
GC_5_722 b_5 NI_5 NS_722 0 7.2276062148210708e-03
GC_5_723 b_5 NI_5 NS_723 0 7.9782887147297667e-03
GC_5_724 b_5 NI_5 NS_724 0 -4.7935801973900908e-03
GC_5_725 b_5 NI_5 NS_725 0 -5.4799474981508502e-04
GC_5_726 b_5 NI_5 NS_726 0 5.0230804901847453e-03
GC_5_727 b_5 NI_5 NS_727 0 2.5034134627312260e-04
GC_5_728 b_5 NI_5 NS_728 0 -4.7520661386946939e-03
GC_5_729 b_5 NI_5 NS_729 0 1.7366272814004955e-09
GC_5_730 b_5 NI_5 NS_730 0 3.2860222505116891e-09
GC_5_731 b_5 NI_5 NS_731 0 -1.4394125008007741e-03
GC_5_732 b_5 NI_5 NS_732 0 7.8706604761739993e-03
GC_5_733 b_5 NI_5 NS_733 0 -1.8574746928498709e-04
GC_5_734 b_5 NI_5 NS_734 0 3.0287972688731223e-03
GC_5_735 b_5 NI_5 NS_735 0 -1.2900533406370399e-04
GC_5_736 b_5 NI_5 NS_736 0 -3.3736684302623529e-03
GC_5_737 b_5 NI_5 NS_737 0 -8.9083181786645915e-04
GC_5_738 b_5 NI_5 NS_738 0 7.5293774121917489e-03
GC_5_739 b_5 NI_5 NS_739 0 3.7906243928354324e-03
GC_5_740 b_5 NI_5 NS_740 0 -6.1490577388279948e-03
GC_5_741 b_5 NI_5 NS_741 0 8.8448813607940954e-08
GC_5_742 b_5 NI_5 NS_742 0 -3.5531433518668937e-07
GC_5_743 b_5 NI_5 NS_743 0 6.7115065628059667e-03
GC_5_744 b_5 NI_5 NS_744 0 -5.3183245754123568e-03
GC_5_745 b_5 NI_5 NS_745 0 -2.6127433872478126e-03
GC_5_746 b_5 NI_5 NS_746 0 6.0487711501957652e-03
GC_5_747 b_5 NI_5 NS_747 0 -4.2945275038195549e-03
GC_5_748 b_5 NI_5 NS_748 0 1.3261562382255842e-05
GC_5_749 b_5 NI_5 NS_749 0 2.7224992724420630e-03
GC_5_750 b_5 NI_5 NS_750 0 -6.1956590818550697e-03
GC_5_751 b_5 NI_5 NS_751 0 2.0898364046733143e-03
GC_5_752 b_5 NI_5 NS_752 0 3.2611136183945248e-03
GC_5_753 b_5 NI_5 NS_753 0 -1.9638287424718617e-03
GC_5_754 b_5 NI_5 NS_754 0 -4.4203348237130367e-03
GC_5_755 b_5 NI_5 NS_755 0 2.8567435015331233e-03
GC_5_756 b_5 NI_5 NS_756 0 8.0017787545880875e-03
GC_5_757 b_5 NI_5 NS_757 0 -3.3198039925024744e-03
GC_5_758 b_5 NI_5 NS_758 0 1.8243968753581004e-09
GC_5_759 b_5 NI_5 NS_759 0 5.5833685855336323e-08
GC_5_760 b_5 NI_5 NS_760 0 1.8994901273373726e-06
GC_5_761 b_5 NI_5 NS_761 0 -9.0391646261060219e-05
GC_5_762 b_5 NI_5 NS_762 0 -5.8816388602288221e-05
GC_5_763 b_5 NI_5 NS_763 0 -1.2620480296526386e-03
GC_5_764 b_5 NI_5 NS_764 0 -3.0052300180571001e-04
GC_5_765 b_5 NI_5 NS_765 0 -1.6884323689189910e-03
GC_5_766 b_5 NI_5 NS_766 0 2.6375240550889274e-03
GC_5_767 b_5 NI_5 NS_767 0 4.9218035302901232e-04
GC_5_768 b_5 NI_5 NS_768 0 5.4232981892436936e-03
GC_5_769 b_5 NI_5 NS_769 0 7.0976984326468900e-03
GC_5_770 b_5 NI_5 NS_770 0 6.5580771105304783e-04
GC_5_771 b_5 NI_5 NS_771 0 6.4693545715985008e-04
GC_5_772 b_5 NI_5 NS_772 0 -6.5981442656357862e-04
GC_5_773 b_5 NI_5 NS_773 0 1.0491635774148079e-03
GC_5_774 b_5 NI_5 NS_774 0 1.5730867844146739e-03
GC_5_775 b_5 NI_5 NS_775 0 1.2639593608042806e-02
GC_5_776 b_5 NI_5 NS_776 0 1.3143543382593282e-02
GC_5_777 b_5 NI_5 NS_777 0 8.7648818791366927e-03
GC_5_778 b_5 NI_5 NS_778 0 -2.0356147037060263e-02
GC_5_779 b_5 NI_5 NS_779 0 8.3908943854833634e-03
GC_5_780 b_5 NI_5 NS_780 0 -2.8818702224687326e-03
GC_5_781 b_5 NI_5 NS_781 0 -1.2619354412556306e-02
GC_5_782 b_5 NI_5 NS_782 0 -3.8807125096877712e-02
GC_5_783 b_5 NI_5 NS_783 0 -7.2444869211372000e-03
GC_5_784 b_5 NI_5 NS_784 0 -2.1485688622041297e-03
GC_5_785 b_5 NI_5 NS_785 0 -5.2275000116047798e-02
GC_5_786 b_5 NI_5 NS_786 0 -1.8767871585090216e-03
GC_5_787 b_5 NI_5 NS_787 0 1.4892259635439470e-02
GC_5_788 b_5 NI_5 NS_788 0 8.6975590071554018e-03
GC_5_789 b_5 NI_5 NS_789 0 -5.9275337103615305e-03
GC_5_790 b_5 NI_5 NS_790 0 4.9905441852537867e-03
GC_5_791 b_5 NI_5 NS_791 0 8.3533718703616578e-03
GC_5_792 b_5 NI_5 NS_792 0 1.1690138985056022e-02
GC_5_793 b_5 NI_5 NS_793 0 4.5590097274008654e-03
GC_5_794 b_5 NI_5 NS_794 0 -2.9247916072175622e-03
GC_5_795 b_5 NI_5 NS_795 0 -7.8932468722468594e-03
GC_5_796 b_5 NI_5 NS_796 0 -8.1501572501387343e-03
GC_5_797 b_5 NI_5 NS_797 0 -5.6782670026900685e-03
GC_5_798 b_5 NI_5 NS_798 0 -6.1945380505947758e-04
GC_5_799 b_5 NI_5 NS_799 0 -1.8070910409072657e-02
GC_5_800 b_5 NI_5 NS_800 0 1.3562270005780287e-02
GC_5_801 b_5 NI_5 NS_801 0 4.7006670363791180e-03
GC_5_802 b_5 NI_5 NS_802 0 4.3832608836261930e-03
GC_5_803 b_5 NI_5 NS_803 0 6.4907980829625501e-04
GC_5_804 b_5 NI_5 NS_804 0 -1.1064122158182963e-04
GC_5_805 b_5 NI_5 NS_805 0 -3.7967884195648990e-03
GC_5_806 b_5 NI_5 NS_806 0 8.8034052685772961e-04
GC_5_807 b_5 NI_5 NS_807 0 -1.1248806791882666e-03
GC_5_808 b_5 NI_5 NS_808 0 1.6693625495463986e-02
GC_5_809 b_5 NI_5 NS_809 0 4.4443841515115498e-03
GC_5_810 b_5 NI_5 NS_810 0 7.1164003236733639e-04
GC_5_811 b_5 NI_5 NS_811 0 -5.2105034486662344e-04
GC_5_812 b_5 NI_5 NS_812 0 -2.2476782286137121e-03
GC_5_813 b_5 NI_5 NS_813 0 -4.9869185765197502e-03
GC_5_814 b_5 NI_5 NS_814 0 2.1058931891973485e-03
GC_5_815 b_5 NI_5 NS_815 0 7.3345854351600246e-03
GC_5_816 b_5 NI_5 NS_816 0 1.4346774371947495e-02
GC_5_817 b_5 NI_5 NS_817 0 4.1867521646059593e-03
GC_5_818 b_5 NI_5 NS_818 0 -1.6800211311655811e-03
GC_5_819 b_5 NI_5 NS_819 0 -3.3979285365229148e-03
GC_5_820 b_5 NI_5 NS_820 0 -2.1020210638149107e-03
GC_5_821 b_5 NI_5 NS_821 0 -5.4224785514777277e-03
GC_5_822 b_5 NI_5 NS_822 0 4.3763691523450027e-03
GC_5_823 b_5 NI_5 NS_823 0 1.3191411507258780e-02
GC_5_824 b_5 NI_5 NS_824 0 8.4408863585243576e-03
GC_5_825 b_5 NI_5 NS_825 0 2.8354700795776245e-03
GC_5_826 b_5 NI_5 NS_826 0 -4.1274251974683816e-03
GC_5_827 b_5 NI_5 NS_827 0 -5.3215591006486431e-03
GC_5_828 b_5 NI_5 NS_828 0 1.1333302092927839e-03
GC_5_829 b_5 NI_5 NS_829 0 -4.4370912591596813e-03
GC_5_830 b_5 NI_5 NS_830 0 8.3056987097559487e-03
GC_5_831 b_5 NI_5 NS_831 0 1.4614310663837527e-02
GC_5_832 b_5 NI_5 NS_832 0 -4.5696925783236212e-04
GC_5_833 b_5 NI_5 NS_833 0 -1.1788295639878674e-03
GC_5_834 b_5 NI_5 NS_834 0 -4.5487508143767525e-03
GC_5_835 b_5 NI_5 NS_835 0 -2.2870885713415106e-03
GC_5_836 b_5 NI_5 NS_836 0 4.3793440719547211e-03
GC_5_837 b_5 NI_5 NS_837 0 1.8255987381408038e-10
GC_5_838 b_5 NI_5 NS_838 0 -1.5799965964392498e-09
GC_5_839 b_5 NI_5 NS_839 0 1.4387717880472554e-03
GC_5_840 b_5 NI_5 NS_840 0 8.2177742617102652e-03
GC_5_841 b_5 NI_5 NS_841 0 -8.7491034135454512e-04
GC_5_842 b_5 NI_5 NS_842 0 -2.2094176122531822e-03
GC_5_843 b_5 NI_5 NS_843 0 -1.4716792699661382e-03
GC_5_844 b_5 NI_5 NS_844 0 2.7485700102958277e-03
GC_5_845 b_5 NI_5 NS_845 0 1.7223950961759811e-03
GC_5_846 b_5 NI_5 NS_846 0 7.6102898186978605e-03
GC_5_847 b_5 NI_5 NS_847 0 7.5930424197294087e-03
GC_5_848 b_5 NI_5 NS_848 0 -3.8216231340066609e-03
GC_5_849 b_5 NI_5 NS_849 0 -4.7008128148994605e-08
GC_5_850 b_5 NI_5 NS_850 0 -2.0170258569992724e-08
GC_5_851 b_5 NI_5 NS_851 0 1.1386078508495318e-02
GC_5_852 b_5 NI_5 NS_852 0 4.4716364341320690e-03
GC_5_853 b_5 NI_5 NS_853 0 -8.6429611410314194e-04
GC_5_854 b_5 NI_5 NS_854 0 6.4881769121089483e-03
GC_5_855 b_5 NI_5 NS_855 0 3.6256398048023632e-03
GC_5_856 b_5 NI_5 NS_856 0 4.0760137287815430e-04
GC_5_857 b_5 NI_5 NS_857 0 6.0652186093334403e-03
GC_5_858 b_5 NI_5 NS_858 0 -4.6566354048473303e-03
GC_5_859 b_5 NI_5 NS_859 0 -3.3846298119627350e-03
GC_5_860 b_5 NI_5 NS_860 0 -1.3607984935558853e-03
GC_5_861 b_5 NI_5 NS_861 0 1.0687130280415729e-04
GC_5_862 b_5 NI_5 NS_862 0 4.4902871968897379e-03
GC_5_863 b_5 NI_5 NS_863 0 7.2784000412120511e-03
GC_5_864 b_5 NI_5 NS_864 0 5.5303118943259661e-03
GC_5_865 b_5 NI_5 NS_865 0 -3.1809050707466072e-05
GC_5_866 b_5 NI_5 NS_866 0 -1.9490390401984754e-12
GC_5_867 b_5 NI_5 NS_867 0 -2.2738569976838423e-10
GC_5_868 b_5 NI_5 NS_868 0 1.0441851732479401e-08
GC_5_869 b_5 NI_5 NS_869 0 6.8674753760868464e-07
GC_5_870 b_5 NI_5 NS_870 0 1.0912849435263397e-07
GC_5_871 b_5 NI_5 NS_871 0 3.1464725378091258e-06
GC_5_872 b_5 NI_5 NS_872 0 -1.3843757425220467e-06
GC_5_873 b_5 NI_5 NS_873 0 -2.7797116731035317e-06
GC_5_874 b_5 NI_5 NS_874 0 -2.8013710424197283e-06
GC_5_875 b_5 NI_5 NS_875 0 4.9066013913795574e-06
GC_5_876 b_5 NI_5 NS_876 0 -5.2640981766404766e-07
GC_5_877 b_5 NI_5 NS_877 0 -7.0388976805970758e-06
GC_5_878 b_5 NI_5 NS_878 0 -8.0734843311859329e-06
GC_5_879 b_5 NI_5 NS_879 0 1.9914092042476401e-08
GC_5_880 b_5 NI_5 NS_880 0 -1.5400079655763619e-06
GC_5_881 b_5 NI_5 NS_881 0 -6.0451837551004206e-06
GC_5_882 b_5 NI_5 NS_882 0 1.9318156784611940e-06
GC_5_883 b_5 NI_5 NS_883 0 5.2997095889031462e-06
GC_5_884 b_5 NI_5 NS_884 0 -5.7096593413725797e-06
GC_5_885 b_5 NI_5 NS_885 0 -1.7020825321890775e-05
GC_5_886 b_5 NI_5 NS_886 0 4.6231739505253500e-06
GC_5_887 b_5 NI_5 NS_887 0 -1.1776749853274284e-06
GC_5_888 b_5 NI_5 NS_888 0 7.0415494665373178e-06
GC_5_889 b_5 NI_5 NS_889 0 -7.1892211460938741e-06
GC_5_890 b_5 NI_5 NS_890 0 -4.5422175065990794e-06
GC_5_891 b_5 NI_5 NS_891 0 -3.3644348848783349e-06
GC_5_892 b_5 NI_5 NS_892 0 7.9554426210622396e-06
GC_5_893 b_5 NI_5 NS_893 0 -2.2172645679678832e-06
GC_5_894 b_5 NI_5 NS_894 0 -4.6363872514452477e-06
GC_5_895 b_5 NI_5 NS_895 0 -3.8558757185374009e-06
GC_5_896 b_5 NI_5 NS_896 0 1.1253137134828167e-05
GC_5_897 b_5 NI_5 NS_897 0 -1.8103182322886142e-07
GC_5_898 b_5 NI_5 NS_898 0 7.1456890704382815e-06
GC_5_899 b_5 NI_5 NS_899 0 -4.1163603098235845e-06
GC_5_900 b_5 NI_5 NS_900 0 1.2239891599612041e-06
GC_5_901 b_5 NI_5 NS_901 0 -6.2986801157470296e-07
GC_5_902 b_5 NI_5 NS_902 0 7.9394007261406871e-06
GC_5_903 b_5 NI_5 NS_903 0 -1.0416947590537041e-06
GC_5_904 b_5 NI_5 NS_904 0 2.1882196166804060e-06
GC_5_905 b_5 NI_5 NS_905 0 -2.4107593993418067e-06
GC_5_906 b_5 NI_5 NS_906 0 8.0524123775358310e-06
GC_5_907 b_5 NI_5 NS_907 0 -1.5236719960058870e-07
GC_5_908 b_5 NI_5 NS_908 0 9.4057513161360350e-06
GC_5_909 b_5 NI_5 NS_909 0 -8.6008111999686094e-07
GC_5_910 b_5 NI_5 NS_910 0 8.6777424917871562e-06
GC_5_911 b_5 NI_5 NS_911 0 -1.3290770441354495e-06
GC_5_912 b_5 NI_5 NS_912 0 3.8594416325902931e-06
GC_5_913 b_5 NI_5 NS_913 0 9.6762987851128415e-07
GC_5_914 b_5 NI_5 NS_914 0 1.1812355584335796e-05
GC_5_915 b_5 NI_5 NS_915 0 1.7367411962011645e-05
GC_5_916 b_5 NI_5 NS_916 0 1.6606439351076272e-05
GC_5_917 b_5 NI_5 NS_917 0 4.7005654356617000e-06
GC_5_918 b_5 NI_5 NS_918 0 7.6012303201727736e-06
GC_5_919 b_5 NI_5 NS_919 0 9.8175726513465718e-06
GC_5_920 b_5 NI_5 NS_920 0 3.8200672239744041e-06
GC_5_921 b_5 NI_5 NS_921 0 6.4427117644219978e-06
GC_5_922 b_5 NI_5 NS_922 0 1.0581086680910590e-05
GC_5_923 b_5 NI_5 NS_923 0 3.1909373780162660e-05
GC_5_924 b_5 NI_5 NS_924 0 -5.8429969212007027e-06
GC_5_925 b_5 NI_5 NS_925 0 7.7884071350338152e-06
GC_5_926 b_5 NI_5 NS_926 0 3.3158520597456623e-06
GC_5_927 b_5 NI_5 NS_927 0 1.1397116905717714e-05
GC_5_928 b_5 NI_5 NS_928 0 -9.9644755546783236e-06
GC_5_929 b_5 NI_5 NS_929 0 1.0344054145509380e-05
GC_5_930 b_5 NI_5 NS_930 0 6.2012168901384595e-06
GC_5_931 b_5 NI_5 NS_931 0 1.5863181650405394e-05
GC_5_932 b_5 NI_5 NS_932 0 -2.9905472214178180e-05
GC_5_933 b_5 NI_5 NS_933 0 7.7033687022619373e-06
GC_5_934 b_5 NI_5 NS_934 0 -2.9069265194729339e-06
GC_5_935 b_5 NI_5 NS_935 0 -3.4527982236542116e-06
GC_5_936 b_5 NI_5 NS_936 0 -1.5725352623950357e-05
GC_5_937 b_5 NI_5 NS_937 0 1.1298999474062330e-05
GC_5_938 b_5 NI_5 NS_938 0 -1.7523101999553523e-06
GC_5_939 b_5 NI_5 NS_939 0 -1.3023508889495958e-05
GC_5_940 b_5 NI_5 NS_940 0 -2.4164323797338041e-05
GC_5_941 b_5 NI_5 NS_941 0 -4.2518814144261436e-07
GC_5_942 b_5 NI_5 NS_942 0 -6.4081584265917462e-06
GC_5_943 b_5 NI_5 NS_943 0 -9.5225953904404882e-06
GC_5_944 b_5 NI_5 NS_944 0 -2.3446767556538479e-06
GC_5_945 b_5 NI_5 NS_945 0 9.7513662028752994e-11
GC_5_946 b_5 NI_5 NS_946 0 5.3586384235852980e-11
GC_5_947 b_5 NI_5 NS_947 0 1.1849077792164896e-06
GC_5_948 b_5 NI_5 NS_948 0 -4.6339012513416611e-06
GC_5_949 b_5 NI_5 NS_949 0 -1.4863761372252775e-06
GC_5_950 b_5 NI_5 NS_950 0 -1.2907052113210419e-06
GC_5_951 b_5 NI_5 NS_951 0 -4.9349921847861124e-06
GC_5_952 b_5 NI_5 NS_952 0 -8.8189364173378315e-07
GC_5_953 b_5 NI_5 NS_953 0 -1.3866100504970447e-06
GC_5_954 b_5 NI_5 NS_954 0 -2.8415046981362699e-06
GC_5_955 b_5 NI_5 NS_955 0 -1.0079602382041263e-05
GC_5_956 b_5 NI_5 NS_956 0 -3.7053039984008183e-06
GC_5_957 b_5 NI_5 NS_957 0 6.6047302988678779e-09
GC_5_958 b_5 NI_5 NS_958 0 5.7466233902049664e-09
GC_5_959 b_5 NI_5 NS_959 0 1.3885986402599670e-06
GC_5_960 b_5 NI_5 NS_960 0 6.7923813461897890e-07
GC_5_961 b_5 NI_5 NS_961 0 -1.7365102029104155e-06
GC_5_962 b_5 NI_5 NS_962 0 3.1379191364764467e-06
GC_5_963 b_5 NI_5 NS_963 0 -9.2489884019493506e-07
GC_5_964 b_5 NI_5 NS_964 0 7.7500977441745498e-07
GC_5_965 b_5 NI_5 NS_965 0 -7.9023121935105756e-06
GC_5_966 b_5 NI_5 NS_966 0 8.1042211466053426e-07
GC_5_967 b_5 NI_5 NS_967 0 -2.4148798686970143e-06
GC_5_968 b_5 NI_5 NS_968 0 2.0815635515205955e-06
GC_5_969 b_5 NI_5 NS_969 0 -2.1260358996063536e-06
GC_5_970 b_5 NI_5 NS_970 0 2.1321344840876506e-06
GC_5_971 b_5 NI_5 NS_971 0 1.1301417882064136e-06
GC_5_972 b_5 NI_5 NS_972 0 2.8148321275733345e-06
GC_5_973 b_5 NI_5 NS_973 0 -1.4324500380219547e-04
GC_5_974 b_5 NI_5 NS_974 0 3.4599473571614782e-11
GC_5_975 b_5 NI_5 NS_975 0 3.0173663891791482e-11
GC_5_976 b_5 NI_5 NS_976 0 9.4206038963802704e-10
GC_5_977 b_5 NI_5 NS_977 0 -2.1091116959165087e-06
GC_5_978 b_5 NI_5 NS_978 0 -1.6534028724614032e-06
GC_5_979 b_5 NI_5 NS_979 0 1.8892523755874762e-06
GC_5_980 b_5 NI_5 NS_980 0 3.8450015283065862e-06
GC_5_981 b_5 NI_5 NS_981 0 3.2880765294835146e-06
GC_5_982 b_5 NI_5 NS_982 0 4.9269026901413863e-06
GC_5_983 b_5 NI_5 NS_983 0 5.8303571902268804e-06
GC_5_984 b_5 NI_5 NS_984 0 -9.0831336686623214e-06
GC_5_985 b_5 NI_5 NS_985 0 -2.5401415892311689e-06
GC_5_986 b_5 NI_5 NS_986 0 -1.3835998140381580e-05
GC_5_987 b_5 NI_5 NS_987 0 -3.5342191349266796e-06
GC_5_988 b_5 NI_5 NS_988 0 2.1965955541030162e-06
GC_5_989 b_5 NI_5 NS_989 0 3.6390210417131202e-06
GC_5_990 b_5 NI_5 NS_990 0 1.2969577615512131e-06
GC_5_991 b_5 NI_5 NS_991 0 7.8997062474368431e-06
GC_5_992 b_5 NI_5 NS_992 0 -3.9683455453607296e-05
GC_5_993 b_5 NI_5 NS_993 0 -4.4005697692644987e-05
GC_5_994 b_5 NI_5 NS_994 0 -8.8267547488270765e-07
GC_5_995 b_5 NI_5 NS_995 0 -1.4766095927885207e-05
GC_5_996 b_5 NI_5 NS_996 0 -8.4725268772861232e-06
GC_5_997 b_5 NI_5 NS_997 0 -7.2348297877387015e-05
GC_5_998 b_5 NI_5 NS_998 0 7.5140020331099233e-05
GC_5_999 b_5 NI_5 NS_999 0 4.6496225986729384e-06
GC_5_1000 b_5 NI_5 NS_1000 0 1.3009889495946494e-05
GC_5_1001 b_5 NI_5 NS_1001 0 6.2664902534681778e-05
GC_5_1002 b_5 NI_5 NS_1002 0 1.2224106210300409e-04
GC_5_1003 b_5 NI_5 NS_1003 0 2.4432197370250135e-07
GC_5_1004 b_5 NI_5 NS_1004 0 -3.6753046295622540e-05
GC_5_1005 b_5 NI_5 NS_1005 0 1.6411265154984306e-05
GC_5_1006 b_5 NI_5 NS_1006 0 3.8870370418552697e-06
GC_5_1007 b_5 NI_5 NS_1007 0 2.4218757552749475e-05
GC_5_1008 b_5 NI_5 NS_1008 0 -3.0243863640212752e-05
GC_5_1009 b_5 NI_5 NS_1009 0 -8.8438563099807464e-06
GC_5_1010 b_5 NI_5 NS_1010 0 -2.2760871431871584e-06
GC_5_1011 b_5 NI_5 NS_1011 0 -8.7280252623841105e-06
GC_5_1012 b_5 NI_5 NS_1012 0 2.5050835882890535e-05
GC_5_1013 b_5 NI_5 NS_1013 0 5.8326426984655712e-06
GC_5_1014 b_5 NI_5 NS_1014 0 8.3787537054273868e-06
GC_5_1015 b_5 NI_5 NS_1015 0 5.5968994772007610e-05
GC_5_1016 b_5 NI_5 NS_1016 0 2.4647283369767361e-05
GC_5_1017 b_5 NI_5 NS_1017 0 3.4490090174253096e-06
GC_5_1018 b_5 NI_5 NS_1018 0 -1.1606186039572972e-05
GC_5_1019 b_5 NI_5 NS_1019 0 -4.0624008989515026e-07
GC_5_1020 b_5 NI_5 NS_1020 0 -1.2992030596488547e-06
GC_5_1021 b_5 NI_5 NS_1021 0 6.7879577288158105e-06
GC_5_1022 b_5 NI_5 NS_1022 0 3.0205385640306798e-06
GC_5_1023 b_5 NI_5 NS_1023 0 4.1591506177496160e-05
GC_5_1024 b_5 NI_5 NS_1024 0 -1.7165542425075311e-05
GC_5_1025 b_5 NI_5 NS_1025 0 -2.5739597184849548e-06
GC_5_1026 b_5 NI_5 NS_1026 0 -7.0282411742968846e-06
GC_5_1027 b_5 NI_5 NS_1027 0 -2.9900893039212231e-06
GC_5_1028 b_5 NI_5 NS_1028 0 1.7603745498449645e-06
GC_5_1029 b_5 NI_5 NS_1029 0 9.5385282655802944e-06
GC_5_1030 b_5 NI_5 NS_1030 0 2.8682641162255170e-06
GC_5_1031 b_5 NI_5 NS_1031 0 2.2731271067177940e-05
GC_5_1032 b_5 NI_5 NS_1032 0 -3.1037336893354611e-05
GC_5_1033 b_5 NI_5 NS_1033 0 -5.6871990009354142e-06
GC_5_1034 b_5 NI_5 NS_1034 0 -3.6245405822499859e-06
GC_5_1035 b_5 NI_5 NS_1035 0 -5.2395264627103735e-07
GC_5_1036 b_5 NI_5 NS_1036 0 5.0176484733036418e-06
GC_5_1037 b_5 NI_5 NS_1037 0 1.2253629391960900e-05
GC_5_1038 b_5 NI_5 NS_1038 0 1.7526939844932501e-07
GC_5_1039 b_5 NI_5 NS_1039 0 1.8081527934614634e-06
GC_5_1040 b_5 NI_5 NS_1040 0 -3.1349647117597911e-05
GC_5_1041 b_5 NI_5 NS_1041 0 -6.7180786310030063e-06
GC_5_1042 b_5 NI_5 NS_1042 0 9.7556402818652511e-07
GC_5_1043 b_5 NI_5 NS_1043 0 4.6118370397777717e-06
GC_5_1044 b_5 NI_5 NS_1044 0 3.8655506612082002e-06
GC_5_1045 b_5 NI_5 NS_1045 0 1.4061774515849650e-05
GC_5_1046 b_5 NI_5 NS_1046 0 -6.0101893326935314e-06
GC_5_1047 b_5 NI_5 NS_1047 0 -1.4015860251487117e-05
GC_5_1048 b_5 NI_5 NS_1048 0 -1.8746808369529216e-05
GC_5_1049 b_5 NI_5 NS_1049 0 -2.5061548171875972e-06
GC_5_1050 b_5 NI_5 NS_1050 0 5.4162611603888574e-06
GC_5_1051 b_5 NI_5 NS_1051 0 4.6576647463596257e-06
GC_5_1052 b_5 NI_5 NS_1052 0 -2.0834586716042294e-06
GC_5_1053 b_5 NI_5 NS_1053 0 -1.4566104014408751e-11
GC_5_1054 b_5 NI_5 NS_1054 0 4.2060567854290715e-12
GC_5_1055 b_5 NI_5 NS_1055 0 5.1979378859549864e-06
GC_5_1056 b_5 NI_5 NS_1056 0 -1.1242581694578139e-05
GC_5_1057 b_5 NI_5 NS_1057 0 -2.6677232273252252e-07
GC_5_1058 b_5 NI_5 NS_1058 0 2.9264734339676127e-06
GC_5_1059 b_5 NI_5 NS_1059 0 2.6444997765484435e-06
GC_5_1060 b_5 NI_5 NS_1060 0 -1.5935804591335003e-06
GC_5_1061 b_5 NI_5 NS_1061 0 2.4075836161090012e-06
GC_5_1062 b_5 NI_5 NS_1062 0 -9.4308013894483517e-06
GC_5_1063 b_5 NI_5 NS_1063 0 -9.9265769593262262e-06
GC_5_1064 b_5 NI_5 NS_1064 0 -3.6883871433070661e-06
GC_5_1065 b_5 NI_5 NS_1065 0 3.1234687508275058e-10
GC_5_1066 b_5 NI_5 NS_1066 0 2.7704382613669457e-10
GC_5_1067 b_5 NI_5 NS_1067 0 -8.5916123125267823e-06
GC_5_1068 b_5 NI_5 NS_1068 0 -5.6864936881821168e-06
GC_5_1069 b_5 NI_5 NS_1069 0 2.2662274440573806e-06
GC_5_1070 b_5 NI_5 NS_1070 0 -6.4520070786707974e-06
GC_5_1071 b_5 NI_5 NS_1071 0 -3.0674012730352132e-06
GC_5_1072 b_5 NI_5 NS_1072 0 -1.3540170638295837e-07
GC_5_1073 b_5 NI_5 NS_1073 0 -7.9220201917139825e-06
GC_5_1074 b_5 NI_5 NS_1074 0 4.8459808285623915e-07
GC_5_1075 b_5 NI_5 NS_1075 0 3.0018508517120846e-06
GC_5_1076 b_5 NI_5 NS_1076 0 2.8730914602888175e-06
GC_5_1077 b_5 NI_5 NS_1077 0 1.2172132117031266e-06
GC_5_1078 b_5 NI_5 NS_1078 0 -3.8814880044022713e-06
GC_5_1079 b_5 NI_5 NS_1079 0 -4.8738054257528034e-06
GC_5_1080 b_5 NI_5 NS_1080 0 -3.9067778766128591e-06
GC_5_1081 b_5 NI_5 NS_1081 0 4.9610769508727464e-05
GC_5_1082 b_5 NI_5 NS_1082 0 3.6353121941747932e-12
GC_5_1083 b_5 NI_5 NS_1083 0 -4.1275403872199043e-12
GC_5_1084 b_5 NI_5 NS_1084 0 9.4606198639672796e-10
GC_5_1085 b_5 NI_5 NS_1085 0 -4.5694206184659050e-08
GC_5_1086 b_5 NI_5 NS_1086 0 2.5276728648265008e-07
GC_5_1087 b_5 NI_5 NS_1087 0 2.5906308305402562e-07
GC_5_1088 b_5 NI_5 NS_1088 0 4.0752866883473338e-07
GC_5_1089 b_5 NI_5 NS_1089 0 -1.3716182147504986e-07
GC_5_1090 b_5 NI_5 NS_1090 0 2.4384810115541381e-07
GC_5_1091 b_5 NI_5 NS_1091 0 7.8139024906597565e-07
GC_5_1092 b_5 NI_5 NS_1092 0 1.4415702305307190e-06
GC_5_1093 b_5 NI_5 NS_1093 0 1.0388733017956534e-06
GC_5_1094 b_5 NI_5 NS_1094 0 -5.2228255958991420e-07
GC_5_1095 b_5 NI_5 NS_1095 0 3.3588430584802711e-07
GC_5_1096 b_5 NI_5 NS_1096 0 8.8677767719493939e-07
GC_5_1097 b_5 NI_5 NS_1097 0 7.3258458483516767e-07
GC_5_1098 b_5 NI_5 NS_1098 0 -3.6895400717544838e-07
GC_5_1099 b_5 NI_5 NS_1099 0 4.3580341521829827e-06
GC_5_1100 b_5 NI_5 NS_1100 0 1.3814609520464018e-06
GC_5_1101 b_5 NI_5 NS_1101 0 -1.6431406325979375e-06
GC_5_1102 b_5 NI_5 NS_1102 0 -3.5781604284357628e-06
GC_5_1103 b_5 NI_5 NS_1103 0 2.3983176289007830e-07
GC_5_1104 b_5 NI_5 NS_1104 0 1.5513164273160372e-06
GC_5_1105 b_5 NI_5 NS_1105 0 2.9719508700035177e-06
GC_5_1106 b_5 NI_5 NS_1106 0 -4.7485563200803433e-06
GC_5_1107 b_5 NI_5 NS_1107 0 -7.7194427121330878e-07
GC_5_1108 b_5 NI_5 NS_1108 0 5.6548804144580451e-07
GC_5_1109 b_5 NI_5 NS_1109 0 5.5722019300009603e-06
GC_5_1110 b_5 NI_5 NS_1110 0 -5.8225124050867622e-06
GC_5_1111 b_5 NI_5 NS_1111 0 -3.3127672387083493e-06
GC_5_1112 b_5 NI_5 NS_1112 0 1.7944209292543809e-06
GC_5_1113 b_5 NI_5 NS_1113 0 8.6215716514200266e-07
GC_5_1114 b_5 NI_5 NS_1114 0 1.2284625509047816e-06
GC_5_1115 b_5 NI_5 NS_1115 0 1.5941346086318947e-06
GC_5_1116 b_5 NI_5 NS_1116 0 -4.1010700697514810e-06
GC_5_1117 b_5 NI_5 NS_1117 0 5.6926932086369470e-07
GC_5_1118 b_5 NI_5 NS_1118 0 1.9922746638593427e-07
GC_5_1119 b_5 NI_5 NS_1119 0 1.7434077086407334e-07
GC_5_1120 b_5 NI_5 NS_1120 0 -4.0363605740056077e-06
GC_5_1121 b_5 NI_5 NS_1121 0 -1.8756594344802056e-07
GC_5_1122 b_5 NI_5 NS_1122 0 1.6761079479975665e-07
GC_5_1123 b_5 NI_5 NS_1123 0 4.6377166523988987e-06
GC_5_1124 b_5 NI_5 NS_1124 0 -6.3334423871300974e-06
GC_5_1125 b_5 NI_5 NS_1125 0 -1.8278214271029545e-06
GC_5_1126 b_5 NI_5 NS_1126 0 -1.2890013763813488e-06
GC_5_1127 b_5 NI_5 NS_1127 0 1.3669191877985715e-06
GC_5_1128 b_5 NI_5 NS_1128 0 -1.1985544267038203e-06
GC_5_1129 b_5 NI_5 NS_1129 0 3.7643259693551039e-07
GC_5_1130 b_5 NI_5 NS_1130 0 -2.0976084981038473e-06
GC_5_1131 b_5 NI_5 NS_1131 0 -1.4875487463781504e-06
GC_5_1132 b_5 NI_5 NS_1132 0 -1.1765894486922943e-05
GC_5_1133 b_5 NI_5 NS_1133 0 -2.2683515217877669e-06
GC_5_1134 b_5 NI_5 NS_1134 0 -1.7024968684475503e-06
GC_5_1135 b_5 NI_5 NS_1135 0 -2.3842940128457256e-06
GC_5_1136 b_5 NI_5 NS_1136 0 -3.9896434497983449e-06
GC_5_1137 b_5 NI_5 NS_1137 0 -1.4876626407255775e-06
GC_5_1138 b_5 NI_5 NS_1138 0 -2.4187941278018903e-06
GC_5_1139 b_5 NI_5 NS_1139 0 -1.0716987004839735e-05
GC_5_1140 b_5 NI_5 NS_1140 0 -7.0850928150889791e-06
GC_5_1141 b_5 NI_5 NS_1141 0 -3.1909448110685312e-06
GC_5_1142 b_5 NI_5 NS_1142 0 -8.5674753336687902e-07
GC_5_1143 b_5 NI_5 NS_1143 0 -5.7476367317748253e-06
GC_5_1144 b_5 NI_5 NS_1144 0 -3.7004872950864556e-07
GC_5_1145 b_5 NI_5 NS_1145 0 -3.1243750307506384e-06
GC_5_1146 b_5 NI_5 NS_1146 0 -1.7461463944176146e-06
GC_5_1147 b_5 NI_5 NS_1147 0 -1.0618663970624777e-05
GC_5_1148 b_5 NI_5 NS_1148 0 3.3753555323240909e-06
GC_5_1149 b_5 NI_5 NS_1149 0 -3.6318005899305165e-06
GC_5_1150 b_5 NI_5 NS_1150 0 8.3009919347028713e-07
GC_5_1151 b_5 NI_5 NS_1151 0 -2.8719522602523983e-06
GC_5_1152 b_5 NI_5 NS_1152 0 3.9430649361726366e-06
GC_5_1153 b_5 NI_5 NS_1153 0 -4.3595838526945594e-06
GC_5_1154 b_5 NI_5 NS_1154 0 1.7264986832051806e-07
GC_5_1155 b_5 NI_5 NS_1155 0 -1.8585267206770095e-06
GC_5_1156 b_5 NI_5 NS_1156 0 7.2740539950004291e-06
GC_5_1157 b_5 NI_5 NS_1157 0 -1.5748460319934688e-06
GC_5_1158 b_5 NI_5 NS_1158 0 2.8115309732277503e-06
GC_5_1159 b_5 NI_5 NS_1159 0 9.3643793900051799e-07
GC_5_1160 b_5 NI_5 NS_1160 0 1.8337161088030159e-06
GC_5_1161 b_5 NI_5 NS_1161 0 -3.0124148066265677e-11
GC_5_1162 b_5 NI_5 NS_1162 0 -3.3889718508537135e-12
GC_5_1163 b_5 NI_5 NS_1163 0 -1.7319002978113763e-06
GC_5_1164 b_5 NI_5 NS_1164 0 2.1529086478862081e-06
GC_5_1165 b_5 NI_5 NS_1165 0 -3.2427999774036517e-07
GC_5_1166 b_5 NI_5 NS_1166 0 1.0583762842791571e-06
GC_5_1167 b_5 NI_5 NS_1167 0 1.4379977511016980e-07
GC_5_1168 b_5 NI_5 NS_1168 0 6.3880009269055626e-07
GC_5_1169 b_5 NI_5 NS_1169 0 -1.0428221756388901e-06
GC_5_1170 b_5 NI_5 NS_1170 0 1.2847611907104427e-06
GC_5_1171 b_5 NI_5 NS_1171 0 9.8816632690318800e-07
GC_5_1172 b_5 NI_5 NS_1172 0 1.8536017681276669e-06
GC_5_1173 b_5 NI_5 NS_1173 0 -1.5199216681472671e-09
GC_5_1174 b_5 NI_5 NS_1174 0 -7.6810688710888625e-10
GC_5_1175 b_5 NI_5 NS_1175 0 -4.6943560189078853e-07
GC_5_1176 b_5 NI_5 NS_1176 0 -2.3372188895553307e-08
GC_5_1177 b_5 NI_5 NS_1177 0 -3.1181061272296796e-07
GC_5_1178 b_5 NI_5 NS_1178 0 1.9126078472445136e-07
GC_5_1179 b_5 NI_5 NS_1179 0 -5.4910130440596450e-07
GC_5_1180 b_5 NI_5 NS_1180 0 1.5141086535733273e-07
GC_5_1181 b_5 NI_5 NS_1181 0 6.6188069255990298e-07
GC_5_1182 b_5 NI_5 NS_1182 0 8.2996733050997711e-07
GC_5_1183 b_5 NI_5 NS_1183 0 2.3288625603947868e-07
GC_5_1184 b_5 NI_5 NS_1184 0 7.0026446212826730e-07
GC_5_1185 b_5 NI_5 NS_1185 0 3.0416342861755592e-09
GC_5_1186 b_5 NI_5 NS_1186 0 -1.3243560290860395e-07
GC_5_1187 b_5 NI_5 NS_1187 0 -3.4705037948412107e-07
GC_5_1188 b_5 NI_5 NS_1188 0 2.9428852748773917e-07
GC_5_1189 b_5 NI_5 NS_1189 0 -9.0232877825115060e-05
GC_5_1190 b_5 NI_5 NS_1190 0 7.1467013071990092e-12
GC_5_1191 b_5 NI_5 NS_1191 0 -5.7273217091038376e-11
GC_5_1192 b_5 NI_5 NS_1192 0 3.3270910391803326e-10
GC_5_1193 b_5 NI_5 NS_1193 0 -1.5775944590719809e-06
GC_5_1194 b_5 NI_5 NS_1194 0 -1.5525971518782960e-06
GC_5_1195 b_5 NI_5 NS_1195 0 9.4591818046387876e-07
GC_5_1196 b_5 NI_5 NS_1196 0 7.1992586496871261e-07
GC_5_1197 b_5 NI_5 NS_1197 0 -2.7042590715342524e-06
GC_5_1198 b_5 NI_5 NS_1198 0 3.0432354429167001e-06
GC_5_1199 b_5 NI_5 NS_1199 0 -3.0477748103264628e-06
GC_5_1200 b_5 NI_5 NS_1200 0 -2.5663673687873772e-06
GC_5_1201 b_5 NI_5 NS_1201 0 1.5140920563295102e-06
GC_5_1202 b_5 NI_5 NS_1202 0 6.0866213157198107e-08
GC_5_1203 b_5 NI_5 NS_1203 0 -1.6616182595846968e-06
GC_5_1204 b_5 NI_5 NS_1204 0 1.7956761153321207e-06
GC_5_1205 b_5 NI_5 NS_1205 0 9.0473692849325610e-07
GC_5_1206 b_5 NI_5 NS_1206 0 4.1356084072413506e-06
GC_5_1207 b_5 NI_5 NS_1207 0 -4.2700433444902418e-06
GC_5_1208 b_5 NI_5 NS_1208 0 -2.0665822122434467e-06
GC_5_1209 b_5 NI_5 NS_1209 0 2.3210734973102237e-06
GC_5_1210 b_5 NI_5 NS_1210 0 -1.9750450209332317e-06
GC_5_1211 b_5 NI_5 NS_1211 0 -1.1664520699678532e-06
GC_5_1212 b_5 NI_5 NS_1212 0 3.2386758377356281e-06
GC_5_1213 b_5 NI_5 NS_1213 0 -8.4927520286743791e-06
GC_5_1214 b_5 NI_5 NS_1214 0 1.1257648125585625e-05
GC_5_1215 b_5 NI_5 NS_1215 0 1.2382783198447869e-06
GC_5_1216 b_5 NI_5 NS_1216 0 -1.6380405557689554e-06
GC_5_1217 b_5 NI_5 NS_1217 0 9.9626673938614572e-06
GC_5_1218 b_5 NI_5 NS_1218 0 1.7510966763208038e-05
GC_5_1219 b_5 NI_5 NS_1219 0 -6.2141837773581737e-07
GC_5_1220 b_5 NI_5 NS_1220 0 -5.7371616893058258e-07
GC_5_1221 b_5 NI_5 NS_1221 0 4.5338160558583943e-07
GC_5_1222 b_5 NI_5 NS_1222 0 -1.3531135909183950e-06
GC_5_1223 b_5 NI_5 NS_1223 0 7.0533203098096421e-06
GC_5_1224 b_5 NI_5 NS_1224 0 -2.6361049632125251e-07
GC_5_1225 b_5 NI_5 NS_1225 0 7.0541848804426509e-07
GC_5_1226 b_5 NI_5 NS_1226 0 2.9816704252497734e-06
GC_5_1227 b_5 NI_5 NS_1227 0 4.2391189212354968e-07
GC_5_1228 b_5 NI_5 NS_1228 0 2.9338682638322837e-06
GC_5_1229 b_5 NI_5 NS_1229 0 1.1537385045309060e-06
GC_5_1230 b_5 NI_5 NS_1230 0 -1.4005640884349448e-06
GC_5_1231 b_5 NI_5 NS_1231 0 9.4429281227096721e-06
GC_5_1232 b_5 NI_5 NS_1232 0 5.2402512330363894e-06
GC_5_1233 b_5 NI_5 NS_1233 0 5.8904321520130972e-07
GC_5_1234 b_5 NI_5 NS_1234 0 1.1278234826042982e-06
GC_5_1235 b_5 NI_5 NS_1235 0 5.5044039198564675e-08
GC_5_1236 b_5 NI_5 NS_1236 0 4.4723215058701425e-07
GC_5_1237 b_5 NI_5 NS_1237 0 1.2859222568804150e-06
GC_5_1238 b_5 NI_5 NS_1238 0 -8.4940917314410593e-07
GC_5_1239 b_5 NI_5 NS_1239 0 9.2174087148623965e-06
GC_5_1240 b_5 NI_5 NS_1240 0 6.4700432272287202e-07
GC_5_1241 b_5 NI_5 NS_1241 0 8.4642396979978098e-07
GC_5_1242 b_5 NI_5 NS_1242 0 1.4278789814611343e-06
GC_5_1243 b_5 NI_5 NS_1243 0 1.0142053963039248e-06
GC_5_1244 b_5 NI_5 NS_1244 0 5.9014676969571083e-07
GC_5_1245 b_5 NI_5 NS_1245 0 1.3671645043380007e-06
GC_5_1246 b_5 NI_5 NS_1246 0 -9.4667621377066751e-07
GC_5_1247 b_5 NI_5 NS_1247 0 8.0330915094369612e-06
GC_5_1248 b_5 NI_5 NS_1248 0 -2.1787314439574020e-06
GC_5_1249 b_5 NI_5 NS_1249 0 1.1742082142122271e-06
GC_5_1250 b_5 NI_5 NS_1250 0 1.5187612756113477e-06
GC_5_1251 b_5 NI_5 NS_1251 0 1.5705996199570524e-06
GC_5_1252 b_5 NI_5 NS_1252 0 -2.4568000382133330e-07
GC_5_1253 b_5 NI_5 NS_1253 0 1.3311045867753754e-06
GC_5_1254 b_5 NI_5 NS_1254 0 -9.9726141044698983e-07
GC_5_1255 b_5 NI_5 NS_1255 0 5.8014304506780170e-06
GC_5_1256 b_5 NI_5 NS_1256 0 -3.9293700911953047e-06
GC_5_1257 b_5 NI_5 NS_1257 0 1.8001462617514058e-06
GC_5_1258 b_5 NI_5 NS_1258 0 1.4046092474634346e-06
GC_5_1259 b_5 NI_5 NS_1259 0 1.0780223406766326e-06
GC_5_1260 b_5 NI_5 NS_1260 0 -1.3987160049828048e-06
GC_5_1261 b_5 NI_5 NS_1261 0 1.4203326975237917e-06
GC_5_1262 b_5 NI_5 NS_1262 0 -1.1295810304691442e-06
GC_5_1263 b_5 NI_5 NS_1263 0 2.9391253217581523e-06
GC_5_1264 b_5 NI_5 NS_1264 0 -4.1900348020136791e-06
GC_5_1265 b_5 NI_5 NS_1265 0 2.2053962291695500e-06
GC_5_1266 b_5 NI_5 NS_1266 0 2.9635278070926982e-07
GC_5_1267 b_5 NI_5 NS_1267 0 -3.3186776888187816e-07
GC_5_1268 b_5 NI_5 NS_1268 0 -1.1800073799302886e-06
GC_5_1269 b_5 NI_5 NS_1269 0 2.4885396467374965e-11
GC_5_1270 b_5 NI_5 NS_1270 0 -4.0917300699322786e-11
GC_5_1271 b_5 NI_5 NS_1271 0 7.9132856034260195e-07
GC_5_1272 b_5 NI_5 NS_1272 0 -1.5907614899351386e-06
GC_5_1273 b_5 NI_5 NS_1273 0 1.2547876777595839e-06
GC_5_1274 b_5 NI_5 NS_1274 0 2.2340461672200087e-07
GC_5_1275 b_5 NI_5 NS_1275 0 1.5908914308320766e-07
GC_5_1276 b_5 NI_5 NS_1276 0 -5.4772244277578070e-07
GC_5_1277 b_5 NI_5 NS_1277 0 5.4957109692567103e-07
GC_5_1278 b_5 NI_5 NS_1278 0 -8.9267217440285703e-07
GC_5_1279 b_5 NI_5 NS_1279 0 1.2802186837889362e-06
GC_5_1280 b_5 NI_5 NS_1280 0 -2.0630237924034743e-06
GC_5_1281 b_5 NI_5 NS_1281 0 4.7395124356503020e-10
GC_5_1282 b_5 NI_5 NS_1282 0 -1.2084264413572410e-09
GC_5_1283 b_5 NI_5 NS_1283 0 5.4791635479142101e-07
GC_5_1284 b_5 NI_5 NS_1284 0 -8.5973170907038488e-07
GC_5_1285 b_5 NI_5 NS_1285 0 7.1441929942668513e-07
GC_5_1286 b_5 NI_5 NS_1286 0 -9.5097395359591102e-07
GC_5_1287 b_5 NI_5 NS_1287 0 8.9079197421095627e-08
GC_5_1288 b_5 NI_5 NS_1288 0 5.0128483930444493e-08
GC_5_1289 b_5 NI_5 NS_1289 0 1.3250939373720850e-06
GC_5_1290 b_5 NI_5 NS_1290 0 -1.2292257183408871e-06
GC_5_1291 b_5 NI_5 NS_1291 0 1.6446054161061553e-06
GC_5_1292 b_5 NI_5 NS_1292 0 -2.9221557614978623e-07
GC_5_1293 b_5 NI_5 NS_1293 0 -2.2768019052200262e-07
GC_5_1294 b_5 NI_5 NS_1294 0 -7.3422400131587217e-07
GC_5_1295 b_5 NI_5 NS_1295 0 7.3335515226528001e-07
GC_5_1296 b_5 NI_5 NS_1296 0 2.8942335427168216e-07
GD_5_1 b_5 NI_5 NA_1 0 3.1568031929873996e-06
GD_5_2 b_5 NI_5 NA_2 0 1.9212503432668103e-05
GD_5_3 b_5 NI_5 NA_3 0 2.2219405014701666e-05
GD_5_4 b_5 NI_5 NA_4 0 1.0510731021863832e-04
GD_5_5 b_5 NI_5 NA_5 0 -1.1040269116041893e-02
GD_5_6 b_5 NI_5 NA_6 0 -4.9039917843811710e-03
GD_5_7 b_5 NI_5 NA_7 0 1.0577033561008323e-02
GD_5_8 b_5 NI_5 NA_8 0 -1.1498023026324552e-03
GD_5_9 b_5 NI_5 NA_9 0 5.7656796858531710e-08
GD_5_10 b_5 NI_5 NA_10 0 1.5903951218009538e-05
GD_5_11 b_5 NI_5 NA_11 0 -3.0002492085413852e-06
GD_5_12 b_5 NI_5 NA_12 0 1.1439017509924456e-05
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 -1.5264055326223407e-04
GC_6_2 b_6 NI_6 NS_2 0 3.6649219803697083e-11
GC_6_3 b_6 NI_6 NS_3 0 1.8927494314323008e-11
GC_6_4 b_6 NI_6 NS_4 0 9.3057798034707992e-10
GC_6_5 b_6 NI_6 NS_5 0 -2.3228432578438686e-06
GC_6_6 b_6 NI_6 NS_6 0 -1.6428402506813695e-06
GC_6_7 b_6 NI_6 NS_7 0 1.4316459214251428e-06
GC_6_8 b_6 NI_6 NS_8 0 3.8987608731532415e-06
GC_6_9 b_6 NI_6 NS_9 0 3.0058872501592151e-06
GC_6_10 b_6 NI_6 NS_10 0 5.4029766610785840e-06
GC_6_11 b_6 NI_6 NS_11 0 5.4599115334325571e-06
GC_6_12 b_6 NI_6 NS_12 0 -8.4815370286447683e-06
GC_6_13 b_6 NI_6 NS_13 0 -2.3141908628278624e-06
GC_6_14 b_6 NI_6 NS_14 0 -1.2723706123326921e-05
GC_6_15 b_6 NI_6 NS_15 0 -3.7422373229155058e-06
GC_6_16 b_6 NI_6 NS_16 0 2.7238948861022121e-06
GC_6_17 b_6 NI_6 NS_17 0 4.5150303792613556e-06
GC_6_18 b_6 NI_6 NS_18 0 1.5307786500822762e-06
GC_6_19 b_6 NI_6 NS_19 0 8.7546485635875665e-06
GC_6_20 b_6 NI_6 NS_20 0 -3.8479440447810489e-05
GC_6_21 b_6 NI_6 NS_21 0 -4.3264344561478150e-05
GC_6_22 b_6 NI_6 NS_22 0 -1.4454256584817443e-06
GC_6_23 b_6 NI_6 NS_23 0 -1.4749708942910464e-05
GC_6_24 b_6 NI_6 NS_24 0 -8.4841759444300327e-06
GC_6_25 b_6 NI_6 NS_25 0 -7.0816020634931421e-05
GC_6_26 b_6 NI_6 NS_26 0 7.5581835459800998e-05
GC_6_27 b_6 NI_6 NS_27 0 4.8531183388139991e-06
GC_6_28 b_6 NI_6 NS_28 0 1.3247715061147525e-05
GC_6_29 b_6 NI_6 NS_29 0 6.5373800829676267e-05
GC_6_30 b_6 NI_6 NS_30 0 1.2307919735115219e-04
GC_6_31 b_6 NI_6 NS_31 0 -1.3648056384514943e-07
GC_6_32 b_6 NI_6 NS_32 0 -3.7823403070185376e-05
GC_6_33 b_6 NI_6 NS_33 0 1.6963540650317057e-05
GC_6_34 b_6 NI_6 NS_34 0 4.3618131817285294e-06
GC_6_35 b_6 NI_6 NS_35 0 2.5306406281669916e-05
GC_6_36 b_6 NI_6 NS_36 0 -3.1223668563984673e-05
GC_6_37 b_6 NI_6 NS_37 0 -8.6240530582695165e-06
GC_6_38 b_6 NI_6 NS_38 0 -2.7321978288785062e-06
GC_6_39 b_6 NI_6 NS_39 0 -8.1952300557998280e-06
GC_6_40 b_6 NI_6 NS_40 0 2.4464289424428995e-05
GC_6_41 b_6 NI_6 NS_41 0 6.0408730816697431e-06
GC_6_42 b_6 NI_6 NS_42 0 8.5944396950360107e-06
GC_6_43 b_6 NI_6 NS_43 0 5.7640097520480125e-05
GC_6_44 b_6 NI_6 NS_44 0 2.4091330709466709e-05
GC_6_45 b_6 NI_6 NS_45 0 3.6448056463085684e-06
GC_6_46 b_6 NI_6 NS_46 0 -1.2427227666394427e-05
GC_6_47 b_6 NI_6 NS_47 0 -7.2855748467425722e-08
GC_6_48 b_6 NI_6 NS_48 0 -1.3777539539239949e-06
GC_6_49 b_6 NI_6 NS_49 0 7.2151384694031405e-06
GC_6_50 b_6 NI_6 NS_50 0 2.9209008531464125e-06
GC_6_51 b_6 NI_6 NS_51 0 4.2719688395613010e-05
GC_6_52 b_6 NI_6 NS_52 0 -1.9006752905723519e-05
GC_6_53 b_6 NI_6 NS_53 0 -2.4853145273174273e-06
GC_6_54 b_6 NI_6 NS_54 0 -7.7712979195929741e-06
GC_6_55 b_6 NI_6 NS_55 0 -2.8170084837633921e-06
GC_6_56 b_6 NI_6 NS_56 0 1.1098380950930774e-06
GC_6_57 b_6 NI_6 NS_57 0 9.8836129831414984e-06
GC_6_58 b_6 NI_6 NS_58 0 2.6878984796884356e-06
GC_6_59 b_6 NI_6 NS_59 0 2.2660344141460226e-05
GC_6_60 b_6 NI_6 NS_60 0 -3.3266185500446366e-05
GC_6_61 b_6 NI_6 NS_61 0 -5.7340514682014511e-06
GC_6_62 b_6 NI_6 NS_62 0 -4.2992031580612423e-06
GC_6_63 b_6 NI_6 NS_63 0 -8.7799528454120592e-07
GC_6_64 b_6 NI_6 NS_64 0 4.2823149494064653e-06
GC_6_65 b_6 NI_6 NS_65 0 1.2543404987341688e-05
GC_6_66 b_6 NI_6 NS_66 0 -1.7550208642716126e-07
GC_6_67 b_6 NI_6 NS_67 0 6.1352852645723629e-07
GC_6_68 b_6 NI_6 NS_68 0 -3.3003904000983482e-05
GC_6_69 b_6 NI_6 NS_69 0 -6.9295725523163948e-06
GC_6_70 b_6 NI_6 NS_70 0 3.5370508800582545e-07
GC_6_71 b_6 NI_6 NS_71 0 3.8626397193917695e-06
GC_6_72 b_6 NI_6 NS_72 0 3.5637552672222811e-06
GC_6_73 b_6 NI_6 NS_73 0 1.4168024987765440e-05
GC_6_74 b_6 NI_6 NS_74 0 -6.6370194185054128e-06
GC_6_75 b_6 NI_6 NS_75 0 -1.5560846421632121e-05
GC_6_76 b_6 NI_6 NS_76 0 -1.9131784917742365e-05
GC_6_77 b_6 NI_6 NS_77 0 -2.9829629257358808e-06
GC_6_78 b_6 NI_6 NS_78 0 5.0701964910700033e-06
GC_6_79 b_6 NI_6 NS_79 0 4.2041749213123217e-06
GC_6_80 b_6 NI_6 NS_80 0 -1.9025757516163620e-06
GC_6_81 b_6 NI_6 NS_81 0 -2.7722125992132913e-11
GC_6_82 b_6 NI_6 NS_82 0 5.4087820899638478e-12
GC_6_83 b_6 NI_6 NS_83 0 4.8942895937900053e-06
GC_6_84 b_6 NI_6 NS_84 0 -1.1671146543794715e-05
GC_6_85 b_6 NI_6 NS_85 0 -5.0227516645649185e-07
GC_6_86 b_6 NI_6 NS_86 0 2.7925975834414354e-06
GC_6_87 b_6 NI_6 NS_87 0 2.3625582144180136e-06
GC_6_88 b_6 NI_6 NS_88 0 -1.5932287151612288e-06
GC_6_89 b_6 NI_6 NS_89 0 2.1702313627834886e-06
GC_6_90 b_6 NI_6 NS_90 0 -9.8796032019875298e-06
GC_6_91 b_6 NI_6 NS_91 0 -1.0601719983688160e-05
GC_6_92 b_6 NI_6 NS_92 0 -3.5478334374594770e-06
GC_6_93 b_6 NI_6 NS_93 0 -2.2615754945366798e-10
GC_6_94 b_6 NI_6 NS_94 0 4.2340218356497706e-10
GC_6_95 b_6 NI_6 NS_95 0 -9.1524871568374543e-06
GC_6_96 b_6 NI_6 NS_96 0 -5.6556579544661693e-06
GC_6_97 b_6 NI_6 NS_97 0 2.0112928704445384e-06
GC_6_98 b_6 NI_6 NS_98 0 -6.6968695379704610e-06
GC_6_99 b_6 NI_6 NS_99 0 -3.3581514623960135e-06
GC_6_100 b_6 NI_6 NS_100 0 -1.8350310502158154e-07
GC_6_101 b_6 NI_6 NS_101 0 -8.5821395414706722e-06
GC_6_102 b_6 NI_6 NS_102 0 5.9057936743777195e-07
GC_6_103 b_6 NI_6 NS_103 0 2.6252870595195957e-06
GC_6_104 b_6 NI_6 NS_104 0 2.8291308595777565e-06
GC_6_105 b_6 NI_6 NS_105 0 1.0192572516621671e-06
GC_6_106 b_6 NI_6 NS_106 0 -3.7248592552942298e-06
GC_6_107 b_6 NI_6 NS_107 0 -5.3998924562925384e-06
GC_6_108 b_6 NI_6 NS_108 0 -4.2209437909207260e-06
GC_6_109 b_6 NI_6 NS_109 0 -5.4772844120695309e-05
GC_6_110 b_6 NI_6 NS_110 0 -6.9629437200645509e-12
GC_6_111 b_6 NI_6 NS_111 0 -2.0817912859138361e-10
GC_6_112 b_6 NI_6 NS_112 0 9.8206144098253359e-09
GC_6_113 b_6 NI_6 NS_113 0 5.4129957677143521e-07
GC_6_114 b_6 NI_6 NS_114 0 4.9187587552106220e-08
GC_6_115 b_6 NI_6 NS_115 0 2.9069068254200984e-06
GC_6_116 b_6 NI_6 NS_116 0 -1.4984891893615365e-06
GC_6_117 b_6 NI_6 NS_117 0 -3.1925349479281577e-06
GC_6_118 b_6 NI_6 NS_118 0 -2.5905350518553044e-06
GC_6_119 b_6 NI_6 NS_119 0 4.5917106068593701e-06
GC_6_120 b_6 NI_6 NS_120 0 -3.9820031445765125e-07
GC_6_121 b_6 NI_6 NS_121 0 -7.4318684383880411e-06
GC_6_122 b_6 NI_6 NS_122 0 -7.4641161902565526e-06
GC_6_123 b_6 NI_6 NS_123 0 -2.5846975908079067e-07
GC_6_124 b_6 NI_6 NS_124 0 -1.3549726422346559e-06
GC_6_125 b_6 NI_6 NS_125 0 -5.8670259208866842e-06
GC_6_126 b_6 NI_6 NS_126 0 2.4876412746608696e-06
GC_6_127 b_6 NI_6 NS_127 0 5.2138883915337892e-06
GC_6_128 b_6 NI_6 NS_128 0 -5.0558572757963265e-06
GC_6_129 b_6 NI_6 NS_129 0 -1.6625735767015013e-05
GC_6_130 b_6 NI_6 NS_130 0 5.0766175329871588e-06
GC_6_131 b_6 NI_6 NS_131 0 -1.1389054443761824e-06
GC_6_132 b_6 NI_6 NS_132 0 7.5150225500193631e-06
GC_6_133 b_6 NI_6 NS_133 0 -6.5962451740772420e-06
GC_6_134 b_6 NI_6 NS_134 0 -4.0226072395498573e-06
GC_6_135 b_6 NI_6 NS_135 0 -3.2518604330029135e-06
GC_6_136 b_6 NI_6 NS_136 0 8.3354888018822377e-06
GC_6_137 b_6 NI_6 NS_137 0 -1.2792490752319117e-06
GC_6_138 b_6 NI_6 NS_138 0 -4.0909169402256802e-06
GC_6_139 b_6 NI_6 NS_139 0 -3.9771512656987145e-06
GC_6_140 b_6 NI_6 NS_140 0 1.1475666952748954e-05
GC_6_141 b_6 NI_6 NS_141 0 -1.4781989710627664e-08
GC_6_142 b_6 NI_6 NS_142 0 7.6669268693975331e-06
GC_6_143 b_6 NI_6 NS_143 0 -3.6189377234133647e-06
GC_6_144 b_6 NI_6 NS_144 0 1.4618089991379339e-06
GC_6_145 b_6 NI_6 NS_145 0 -3.4651571657334917e-07
GC_6_146 b_6 NI_6 NS_146 0 8.4080178150468161e-06
GC_6_147 b_6 NI_6 NS_147 0 -5.5944460371679973e-07
GC_6_148 b_6 NI_6 NS_148 0 2.1381468703751423e-06
GC_6_149 b_6 NI_6 NS_149 0 -2.2883710658551187e-06
GC_6_150 b_6 NI_6 NS_150 0 8.4915537563568657e-06
GC_6_151 b_6 NI_6 NS_151 0 7.3273015304509391e-07
GC_6_152 b_6 NI_6 NS_152 0 9.9252263218135145e-06
GC_6_153 b_6 NI_6 NS_153 0 -7.0096484037387217e-07
GC_6_154 b_6 NI_6 NS_154 0 8.9537435601072310e-06
GC_6_155 b_6 NI_6 NS_155 0 -1.2260745285754294e-06
GC_6_156 b_6 NI_6 NS_156 0 4.0765953371153705e-06
GC_6_157 b_6 NI_6 NS_157 0 1.3021507529876134e-06
GC_6_158 b_6 NI_6 NS_158 0 1.2333188303515230e-05
GC_6_159 b_6 NI_6 NS_159 0 1.8798613922335710e-05
GC_6_160 b_6 NI_6 NS_160 0 1.7017275247839715e-05
GC_6_161 b_6 NI_6 NS_161 0 5.0479537448427585e-06
GC_6_162 b_6 NI_6 NS_162 0 7.8839365838292269e-06
GC_6_163 b_6 NI_6 NS_163 0 1.0389989274283236e-05
GC_6_164 b_6 NI_6 NS_164 0 3.8923638936471031e-06
GC_6_165 b_6 NI_6 NS_165 0 6.8759109014526046e-06
GC_6_166 b_6 NI_6 NS_166 0 1.1069323429494128e-05
GC_6_167 b_6 NI_6 NS_167 0 3.3658578081514531e-05
GC_6_168 b_6 NI_6 NS_168 0 -6.2040446915443295e-06
GC_6_169 b_6 NI_6 NS_169 0 8.2351361031573562e-06
GC_6_170 b_6 NI_6 NS_170 0 3.4806557640994637e-06
GC_6_171 b_6 NI_6 NS_171 0 1.2053460701628581e-05
GC_6_172 b_6 NI_6 NS_172 0 -1.0358836390149264e-05
GC_6_173 b_6 NI_6 NS_173 0 1.0858559160024193e-05
GC_6_174 b_6 NI_6 NS_174 0 6.5736103075053291e-06
GC_6_175 b_6 NI_6 NS_175 0 1.7121023609543903e-05
GC_6_176 b_6 NI_6 NS_176 0 -3.0993299684994132e-05
GC_6_177 b_6 NI_6 NS_177 0 8.1831186676494554e-06
GC_6_178 b_6 NI_6 NS_178 0 -2.9223707986273811e-06
GC_6_179 b_6 NI_6 NS_179 0 -3.1851996427976511e-06
GC_6_180 b_6 NI_6 NS_180 0 -1.6372769431268230e-05
GC_6_181 b_6 NI_6 NS_181 0 1.1876730642203001e-05
GC_6_182 b_6 NI_6 NS_182 0 -1.5556616531573666e-06
GC_6_183 b_6 NI_6 NS_183 0 -1.2637532357685594e-05
GC_6_184 b_6 NI_6 NS_184 0 -2.5277366029824179e-05
GC_6_185 b_6 NI_6 NS_185 0 -1.0768074212464627e-07
GC_6_186 b_6 NI_6 NS_186 0 -6.6428262826827158e-06
GC_6_187 b_6 NI_6 NS_187 0 -9.5779958521991351e-06
GC_6_188 b_6 NI_6 NS_188 0 -2.6885578329866993e-06
GC_6_189 b_6 NI_6 NS_189 0 1.0207143126925955e-10
GC_6_190 b_6 NI_6 NS_190 0 4.5675821892604927e-11
GC_6_191 b_6 NI_6 NS_191 0 1.5500865529281238e-06
GC_6_192 b_6 NI_6 NS_192 0 -4.7010659228057024e-06
GC_6_193 b_6 NI_6 NS_193 0 -1.3389448841447365e-06
GC_6_194 b_6 NI_6 NS_194 0 -1.3668614568019745e-06
GC_6_195 b_6 NI_6 NS_195 0 -4.8399313763360886e-06
GC_6_196 b_6 NI_6 NS_196 0 -1.0276602110663776e-06
GC_6_197 b_6 NI_6 NS_197 0 -1.0646410860870592e-06
GC_6_198 b_6 NI_6 NS_198 0 -2.7378262741847625e-06
GC_6_199 b_6 NI_6 NS_199 0 -9.9890614160465737e-06
GC_6_200 b_6 NI_6 NS_200 0 -4.1192124164004082e-06
GC_6_201 b_6 NI_6 NS_201 0 6.6959739008716804e-09
GC_6_202 b_6 NI_6 NS_202 0 5.4073950215518974e-09
GC_6_203 b_6 NI_6 NS_203 0 1.7777237136199191e-06
GC_6_204 b_6 NI_6 NS_204 0 4.4395341240508439e-07
GC_6_205 b_6 NI_6 NS_205 0 -1.5869734192722623e-06
GC_6_206 b_6 NI_6 NS_206 0 3.2264935079944614e-06
GC_6_207 b_6 NI_6 NS_207 0 -8.2721059307802136e-07
GC_6_208 b_6 NI_6 NS_208 0 6.9325931935675971e-07
GC_6_209 b_6 NI_6 NS_209 0 -7.6673735587582635e-06
GC_6_210 b_6 NI_6 NS_210 0 4.7218365551631365e-07
GC_6_211 b_6 NI_6 NS_211 0 -2.2070926830037886e-06
GC_6_212 b_6 NI_6 NS_212 0 1.9527358638013687e-06
GC_6_213 b_6 NI_6 NS_213 0 -2.0870472355755708e-06
GC_6_214 b_6 NI_6 NS_214 0 1.9632476078778956e-06
GC_6_215 b_6 NI_6 NS_215 0 1.2949331350686769e-06
GC_6_216 b_6 NI_6 NS_216 0 2.8398323240101710e-06
GC_6_217 b_6 NI_6 NS_217 0 -6.4105861506774350e-04
GC_6_218 b_6 NI_6 NS_218 0 -9.7197848733164243e-11
GC_6_219 b_6 NI_6 NS_219 0 3.8858264524741188e-09
GC_6_220 b_6 NI_6 NS_220 0 -6.7399748993742727e-08
GC_6_221 b_6 NI_6 NS_221 0 -1.1325349374590708e-05
GC_6_222 b_6 NI_6 NS_222 0 -9.3599508361932634e-06
GC_6_223 b_6 NI_6 NS_223 0 -2.2402057161078846e-06
GC_6_224 b_6 NI_6 NS_224 0 1.9787863310358243e-07
GC_6_225 b_6 NI_6 NS_225 0 -3.0414370435521898e-05
GC_6_226 b_6 NI_6 NS_226 0 2.7141390509978107e-05
GC_6_227 b_6 NI_6 NS_227 0 -3.3444217399673500e-05
GC_6_228 b_6 NI_6 NS_228 0 8.1131392889947043e-06
GC_6_229 b_6 NI_6 NS_229 0 3.1774137748961086e-05
GC_6_230 b_6 NI_6 NS_230 0 2.7463320156026254e-05
GC_6_231 b_6 NI_6 NS_231 0 -9.1036112123762495e-06
GC_6_232 b_6 NI_6 NS_232 0 1.4796418004090470e-05
GC_6_233 b_6 NI_6 NS_233 0 1.2667859729246203e-05
GC_6_234 b_6 NI_6 NS_234 0 3.7134956782147278e-05
GC_6_235 b_6 NI_6 NS_235 0 -1.1026764730346091e-05
GC_6_236 b_6 NI_6 NS_236 0 6.8453885502915300e-05
GC_6_237 b_6 NI_6 NS_237 0 9.5993858814715253e-05
GC_6_238 b_6 NI_6 NS_238 0 -6.6259870461554226e-05
GC_6_239 b_6 NI_6 NS_239 0 2.7201064731113508e-05
GC_6_240 b_6 NI_6 NS_240 0 3.2003867205384785e-05
GC_6_241 b_6 NI_6 NS_241 0 -7.0531925239586030e-06
GC_6_242 b_6 NI_6 NS_242 0 -7.2616518322595453e-05
GC_6_243 b_6 NI_6 NS_243 0 -9.8456931535958475e-06
GC_6_244 b_6 NI_6 NS_244 0 -3.4285202543218303e-05
GC_6_245 b_6 NI_6 NS_245 0 -7.6897131390768632e-05
GC_6_246 b_6 NI_6 NS_246 0 1.8745808828705365e-05
GC_6_247 b_6 NI_6 NS_247 0 2.4874720629934380e-05
GC_6_248 b_6 NI_6 NS_248 0 5.1393202484541850e-05
GC_6_249 b_6 NI_6 NS_249 0 -2.3342748917890293e-05
GC_6_250 b_6 NI_6 NS_250 0 -3.7551236393181415e-06
GC_6_251 b_6 NI_6 NS_251 0 7.0090143658303733e-05
GC_6_252 b_6 NI_6 NS_252 0 4.4926280941638859e-05
GC_6_253 b_6 NI_6 NS_253 0 2.9399647549506764e-05
GC_6_254 b_6 NI_6 NS_254 0 1.9985842113520886e-05
GC_6_255 b_6 NI_6 NS_255 0 -7.2378854546753111e-06
GC_6_256 b_6 NI_6 NS_256 0 -2.5815194601862029e-05
GC_6_257 b_6 NI_6 NS_257 0 -7.5769884773068691e-06
GC_6_258 b_6 NI_6 NS_258 0 -2.5457578469617094e-05
GC_6_259 b_6 NI_6 NS_259 0 6.9370843825887060e-06
GC_6_260 b_6 NI_6 NS_260 0 4.9224246814201206e-05
GC_6_261 b_6 NI_6 NS_261 0 1.2889452021389758e-05
GC_6_262 b_6 NI_6 NS_262 0 2.7625570774978338e-05
GC_6_263 b_6 NI_6 NS_263 0 5.8786692777324865e-06
GC_6_264 b_6 NI_6 NS_264 0 2.1442877179698809e-06
GC_6_265 b_6 NI_6 NS_265 0 -6.1844722745396538e-07
GC_6_266 b_6 NI_6 NS_266 0 -1.5585956418825055e-05
GC_6_267 b_6 NI_6 NS_267 0 5.6423026127808486e-05
GC_6_268 b_6 NI_6 NS_268 0 3.8203674322081544e-05
GC_6_269 b_6 NI_6 NS_269 0 1.9996580966128683e-05
GC_6_270 b_6 NI_6 NS_270 0 1.5002575526345202e-05
GC_6_271 b_6 NI_6 NS_271 0 8.4325587532217153e-06
GC_6_272 b_6 NI_6 NS_272 0 -1.2893614736196838e-05
GC_6_273 b_6 NI_6 NS_273 0 -5.6500652378529032e-06
GC_6_274 b_6 NI_6 NS_274 0 -1.4195065471457969e-05
GC_6_275 b_6 NI_6 NS_275 0 6.6301826291428496e-05
GC_6_276 b_6 NI_6 NS_276 0 1.2978543121911713e-05
GC_6_277 b_6 NI_6 NS_277 0 2.2841948169633930e-05
GC_6_278 b_6 NI_6 NS_278 0 5.0487029290596485e-06
GC_6_279 b_6 NI_6 NS_279 0 -5.5524465592330971e-06
GC_6_280 b_6 NI_6 NS_280 0 -2.2079790260345179e-05
GC_6_281 b_6 NI_6 NS_281 0 -9.1403127087109752e-06
GC_6_282 b_6 NI_6 NS_282 0 -7.2135316698886164e-06
GC_6_283 b_6 NI_6 NS_283 0 6.0763587252473918e-05
GC_6_284 b_6 NI_6 NS_284 0 -9.5420678370480528e-06
GC_6_285 b_6 NI_6 NS_285 0 2.1478227851639046e-05
GC_6_286 b_6 NI_6 NS_286 0 -7.3421543121298824e-06
GC_6_287 b_6 NI_6 NS_287 0 -2.3108195879337222e-05
GC_6_288 b_6 NI_6 NS_288 0 -1.3186405294402354e-05
GC_6_289 b_6 NI_6 NS_289 0 -8.6384546345367918e-06
GC_6_290 b_6 NI_6 NS_290 0 4.3948700661476587e-06
GC_6_291 b_6 NI_6 NS_291 0 4.5484339018437442e-05
GC_6_292 b_6 NI_6 NS_292 0 -2.5717089267822055e-05
GC_6_293 b_6 NI_6 NS_293 0 6.0380911352361642e-06
GC_6_294 b_6 NI_6 NS_294 0 -1.6494070546845589e-05
GC_6_295 b_6 NI_6 NS_295 0 -1.8737711427559523e-05
GC_6_296 b_6 NI_6 NS_296 0 8.6024235234489824e-06
GC_6_297 b_6 NI_6 NS_297 0 -4.6784477276804164e-11
GC_6_298 b_6 NI_6 NS_298 0 -1.7807466738014455e-10
GC_6_299 b_6 NI_6 NS_299 0 1.7771662742622918e-06
GC_6_300 b_6 NI_6 NS_300 0 8.7585030565030666e-06
GC_6_301 b_6 NI_6 NS_301 0 2.2074348799744727e-06
GC_6_302 b_6 NI_6 NS_302 0 -7.0114804648016692e-06
GC_6_303 b_6 NI_6 NS_303 0 -9.0081319052681285e-06
GC_6_304 b_6 NI_6 NS_304 0 5.7591249128966879e-06
GC_6_305 b_6 NI_6 NS_305 0 4.7915722625420456e-06
GC_6_306 b_6 NI_6 NS_306 0 1.1558577380103885e-05
GC_6_307 b_6 NI_6 NS_307 0 2.4562418340236008e-05
GC_6_308 b_6 NI_6 NS_308 0 -2.1173228122305516e-05
GC_6_309 b_6 NI_6 NS_309 0 -5.7146444857208379e-09
GC_6_310 b_6 NI_6 NS_310 0 -5.6481292434687078e-09
GC_6_311 b_6 NI_6 NS_311 0 3.0658431378985196e-05
GC_6_312 b_6 NI_6 NS_312 0 7.4840761090345332e-06
GC_6_313 b_6 NI_6 NS_313 0 -2.6776559877564490e-06
GC_6_314 b_6 NI_6 NS_314 0 1.1046091148907756e-05
GC_6_315 b_6 NI_6 NS_315 0 8.0413961888927921e-06
GC_6_316 b_6 NI_6 NS_316 0 1.1940897562848157e-06
GC_6_317 b_6 NI_6 NS_317 0 1.9118667233523270e-05
GC_6_318 b_6 NI_6 NS_318 0 -2.1563824578677328e-05
GC_6_319 b_6 NI_6 NS_319 0 -6.5506355132872060e-06
GC_6_320 b_6 NI_6 NS_320 0 -7.4600009908265993e-06
GC_6_321 b_6 NI_6 NS_321 0 -5.3917913583534550e-06
GC_6_322 b_6 NI_6 NS_322 0 1.2485350877305975e-05
GC_6_323 b_6 NI_6 NS_323 0 1.6112330214245082e-05
GC_6_324 b_6 NI_6 NS_324 0 7.3766610488005514e-06
GC_6_325 b_6 NI_6 NS_325 0 7.9288748106353209e-05
GC_6_326 b_6 NI_6 NS_326 0 -1.2174291277099575e-10
GC_6_327 b_6 NI_6 NS_327 0 -2.0288821250974514e-09
GC_6_328 b_6 NI_6 NS_328 0 3.4022340935787456e-08
GC_6_329 b_6 NI_6 NS_329 0 -3.3983706979251914e-07
GC_6_330 b_6 NI_6 NS_330 0 -3.3574283695044813e-07
GC_6_331 b_6 NI_6 NS_331 0 -5.7584242004036873e-07
GC_6_332 b_6 NI_6 NS_332 0 9.6675315570907827e-06
GC_6_333 b_6 NI_6 NS_333 0 1.3105676026046349e-05
GC_6_334 b_6 NI_6 NS_334 0 -1.2342181871068711e-05
GC_6_335 b_6 NI_6 NS_335 0 -1.7112606855796874e-05
GC_6_336 b_6 NI_6 NS_336 0 8.5764476714018057e-06
GC_6_337 b_6 NI_6 NS_337 0 2.8663170608251613e-05
GC_6_338 b_6 NI_6 NS_338 0 -7.4194702283476501e-06
GC_6_339 b_6 NI_6 NS_339 0 -2.8956659508489905e-06
GC_6_340 b_6 NI_6 NS_340 0 -3.4130742210846956e-06
GC_6_341 b_6 NI_6 NS_341 0 -3.2449804147242011e-06
GC_6_342 b_6 NI_6 NS_342 0 -1.5090311596072427e-05
GC_6_343 b_6 NI_6 NS_343 0 -2.4828337472517017e-05
GC_6_344 b_6 NI_6 NS_344 0 3.9221721286812920e-05
GC_6_345 b_6 NI_6 NS_345 0 3.6987644414638259e-05
GC_6_346 b_6 NI_6 NS_346 0 -4.7225340811290426e-05
GC_6_347 b_6 NI_6 NS_347 0 -3.0518339461971297e-05
GC_6_348 b_6 NI_6 NS_348 0 -2.1425302161267035e-05
GC_6_349 b_6 NI_6 NS_349 0 3.2014658244159357e-05
GC_6_350 b_6 NI_6 NS_350 0 2.6387854860634392e-05
GC_6_351 b_6 NI_6 NS_351 0 -1.8545633806795780e-05
GC_6_352 b_6 NI_6 NS_352 0 -2.9076395143778122e-05
GC_6_353 b_6 NI_6 NS_353 0 2.0026492942475261e-05
GC_6_354 b_6 NI_6 NS_354 0 5.9804793797451665e-05
GC_6_355 b_6 NI_6 NS_355 0 -2.0977330629786661e-05
GC_6_356 b_6 NI_6 NS_356 0 -5.5613753236292245e-05
GC_6_357 b_6 NI_6 NS_357 0 -3.1646152877055207e-05
GC_6_358 b_6 NI_6 NS_358 0 -1.2116541199858885e-05
GC_6_359 b_6 NI_6 NS_359 0 1.9561870496163475e-05
GC_6_360 b_6 NI_6 NS_360 0 1.3806626329972756e-05
GC_6_361 b_6 NI_6 NS_361 0 -2.4957198274251179e-05
GC_6_362 b_6 NI_6 NS_362 0 -1.1262318012278381e-05
GC_6_363 b_6 NI_6 NS_363 0 2.0179937023939578e-05
GC_6_364 b_6 NI_6 NS_364 0 1.0341639104802652e-05
GC_6_365 b_6 NI_6 NS_365 0 -1.8434218523731557e-05
GC_6_366 b_6 NI_6 NS_366 0 -2.1152540732363728e-05
GC_6_367 b_6 NI_6 NS_367 0 4.2957737175938267e-06
GC_6_368 b_6 NI_6 NS_368 0 3.1958082300697624e-05
GC_6_369 b_6 NI_6 NS_369 0 -8.4065272336609101e-06
GC_6_370 b_6 NI_6 NS_370 0 -2.6582396538829059e-05
GC_6_371 b_6 NI_6 NS_371 0 -2.0402888452019782e-06
GC_6_372 b_6 NI_6 NS_372 0 1.5416009959469692e-06
GC_6_373 b_6 NI_6 NS_373 0 -1.9679904102930060e-05
GC_6_374 b_6 NI_6 NS_374 0 -1.2198708820999917e-05
GC_6_375 b_6 NI_6 NS_375 0 5.5390028033574826e-06
GC_6_376 b_6 NI_6 NS_376 0 2.1304113305830235e-05
GC_6_377 b_6 NI_6 NS_377 0 -1.6263704313578511e-05
GC_6_378 b_6 NI_6 NS_378 0 -1.4842861964442205e-05
GC_6_379 b_6 NI_6 NS_379 0 9.0210300899564892e-07
GC_6_380 b_6 NI_6 NS_380 0 5.5179726163849487e-06
GC_6_381 b_6 NI_6 NS_381 0 -2.5230906358176399e-05
GC_6_382 b_6 NI_6 NS_382 0 -1.0007044512823751e-05
GC_6_383 b_6 NI_6 NS_383 0 7.5032628472194224e-06
GC_6_384 b_6 NI_6 NS_384 0 2.3878270286146259e-05
GC_6_385 b_6 NI_6 NS_385 0 -2.0944113393119213e-05
GC_6_386 b_6 NI_6 NS_386 0 -5.6385641211324178e-06
GC_6_387 b_6 NI_6 NS_387 0 5.9392830426240017e-06
GC_6_388 b_6 NI_6 NS_388 0 7.9059439636107839e-06
GC_6_389 b_6 NI_6 NS_389 0 -3.0918933999592312e-05
GC_6_390 b_6 NI_6 NS_390 0 -2.7455169659095074e-06
GC_6_391 b_6 NI_6 NS_391 0 1.8051693568372104e-05
GC_6_392 b_6 NI_6 NS_392 0 2.6172446386126890e-05
GC_6_393 b_6 NI_6 NS_393 0 -2.2120772812827755e-05
GC_6_394 b_6 NI_6 NS_394 0 6.9971042661228870e-06
GC_6_395 b_6 NI_6 NS_395 0 1.5076744121767528e-05
GC_6_396 b_6 NI_6 NS_396 0 4.4857565844525819e-06
GC_6_397 b_6 NI_6 NS_397 0 -3.5006192715710492e-05
GC_6_398 b_6 NI_6 NS_398 0 1.3594831664631521e-05
GC_6_399 b_6 NI_6 NS_399 0 3.7185055201395230e-05
GC_6_400 b_6 NI_6 NS_400 0 1.3344808458994698e-05
GC_6_401 b_6 NI_6 NS_401 0 -7.9971577182544669e-06
GC_6_402 b_6 NI_6 NS_402 0 1.9077538438475928e-05
GC_6_403 b_6 NI_6 NS_403 0 1.2877244190563973e-05
GC_6_404 b_6 NI_6 NS_404 0 -1.0947056129820303e-05
GC_6_405 b_6 NI_6 NS_405 0 1.1098889656200731e-10
GC_6_406 b_6 NI_6 NS_406 0 4.4127826136394625e-11
GC_6_407 b_6 NI_6 NS_407 0 -1.3992975398868235e-05
GC_6_408 b_6 NI_6 NS_408 0 2.6116738196756830e-05
GC_6_409 b_6 NI_6 NS_409 0 -2.1466198241331191e-06
GC_6_410 b_6 NI_6 NS_410 0 1.0636847819256651e-05
GC_6_411 b_6 NI_6 NS_411 0 6.1623438723870680e-06
GC_6_412 b_6 NI_6 NS_412 0 -8.3666724758380773e-06
GC_6_413 b_6 NI_6 NS_413 0 -8.3609167002666577e-06
GC_6_414 b_6 NI_6 NS_414 0 2.5491814167152571e-05
GC_6_415 b_6 NI_6 NS_415 0 2.5015772726253701e-05
GC_6_416 b_6 NI_6 NS_416 0 -9.9981301841886497e-06
GC_6_417 b_6 NI_6 NS_417 0 4.8733519911353127e-09
GC_6_418 b_6 NI_6 NS_418 0 -1.1063138925369404e-09
GC_6_419 b_6 NI_6 NS_419 0 2.6321680396746009e-05
GC_6_420 b_6 NI_6 NS_420 0 -1.2477251478641133e-05
GC_6_421 b_6 NI_6 NS_421 0 -8.3190506966046506e-06
GC_6_422 b_6 NI_6 NS_422 0 1.8150061776724023e-05
GC_6_423 b_6 NI_6 NS_423 0 -1.0398845374974583e-05
GC_6_424 b_6 NI_6 NS_424 0 -2.8340374495061405e-07
GC_6_425 b_6 NI_6 NS_425 0 1.9410927993698879e-05
GC_6_426 b_6 NI_6 NS_426 0 -1.4077514439135026e-05
GC_6_427 b_6 NI_6 NS_427 0 7.1590822029446791e-06
GC_6_428 b_6 NI_6 NS_428 0 1.1754924684312183e-05
GC_6_429 b_6 NI_6 NS_429 0 -1.8100738648006720e-07
GC_6_430 b_6 NI_6 NS_430 0 -1.4547290086435440e-05
GC_6_431 b_6 NI_6 NS_431 0 1.3082934427983040e-05
GC_6_432 b_6 NI_6 NS_432 0 2.7942030069395410e-05
GC_6_433 b_6 NI_6 NS_433 0 -1.0963073147016847e-02
GC_6_434 b_6 NI_6 NS_434 0 8.3276069722895560e-09
GC_6_435 b_6 NI_6 NS_435 0 9.8608101381736882e-07
GC_6_436 b_6 NI_6 NS_436 0 3.6177580657623515e-05
GC_6_437 b_6 NI_6 NS_437 0 4.3739141969593720e-03
GC_6_438 b_6 NI_6 NS_438 0 -3.4750185261802238e-03
GC_6_439 b_6 NI_6 NS_439 0 -3.7382622061470738e-03
GC_6_440 b_6 NI_6 NS_440 0 6.2463727604606884e-03
GC_6_441 b_6 NI_6 NS_441 0 -8.7586386078073904e-03
GC_6_442 b_6 NI_6 NS_442 0 -5.9567971569784864e-03
GC_6_443 b_6 NI_6 NS_443 0 9.2115215452220987e-03
GC_6_444 b_6 NI_6 NS_444 0 -5.9461495188750596e-03
GC_6_445 b_6 NI_6 NS_445 0 7.1478634000118110e-03
GC_6_446 b_6 NI_6 NS_446 0 1.1907369213458625e-02
GC_6_447 b_6 NI_6 NS_447 0 -4.2314323917051260e-03
GC_6_448 b_6 NI_6 NS_448 0 -1.1324268691774123e-03
GC_6_449 b_6 NI_6 NS_449 0 -8.8598487071688582e-03
GC_6_450 b_6 NI_6 NS_450 0 -4.7418026353755960e-04
GC_6_451 b_6 NI_6 NS_451 0 1.4618444174231637e-02
GC_6_452 b_6 NI_6 NS_452 0 -1.0343815087950731e-02
GC_6_453 b_6 NI_6 NS_453 0 1.6441826489045835e-02
GC_6_454 b_6 NI_6 NS_454 0 4.0225060997904610e-03
GC_6_455 b_6 NI_6 NS_455 0 -1.1482358850963490e-02
GC_6_456 b_6 NI_6 NS_456 0 -2.4511033559305225e-04
GC_6_457 b_6 NI_6 NS_457 0 -1.6636877553690095e-02
GC_6_458 b_6 NI_6 NS_458 0 -4.4573846014270530e-02
GC_6_459 b_6 NI_6 NS_459 0 1.0652634812358328e-02
GC_6_460 b_6 NI_6 NS_460 0 1.1245756323394127e-03
GC_6_461 b_6 NI_6 NS_461 0 -4.8294088772321782e-02
GC_6_462 b_6 NI_6 NS_462 0 1.1061721686025391e-02
GC_6_463 b_6 NI_6 NS_463 0 -1.0433755509328260e-02
GC_6_464 b_6 NI_6 NS_464 0 4.8882535113729526e-04
GC_6_465 b_6 NI_6 NS_465 0 9.7769909733484133e-03
GC_6_466 b_6 NI_6 NS_466 0 -5.7680085209487560e-04
GC_6_467 b_6 NI_6 NS_467 0 4.6095816845729137e-03
GC_6_468 b_6 NI_6 NS_468 0 2.4174009226847384e-02
GC_6_469 b_6 NI_6 NS_469 0 -1.0735352775947357e-02
GC_6_470 b_6 NI_6 NS_470 0 1.9692039622511695e-03
GC_6_471 b_6 NI_6 NS_471 0 -8.4727284429668773e-03
GC_6_472 b_6 NI_6 NS_472 0 -1.3537883051804839e-02
GC_6_473 b_6 NI_6 NS_473 0 1.0150133997969334e-02
GC_6_474 b_6 NI_6 NS_474 0 9.8140819990987687e-04
GC_6_475 b_6 NI_6 NS_475 0 -1.9163126575998338e-02
GC_6_476 b_6 NI_6 NS_476 0 2.8679169992180634e-02
GC_6_477 b_6 NI_6 NS_477 0 -9.6128537817313578e-03
GC_6_478 b_6 NI_6 NS_478 0 -9.6554886553448782e-04
GC_6_479 b_6 NI_6 NS_479 0 1.8914227750156008e-03
GC_6_480 b_6 NI_6 NS_480 0 -1.3780560531005629e-03
GC_6_481 b_6 NI_6 NS_481 0 9.4683001348545206e-03
GC_6_482 b_6 NI_6 NS_482 0 -2.4741908635168776e-04
GC_6_483 b_6 NI_6 NS_483 0 -1.4945599432234766e-04
GC_6_484 b_6 NI_6 NS_484 0 3.0270093038688682e-02
GC_6_485 b_6 NI_6 NS_485 0 -8.5288668240693418e-03
GC_6_486 b_6 NI_6 NS_486 0 1.5478406748744460e-04
GC_6_487 b_6 NI_6 NS_487 0 2.1681617412530230e-04
GC_6_488 b_6 NI_6 NS_488 0 -5.4812575122660133e-03
GC_6_489 b_6 NI_6 NS_489 0 1.0036165885359011e-02
GC_6_490 b_6 NI_6 NS_490 0 -3.3857706452001602e-04
GC_6_491 b_6 NI_6 NS_491 0 8.9341636430440782e-03
GC_6_492 b_6 NI_6 NS_492 0 2.6365820291616292e-02
GC_6_493 b_6 NI_6 NS_493 0 -8.3555392460473894e-03
GC_6_494 b_6 NI_6 NS_494 0 1.3766456076561245e-03
GC_6_495 b_6 NI_6 NS_495 0 -2.5869084462321105e-03
GC_6_496 b_6 NI_6 NS_496 0 -7.3539563271986510e-03
GC_6_497 b_6 NI_6 NS_497 0 1.0553563516664911e-02
GC_6_498 b_6 NI_6 NS_498 0 -8.2348946291138680e-04
GC_6_499 b_6 NI_6 NS_499 0 1.4439011337467701e-02
GC_6_500 b_6 NI_6 NS_500 0 1.9950606833564841e-02
GC_6_501 b_6 NI_6 NS_501 0 -8.2760873029916523e-03
GC_6_502 b_6 NI_6 NS_502 0 2.9305066323063169e-03
GC_6_503 b_6 NI_6 NS_503 0 -5.5941949006485378e-03
GC_6_504 b_6 NI_6 NS_504 0 -6.9177103658684680e-03
GC_6_505 b_6 NI_6 NS_505 0 1.1244063171655163e-02
GC_6_506 b_6 NI_6 NS_506 0 -1.3754145456894129e-03
GC_6_507 b_6 NI_6 NS_507 0 1.5700530230488351e-02
GC_6_508 b_6 NI_6 NS_508 0 1.2945594351200738e-02
GC_6_509 b_6 NI_6 NS_509 0 -7.1893616670266622e-03
GC_6_510 b_6 NI_6 NS_510 0 5.1106079498219057e-03
GC_6_511 b_6 NI_6 NS_511 0 -6.8765833538458115e-03
GC_6_512 b_6 NI_6 NS_512 0 -4.8360425887050765e-03
GC_6_513 b_6 NI_6 NS_513 0 4.7734485803383725e-09
GC_6_514 b_6 NI_6 NS_514 0 4.4199393938065769e-08
GC_6_515 b_6 NI_6 NS_515 0 1.2004105139439270e-02
GC_6_516 b_6 NI_6 NS_516 0 -2.5766627533470852e-03
GC_6_517 b_6 NI_6 NS_517 0 -5.2510753379389711e-03
GC_6_518 b_6 NI_6 NS_518 0 4.7015459439890507e-03
GC_6_519 b_6 NI_6 NS_519 0 -6.1588970358766003e-03
GC_6_520 b_6 NI_6 NS_520 0 -4.3232024915841874e-03
GC_6_521 b_6 NI_6 NS_521 0 1.1774219578108109e-02
GC_6_522 b_6 NI_6 NS_522 0 -3.7297221701913861e-03
GC_6_523 b_6 NI_6 NS_523 0 1.2978428111063235e-02
GC_6_524 b_6 NI_6 NS_524 0 9.4653978068943434e-03
GC_6_525 b_6 NI_6 NS_525 0 3.9180870903957171e-06
GC_6_526 b_6 NI_6 NS_526 0 -9.4184451040016613e-07
GC_6_527 b_6 NI_6 NS_527 0 1.6087880742317859e-02
GC_6_528 b_6 NI_6 NS_528 0 1.6769945833813547e-02
GC_6_529 b_6 NI_6 NS_529 0 1.2047068377842014e-02
GC_6_530 b_6 NI_6 NS_530 0 -2.4806928004426528e-03
GC_6_531 b_6 NI_6 NS_531 0 -8.3607713536286744e-03
GC_6_532 b_6 NI_6 NS_532 0 7.9691329515188186e-05
GC_6_533 b_6 NI_6 NS_533 0 1.1309400927670469e-02
GC_6_534 b_6 NI_6 NS_534 0 7.3306470967411516e-03
GC_6_535 b_6 NI_6 NS_535 0 -4.6732526078708432e-03
GC_6_536 b_6 NI_6 NS_536 0 7.3569228915685413e-03
GC_6_537 b_6 NI_6 NS_537 0 -8.0809725622685586e-03
GC_6_538 b_6 NI_6 NS_538 0 -3.7224018493389032e-03
GC_6_539 b_6 NI_6 NS_539 0 1.5958293637794708e-02
GC_6_540 b_6 NI_6 NS_540 0 -7.7554803149061310e-03
GC_6_541 b_6 NI_6 NS_541 0 -1.3590038758595054e-02
GC_6_542 b_6 NI_6 NS_542 0 5.7574113574498685e-09
GC_6_543 b_6 NI_6 NS_543 0 -1.0755251955003728e-06
GC_6_544 b_6 NI_6 NS_544 0 -2.3265200914775897e-05
GC_6_545 b_6 NI_6 NS_545 0 3.4981851747790032e-04
GC_6_546 b_6 NI_6 NS_546 0 -1.9740598410816467e-04
GC_6_547 b_6 NI_6 NS_547 0 -1.5437483444288376e-03
GC_6_548 b_6 NI_6 NS_548 0 -2.3356983122441903e-03
GC_6_549 b_6 NI_6 NS_549 0 -5.1340364113436742e-05
GC_6_550 b_6 NI_6 NS_550 0 4.3605120496331114e-03
GC_6_551 b_6 NI_6 NS_551 0 1.6175824927349754e-03
GC_6_552 b_6 NI_6 NS_552 0 -5.9520405602870577e-03
GC_6_553 b_6 NI_6 NS_553 0 -4.9853593163292978e-03
GC_6_554 b_6 NI_6 NS_554 0 6.4563571009631851e-03
GC_6_555 b_6 NI_6 NS_555 0 1.1341380715635613e-03
GC_6_556 b_6 NI_6 NS_556 0 -5.0675425946496893e-04
GC_6_557 b_6 NI_6 NS_557 0 2.7871014128825308e-03
GC_6_558 b_6 NI_6 NS_558 0 2.3388044429881205e-03
GC_6_559 b_6 NI_6 NS_559 0 -4.3321682726311884e-03
GC_6_560 b_6 NI_6 NS_560 0 -1.3583565618000427e-02
GC_6_561 b_6 NI_6 NS_561 0 1.5695038276341802e-03
GC_6_562 b_6 NI_6 NS_562 0 1.7683041197579623e-02
GC_6_563 b_6 NI_6 NS_563 0 9.8323126131528195e-03
GC_6_564 b_6 NI_6 NS_564 0 -2.3109432708630214e-03
GC_6_565 b_6 NI_6 NS_565 0 -1.3157073609238679e-02
GC_6_566 b_6 NI_6 NS_566 0 2.2142408000817393e-03
GC_6_567 b_6 NI_6 NS_567 0 9.1925784034046741e-03
GC_6_568 b_6 NI_6 NS_568 0 1.9425112077200561e-03
GC_6_569 b_6 NI_6 NS_569 0 -1.8069422469017639e-02
GC_6_570 b_6 NI_6 NS_570 0 -6.4922283942859104e-03
GC_6_571 b_6 NI_6 NS_571 0 1.5725028675783206e-02
GC_6_572 b_6 NI_6 NS_572 0 6.4951447484252823e-03
GC_6_573 b_6 NI_6 NS_573 0 8.1032003105175002e-03
GC_6_574 b_6 NI_6 NS_574 0 -4.2110876475473565e-03
GC_6_575 b_6 NI_6 NS_575 0 -7.5660795372930563e-03
GC_6_576 b_6 NI_6 NS_576 0 2.0432100992717203e-03
GC_6_577 b_6 NI_6 NS_577 0 6.6854379760948428e-03
GC_6_578 b_6 NI_6 NS_578 0 -2.7541177502803087e-03
GC_6_579 b_6 NI_6 NS_579 0 -6.6055144911247102e-03
GC_6_580 b_6 NI_6 NS_580 0 2.9142121005511037e-03
GC_6_581 b_6 NI_6 NS_581 0 7.6544557708656535e-03
GC_6_582 b_6 NI_6 NS_582 0 4.7732052876357447e-04
GC_6_583 b_6 NI_6 NS_583 0 -9.4088268642746591e-03
GC_6_584 b_6 NI_6 NS_584 0 -5.1695959250246722e-03
GC_6_585 b_6 NI_6 NS_585 0 6.8169842482273622e-03
GC_6_586 b_6 NI_6 NS_586 0 4.1131794029751669e-03
GC_6_587 b_6 NI_6 NS_587 0 -3.9574846280544991e-04
GC_6_588 b_6 NI_6 NS_588 0 -9.3604180763582647e-04
GC_6_589 b_6 NI_6 NS_589 0 5.6653317207762156e-03
GC_6_590 b_6 NI_6 NS_590 0 -1.3801820683056131e-03
GC_6_591 b_6 NI_6 NS_591 0 -9.2023184182151892e-03
GC_6_592 b_6 NI_6 NS_592 0 -1.2456050726622463e-03
GC_6_593 b_6 NI_6 NS_593 0 5.9915313907572361e-03
GC_6_594 b_6 NI_6 NS_594 0 7.3808348578695889e-04
GC_6_595 b_6 NI_6 NS_595 0 -2.6544549900193470e-03
GC_6_596 b_6 NI_6 NS_596 0 2.4842222125170282e-04
GC_6_597 b_6 NI_6 NS_597 0 6.6958828091666115e-03
GC_6_598 b_6 NI_6 NS_598 0 -2.2582329946150025e-03
GC_6_599 b_6 NI_6 NS_599 0 -9.3158089924144406e-03
GC_6_600 b_6 NI_6 NS_600 0 1.5268648283372664e-03
GC_6_601 b_6 NI_6 NS_601 0 5.7300536260806939e-03
GC_6_602 b_6 NI_6 NS_602 0 -1.5007448373695143e-03
GC_6_603 b_6 NI_6 NS_603 0 -3.3211781925184011e-03
GC_6_604 b_6 NI_6 NS_604 0 2.4082389398277226e-03
GC_6_605 b_6 NI_6 NS_605 0 7.2643742621708038e-03
GC_6_606 b_6 NI_6 NS_606 0 -4.0966037542831601e-03
GC_6_607 b_6 NI_6 NS_607 0 -8.5936681109158360e-03
GC_6_608 b_6 NI_6 NS_608 0 4.2025452154413855e-03
GC_6_609 b_6 NI_6 NS_609 0 4.8158705784497602e-03
GC_6_610 b_6 NI_6 NS_610 0 -3.8696540515473659e-03
GC_6_611 b_6 NI_6 NS_611 0 -2.4037860168783709e-03
GC_6_612 b_6 NI_6 NS_612 0 4.7598874104289694e-03
GC_6_613 b_6 NI_6 NS_613 0 7.0540631349610477e-03
GC_6_614 b_6 NI_6 NS_614 0 -7.3479437791381472e-03
GC_6_615 b_6 NI_6 NS_615 0 -7.1271032067402847e-03
GC_6_616 b_6 NI_6 NS_616 0 6.8936503102673928e-03
GC_6_617 b_6 NI_6 NS_617 0 1.6683514128539600e-03
GC_6_618 b_6 NI_6 NS_618 0 -5.2972255960429416e-03
GC_6_619 b_6 NI_6 NS_619 0 5.9423078355028353e-04
GC_6_620 b_6 NI_6 NS_620 0 5.4734770636632752e-03
GC_6_621 b_6 NI_6 NS_621 0 -4.1996224591138842e-09
GC_6_622 b_6 NI_6 NS_622 0 -1.3215473074977930e-08
GC_6_623 b_6 NI_6 NS_623 0 2.7118324802205287e-03
GC_6_624 b_6 NI_6 NS_624 0 -8.5806166158299748e-03
GC_6_625 b_6 NI_6 NS_625 0 8.7189105151600345e-04
GC_6_626 b_6 NI_6 NS_626 0 -3.4318678539232116e-03
GC_6_627 b_6 NI_6 NS_627 0 6.2897431415985582e-04
GC_6_628 b_6 NI_6 NS_628 0 4.0346894477519815e-03
GC_6_629 b_6 NI_6 NS_629 0 2.1766535629689668e-03
GC_6_630 b_6 NI_6 NS_630 0 -8.1586516493606497e-03
GC_6_631 b_6 NI_6 NS_631 0 -3.4870480262387043e-03
GC_6_632 b_6 NI_6 NS_632 0 7.0184773261584912e-03
GC_6_633 b_6 NI_6 NS_633 0 -9.0338470132873869e-08
GC_6_634 b_6 NI_6 NS_634 0 -3.0340980818071843e-07
GC_6_635 b_6 NI_6 NS_635 0 -8.0011233891473365e-03
GC_6_636 b_6 NI_6 NS_636 0 5.3809331600616185e-03
GC_6_637 b_6 NI_6 NS_637 0 4.1753794557670629e-03
GC_6_638 b_6 NI_6 NS_638 0 -6.8471564425540378e-03
GC_6_639 b_6 NI_6 NS_639 0 5.3267679624766171e-03
GC_6_640 b_6 NI_6 NS_640 0 7.4221568060223826e-04
GC_6_641 b_6 NI_6 NS_641 0 -2.3672765884588920e-03
GC_6_642 b_6 NI_6 NS_642 0 6.8575175439451489e-03
GC_6_643 b_6 NI_6 NS_643 0 -1.4866281827221163e-03
GC_6_644 b_6 NI_6 NS_644 0 -4.2154555137041061e-03
GC_6_645 b_6 NI_6 NS_645 0 2.3568558413644305e-03
GC_6_646 b_6 NI_6 NS_646 0 5.0372669558085732e-03
GC_6_647 b_6 NI_6 NS_647 0 -1.9997035533974648e-03
GC_6_648 b_6 NI_6 NS_648 0 -8.9736637719760037e-03
GC_6_649 b_6 NI_6 NS_649 0 -3.3197615077371393e-03
GC_6_650 b_6 NI_6 NS_650 0 1.8243968467886715e-09
GC_6_651 b_6 NI_6 NS_651 0 5.5833686493646005e-08
GC_6_652 b_6 NI_6 NS_652 0 1.8994900695613252e-06
GC_6_653 b_6 NI_6 NS_653 0 -9.0391575333653381e-05
GC_6_654 b_6 NI_6 NS_654 0 -5.8816093922433504e-05
GC_6_655 b_6 NI_6 NS_655 0 -1.2620478087099348e-03
GC_6_656 b_6 NI_6 NS_656 0 -3.0052236560350185e-04
GC_6_657 b_6 NI_6 NS_657 0 -1.6884314959624673e-03
GC_6_658 b_6 NI_6 NS_658 0 2.6375243457915395e-03
GC_6_659 b_6 NI_6 NS_659 0 4.9218123318524483e-04
GC_6_660 b_6 NI_6 NS_660 0 5.4232987542358561e-03
GC_6_661 b_6 NI_6 NS_661 0 7.0977003071706927e-03
GC_6_662 b_6 NI_6 NS_662 0 6.5580733311810439e-04
GC_6_663 b_6 NI_6 NS_663 0 6.4693661373059930e-04
GC_6_664 b_6 NI_6 NS_664 0 -6.5981382850546311e-04
GC_6_665 b_6 NI_6 NS_665 0 1.0491643622529390e-03
GC_6_666 b_6 NI_6 NS_666 0 1.5730848825159097e-03
GC_6_667 b_6 NI_6 NS_667 0 1.2639596499611553e-02
GC_6_668 b_6 NI_6 NS_668 0 1.3143541779153981e-02
GC_6_669 b_6 NI_6 NS_669 0 8.7648802086294567e-03
GC_6_670 b_6 NI_6 NS_670 0 -2.0356149451787115e-02
GC_6_671 b_6 NI_6 NS_671 0 8.3908950576274833e-03
GC_6_672 b_6 NI_6 NS_672 0 -2.8818704505459126e-03
GC_6_673 b_6 NI_6 NS_673 0 -1.2619354463849200e-02
GC_6_674 b_6 NI_6 NS_674 0 -3.8807130047445175e-02
GC_6_675 b_6 NI_6 NS_675 0 -7.2444872565977517e-03
GC_6_676 b_6 NI_6 NS_676 0 -2.1485695287403739e-03
GC_6_677 b_6 NI_6 NS_677 0 -5.2275002091240481e-02
GC_6_678 b_6 NI_6 NS_678 0 -1.8767942545637238e-03
GC_6_679 b_6 NI_6 NS_679 0 1.4892258823857646e-02
GC_6_680 b_6 NI_6 NS_680 0 8.6975609016729238e-03
GC_6_681 b_6 NI_6 NS_681 0 -5.9275334219090819e-03
GC_6_682 b_6 NI_6 NS_682 0 4.9905430455346005e-03
GC_6_683 b_6 NI_6 NS_683 0 8.3533688017791603e-03
GC_6_684 b_6 NI_6 NS_684 0 1.1690136307630480e-02
GC_6_685 b_6 NI_6 NS_685 0 4.5590086452298641e-03
GC_6_686 b_6 NI_6 NS_686 0 -2.9247924675726510e-03
GC_6_687 b_6 NI_6 NS_687 0 -7.8932497667644451e-03
GC_6_688 b_6 NI_6 NS_688 0 -8.1501573080331458e-03
GC_6_689 b_6 NI_6 NS_689 0 -5.6782675818707129e-03
GC_6_690 b_6 NI_6 NS_690 0 -6.1945400958757571e-04
GC_6_691 b_6 NI_6 NS_691 0 -1.8070913512836042e-02
GC_6_692 b_6 NI_6 NS_692 0 1.3562267899791666e-02
GC_6_693 b_6 NI_6 NS_693 0 4.7006660093112254e-03
GC_6_694 b_6 NI_6 NS_694 0 4.3832612388289560e-03
GC_6_695 b_6 NI_6 NS_695 0 6.4907931484364063e-04
GC_6_696 b_6 NI_6 NS_696 0 -1.1064190397599845e-04
GC_6_697 b_6 NI_6 NS_697 0 -3.7967898148101825e-03
GC_6_698 b_6 NI_6 NS_698 0 8.8034002846069839e-04
GC_6_699 b_6 NI_6 NS_699 0 -1.1248852084006782e-03
GC_6_700 b_6 NI_6 NS_700 0 1.6693626560781577e-02
GC_6_701 b_6 NI_6 NS_701 0 4.4443837140775008e-03
GC_6_702 b_6 NI_6 NS_702 0 7.1164090448535568e-04
GC_6_703 b_6 NI_6 NS_703 0 -5.2105051454657723e-04
GC_6_704 b_6 NI_6 NS_704 0 -2.2476775716620263e-03
GC_6_705 b_6 NI_6 NS_705 0 -4.9869184167121708e-03
GC_6_706 b_6 NI_6 NS_706 0 2.1058932026494859e-03
GC_6_707 b_6 NI_6 NS_707 0 7.3345843717240568e-03
GC_6_708 b_6 NI_6 NS_708 0 1.4346772732864417e-02
GC_6_709 b_6 NI_6 NS_709 0 4.1867517342199746e-03
GC_6_710 b_6 NI_6 NS_710 0 -1.6800221464430519e-03
GC_6_711 b_6 NI_6 NS_711 0 -3.3979308305906756e-03
GC_6_712 b_6 NI_6 NS_712 0 -2.1020221578788379e-03
GC_6_713 b_6 NI_6 NS_713 0 -5.4224795890380649e-03
GC_6_714 b_6 NI_6 NS_714 0 4.3763674871928849e-03
GC_6_715 b_6 NI_6 NS_715 0 1.3191405138688292e-02
GC_6_716 b_6 NI_6 NS_716 0 8.4408875034005966e-03
GC_6_717 b_6 NI_6 NS_717 0 2.8354678435269487e-03
GC_6_718 b_6 NI_6 NS_718 0 -4.1274253349564928e-03
GC_6_719 b_6 NI_6 NS_719 0 -5.3215613230191989e-03
GC_6_720 b_6 NI_6 NS_720 0 1.1333329869811901e-03
GC_6_721 b_6 NI_6 NS_721 0 -4.4370944731840483e-03
GC_6_722 b_6 NI_6 NS_722 0 8.3056983000051668e-03
GC_6_723 b_6 NI_6 NS_723 0 1.4614309671753456e-02
GC_6_724 b_6 NI_6 NS_724 0 -4.5696282958441082e-04
GC_6_725 b_6 NI_6 NS_725 0 -1.1788303179580354e-03
GC_6_726 b_6 NI_6 NS_726 0 -4.5487487054969933e-03
GC_6_727 b_6 NI_6 NS_727 0 -2.2870873693035488e-03
GC_6_728 b_6 NI_6 NS_728 0 4.3793455117554763e-03
GC_6_729 b_6 NI_6 NS_729 0 1.8266346737059817e-10
GC_6_730 b_6 NI_6 NS_730 0 -1.5798165184135557e-09
GC_6_731 b_6 NI_6 NS_731 0 1.4387706854717410e-03
GC_6_732 b_6 NI_6 NS_732 0 8.2177758807261293e-03
GC_6_733 b_6 NI_6 NS_733 0 -8.7491003055263812e-04
GC_6_734 b_6 NI_6 NS_734 0 -2.2094167279667330e-03
GC_6_735 b_6 NI_6 NS_735 0 -1.4716785383786283e-03
GC_6_736 b_6 NI_6 NS_736 0 2.7485704243204539e-03
GC_6_737 b_6 NI_6 NS_737 0 1.7223951665452245e-03
GC_6_738 b_6 NI_6 NS_738 0 7.6102907946191418e-03
GC_6_739 b_6 NI_6 NS_739 0 7.5930439282542624e-03
GC_6_740 b_6 NI_6 NS_740 0 -3.8216212223072346e-03
GC_6_741 b_6 NI_6 NS_741 0 -4.7008113716645724e-08
GC_6_742 b_6 NI_6 NS_742 0 -2.0170175914234259e-08
GC_6_743 b_6 NI_6 NS_743 0 1.1386078511073686e-02
GC_6_744 b_6 NI_6 NS_744 0 4.4716365186098176e-03
GC_6_745 b_6 NI_6 NS_745 0 -8.6429611106540012e-04
GC_6_746 b_6 NI_6 NS_746 0 6.4881769365568095e-03
GC_6_747 b_6 NI_6 NS_747 0 3.6256397905606191e-03
GC_6_748 b_6 NI_6 NS_748 0 4.0760139183517244e-04
GC_6_749 b_6 NI_6 NS_749 0 6.0652196136472018e-03
GC_6_750 b_6 NI_6 NS_750 0 -4.6566352533464516e-03
GC_6_751 b_6 NI_6 NS_751 0 -3.3846294272665486e-03
GC_6_752 b_6 NI_6 NS_752 0 -1.3607984535455012e-03
GC_6_753 b_6 NI_6 NS_753 0 1.0687140882699213e-04
GC_6_754 b_6 NI_6 NS_754 0 4.4902870768153092e-03
GC_6_755 b_6 NI_6 NS_755 0 7.2783999813534547e-03
GC_6_756 b_6 NI_6 NS_756 0 5.5303118665771152e-03
GC_6_757 b_6 NI_6 NS_757 0 1.4425741233363850e-03
GC_6_758 b_6 NI_6 NS_758 0 -3.5904351747149312e-09
GC_6_759 b_6 NI_6 NS_759 0 -4.7342043128150009e-08
GC_6_760 b_6 NI_6 NS_760 0 -3.5032371832118765e-06
GC_6_761 b_6 NI_6 NS_761 0 -3.6675402607324649e-04
GC_6_762 b_6 NI_6 NS_762 0 1.3531649500525661e-04
GC_6_763 b_6 NI_6 NS_763 0 1.1270906314471171e-03
GC_6_764 b_6 NI_6 NS_764 0 1.9466317752188215e-03
GC_6_765 b_6 NI_6 NS_765 0 -5.2133213260549001e-05
GC_6_766 b_6 NI_6 NS_766 0 -3.4959654435807565e-03
GC_6_767 b_6 NI_6 NS_767 0 -1.5728294785790976e-03
GC_6_768 b_6 NI_6 NS_768 0 5.0835060984192465e-03
GC_6_769 b_6 NI_6 NS_769 0 4.2660496763269884e-03
GC_6_770 b_6 NI_6 NS_770 0 -4.9897929070205401e-03
GC_6_771 b_6 NI_6 NS_771 0 -1.0071498745518562e-03
GC_6_772 b_6 NI_6 NS_772 0 5.5941858275031339e-04
GC_6_773 b_6 NI_6 NS_773 0 -2.0791293775649241e-03
GC_6_774 b_6 NI_6 NS_774 0 -1.8719560941386167e-03
GC_6_775 b_6 NI_6 NS_775 0 3.6235024008862251e-03
GC_6_776 b_6 NI_6 NS_776 0 1.1644121681272452e-02
GC_6_777 b_6 NI_6 NS_777 0 -8.7672702084263675e-04
GC_6_778 b_6 NI_6 NS_778 0 -1.4855229418282772e-02
GC_6_779 b_6 NI_6 NS_779 0 -8.1250075384111456e-03
GC_6_780 b_6 NI_6 NS_780 0 1.9028461816925661e-03
GC_6_781 b_6 NI_6 NS_781 0 1.1255574803279393e-02
GC_6_782 b_6 NI_6 NS_782 0 -1.8013331256157784e-03
GC_6_783 b_6 NI_6 NS_783 0 -7.5649379463101690e-03
GC_6_784 b_6 NI_6 NS_784 0 -1.6931181032836292e-03
GC_6_785 b_6 NI_6 NS_785 0 1.5263484753164563e-02
GC_6_786 b_6 NI_6 NS_786 0 5.3089269962557119e-03
GC_6_787 b_6 NI_6 NS_787 0 -1.3074208628142386e-02
GC_6_788 b_6 NI_6 NS_788 0 -5.4740974161817078e-03
GC_6_789 b_6 NI_6 NS_789 0 -6.6401727829745278e-03
GC_6_790 b_6 NI_6 NS_790 0 3.4469264645533102e-03
GC_6_791 b_6 NI_6 NS_791 0 6.3571562313446267e-03
GC_6_792 b_6 NI_6 NS_792 0 -1.8769366072077583e-03
GC_6_793 b_6 NI_6 NS_793 0 -5.4767784441416244e-03
GC_6_794 b_6 NI_6 NS_794 0 2.1761634539402015e-03
GC_6_795 b_6 NI_6 NS_795 0 5.3904708368408541e-03
GC_6_796 b_6 NI_6 NS_796 0 -2.6291409730218114e-03
GC_6_797 b_6 NI_6 NS_797 0 -6.3068613300950385e-03
GC_6_798 b_6 NI_6 NS_798 0 -4.8944546422454794e-04
GC_6_799 b_6 NI_6 NS_799 0 7.6383029102316431e-03
GC_6_800 b_6 NI_6 NS_800 0 3.6283278334162559e-03
GC_6_801 b_6 NI_6 NS_801 0 -5.8333235006030430e-03
GC_6_802 b_6 NI_6 NS_802 0 -3.4684301765322894e-03
GC_6_803 b_6 NI_6 NS_803 0 2.9592188619425685e-04
GC_6_804 b_6 NI_6 NS_804 0 5.5702924793220364e-04
GC_6_805 b_6 NI_6 NS_805 0 -4.9284028867594898e-03
GC_6_806 b_6 NI_6 NS_806 0 8.8733927007926192e-04
GC_6_807 b_6 NI_6 NS_807 0 6.2016450885671775e-03
GC_6_808 b_6 NI_6 NS_808 0 6.8248096800231899e-04
GC_6_809 b_6 NI_6 NS_809 0 -5.3226827419087528e-03
GC_6_810 b_6 NI_6 NS_810 0 -4.8918921539248044e-04
GC_6_811 b_6 NI_6 NS_811 0 1.5482735936977537e-03
GC_6_812 b_6 NI_6 NS_812 0 -4.6609097844113840e-05
GC_6_813 b_6 NI_6 NS_813 0 -6.0242735565756373e-03
GC_6_814 b_6 NI_6 NS_814 0 1.9161516125140510e-03
GC_6_815 b_6 NI_6 NS_815 0 6.2494033703015981e-03
GC_6_816 b_6 NI_6 NS_816 0 2.0850497458901803e-04
GC_6_817 b_6 NI_6 NS_817 0 -5.0636589476607090e-03
GC_6_818 b_6 NI_6 NS_818 0 1.6954532766883591e-03
GC_6_819 b_6 NI_6 NS_819 0 2.4806588151513086e-03
GC_6_820 b_6 NI_6 NS_820 0 -9.6015728238764875e-04
GC_6_821 b_6 NI_6 NS_821 0 -6.5381320997607217e-03
GC_6_822 b_6 NI_6 NS_822 0 3.8750074877559556e-03
GC_6_823 b_6 NI_6 NS_823 0 7.4722547471554072e-03
GC_6_824 b_6 NI_6 NS_824 0 -1.0944729982741304e-03
GC_6_825 b_6 NI_6 NS_825 0 -3.9943218502332123e-03
GC_6_826 b_6 NI_6 NS_826 0 4.0357752359328229e-03
GC_6_827 b_6 NI_6 NS_827 0 2.8552014001051273e-03
GC_6_828 b_6 NI_6 NS_828 0 -3.0472625143400278e-03
GC_6_829 b_6 NI_6 NS_829 0 -6.0351388735177666e-03
GC_6_830 b_6 NI_6 NS_830 0 7.2276062239162477e-03
GC_6_831 b_6 NI_6 NS_831 0 7.9782887395805496e-03
GC_6_832 b_6 NI_6 NS_832 0 -4.7935802390633867e-03
GC_6_833 b_6 NI_6 NS_833 0 -5.4799473742592544e-04
GC_6_834 b_6 NI_6 NS_834 0 5.0230804803337659e-03
GC_6_835 b_6 NI_6 NS_835 0 2.5034134498541210e-04
GC_6_836 b_6 NI_6 NS_836 0 -4.7520661524518056e-03
GC_6_837 b_6 NI_6 NS_837 0 1.7366273020420207e-09
GC_6_838 b_6 NI_6 NS_838 0 3.2860219100722032e-09
GC_6_839 b_6 NI_6 NS_839 0 -1.4394124885463602e-03
GC_6_840 b_6 NI_6 NS_840 0 7.8706604719082068e-03
GC_6_841 b_6 NI_6 NS_841 0 -1.8574746552919573e-04
GC_6_842 b_6 NI_6 NS_842 0 3.0287972650494101e-03
GC_6_843 b_6 NI_6 NS_843 0 -1.2900533253323610e-04
GC_6_844 b_6 NI_6 NS_844 0 -3.3736684356684204e-03
GC_6_845 b_6 NI_6 NS_845 0 -8.9083180904216965e-04
GC_6_846 b_6 NI_6 NS_846 0 7.5293774109586944e-03
GC_6_847 b_6 NI_6 NS_847 0 3.7906243942544358e-03
GC_6_848 b_6 NI_6 NS_848 0 -6.1490577537347806e-03
GC_6_849 b_6 NI_6 NS_849 0 8.8448812800164688e-08
GC_6_850 b_6 NI_6 NS_850 0 -3.5531433930158850e-07
GC_6_851 b_6 NI_6 NS_851 0 6.7115065644237299e-03
GC_6_852 b_6 NI_6 NS_852 0 -5.3183245801309833e-03
GC_6_853 b_6 NI_6 NS_853 0 -2.6127433844451969e-03
GC_6_854 b_6 NI_6 NS_854 0 6.0487711490434552e-03
GC_6_855 b_6 NI_6 NS_855 0 -4.2945275031913326e-03
GC_6_856 b_6 NI_6 NS_856 0 1.3261561751562693e-05
GC_6_857 b_6 NI_6 NS_857 0 2.7224992743036238e-03
GC_6_858 b_6 NI_6 NS_858 0 -6.1956590921680354e-03
GC_6_859 b_6 NI_6 NS_859 0 2.0898364070663007e-03
GC_6_860 b_6 NI_6 NS_860 0 3.2611136133748951e-03
GC_6_861 b_6 NI_6 NS_861 0 -1.9638287434536657e-03
GC_6_862 b_6 NI_6 NS_862 0 -4.4203348271417177e-03
GC_6_863 b_6 NI_6 NS_863 0 2.8567435038813417e-03
GC_6_864 b_6 NI_6 NS_864 0 8.0017787559365054e-03
GC_6_865 b_6 NI_6 NS_865 0 -1.4324864070388216e-04
GC_6_866 b_6 NI_6 NS_866 0 3.4599467632020393e-11
GC_6_867 b_6 NI_6 NS_867 0 3.0174581320017198e-11
GC_6_868 b_6 NI_6 NS_868 0 9.4202339998135707e-10
GC_6_869 b_6 NI_6 NS_869 0 -2.1091457317140727e-06
GC_6_870 b_6 NI_6 NS_870 0 -1.6534096847357484e-06
GC_6_871 b_6 NI_6 NS_871 0 1.8892051209049264e-06
GC_6_872 b_6 NI_6 NS_872 0 3.8449850343838746e-06
GC_6_873 b_6 NI_6 NS_873 0 3.2880567322659333e-06
GC_6_874 b_6 NI_6 NS_874 0 4.9269638868930100e-06
GC_6_875 b_6 NI_6 NS_875 0 5.8302987679642168e-06
GC_6_876 b_6 NI_6 NS_876 0 -9.0830944448677718e-06
GC_6_877 b_6 NI_6 NS_877 0 -2.5402013598986857e-06
GC_6_878 b_6 NI_6 NS_878 0 -1.3835961776218204e-05
GC_6_879 b_6 NI_6 NS_879 0 -3.5342732938184657e-06
GC_6_880 b_6 NI_6 NS_880 0 2.1966333005944464e-06
GC_6_881 b_6 NI_6 NS_881 0 3.6391305956678683e-06
GC_6_882 b_6 NI_6 NS_882 0 1.2970513585538672e-06
GC_6_883 b_6 NI_6 NS_883 0 7.8997729679709276e-06
GC_6_884 b_6 NI_6 NS_884 0 -3.9683335078830703e-05
GC_6_885 b_6 NI_6 NS_885 0 -4.4005792825484432e-05
GC_6_886 b_6 NI_6 NS_886 0 -8.8282327276510609e-07
GC_6_887 b_6 NI_6 NS_887 0 -1.4766050615859493e-05
GC_6_888 b_6 NI_6 NS_888 0 -8.4725925754117908e-06
GC_6_889 b_6 NI_6 NS_889 0 -7.2348590426860566e-05
GC_6_890 b_6 NI_6 NS_890 0 7.5140396584880769e-05
GC_6_891 b_6 NI_6 NS_891 0 4.6495319187927653e-06
GC_6_892 b_6 NI_6 NS_892 0 1.3009967517210407e-05
GC_6_893 b_6 NI_6 NS_893 0 6.2665097400042415e-05
GC_6_894 b_6 NI_6 NS_894 0 1.2224194269646658e-04
GC_6_895 b_6 NI_6 NS_895 0 2.4457335768479032e-07
GC_6_896 b_6 NI_6 NS_896 0 -3.6753277840645116e-05
GC_6_897 b_6 NI_6 NS_897 0 1.6411258782030658e-05
GC_6_898 b_6 NI_6 NS_898 0 3.8871919102622316e-06
GC_6_899 b_6 NI_6 NS_899 0 2.4219128417047415e-05
GC_6_900 b_6 NI_6 NS_900 0 -3.0244018059555093e-05
GC_6_901 b_6 NI_6 NS_901 0 -8.8437631769636924e-06
GC_6_902 b_6 NI_6 NS_902 0 -2.2761552315330025e-06
GC_6_903 b_6 NI_6 NS_903 0 -8.7280491673389642e-06
GC_6_904 b_6 NI_6 NS_904 0 2.5050975032957038e-05
GC_6_905 b_6 NI_6 NS_905 0 5.8325735593331687e-06
GC_6_906 b_6 NI_6 NS_906 0 8.3788316390864721e-06
GC_6_907 b_6 NI_6 NS_907 0 5.5969447649002548e-05
GC_6_908 b_6 NI_6 NS_908 0 2.4647593554246866e-05
GC_6_909 b_6 NI_6 NS_909 0 3.4492085952306533e-06
GC_6_910 b_6 NI_6 NS_910 0 -1.1606262499177152e-05
GC_6_911 b_6 NI_6 NS_911 0 -4.0620355742236124e-07
GC_6_912 b_6 NI_6 NS_912 0 -1.2991929005260041e-06
GC_6_913 b_6 NI_6 NS_913 0 6.7879721140405351e-06
GC_6_914 b_6 NI_6 NS_914 0 3.0205805034449130e-06
GC_6_915 b_6 NI_6 NS_915 0 4.1592022079281475e-05
GC_6_916 b_6 NI_6 NS_916 0 -1.7165656659661355e-05
GC_6_917 b_6 NI_6 NS_917 0 -2.5738414942771147e-06
GC_6_918 b_6 NI_6 NS_918 0 -7.0283371096076546e-06
GC_6_919 b_6 NI_6 NS_919 0 -2.9900618733030672e-06
GC_6_920 b_6 NI_6 NS_920 0 1.7603142920091398e-06
GC_6_921 b_6 NI_6 NS_921 0 9.5385441624539742e-06
GC_6_922 b_6 NI_6 NS_922 0 2.8682883723567672e-06
GC_6_923 b_6 NI_6 NS_923 0 2.2731559503514391e-05
GC_6_924 b_6 NI_6 NS_924 0 -3.1037614858118868e-05
GC_6_925 b_6 NI_6 NS_925 0 -5.6871533623039327e-06
GC_6_926 b_6 NI_6 NS_926 0 -3.6246179722499213e-06
GC_6_927 b_6 NI_6 NS_927 0 -5.2395965286833206e-07
GC_6_928 b_6 NI_6 NS_928 0 5.0176248988801396e-06
GC_6_929 b_6 NI_6 NS_929 0 1.2253679910732575e-05
GC_6_930 b_6 NI_6 NS_930 0 1.7531652179123602e-07
GC_6_931 b_6 NI_6 NS_931 0 1.8083170695188806e-06
GC_6_932 b_6 NI_6 NS_932 0 -3.1349940458809069e-05
GC_6_933 b_6 NI_6 NS_933 0 -6.7180468929919325e-06
GC_6_934 b_6 NI_6 NS_934 0 9.7548984033982666e-07
GC_6_935 b_6 NI_6 NS_935 0 4.6118149147777729e-06
GC_6_936 b_6 NI_6 NS_936 0 3.8655024353917893e-06
GC_6_937 b_6 NI_6 NS_937 0 1.4061852739223348e-05
GC_6_938 b_6 NI_6 NS_938 0 -6.0101949940870876e-06
GC_6_939 b_6 NI_6 NS_939 0 -1.4015897413645019e-05
GC_6_940 b_6 NI_6 NS_940 0 -1.8747008544404041e-05
GC_6_941 b_6 NI_6 NS_941 0 -2.5061617140895530e-06
GC_6_942 b_6 NI_6 NS_942 0 5.4162182926779556e-06
GC_6_943 b_6 NI_6 NS_943 0 4.6576524122395444e-06
GC_6_944 b_6 NI_6 NS_944 0 -2.0834711745067344e-06
GC_6_945 b_6 NI_6 NS_945 0 -1.4565769591338177e-11
GC_6_946 b_6 NI_6 NS_946 0 4.2046046964607029e-12
GC_6_947 b_6 NI_6 NS_947 0 5.1979791464288049e-06
GC_6_948 b_6 NI_6 NS_948 0 -1.1242606331306605e-05
GC_6_949 b_6 NI_6 NS_949 0 -2.6676589020784989e-07
GC_6_950 b_6 NI_6 NS_950 0 2.9264564739919444e-06
GC_6_951 b_6 NI_6 NS_951 0 2.6445021056645551e-06
GC_6_952 b_6 NI_6 NS_952 0 -1.5935958540201036e-06
GC_6_953 b_6 NI_6 NS_953 0 2.4076268287215001e-06
GC_6_954 b_6 NI_6 NS_954 0 -9.4308107605498062e-06
GC_6_955 b_6 NI_6 NS_955 0 -9.9265954482454993e-06
GC_6_956 b_6 NI_6 NS_956 0 -3.6884528492557378e-06
GC_6_957 b_6 NI_6 NS_957 0 3.1234824120851768e-10
GC_6_958 b_6 NI_6 NS_958 0 2.7697760132315182e-10
GC_6_959 b_6 NI_6 NS_959 0 -8.5916096677855126e-06
GC_6_960 b_6 NI_6 NS_960 0 -5.6865018401105187e-06
GC_6_961 b_6 NI_6 NS_961 0 2.2662363177774279e-06
GC_6_962 b_6 NI_6 NS_962 0 -6.4520167074772378e-06
GC_6_963 b_6 NI_6 NS_963 0 -3.0673941811149788e-06
GC_6_964 b_6 NI_6 NS_964 0 -1.3540707208082387e-07
GC_6_965 b_6 NI_6 NS_965 0 -7.9220182963082988e-06
GC_6_966 b_6 NI_6 NS_966 0 4.8453491833371352e-07
GC_6_967 b_6 NI_6 NS_967 0 3.0018482516193619e-06
GC_6_968 b_6 NI_6 NS_968 0 2.8730585708417800e-06
GC_6_969 b_6 NI_6 NS_969 0 1.2171961224846272e-06
GC_6_970 b_6 NI_6 NS_970 0 -3.8814955134215981e-06
GC_6_971 b_6 NI_6 NS_971 0 -4.8737987917712779e-06
GC_6_972 b_6 NI_6 NS_972 0 -3.9067803325292269e-06
GC_6_973 b_6 NI_6 NS_973 0 -3.0637392627561084e-05
GC_6_974 b_6 NI_6 NS_974 0 -1.9701788900989091e-12
GC_6_975 b_6 NI_6 NS_975 0 -2.2726002432827514e-10
GC_6_976 b_6 NI_6 NS_976 0 1.0440684633505415e-08
GC_6_977 b_6 NI_6 NS_977 0 6.9327075003054653e-07
GC_6_978 b_6 NI_6 NS_978 0 1.0332693288744298e-07
GC_6_979 b_6 NI_6 NS_979 0 3.1648136438565568e-06
GC_6_980 b_6 NI_6 NS_980 0 -1.3944687702703775e-06
GC_6_981 b_6 NI_6 NS_981 0 -2.7897599646584512e-06
GC_6_982 b_6 NI_6 NS_982 0 -2.8314313832247718e-06
GC_6_983 b_6 NI_6 NS_983 0 4.9208217028607224e-06
GC_6_984 b_6 NI_6 NS_984 0 -5.3538933989723200e-07
GC_6_985 b_6 NI_6 NS_985 0 -7.0691797507249311e-06
GC_6_986 b_6 NI_6 NS_986 0 -8.1237002541663642e-06
GC_6_987 b_6 NI_6 NS_987 0 1.8605993430755484e-08
GC_6_988 b_6 NI_6 NS_988 0 -1.5534374209472310e-06
GC_6_989 b_6 NI_6 NS_989 0 -6.0814386714532330e-06
GC_6_990 b_6 NI_6 NS_990 0 1.9319036551972675e-06
GC_6_991 b_6 NI_6 NS_991 0 5.3119887789057661e-06
GC_6_992 b_6 NI_6 NS_992 0 -5.7335801442955760e-06
GC_6_993 b_6 NI_6 NS_993 0 -1.7096906077749549e-05
GC_6_994 b_6 NI_6 NS_994 0 4.6242225665948065e-06
GC_6_995 b_6 NI_6 NS_995 0 -1.1944686918143934e-06
GC_6_996 b_6 NI_6 NS_996 0 7.0592835588547843e-06
GC_6_997 b_6 NI_6 NS_997 0 -7.2285772523319732e-06
GC_6_998 b_6 NI_6 NS_998 0 -4.5688870227889859e-06
GC_6_999 b_6 NI_6 NS_999 0 -3.3893053275519803e-06
GC_6_1000 b_6 NI_6 NS_1000 0 7.9766987733916595e-06
GC_6_1001 b_6 NI_6 NS_1001 0 -2.2427659551997014e-06
GC_6_1002 b_6 NI_6 NS_1002 0 -4.6664999979183040e-06
GC_6_1003 b_6 NI_6 NS_1003 0 -3.8807669960726156e-06
GC_6_1004 b_6 NI_6 NS_1004 0 1.1289712256580433e-05
GC_6_1005 b_6 NI_6 NS_1005 0 -1.9128083374255178e-07
GC_6_1006 b_6 NI_6 NS_1006 0 7.1636505735151789e-06
GC_6_1007 b_6 NI_6 NS_1007 0 -4.1441824359101055e-06
GC_6_1008 b_6 NI_6 NS_1008 0 1.2150894653025325e-06
GC_6_1009 b_6 NI_6 NS_1009 0 -6.4403623064902790e-07
GC_6_1010 b_6 NI_6 NS_1010 0 7.9591241419361221e-06
GC_6_1011 b_6 NI_6 NS_1011 0 -1.0603801532821055e-06
GC_6_1012 b_6 NI_6 NS_1012 0 2.1884897969850647e-06
GC_6_1013 b_6 NI_6 NS_1013 0 -2.4285512394424080e-06
GC_6_1014 b_6 NI_6 NS_1014 0 8.0706353141039482e-06
GC_6_1015 b_6 NI_6 NS_1015 0 -1.7503981933420986e-07
GC_6_1016 b_6 NI_6 NS_1016 0 9.4003707188776012e-06
GC_6_1017 b_6 NI_6 NS_1017 0 -8.8143844632507627e-07
GC_6_1018 b_6 NI_6 NS_1018 0 8.6988676679423796e-06
GC_6_1019 b_6 NI_6 NS_1019 0 -1.3355222536180013e-06
GC_6_1020 b_6 NI_6 NS_1020 0 3.8589146292692184e-06
GC_6_1021 b_6 NI_6 NS_1021 0 9.5135043942930140e-07
GC_6_1022 b_6 NI_6 NS_1022 0 1.1830488743677764e-05
GC_6_1023 b_6 NI_6 NS_1023 0 1.7339678181432823e-05
GC_6_1024 b_6 NI_6 NS_1024 0 1.6620957406980684e-05
GC_6_1025 b_6 NI_6 NS_1025 0 4.6876734722830669e-06
GC_6_1026 b_6 NI_6 NS_1026 0 7.6215654801057031e-06
GC_6_1027 b_6 NI_6 NS_1027 0 9.8092198845097941e-06
GC_6_1028 b_6 NI_6 NS_1028 0 3.8277643400692211e-06
GC_6_1029 b_6 NI_6 NS_1029 0 6.4308508352105446e-06
GC_6_1030 b_6 NI_6 NS_1030 0 1.0600263312473105e-05
GC_6_1031 b_6 NI_6 NS_1031 0 3.1894622562952962e-05
GC_6_1032 b_6 NI_6 NS_1032 0 -5.8207799226560567e-06
GC_6_1033 b_6 NI_6 NS_1033 0 7.7815651621449348e-06
GC_6_1034 b_6 NI_6 NS_1034 0 3.3341158985119182e-06
GC_6_1035 b_6 NI_6 NS_1035 0 1.1392291394593068e-05
GC_6_1036 b_6 NI_6 NS_1036 0 -9.9543851766476265e-06
GC_6_1037 b_6 NI_6 NS_1037 0 1.0335938050039953e-05
GC_6_1038 b_6 NI_6 NS_1038 0 6.2186471320492545e-06
GC_6_1039 b_6 NI_6 NS_1039 0 1.5858030353626564e-05
GC_6_1040 b_6 NI_6 NS_1040 0 -2.9884766593588657e-05
GC_6_1041 b_6 NI_6 NS_1041 0 7.7006040529127063e-06
GC_6_1042 b_6 NI_6 NS_1042 0 -2.8908264810862044e-06
GC_6_1043 b_6 NI_6 NS_1043 0 -3.4539415772998637e-06
GC_6_1044 b_6 NI_6 NS_1044 0 -1.5715634433190754e-05
GC_6_1045 b_6 NI_6 NS_1045 0 1.1293336763338488e-05
GC_6_1046 b_6 NI_6 NS_1046 0 -1.7359447111238037e-06
GC_6_1047 b_6 NI_6 NS_1047 0 -1.3020290064558145e-05
GC_6_1048 b_6 NI_6 NS_1048 0 -2.4148618036394421e-05
GC_6_1049 b_6 NI_6 NS_1049 0 -4.2214977119029767e-07
GC_6_1050 b_6 NI_6 NS_1050 0 -6.3952475510301904e-06
GC_6_1051 b_6 NI_6 NS_1051 0 -9.5214715151193812e-06
GC_6_1052 b_6 NI_6 NS_1052 0 -2.3393117943722041e-06
GC_6_1053 b_6 NI_6 NS_1053 0 9.7737469529915419e-11
GC_6_1054 b_6 NI_6 NS_1054 0 5.3682970592318579e-11
GC_6_1055 b_6 NI_6 NS_1055 0 1.1864487993221074e-06
GC_6_1056 b_6 NI_6 NS_1056 0 -4.6217717348696747e-06
GC_6_1057 b_6 NI_6 NS_1057 0 -1.4846152847397040e-06
GC_6_1058 b_6 NI_6 NS_1058 0 -1.2851849410326793e-06
GC_6_1059 b_6 NI_6 NS_1059 0 -4.9361111558349093e-06
GC_6_1060 b_6 NI_6 NS_1060 0 -8.7754694675992366e-07
GC_6_1061 b_6 NI_6 NS_1061 0 -1.3873432084914194e-06
GC_6_1062 b_6 NI_6 NS_1062 0 -2.8331812727207967e-06
GC_6_1063 b_6 NI_6 NS_1063 0 -1.0078501125690919e-05
GC_6_1064 b_6 NI_6 NS_1064 0 -3.6998807613256413e-06
GC_6_1065 b_6 NI_6 NS_1065 0 6.6046400030560755e-09
GC_6_1066 b_6 NI_6 NS_1066 0 5.7462999558495321e-09
GC_6_1067 b_6 NI_6 NS_1067 0 1.3894890386921221e-06
GC_6_1068 b_6 NI_6 NS_1068 0 6.7846014562375019e-07
GC_6_1069 b_6 NI_6 NS_1069 0 -1.7344558258936674e-06
GC_6_1070 b_6 NI_6 NS_1070 0 3.1417316060333096e-06
GC_6_1071 b_6 NI_6 NS_1071 0 -9.2518097978972977e-07
GC_6_1072 b_6 NI_6 NS_1072 0 7.7635650409730743e-07
GC_6_1073 b_6 NI_6 NS_1073 0 -7.9006813972920457e-06
GC_6_1074 b_6 NI_6 NS_1074 0 8.1641422599338337e-07
GC_6_1075 b_6 NI_6 NS_1075 0 -2.4105961034727568e-06
GC_6_1076 b_6 NI_6 NS_1076 0 2.0859203667112411e-06
GC_6_1077 b_6 NI_6 NS_1077 0 -2.1253693848796860e-06
GC_6_1078 b_6 NI_6 NS_1078 0 2.1337375380059271e-06
GC_6_1079 b_6 NI_6 NS_1079 0 1.1308769262448768e-06
GC_6_1080 b_6 NI_6 NS_1080 0 2.8161633841349760e-06
GC_6_1081 b_6 NI_6 NS_1081 0 -9.0136324675633118e-05
GC_6_1082 b_6 NI_6 NS_1082 0 7.1502555862506125e-12
GC_6_1083 b_6 NI_6 NS_1083 0 -5.7297248174278353e-11
GC_6_1084 b_6 NI_6 NS_1084 0 3.3361295279621262e-10
GC_6_1085 b_6 NI_6 NS_1085 0 -1.5721767629538323e-06
GC_6_1086 b_6 NI_6 NS_1086 0 -1.5573912424820836e-06
GC_6_1087 b_6 NI_6 NS_1087 0 9.4297753429023430e-07
GC_6_1088 b_6 NI_6 NS_1088 0 7.2566254607475550e-07
GC_6_1089 b_6 NI_6 NS_1089 0 -2.7196303334875077e-06
GC_6_1090 b_6 NI_6 NS_1090 0 3.0307848496909001e-06
GC_6_1091 b_6 NI_6 NS_1091 0 -3.0496638824230564e-06
GC_6_1092 b_6 NI_6 NS_1092 0 -2.5769713216498874e-06
GC_6_1093 b_6 NI_6 NS_1093 0 1.5158968923593623e-06
GC_6_1094 b_6 NI_6 NS_1094 0 9.0893433349421315e-08
GC_6_1095 b_6 NI_6 NS_1095 0 -1.6657821916929438e-06
GC_6_1096 b_6 NI_6 NS_1096 0 1.7972653937360592e-06
GC_6_1097 b_6 NI_6 NS_1097 0 8.9123525014313650e-07
GC_6_1098 b_6 NI_6 NS_1098 0 4.1366205450534416e-06
GC_6_1099 b_6 NI_6 NS_1099 0 -4.2927672867884478e-06
GC_6_1100 b_6 NI_6 NS_1100 0 -2.0599997759971169e-06
GC_6_1101 b_6 NI_6 NS_1101 0 2.3787683629134253e-06
GC_6_1102 b_6 NI_6 NS_1102 0 -1.9358839831990853e-06
GC_6_1103 b_6 NI_6 NS_1103 0 -1.1788210641087254e-06
GC_6_1104 b_6 NI_6 NS_1104 0 3.2601431197261090e-06
GC_6_1105 b_6 NI_6 NS_1105 0 -8.4124102124693396e-06
GC_6_1106 b_6 NI_6 NS_1106 0 1.1213008488202299e-05
GC_6_1107 b_6 NI_6 NS_1107 0 1.2598096429606961e-06
GC_6_1108 b_6 NI_6 NS_1108 0 -1.6518673655730096e-06
GC_6_1109 b_6 NI_6 NS_1109 0 9.9604694056384736e-06
GC_6_1110 b_6 NI_6 NS_1110 0 1.7407374017860053e-05
GC_6_1111 b_6 NI_6 NS_1111 0 -6.6234898443768555e-07
GC_6_1112 b_6 NI_6 NS_1112 0 -5.4666971754082105e-07
GC_6_1113 b_6 NI_6 NS_1113 0 4.5572771096953712e-07
GC_6_1114 b_6 NI_6 NS_1114 0 -1.3700998658097223e-06
GC_6_1115 b_6 NI_6 NS_1115 0 7.0273615567041306e-06
GC_6_1116 b_6 NI_6 NS_1116 0 -2.3133395482826009e-07
GC_6_1117 b_6 NI_6 NS_1117 0 6.9999672531334962e-07
GC_6_1118 b_6 NI_6 NS_1118 0 2.9955126122386900e-06
GC_6_1119 b_6 NI_6 NS_1119 0 4.4108793973868417e-07
GC_6_1120 b_6 NI_6 NS_1120 0 2.9100613166788581e-06
GC_6_1121 b_6 NI_6 NS_1121 0 1.1671201397215561e-06
GC_6_1122 b_6 NI_6 NS_1122 0 -1.4115770154417524e-06
GC_6_1123 b_6 NI_6 NS_1123 0 9.4124669791332229e-06
GC_6_1124 b_6 NI_6 NS_1124 0 5.2153716915289170e-06
GC_6_1125 b_6 NI_6 NS_1125 0 5.7060076692084278e-07
GC_6_1126 b_6 NI_6 NS_1126 0 1.1337175239046775e-06
GC_6_1127 b_6 NI_6 NS_1127 0 5.6635657211078908e-08
GC_6_1128 b_6 NI_6 NS_1128 0 4.4780048583390847e-07
GC_6_1129 b_6 NI_6 NS_1129 0 1.2930173453017109e-06
GC_6_1130 b_6 NI_6 NS_1130 0 -8.5758344478152843e-07
GC_6_1131 b_6 NI_6 NS_1131 0 9.1863075729678575e-06
GC_6_1132 b_6 NI_6 NS_1132 0 6.5375039287412692e-07
GC_6_1133 b_6 NI_6 NS_1133 0 8.3834867855354149e-07
GC_6_1134 b_6 NI_6 NS_1134 0 1.4354668713502649e-06
GC_6_1135 b_6 NI_6 NS_1135 0 1.0193399835208624e-06
GC_6_1136 b_6 NI_6 NS_1136 0 5.8698357721206326e-07
GC_6_1137 b_6 NI_6 NS_1137 0 1.3710352364329224e-06
GC_6_1138 b_6 NI_6 NS_1138 0 -9.5622299128214045e-07
GC_6_1139 b_6 NI_6 NS_1139 0 8.0098262742061443e-06
GC_6_1140 b_6 NI_6 NS_1140 0 -2.1610484136729379e-06
GC_6_1141 b_6 NI_6 NS_1141 0 1.1721236843559445e-06
GC_6_1142 b_6 NI_6 NS_1142 0 1.5263103790329470e-06
GC_6_1143 b_6 NI_6 NS_1143 0 1.5749311925884211e-06
GC_6_1144 b_6 NI_6 NS_1144 0 -2.5367781262157637e-07
GC_6_1145 b_6 NI_6 NS_1145 0 1.3308042121153192e-06
GC_6_1146 b_6 NI_6 NS_1146 0 -1.0066157831291740e-06
GC_6_1147 b_6 NI_6 NS_1147 0 5.7892180576794180e-06
GC_6_1148 b_6 NI_6 NS_1148 0 -3.9086683510452168e-06
GC_6_1149 b_6 NI_6 NS_1149 0 1.8024603896025247e-06
GC_6_1150 b_6 NI_6 NS_1150 0 1.4095139378120783e-06
GC_6_1151 b_6 NI_6 NS_1151 0 1.0763959891285198e-06
GC_6_1152 b_6 NI_6 NS_1152 0 -1.4081557091405275e-06
GC_6_1153 b_6 NI_6 NS_1153 0 1.4146271252184701e-06
GC_6_1154 b_6 NI_6 NS_1154 0 -1.1369767640502012e-06
GC_6_1155 b_6 NI_6 NS_1155 0 2.9379344018858220e-06
GC_6_1156 b_6 NI_6 NS_1156 0 -4.1714633763493070e-06
GC_6_1157 b_6 NI_6 NS_1157 0 2.2085081851629802e-06
GC_6_1158 b_6 NI_6 NS_1158 0 2.9634104900437647e-07
GC_6_1159 b_6 NI_6 NS_1159 0 -3.3704622656083913e-07
GC_6_1160 b_6 NI_6 NS_1160 0 -1.1837401272903804e-06
GC_6_1161 b_6 NI_6 NS_1161 0 2.4875083328704189e-11
GC_6_1162 b_6 NI_6 NS_1162 0 -4.0913108544532353e-11
GC_6_1163 b_6 NI_6 NS_1163 0 7.8538972831461179e-07
GC_6_1164 b_6 NI_6 NS_1164 0 -1.5911479702283517e-06
GC_6_1165 b_6 NI_6 NS_1165 0 1.2557723578829168e-06
GC_6_1166 b_6 NI_6 NS_1166 0 2.2315376579670528e-07
GC_6_1167 b_6 NI_6 NS_1167 0 1.5659218838254300e-07
GC_6_1168 b_6 NI_6 NS_1168 0 -5.4948818560856513e-07
GC_6_1169 b_6 NI_6 NS_1169 0 5.4537121389050551e-07
GC_6_1170 b_6 NI_6 NS_1170 0 -8.9276718239199553e-07
GC_6_1171 b_6 NI_6 NS_1171 0 1.2830273724135556e-06
GC_6_1172 b_6 NI_6 NS_1172 0 -2.0549369121533973e-06
GC_6_1173 b_6 NI_6 NS_1173 0 4.7366134917157180e-10
GC_6_1174 b_6 NI_6 NS_1174 0 -1.2085642547890880e-09
GC_6_1175 b_6 NI_6 NS_1175 0 5.4539170274125565e-07
GC_6_1176 b_6 NI_6 NS_1176 0 -8.5655969664391391e-07
GC_6_1177 b_6 NI_6 NS_1177 0 7.1232733492307373e-07
GC_6_1178 b_6 NI_6 NS_1178 0 -9.5180807724037970e-07
GC_6_1179 b_6 NI_6 NS_1179 0 8.8751985551023756e-08
GC_6_1180 b_6 NI_6 NS_1180 0 5.0688941439428539e-08
GC_6_1181 b_6 NI_6 NS_1181 0 1.3271496873867863e-06
GC_6_1182 b_6 NI_6 NS_1182 0 -1.2248142507374969e-06
GC_6_1183 b_6 NI_6 NS_1183 0 1.6449395225540219e-06
GC_6_1184 b_6 NI_6 NS_1184 0 -2.9372095525334584e-07
GC_6_1185 b_6 NI_6 NS_1185 0 -2.3012991323750509e-07
GC_6_1186 b_6 NI_6 NS_1186 0 -7.3458670407458323e-07
GC_6_1187 b_6 NI_6 NS_1187 0 7.3260767551048154e-07
GC_6_1188 b_6 NI_6 NS_1188 0 2.8937258575640461e-07
GC_6_1189 b_6 NI_6 NS_1189 0 4.9622892078738299e-05
GC_6_1190 b_6 NI_6 NS_1190 0 3.6303232873700738e-12
GC_6_1191 b_6 NI_6 NS_1191 0 -4.1065119835124740e-12
GC_6_1192 b_6 NI_6 NS_1192 0 9.4552646741476397e-10
GC_6_1193 b_6 NI_6 NS_1193 0 -4.5592729239358077e-08
GC_6_1194 b_6 NI_6 NS_1194 0 2.5302102935711645e-07
GC_6_1195 b_6 NI_6 NS_1195 0 2.5930072744228142e-07
GC_6_1196 b_6 NI_6 NS_1196 0 4.0791660376520017e-07
GC_6_1197 b_6 NI_6 NS_1197 0 -1.3649523336941601e-07
GC_6_1198 b_6 NI_6 NS_1198 0 2.4393638864996197e-07
GC_6_1199 b_6 NI_6 NS_1199 0 7.8203514142467763e-07
GC_6_1200 b_6 NI_6 NS_1200 0 1.4417034245792251e-06
GC_6_1201 b_6 NI_6 NS_1201 0 1.0397084214724829e-06
GC_6_1202 b_6 NI_6 NS_1202 0 -5.2292443105339315e-07
GC_6_1203 b_6 NI_6 NS_1203 0 3.3637638265764777e-07
GC_6_1204 b_6 NI_6 NS_1204 0 8.8673923929050186e-07
GC_6_1205 b_6 NI_6 NS_1205 0 7.3264031448761284e-07
GC_6_1206 b_6 NI_6 NS_1206 0 -3.6972329301733256e-07
GC_6_1207 b_6 NI_6 NS_1207 0 4.3588550018348819e-06
GC_6_1208 b_6 NI_6 NS_1208 0 1.3805937882958914e-06
GC_6_1209 b_6 NI_6 NS_1209 0 -1.6438411660936222e-06
GC_6_1210 b_6 NI_6 NS_1210 0 -3.5789182254246461e-06
GC_6_1211 b_6 NI_6 NS_1211 0 2.4006573946843829e-07
GC_6_1212 b_6 NI_6 NS_1212 0 1.5509787143483403e-06
GC_6_1213 b_6 NI_6 NS_1213 0 2.9713807086122570e-06
GC_6_1214 b_6 NI_6 NS_1214 0 -4.7497997904785026e-06
GC_6_1215 b_6 NI_6 NS_1215 0 -7.7198179823281751e-07
GC_6_1216 b_6 NI_6 NS_1216 0 5.6526085814021255e-07
GC_6_1217 b_6 NI_6 NS_1217 0 5.5714203379849249e-06
GC_6_1218 b_6 NI_6 NS_1218 0 -5.8239761940734889e-06
GC_6_1219 b_6 NI_6 NS_1219 0 -3.3126924551666642e-06
GC_6_1220 b_6 NI_6 NS_1220 0 1.7946939167787273e-06
GC_6_1221 b_6 NI_6 NS_1221 0 8.6225856884913098e-07
GC_6_1222 b_6 NI_6 NS_1222 0 1.2280691633840723e-06
GC_6_1223 b_6 NI_6 NS_1223 0 1.5935580397522229e-06
GC_6_1224 b_6 NI_6 NS_1224 0 -4.1016196624991178e-06
GC_6_1225 b_6 NI_6 NS_1225 0 5.6918432674550418e-07
GC_6_1226 b_6 NI_6 NS_1226 0 1.9886999347009612e-07
GC_6_1227 b_6 NI_6 NS_1227 0 1.7374832420059089e-07
GC_6_1228 b_6 NI_6 NS_1228 0 -4.0365325732244473e-06
GC_6_1229 b_6 NI_6 NS_1229 0 -1.8756568232188815e-07
GC_6_1230 b_6 NI_6 NS_1230 0 1.6738459329504198e-07
GC_6_1231 b_6 NI_6 NS_1231 0 4.6371532258191252e-06
GC_6_1232 b_6 NI_6 NS_1232 0 -6.3342163801214933e-06
GC_6_1233 b_6 NI_6 NS_1233 0 -1.8279082401390849e-06
GC_6_1234 b_6 NI_6 NS_1234 0 -1.2891003720581293e-06
GC_6_1235 b_6 NI_6 NS_1235 0 1.3669285990901595e-06
GC_6_1236 b_6 NI_6 NS_1236 0 -1.1987254571348222e-06
GC_6_1237 b_6 NI_6 NS_1237 0 3.7640843439794355e-07
GC_6_1238 b_6 NI_6 NS_1238 0 -2.0979974752339792e-06
GC_6_1239 b_6 NI_6 NS_1239 0 -1.4883372607250101e-06
GC_6_1240 b_6 NI_6 NS_1240 0 -1.1766922742026087e-05
GC_6_1241 b_6 NI_6 NS_1241 0 -2.2685261424277725e-06
GC_6_1242 b_6 NI_6 NS_1242 0 -1.7028017088373762e-06
GC_6_1243 b_6 NI_6 NS_1243 0 -2.3846885058590163e-06
GC_6_1244 b_6 NI_6 NS_1244 0 -3.9900409387181535e-06
GC_6_1245 b_6 NI_6 NS_1245 0 -1.4877942972785012e-06
GC_6_1246 b_6 NI_6 NS_1246 0 -2.4193237709239337e-06
GC_6_1247 b_6 NI_6 NS_1247 0 -1.0718666974195810e-05
GC_6_1248 b_6 NI_6 NS_1248 0 -7.0858396828241823e-06
GC_6_1249 b_6 NI_6 NS_1249 0 -3.1913008936794725e-06
GC_6_1250 b_6 NI_6 NS_1250 0 -8.5705636285714992e-07
GC_6_1251 b_6 NI_6 NS_1251 0 -5.7484893235574218e-06
GC_6_1252 b_6 NI_6 NS_1252 0 -3.7009189415087604e-07
GC_6_1253 b_6 NI_6 NS_1253 0 -3.1247011179236963e-06
GC_6_1254 b_6 NI_6 NS_1254 0 -1.7467010566624070e-06
GC_6_1255 b_6 NI_6 NS_1255 0 -1.0620563759525155e-05
GC_6_1256 b_6 NI_6 NS_1256 0 3.3757026877594932e-06
GC_6_1257 b_6 NI_6 NS_1257 0 -3.6323502073644157e-06
GC_6_1258 b_6 NI_6 NS_1258 0 8.2990738611260243e-07
GC_6_1259 b_6 NI_6 NS_1259 0 -2.8726621383215847e-06
GC_6_1260 b_6 NI_6 NS_1260 0 3.9436371965494403e-06
GC_6_1261 b_6 NI_6 NS_1261 0 -4.3602282324877581e-06
GC_6_1262 b_6 NI_6 NS_1262 0 1.7215241685347608e-07
GC_6_1263 b_6 NI_6 NS_1263 0 -1.8596080451781374e-06
GC_6_1264 b_6 NI_6 NS_1264 0 7.2753449785330666e-06
GC_6_1265 b_6 NI_6 NS_1265 0 -1.5754115319638849e-06
GC_6_1266 b_6 NI_6 NS_1266 0 2.8117901487297631e-06
GC_6_1267 b_6 NI_6 NS_1267 0 9.3640963896643502e-07
GC_6_1268 b_6 NI_6 NS_1268 0 1.8342904809091011e-06
GC_6_1269 b_6 NI_6 NS_1269 0 -3.0126840328697078e-11
GC_6_1270 b_6 NI_6 NS_1270 0 -3.3795089032961796e-12
GC_6_1271 b_6 NI_6 NS_1271 0 -1.7324948658585524e-06
GC_6_1272 b_6 NI_6 NS_1272 0 2.1530116127260925e-06
GC_6_1273 b_6 NI_6 NS_1273 0 -3.2447816939980742e-07
GC_6_1274 b_6 NI_6 NS_1274 0 1.0585500720462542e-06
GC_6_1275 b_6 NI_6 NS_1275 0 1.4373499792284570e-07
GC_6_1276 b_6 NI_6 NS_1276 0 6.3907925419538792e-07
GC_6_1277 b_6 NI_6 NS_1277 0 -1.0432330340681828e-06
GC_6_1278 b_6 NI_6 NS_1278 0 1.2848488860883879e-06
GC_6_1279 b_6 NI_6 NS_1279 0 9.8805433356664043e-07
GC_6_1280 b_6 NI_6 NS_1280 0 1.8543072421426810e-06
GC_6_1281 b_6 NI_6 NS_1281 0 -1.5200215646202955e-09
GC_6_1282 b_6 NI_6 NS_1282 0 -7.6813243270803659e-10
GC_6_1283 b_6 NI_6 NS_1283 0 -4.6961262362619734e-07
GC_6_1284 b_6 NI_6 NS_1284 0 -2.3333645960305183e-08
GC_6_1285 b_6 NI_6 NS_1285 0 -3.1184768883712145e-07
GC_6_1286 b_6 NI_6 NS_1286 0 1.9127777368944800e-07
GC_6_1287 b_6 NI_6 NS_1287 0 -5.4919344556834409e-07
GC_6_1288 b_6 NI_6 NS_1288 0 1.5141538437307524e-07
GC_6_1289 b_6 NI_6 NS_1289 0 6.6185625258998342e-07
GC_6_1290 b_6 NI_6 NS_1290 0 8.3046390744418850e-07
GC_6_1291 b_6 NI_6 NS_1291 0 2.3283649306679413e-07
GC_6_1292 b_6 NI_6 NS_1292 0 7.0047503798867483e-07
GC_6_1293 b_6 NI_6 NS_1293 0 3.0951615143653210e-09
GC_6_1294 b_6 NI_6 NS_1294 0 -1.3231310667077663e-07
GC_6_1295 b_6 NI_6 NS_1295 0 -3.4727150870241052e-07
GC_6_1296 b_6 NI_6 NS_1296 0 2.9413059095663639e-07
GD_6_1 b_6 NI_6 NA_1 0 1.9211926466556270e-05
GD_6_2 b_6 NI_6 NA_2 0 3.5826268307878507e-06
GD_6_3 b_6 NI_6 NA_3 0 1.0511509584810319e-04
GD_6_4 b_6 NI_6 NA_4 0 2.2219274622720857e-05
GD_6_5 b_6 NI_6 NA_5 0 -4.9039972962224843e-03
GD_6_6 b_6 NI_6 NA_6 0 -1.1040269116042035e-02
GD_6_7 b_6 NI_6 NA_7 0 -1.1498071994794749e-03
GD_6_8 b_6 NI_6 NA_8 0 1.0577033559931812e-02
GD_6_9 b_6 NI_6 NA_9 0 1.5904542451315317e-05
GD_6_10 b_6 NI_6 NA_10 0 -3.7841718931773767e-07
GD_6_11 b_6 NI_6 NA_11 0 1.1430787472871246e-05
GD_6_12 b_6 NI_6 NA_12 0 -2.9989191181763534e-06
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 4.7631966946558960e-05
GC_7_2 b_7 NI_7 NS_2 0 7.4845515681842993e-12
GC_7_3 b_7 NI_7 NS_3 0 -1.8841447336015248e-11
GC_7_4 b_7 NI_7 NS_4 0 9.9252817843023913e-10
GC_7_5 b_7 NI_7 NS_5 0 -6.5468925148042918e-08
GC_7_6 b_7 NI_7 NS_6 0 2.4788334776608618e-07
GC_7_7 b_7 NI_7 NS_7 0 2.2310536449618617e-07
GC_7_8 b_7 NI_7 NS_8 0 4.0419326477214767e-07
GC_7_9 b_7 NI_7 NS_9 0 -1.7538227153262589e-07
GC_7_10 b_7 NI_7 NS_10 0 2.7605818803192090e-07
GC_7_11 b_7 NI_7 NS_11 0 7.2646978815622828e-07
GC_7_12 b_7 NI_7 NS_12 0 1.4718717698435661e-06
GC_7_13 b_7 NI_7 NS_13 0 1.0323109306589985e-06
GC_7_14 b_7 NI_7 NS_14 0 -4.2531103623850424e-07
GC_7_15 b_7 NI_7 NS_15 0 3.0287118581505716e-07
GC_7_16 b_7 NI_7 NS_16 0 9.1872026082369899e-07
GC_7_17 b_7 NI_7 NS_17 0 7.8010433989347938e-07
GC_7_18 b_7 NI_7 NS_18 0 -3.1455706660929672e-07
GC_7_19 b_7 NI_7 NS_19 0 4.3375164436419900e-06
GC_7_20 b_7 NI_7 NS_20 0 1.5052412278201375e-06
GC_7_21 b_7 NI_7 NS_21 0 -1.5165559971160282e-06
GC_7_22 b_7 NI_7 NS_22 0 -3.5706885286041766e-06
GC_7_23 b_7 NI_7 NS_23 0 2.4327995990603282e-07
GC_7_24 b_7 NI_7 NS_24 0 1.5795052291293579e-06
GC_7_25 b_7 NI_7 NS_25 0 3.1040272062315899e-06
GC_7_26 b_7 NI_7 NS_26 0 -4.6709509700649332e-06
GC_7_27 b_7 NI_7 NS_27 0 -7.4669659896911298e-07
GC_7_28 b_7 NI_7 NS_28 0 5.6972902333467199e-07
GC_7_29 b_7 NI_7 NS_29 0 5.7308733202838435e-06
GC_7_30 b_7 NI_7 NS_30 0 -5.7318870497247155e-06
GC_7_31 b_7 NI_7 NS_31 0 -3.3217238132258408e-06
GC_7_32 b_7 NI_7 NS_32 0 1.7569737156884520e-06
GC_7_33 b_7 NI_7 NS_33 0 8.8313630992013375e-07
GC_7_34 b_7 NI_7 NS_34 0 1.2588766400538333e-06
GC_7_35 b_7 NI_7 NS_35 0 1.6940415842696759e-06
GC_7_36 b_7 NI_7 NS_36 0 -4.0841762498991572e-06
GC_7_37 b_7 NI_7 NS_37 0 6.1060207350846576e-07
GC_7_38 b_7 NI_7 NS_38 0 2.1519047006854608e-07
GC_7_39 b_7 NI_7 NS_39 0 2.5345205669648764e-07
GC_7_40 b_7 NI_7 NS_40 0 -4.0636606604625441e-06
GC_7_41 b_7 NI_7 NS_41 0 -1.5617930065341380e-07
GC_7_42 b_7 NI_7 NS_42 0 1.7811620600145741e-07
GC_7_43 b_7 NI_7 NS_43 0 4.7913306474094295e-06
GC_7_44 b_7 NI_7 NS_44 0 -6.3202229633087762e-06
GC_7_45 b_7 NI_7 NS_45 0 -1.7962215414410845e-06
GC_7_46 b_7 NI_7 NS_46 0 -1.3136347779657275e-06
GC_7_47 b_7 NI_7 NS_47 0 1.4000599993834882e-06
GC_7_48 b_7 NI_7 NS_48 0 -1.1889560269279738e-06
GC_7_49 b_7 NI_7 NS_49 0 4.3422443417980876e-07
GC_7_50 b_7 NI_7 NS_50 0 -2.1045341782058328e-06
GC_7_51 b_7 NI_7 NS_51 0 -1.3395088127396419e-06
GC_7_52 b_7 NI_7 NS_52 0 -1.1872484490482143e-05
GC_7_53 b_7 NI_7 NS_53 0 -2.2432648860900503e-06
GC_7_54 b_7 NI_7 NS_54 0 -1.7314842309367918e-06
GC_7_55 b_7 NI_7 NS_55 0 -2.3524775701491194e-06
GC_7_56 b_7 NI_7 NS_56 0 -4.0390075982651929e-06
GC_7_57 b_7 NI_7 NS_57 0 -1.4499764003193982e-06
GC_7_58 b_7 NI_7 NS_58 0 -2.4370092964593722e-06
GC_7_59 b_7 NI_7 NS_59 0 -1.0683069533826621e-05
GC_7_60 b_7 NI_7 NS_60 0 -7.2200572148090000e-06
GC_7_61 b_7 NI_7 NS_61 0 -3.1781716401460233e-06
GC_7_62 b_7 NI_7 NS_62 0 -8.7729187697377620e-07
GC_7_63 b_7 NI_7 NS_63 0 -5.7541058597961405e-06
GC_7_64 b_7 NI_7 NS_64 0 -4.1607484423600735e-07
GC_7_65 b_7 NI_7 NS_65 0 -3.0997357383233849e-06
GC_7_66 b_7 NI_7 NS_66 0 -1.7555840722633963e-06
GC_7_67 b_7 NI_7 NS_67 0 -1.0627585100815261e-05
GC_7_68 b_7 NI_7 NS_68 0 3.2953774205070929e-06
GC_7_69 b_7 NI_7 NS_69 0 -3.6183712820320184e-06
GC_7_70 b_7 NI_7 NS_70 0 8.1870306375441761e-07
GC_7_71 b_7 NI_7 NS_71 0 -2.8814465509304798e-06
GC_7_72 b_7 NI_7 NS_72 0 3.9140066272928724e-06
GC_7_73 b_7 NI_7 NS_73 0 -4.3309334795739549e-06
GC_7_74 b_7 NI_7 NS_74 0 1.7127381880754197e-07
GC_7_75 b_7 NI_7 NS_75 0 -1.8671475615398519e-06
GC_7_76 b_7 NI_7 NS_76 0 7.2126071725172817e-06
GC_7_77 b_7 NI_7 NS_77 0 -1.5633432353133259e-06
GC_7_78 b_7 NI_7 NS_78 0 2.7935666271467218e-06
GC_7_79 b_7 NI_7 NS_79 0 9.2396491029579401e-07
GC_7_80 b_7 NI_7 NS_80 0 1.8140039662102593e-06
GC_7_81 b_7 NI_7 NS_81 0 -3.0213685789724924e-11
GC_7_82 b_7 NI_7 NS_82 0 -3.9931475956168604e-12
GC_7_83 b_7 NI_7 NS_83 0 -1.7134382599510951e-06
GC_7_84 b_7 NI_7 NS_84 0 2.1404403455519030e-06
GC_7_85 b_7 NI_7 NS_85 0 -3.2436353778035551e-07
GC_7_86 b_7 NI_7 NS_86 0 1.0487453848481990e-06
GC_7_87 b_7 NI_7 NS_87 0 1.4400256463229223e-07
GC_7_88 b_7 NI_7 NS_88 0 6.2111542664577477e-07
GC_7_89 b_7 NI_7 NS_89 0 -1.0462324686081481e-06
GC_7_90 b_7 NI_7 NS_90 0 1.2710919853041630e-06
GC_7_91 b_7 NI_7 NS_91 0 9.7965191833771816e-07
GC_7_92 b_7 NI_7 NS_92 0 1.8189635595557154e-06
GC_7_93 b_7 NI_7 NS_93 0 -1.5165334427340345e-09
GC_7_94 b_7 NI_7 NS_94 0 -7.8078233781151703e-10
GC_7_95 b_7 NI_7 NS_95 0 -4.8470522465135096e-07
GC_7_96 b_7 NI_7 NS_96 0 -2.7510766463683923e-08
GC_7_97 b_7 NI_7 NS_97 0 -3.1050735924549243e-07
GC_7_98 b_7 NI_7 NS_98 0 1.7476029169890767e-07
GC_7_99 b_7 NI_7 NS_99 0 -5.5079987921206176e-07
GC_7_100 b_7 NI_7 NS_100 0 1.5190555443158876e-07
GC_7_101 b_7 NI_7 NS_101 0 6.6424926825704255e-07
GC_7_102 b_7 NI_7 NS_102 0 8.1076600609659581e-07
GC_7_103 b_7 NI_7 NS_103 0 2.1776781220687560e-07
GC_7_104 b_7 NI_7 NS_104 0 6.9571010181021462e-07
GC_7_105 b_7 NI_7 NS_105 0 1.0940213103610424e-08
GC_7_106 b_7 NI_7 NS_106 0 -1.3810919825212781e-07
GC_7_107 b_7 NI_7 NS_107 0 -3.4771245244287973e-07
GC_7_108 b_7 NI_7 NS_108 0 2.9453641711061325e-07
GC_7_109 b_7 NI_7 NS_109 0 -8.9925137525303784e-05
GC_7_110 b_7 NI_7 NS_110 0 3.3207015404536118e-12
GC_7_111 b_7 NI_7 NS_111 0 -4.3128817098512642e-11
GC_7_112 b_7 NI_7 NS_112 0 3.0190792527993700e-10
GC_7_113 b_7 NI_7 NS_113 0 -1.5707266998279248e-06
GC_7_114 b_7 NI_7 NS_114 0 -1.5515332936728513e-06
GC_7_115 b_7 NI_7 NS_115 0 9.5011122046084813e-07
GC_7_116 b_7 NI_7 NS_116 0 7.0859746109594679e-07
GC_7_117 b_7 NI_7 NS_117 0 -2.7109495454425127e-06
GC_7_118 b_7 NI_7 NS_118 0 3.0183037772233092e-06
GC_7_119 b_7 NI_7 NS_119 0 -3.0631390801589227e-06
GC_7_120 b_7 NI_7 NS_120 0 -2.5681861474502426e-06
GC_7_121 b_7 NI_7 NS_121 0 1.4917516300875810e-06
GC_7_122 b_7 NI_7 NS_122 0 8.4631729107066178e-08
GC_7_123 b_7 NI_7 NS_123 0 -1.6569922646023009e-06
GC_7_124 b_7 NI_7 NS_124 0 1.7806155863648009e-06
GC_7_125 b_7 NI_7 NS_125 0 8.7351325963540654e-07
GC_7_126 b_7 NI_7 NS_126 0 4.1342407457068660e-06
GC_7_127 b_7 NI_7 NS_127 0 -4.3581708274511181e-06
GC_7_128 b_7 NI_7 NS_128 0 -1.9912099995526725e-06
GC_7_129 b_7 NI_7 NS_129 0 2.4348194737448496e-06
GC_7_130 b_7 NI_7 NS_130 0 -1.8849490996909452e-06
GC_7_131 b_7 NI_7 NS_131 0 -1.1509987502288401e-06
GC_7_132 b_7 NI_7 NS_132 0 3.2760392892900912e-06
GC_7_133 b_7 NI_7 NS_133 0 -8.2168044855203814e-06
GC_7_134 b_7 NI_7 NS_134 0 1.1138771452891388e-05
GC_7_135 b_7 NI_7 NS_135 0 1.2480511957103064e-06
GC_7_136 b_7 NI_7 NS_136 0 -1.6722623696503041e-06
GC_7_137 b_7 NI_7 NS_137 0 9.8795690249265224e-06
GC_7_138 b_7 NI_7 NS_138 0 1.7077759120098524e-05
GC_7_139 b_7 NI_7 NS_139 0 -6.7063777910880669e-07
GC_7_140 b_7 NI_7 NS_140 0 -4.6941551841482848e-07
GC_7_141 b_7 NI_7 NS_141 0 4.0634682689216991e-07
GC_7_142 b_7 NI_7 NS_142 0 -1.3870420170537907e-06
GC_7_143 b_7 NI_7 NS_143 0 6.8974674890354218e-06
GC_7_144 b_7 NI_7 NS_144 0 -1.5805647125497159e-07
GC_7_145 b_7 NI_7 NS_145 0 7.1137371993578584e-07
GC_7_146 b_7 NI_7 NS_146 0 3.0107754439086927e-06
GC_7_147 b_7 NI_7 NS_147 0 5.0116847832179911e-07
GC_7_148 b_7 NI_7 NS_148 0 2.8944302541545382e-06
GC_7_149 b_7 NI_7 NS_149 0 1.1551642732096831e-06
GC_7_150 b_7 NI_7 NS_150 0 -1.4201311040104945e-06
GC_7_151 b_7 NI_7 NS_151 0 9.2615647686842507e-06
GC_7_152 b_7 NI_7 NS_152 0 5.1119617725432236e-06
GC_7_153 b_7 NI_7 NS_153 0 5.5744833193432640e-07
GC_7_154 b_7 NI_7 NS_154 0 1.1628096368159025e-06
GC_7_155 b_7 NI_7 NS_155 0 4.5595150036943773e-08
GC_7_156 b_7 NI_7 NS_156 0 4.6106139588891227e-07
GC_7_157 b_7 NI_7 NS_157 0 1.2710005409115873e-06
GC_7_158 b_7 NI_7 NS_158 0 -8.4419934977842505e-07
GC_7_159 b_7 NI_7 NS_159 0 9.0349148585355095e-06
GC_7_160 b_7 NI_7 NS_160 0 7.0641231338948312e-07
GC_7_161 b_7 NI_7 NS_161 0 8.3856109355462797e-07
GC_7_162 b_7 NI_7 NS_162 0 1.4664546274636352e-06
GC_7_163 b_7 NI_7 NS_163 0 1.0338744731259049e-06
GC_7_164 b_7 NI_7 NS_164 0 6.2486116777460570e-07
GC_7_165 b_7 NI_7 NS_165 0 1.3512302282790773e-06
GC_7_166 b_7 NI_7 NS_166 0 -9.4050027863084281e-07
GC_7_167 b_7 NI_7 NS_167 0 7.9401787568099950e-06
GC_7_168 b_7 NI_7 NS_168 0 -2.0574336692606511e-06
GC_7_169 b_7 NI_7 NS_169 0 1.1774868207139395e-06
GC_7_170 b_7 NI_7 NS_170 0 1.5557215510933050e-06
GC_7_171 b_7 NI_7 NS_171 0 1.6144416346318521e-06
GC_7_172 b_7 NI_7 NS_172 0 -2.1447334196261452e-07
GC_7_173 b_7 NI_7 NS_173 0 1.3152795445498034e-06
GC_7_174 b_7 NI_7 NS_174 0 -9.8120406898038024e-07
GC_7_175 b_7 NI_7 NS_175 0 5.8097268139479410e-06
GC_7_176 b_7 NI_7 NS_176 0 -3.8284853859855166e-06
GC_7_177 b_7 NI_7 NS_177 0 1.8107763242422285e-06
GC_7_178 b_7 NI_7 NS_178 0 1.4375766988104311e-06
GC_7_179 b_7 NI_7 NS_179 0 1.1299062145066183e-06
GC_7_180 b_7 NI_7 NS_180 0 -1.3882895137721936e-06
GC_7_181 b_7 NI_7 NS_181 0 1.4160170134936263e-06
GC_7_182 b_7 NI_7 NS_182 0 -1.0986919513817648e-06
GC_7_183 b_7 NI_7 NS_183 0 2.9955763893206041e-06
GC_7_184 b_7 NI_7 NS_184 0 -4.1669843017254318e-06
GC_7_185 b_7 NI_7 NS_185 0 2.2265255120263448e-06
GC_7_186 b_7 NI_7 NS_186 0 3.1296203494060254e-07
GC_7_187 b_7 NI_7 NS_187 0 -3.0639562821957853e-07
GC_7_188 b_7 NI_7 NS_188 0 -1.1888571372685726e-06
GC_7_189 b_7 NI_7 NS_189 0 2.5432671247243125e-11
GC_7_190 b_7 NI_7 NS_190 0 -4.1105506091219085e-11
GC_7_191 b_7 NI_7 NS_191 0 8.0940173594058295e-07
GC_7_192 b_7 NI_7 NS_192 0 -1.5691564293716276e-06
GC_7_193 b_7 NI_7 NS_193 0 1.2651493716373758e-06
GC_7_194 b_7 NI_7 NS_194 0 2.2094680681391598e-07
GC_7_195 b_7 NI_7 NS_195 0 1.6270285684478959e-07
GC_7_196 b_7 NI_7 NS_196 0 -5.4918374177207124e-07
GC_7_197 b_7 NI_7 NS_197 0 5.5453372486212388e-07
GC_7_198 b_7 NI_7 NS_198 0 -8.6155709493891055e-07
GC_7_199 b_7 NI_7 NS_199 0 1.3101220080844703e-06
GC_7_200 b_7 NI_7 NS_200 0 -2.0776519945388766e-06
GC_7_201 b_7 NI_7 NS_201 0 4.9004256053118770e-10
GC_7_202 b_7 NI_7 NS_202 0 -1.2286548743533631e-09
GC_7_203 b_7 NI_7 NS_203 0 5.5269533022176542e-07
GC_7_204 b_7 NI_7 NS_204 0 -8.6347619060784736e-07
GC_7_205 b_7 NI_7 NS_205 0 7.1657187060196998e-07
GC_7_206 b_7 NI_7 NS_206 0 -9.5174159257651988e-07
GC_7_207 b_7 NI_7 NS_207 0 9.1484167548771759e-08
GC_7_208 b_7 NI_7 NS_208 0 4.9336905657722897e-08
GC_7_209 b_7 NI_7 NS_209 0 1.3737752544353467e-06
GC_7_210 b_7 NI_7 NS_210 0 -1.2452351870806522e-06
GC_7_211 b_7 NI_7 NS_211 0 1.6627819059840762e-06
GC_7_212 b_7 NI_7 NS_212 0 -3.1746238572373524e-07
GC_7_213 b_7 NI_7 NS_213 0 -2.3880345920376409e-07
GC_7_214 b_7 NI_7 NS_214 0 -7.4466902694736191e-07
GC_7_215 b_7 NI_7 NS_215 0 7.3884951276105620e-07
GC_7_216 b_7 NI_7 NS_216 0 2.9287388822209100e-07
GC_7_217 b_7 NI_7 NS_217 0 -2.8450109010455024e-05
GC_7_218 b_7 NI_7 NS_218 0 -9.0137019991392671e-13
GC_7_219 b_7 NI_7 NS_219 0 -2.3532354983913329e-10
GC_7_220 b_7 NI_7 NS_220 0 1.0469898403828317e-08
GC_7_221 b_7 NI_7 NS_221 0 7.2361377555210130e-07
GC_7_222 b_7 NI_7 NS_222 0 1.1682418614927328e-07
GC_7_223 b_7 NI_7 NS_223 0 3.2158789041487332e-06
GC_7_224 b_7 NI_7 NS_224 0 -1.3848969882192265e-06
GC_7_225 b_7 NI_7 NS_225 0 -2.7214326435008593e-06
GC_7_226 b_7 NI_7 NS_226 0 -2.8594433451887567e-06
GC_7_227 b_7 NI_7 NS_227 0 5.0260142923809230e-06
GC_7_228 b_7 NI_7 NS_228 0 -5.8504264544669851e-07
GC_7_229 b_7 NI_7 NS_229 0 -7.0572386582488509e-06
GC_7_230 b_7 NI_7 NS_230 0 -8.2657447345377763e-06
GC_7_231 b_7 NI_7 NS_231 0 8.4163795005262638e-08
GC_7_232 b_7 NI_7 NS_232 0 -1.5979811135919314e-06
GC_7_233 b_7 NI_7 NS_233 0 -6.1458564384684910e-06
GC_7_234 b_7 NI_7 NS_234 0 1.8452524766470391e-06
GC_7_235 b_7 NI_7 NS_235 0 5.3927004264957291e-06
GC_7_236 b_7 NI_7 NS_236 0 -5.9846569934136712e-06
GC_7_237 b_7 NI_7 NS_237 0 -1.7353900743671204e-05
GC_7_238 b_7 NI_7 NS_238 0 4.6493306406104387e-06
GC_7_239 b_7 NI_7 NS_239 0 -1.1603762174071007e-06
GC_7_240 b_7 NI_7 NS_240 0 7.0453709479424970e-06
GC_7_241 b_7 NI_7 NS_241 0 -7.4845948325220003e-06
GC_7_242 b_7 NI_7 NS_242 0 -4.7597379235542805e-06
GC_7_243 b_7 NI_7 NS_243 0 -3.4153040762122801e-06
GC_7_244 b_7 NI_7 NS_244 0 8.0176902728308036e-06
GC_7_245 b_7 NI_7 NS_245 0 -2.5103464023047247e-06
GC_7_246 b_7 NI_7 NS_246 0 -4.9392785167785019e-06
GC_7_247 b_7 NI_7 NS_247 0 -3.8632871770144922e-06
GC_7_248 b_7 NI_7 NS_248 0 1.1456367727594994e-05
GC_7_249 b_7 NI_7 NS_249 0 -1.7994811476379881e-07
GC_7_250 b_7 NI_7 NS_250 0 7.1537422215474852e-06
GC_7_251 b_7 NI_7 NS_251 0 -4.3372987496911446e-06
GC_7_252 b_7 NI_7 NS_252 0 1.1467067961473793e-06
GC_7_253 b_7 NI_7 NS_253 0 -6.7842101007949110e-07
GC_7_254 b_7 NI_7 NS_254 0 7.9730691507698692e-06
GC_7_255 b_7 NI_7 NS_255 0 -1.2189492604492117e-06
GC_7_256 b_7 NI_7 NS_256 0 2.1994255094585245e-06
GC_7_257 b_7 NI_7 NS_257 0 -2.4670330842175054e-06
GC_7_258 b_7 NI_7 NS_258 0 8.1096126488037533e-06
GC_7_259 b_7 NI_7 NS_259 0 -3.9818466661294583e-07
GC_7_260 b_7 NI_7 NS_260 0 9.3212490244348546e-06
GC_7_261 b_7 NI_7 NS_261 0 -9.4389218110021648e-07
GC_7_262 b_7 NI_7 NS_262 0 8.7939545351285855e-06
GC_7_263 b_7 NI_7 NS_263 0 -1.3825917461186113e-06
GC_7_264 b_7 NI_7 NS_264 0 3.8436288294467254e-06
GC_7_265 b_7 NI_7 NS_265 0 8.7890300118402039e-07
GC_7_266 b_7 NI_7 NS_266 0 1.1882942069115950e-05
GC_7_267 b_7 NI_7 NS_267 0 1.7118689258311150e-05
GC_7_268 b_7 NI_7 NS_268 0 1.6747351739254846e-05
GC_7_269 b_7 NI_7 NS_269 0 4.6531239620865810e-06
GC_7_270 b_7 NI_7 NS_270 0 7.7083933880062519e-06
GC_7_271 b_7 NI_7 NS_271 0 9.7617617756947417e-06
GC_7_272 b_7 NI_7 NS_272 0 3.8979688816289244e-06
GC_7_273 b_7 NI_7 NS_273 0 6.3871972959350766e-06
GC_7_274 b_7 NI_7 NS_274 0 1.0670549943454131e-05
GC_7_275 b_7 NI_7 NS_275 0 3.1859678126256064e-05
GC_7_276 b_7 NI_7 NS_276 0 -5.6286006589521356e-06
GC_7_277 b_7 NI_7 NS_277 0 7.7729849699531212e-06
GC_7_278 b_7 NI_7 NS_278 0 3.3978521648350320e-06
GC_7_279 b_7 NI_7 NS_279 0 1.1412307183718587e-05
GC_7_280 b_7 NI_7 NS_280 0 -9.8828256412099411e-06
GC_7_281 b_7 NI_7 NS_281 0 1.0308208970263038e-05
GC_7_282 b_7 NI_7 NS_282 0 6.2712889959454467e-06
GC_7_283 b_7 NI_7 NS_283 0 1.5926514842468387e-05
GC_7_284 b_7 NI_7 NS_284 0 -2.9763092896633639e-05
GC_7_285 b_7 NI_7 NS_285 0 7.6989670181538355e-06
GC_7_286 b_7 NI_7 NS_286 0 -2.8503570682419964e-06
GC_7_287 b_7 NI_7 NS_287 0 -3.4066363400809783e-06
GC_7_288 b_7 NI_7 NS_288 0 -1.5683575741775546e-05
GC_7_289 b_7 NI_7 NS_289 0 1.1265212055601548e-05
GC_7_290 b_7 NI_7 NS_290 0 -1.7001882135937927e-06
GC_7_291 b_7 NI_7 NS_291 0 -1.2934679513111400e-05
GC_7_292 b_7 NI_7 NS_292 0 -2.4095960897216839e-05
GC_7_293 b_7 NI_7 NS_293 0 -4.1482501424851214e-07
GC_7_294 b_7 NI_7 NS_294 0 -6.3721083492295655e-06
GC_7_295 b_7 NI_7 NS_295 0 -9.4862697462526194e-06
GC_7_296 b_7 NI_7 NS_296 0 -2.3404463473477483e-06
GC_7_297 b_7 NI_7 NS_297 0 9.7943009146926326e-11
GC_7_298 b_7 NI_7 NS_298 0 5.4145733933964428e-11
GC_7_299 b_7 NI_7 NS_299 0 1.1788424826391243e-06
GC_7_300 b_7 NI_7 NS_300 0 -4.6057062340473968e-06
GC_7_301 b_7 NI_7 NS_301 0 -1.4797996487510218e-06
GC_7_302 b_7 NI_7 NS_302 0 -1.2848527597536336e-06
GC_7_303 b_7 NI_7 NS_303 0 -4.9236175031598049e-06
GC_7_304 b_7 NI_7 NS_304 0 -8.7275585094081344e-07
GC_7_305 b_7 NI_7 NS_305 0 -1.3800578692018385e-06
GC_7_306 b_7 NI_7 NS_306 0 -2.8436550596928210e-06
GC_7_307 b_7 NI_7 NS_307 0 -1.0040390018300259e-05
GC_7_308 b_7 NI_7 NS_308 0 -3.6858172576700502e-06
GC_7_309 b_7 NI_7 NS_309 0 6.6581509786374768e-09
GC_7_310 b_7 NI_7 NS_310 0 5.7685224972499398e-09
GC_7_311 b_7 NI_7 NS_311 0 1.3973574957490061e-06
GC_7_312 b_7 NI_7 NS_312 0 6.7929616614619743e-07
GC_7_313 b_7 NI_7 NS_313 0 -1.7307673991845331e-06
GC_7_314 b_7 NI_7 NS_314 0 3.1503399720393280e-06
GC_7_315 b_7 NI_7 NS_315 0 -9.2380473746603920e-07
GC_7_316 b_7 NI_7 NS_316 0 7.7445358092014356e-07
GC_7_317 b_7 NI_7 NS_317 0 -7.9050294315926557e-06
GC_7_318 b_7 NI_7 NS_318 0 8.2698605361166494e-07
GC_7_319 b_7 NI_7 NS_319 0 -2.4152010232526735e-06
GC_7_320 b_7 NI_7 NS_320 0 2.0790177153280299e-06
GC_7_321 b_7 NI_7 NS_321 0 -2.1277774428300464e-06
GC_7_322 b_7 NI_7 NS_322 0 2.1503900805953420e-06
GC_7_323 b_7 NI_7 NS_323 0 1.1274193112787230e-06
GC_7_324 b_7 NI_7 NS_324 0 2.8111017592281511e-06
GC_7_325 b_7 NI_7 NS_325 0 -1.4436373535033298e-04
GC_7_326 b_7 NI_7 NS_326 0 3.3291387303585096e-11
GC_7_327 b_7 NI_7 NS_327 0 3.9882099425946800e-11
GC_7_328 b_7 NI_7 NS_328 0 9.0903672101921779e-10
GC_7_329 b_7 NI_7 NS_329 0 -2.1100782333540289e-06
GC_7_330 b_7 NI_7 NS_330 0 -1.6555674177524564e-06
GC_7_331 b_7 NI_7 NS_331 0 1.8947205468173026e-06
GC_7_332 b_7 NI_7 NS_332 0 3.8512917976862835e-06
GC_7_333 b_7 NI_7 NS_333 0 3.3113005804393602e-06
GC_7_334 b_7 NI_7 NS_334 0 4.9314150887762951e-06
GC_7_335 b_7 NI_7 NS_335 0 5.8708136782200842e-06
GC_7_336 b_7 NI_7 NS_336 0 -9.1115745743130765e-06
GC_7_337 b_7 NI_7 NS_337 0 -2.5609916430641102e-06
GC_7_338 b_7 NI_7 NS_338 0 -1.3919625909142548e-05
GC_7_339 b_7 NI_7 NS_339 0 -3.5429293493742383e-06
GC_7_340 b_7 NI_7 NS_340 0 2.1898054511600127e-06
GC_7_341 b_7 NI_7 NS_341 0 3.6501936456946169e-06
GC_7_342 b_7 NI_7 NS_342 0 1.2869481938549338e-06
GC_7_343 b_7 NI_7 NS_343 0 8.0000493802760078e-06
GC_7_344 b_7 NI_7 NS_344 0 -3.9897559259689219e-05
GC_7_345 b_7 NI_7 NS_345 0 -4.4313711733608574e-05
GC_7_346 b_7 NI_7 NS_346 0 -9.3697111382649157e-07
GC_7_347 b_7 NI_7 NS_347 0 -1.4827741601983220e-05
GC_7_348 b_7 NI_7 NS_348 0 -8.5761184048024682e-06
GC_7_349 b_7 NI_7 NS_349 0 -7.2939514799192899e-05
GC_7_350 b_7 NI_7 NS_350 0 7.5520238143228006e-05
GC_7_351 b_7 NI_7 NS_351 0 4.6289617882119877e-06
GC_7_352 b_7 NI_7 NS_352 0 1.3120054226334590e-05
GC_7_353 b_7 NI_7 NS_353 0 6.2840275979586218e-05
GC_7_354 b_7 NI_7 NS_354 0 1.2319963875398379e-04
GC_7_355 b_7 NI_7 NS_355 0 3.6327008844696044e-07
GC_7_356 b_7 NI_7 NS_356 0 -3.7019876311510890e-05
GC_7_357 b_7 NI_7 NS_357 0 1.6508676241033001e-05
GC_7_358 b_7 NI_7 NS_358 0 3.9672167862995570e-06
GC_7_359 b_7 NI_7 NS_359 0 2.4447788536671013e-05
GC_7_360 b_7 NI_7 NS_360 0 -3.0457955770084245e-05
GC_7_361 b_7 NI_7 NS_361 0 -8.8967721333999483e-06
GC_7_362 b_7 NI_7 NS_362 0 -2.3402098735877741e-06
GC_7_363 b_7 NI_7 NS_363 0 -8.8832850311499966e-06
GC_7_364 b_7 NI_7 NS_364 0 2.5237311700210069e-05
GC_7_365 b_7 NI_7 NS_365 0 5.8267217080779025e-06
GC_7_366 b_7 NI_7 NS_366 0 8.4670740135772346e-06
GC_7_367 b_7 NI_7 NS_367 0 5.6328294959376077e-05
GC_7_368 b_7 NI_7 NS_368 0 2.4970035889554806e-05
GC_7_369 b_7 NI_7 NS_369 0 3.5271362125614106e-06
GC_7_370 b_7 NI_7 NS_370 0 -1.1687102201658606e-05
GC_7_371 b_7 NI_7 NS_371 0 -4.0893620230356692e-07
GC_7_372 b_7 NI_7 NS_372 0 -1.3155525017791929e-06
GC_7_373 b_7 NI_7 NS_373 0 6.8059515917161994e-06
GC_7_374 b_7 NI_7 NS_374 0 3.0643177200443256e-06
GC_7_375 b_7 NI_7 NS_375 0 4.1947345442178175e-05
GC_7_376 b_7 NI_7 NS_376 0 -1.7198851167711414e-05
GC_7_377 b_7 NI_7 NS_377 0 -2.5587325623490220e-06
GC_7_378 b_7 NI_7 NS_378 0 -7.0969114422461084e-06
GC_7_379 b_7 NI_7 NS_379 0 -3.0311216968808503e-06
GC_7_380 b_7 NI_7 NS_380 0 1.7555079664938645e-06
GC_7_381 b_7 NI_7 NS_381 0 9.5694253140783602e-06
GC_7_382 b_7 NI_7 NS_382 0 2.9161001707619077e-06
GC_7_383 b_7 NI_7 NS_383 0 2.2975733315351055e-05
GC_7_384 b_7 NI_7 NS_384 0 -3.1187552552219614e-05
GC_7_385 b_7 NI_7 NS_385 0 -5.6937409793793131e-06
GC_7_386 b_7 NI_7 NS_386 0 -3.6756843403623617e-06
GC_7_387 b_7 NI_7 NS_387 0 -5.6140290206715984e-07
GC_7_388 b_7 NI_7 NS_388 0 5.0284604168137977e-06
GC_7_389 b_7 NI_7 NS_389 0 1.2292599722114543e-05
GC_7_390 b_7 NI_7 NS_390 0 2.0420805557735008e-07
GC_7_391 b_7 NI_7 NS_391 0 1.9184400593438847e-06
GC_7_392 b_7 NI_7 NS_392 0 -3.1503455546282967e-05
GC_7_393 b_7 NI_7 NS_393 0 -6.7231151650604399e-06
GC_7_394 b_7 NI_7 NS_394 0 9.4627462512202167e-07
GC_7_395 b_7 NI_7 NS_395 0 4.5912590890620542e-06
GC_7_396 b_7 NI_7 NS_396 0 3.8667896211982772e-06
GC_7_397 b_7 NI_7 NS_397 0 1.4096550353693015e-05
GC_7_398 b_7 NI_7 NS_398 0 -6.0052051202605487e-06
GC_7_399 b_7 NI_7 NS_399 0 -1.3991415688155794e-05
GC_7_400 b_7 NI_7 NS_400 0 -1.8834210417608704e-05
GC_7_401 b_7 NI_7 NS_401 0 -2.5005394032594012e-06
GC_7_402 b_7 NI_7 NS_402 0 5.3959386522720470e-06
GC_7_403 b_7 NI_7 NS_403 0 4.6402339650707107e-06
GC_7_404 b_7 NI_7 NS_404 0 -2.0953515482236344e-06
GC_7_405 b_7 NI_7 NS_405 0 -1.4466712168479286e-11
GC_7_406 b_7 NI_7 NS_406 0 3.9863998002107105e-12
GC_7_407 b_7 NI_7 NS_407 0 5.2050436760924432e-06
GC_7_408 b_7 NI_7 NS_408 0 -1.1255637506104323e-05
GC_7_409 b_7 NI_7 NS_409 0 -2.6207805365397699e-07
GC_7_410 b_7 NI_7 NS_410 0 2.9240741721436538e-06
GC_7_411 b_7 NI_7 NS_411 0 2.6491364981996882e-06
GC_7_412 b_7 NI_7 NS_412 0 -1.6106156442507593e-06
GC_7_413 b_7 NI_7 NS_413 0 2.4311195868717799e-06
GC_7_414 b_7 NI_7 NS_414 0 -9.4257144225246813e-06
GC_7_415 b_7 NI_7 NS_415 0 -9.9191023744807521e-06
GC_7_416 b_7 NI_7 NS_416 0 -3.6952523716666837e-06
GC_7_417 b_7 NI_7 NS_417 0 3.1959673367626157e-10
GC_7_418 b_7 NI_7 NS_418 0 2.6406121421726251e-10
GC_7_419 b_7 NI_7 NS_419 0 -8.5810808272950858e-06
GC_7_420 b_7 NI_7 NS_420 0 -5.7196666115889418e-06
GC_7_421 b_7 NI_7 NS_421 0 2.2759088243607779e-06
GC_7_422 b_7 NI_7 NS_422 0 -6.4442872801461139e-06
GC_7_423 b_7 NI_7 NS_423 0 -3.0692758063640964e-06
GC_7_424 b_7 NI_7 NS_424 0 -1.3767141828140062e-07
GC_7_425 b_7 NI_7 NS_425 0 -7.9175943952123413e-06
GC_7_426 b_7 NI_7 NS_426 0 4.8805512885631643e-07
GC_7_427 b_7 NI_7 NS_427 0 3.0157381949114486e-06
GC_7_428 b_7 NI_7 NS_428 0 2.8670369036843247e-06
GC_7_429 b_7 NI_7 NS_429 0 1.2342980748281233e-06
GC_7_430 b_7 NI_7 NS_430 0 -3.9109811129983600e-06
GC_7_431 b_7 NI_7 NS_431 0 -4.8692444772841975e-06
GC_7_432 b_7 NI_7 NS_432 0 -3.9053550416086599e-06
GC_7_433 b_7 NI_7 NS_433 0 1.4425741233361886e-03
GC_7_434 b_7 NI_7 NS_434 0 -3.5904351747023481e-09
GC_7_435 b_7 NI_7 NS_435 0 -4.7342043128233263e-08
GC_7_436 b_7 NI_7 NS_436 0 -3.5032371832117494e-06
GC_7_437 b_7 NI_7 NS_437 0 -3.6675402607323326e-04
GC_7_438 b_7 NI_7 NS_438 0 1.3531649500526485e-04
GC_7_439 b_7 NI_7 NS_439 0 1.1270906314471225e-03
GC_7_440 b_7 NI_7 NS_440 0 1.9466317752188139e-03
GC_7_441 b_7 NI_7 NS_441 0 -5.2133213260550092e-05
GC_7_442 b_7 NI_7 NS_442 0 -3.4959654435807886e-03
GC_7_443 b_7 NI_7 NS_443 0 -1.5728294785791698e-03
GC_7_444 b_7 NI_7 NS_444 0 5.0835060984192309e-03
GC_7_445 b_7 NI_7 NS_445 0 4.2660496763269598e-03
GC_7_446 b_7 NI_7 NS_446 0 -4.9897929070204586e-03
GC_7_447 b_7 NI_7 NS_447 0 -1.0071498745518805e-03
GC_7_448 b_7 NI_7 NS_448 0 5.5941858275035589e-04
GC_7_449 b_7 NI_7 NS_449 0 -2.0791293775648707e-03
GC_7_450 b_7 NI_7 NS_450 0 -1.8719560941385857e-03
GC_7_451 b_7 NI_7 NS_451 0 3.6235024008862845e-03
GC_7_452 b_7 NI_7 NS_452 0 1.1644121681272544e-02
GC_7_453 b_7 NI_7 NS_453 0 -8.7672702084257549e-04
GC_7_454 b_7 NI_7 NS_454 0 -1.4855229418282824e-02
GC_7_455 b_7 NI_7 NS_455 0 -8.1250075384110953e-03
GC_7_456 b_7 NI_7 NS_456 0 1.9028461816925867e-03
GC_7_457 b_7 NI_7 NS_457 0 1.1255574803279458e-02
GC_7_458 b_7 NI_7 NS_458 0 -1.8013331256158493e-03
GC_7_459 b_7 NI_7 NS_459 0 -7.5649379463101586e-03
GC_7_460 b_7 NI_7 NS_460 0 -1.6931181032836427e-03
GC_7_461 b_7 NI_7 NS_461 0 1.5263484753164743e-02
GC_7_462 b_7 NI_7 NS_462 0 5.3089269962556156e-03
GC_7_463 b_7 NI_7 NS_463 0 -1.3074208628142452e-02
GC_7_464 b_7 NI_7 NS_464 0 -5.4740974161817165e-03
GC_7_465 b_7 NI_7 NS_465 0 -6.6401727829744819e-03
GC_7_466 b_7 NI_7 NS_466 0 3.4469264645533054e-03
GC_7_467 b_7 NI_7 NS_467 0 6.3571562313446449e-03
GC_7_468 b_7 NI_7 NS_468 0 -1.8769366072078938e-03
GC_7_469 b_7 NI_7 NS_469 0 -5.4767784441415923e-03
GC_7_470 b_7 NI_7 NS_470 0 2.1761634539401546e-03
GC_7_471 b_7 NI_7 NS_471 0 5.3904708368407890e-03
GC_7_472 b_7 NI_7 NS_472 0 -2.6291409730219281e-03
GC_7_473 b_7 NI_7 NS_473 0 -6.3068613300950194e-03
GC_7_474 b_7 NI_7 NS_474 0 -4.8944546422459130e-04
GC_7_475 b_7 NI_7 NS_475 0 7.6383029102315243e-03
GC_7_476 b_7 NI_7 NS_476 0 3.6283278334159554e-03
GC_7_477 b_7 NI_7 NS_477 0 -5.8333235006031350e-03
GC_7_478 b_7 NI_7 NS_478 0 -3.4684301765323076e-03
GC_7_479 b_7 NI_7 NS_479 0 2.9592188619419760e-04
GC_7_480 b_7 NI_7 NS_480 0 5.5702924793212384e-04
GC_7_481 b_7 NI_7 NS_481 0 -4.9284028867596103e-03
GC_7_482 b_7 NI_7 NS_482 0 8.8733927007922484e-04
GC_7_483 b_7 NI_7 NS_483 0 6.2016450885667542e-03
GC_7_484 b_7 NI_7 NS_484 0 6.8248096800240952e-04
GC_7_485 b_7 NI_7 NS_485 0 -5.3226827419088144e-03
GC_7_486 b_7 NI_7 NS_486 0 -4.8918921539239956e-04
GC_7_487 b_7 NI_7 NS_487 0 1.5482735936976748e-03
GC_7_488 b_7 NI_7 NS_488 0 -4.6609097843995798e-05
GC_7_489 b_7 NI_7 NS_489 0 -6.0242735565756798e-03
GC_7_490 b_7 NI_7 NS_490 0 1.9161516125141217e-03
GC_7_491 b_7 NI_7 NS_491 0 6.2494033703015947e-03
GC_7_492 b_7 NI_7 NS_492 0 2.0850497458923365e-04
GC_7_493 b_7 NI_7 NS_493 0 -5.0636589476606986e-03
GC_7_494 b_7 NI_7 NS_494 0 1.6954532766883816e-03
GC_7_495 b_7 NI_7 NS_495 0 2.4806588151512817e-03
GC_7_496 b_7 NI_7 NS_496 0 -9.6015728238761991e-04
GC_7_497 b_7 NI_7 NS_497 0 -6.5381320997607729e-03
GC_7_498 b_7 NI_7 NS_498 0 3.8750074877559469e-03
GC_7_499 b_7 NI_7 NS_499 0 7.4722547471553049e-03
GC_7_500 b_7 NI_7 NS_500 0 -1.0944729982738822e-03
GC_7_501 b_7 NI_7 NS_501 0 -3.9943218502332513e-03
GC_7_502 b_7 NI_7 NS_502 0 4.0357752359329174e-03
GC_7_503 b_7 NI_7 NS_503 0 2.8552014001052097e-03
GC_7_504 b_7 NI_7 NS_504 0 -3.0472625143398886e-03
GC_7_505 b_7 NI_7 NS_505 0 -6.0351388735178342e-03
GC_7_506 b_7 NI_7 NS_506 0 7.2276062239163726e-03
GC_7_507 b_7 NI_7 NS_507 0 7.9782887395807960e-03
GC_7_508 b_7 NI_7 NS_508 0 -4.7935802390632254e-03
GC_7_509 b_7 NI_7 NS_509 0 -5.4799473742584033e-04
GC_7_510 b_7 NI_7 NS_510 0 5.0230804803338596e-03
GC_7_511 b_7 NI_7 NS_511 0 2.5034134498552686e-04
GC_7_512 b_7 NI_7 NS_512 0 -4.7520661524518403e-03
GC_7_513 b_7 NI_7 NS_513 0 1.7366273020438390e-09
GC_7_514 b_7 NI_7 NS_514 0 3.2860219100700802e-09
GC_7_515 b_7 NI_7 NS_515 0 -1.4394124885462700e-03
GC_7_516 b_7 NI_7 NS_516 0 7.8706604719082883e-03
GC_7_517 b_7 NI_7 NS_517 0 -1.8574746552913943e-04
GC_7_518 b_7 NI_7 NS_518 0 3.0287972650494062e-03
GC_7_519 b_7 NI_7 NS_519 0 -1.2900533253319585e-04
GC_7_520 b_7 NI_7 NS_520 0 -3.3736684356684603e-03
GC_7_521 b_7 NI_7 NS_521 0 -8.9083180904211067e-04
GC_7_522 b_7 NI_7 NS_522 0 7.5293774109587040e-03
GC_7_523 b_7 NI_7 NS_523 0 3.7906243942545602e-03
GC_7_524 b_7 NI_7 NS_524 0 -6.1490577537348500e-03
GC_7_525 b_7 NI_7 NS_525 0 8.8448812800010409e-08
GC_7_526 b_7 NI_7 NS_526 0 -3.5531433930165664e-07
GC_7_527 b_7 NI_7 NS_527 0 6.7115065644237594e-03
GC_7_528 b_7 NI_7 NS_528 0 -5.3183245801310293e-03
GC_7_529 b_7 NI_7 NS_529 0 -2.6127433844451622e-03
GC_7_530 b_7 NI_7 NS_530 0 6.0487711490434587e-03
GC_7_531 b_7 NI_7 NS_531 0 -4.2945275031913274e-03
GC_7_532 b_7 NI_7 NS_532 0 1.3261561751555217e-05
GC_7_533 b_7 NI_7 NS_533 0 2.7224992743036520e-03
GC_7_534 b_7 NI_7 NS_534 0 -6.1956590921680823e-03
GC_7_535 b_7 NI_7 NS_535 0 2.0898364070663384e-03
GC_7_536 b_7 NI_7 NS_536 0 3.2611136133748864e-03
GC_7_537 b_7 NI_7 NS_537 0 -1.9638287434536519e-03
GC_7_538 b_7 NI_7 NS_538 0 -4.4203348271417446e-03
GC_7_539 b_7 NI_7 NS_539 0 2.8567435038813586e-03
GC_7_540 b_7 NI_7 NS_540 0 8.0017787559365106e-03
GC_7_541 b_7 NI_7 NS_541 0 -3.3198038956681582e-03
GC_7_542 b_7 NI_7 NS_542 0 1.8243969736365533e-09
GC_7_543 b_7 NI_7 NS_543 0 5.5833684882506317e-08
GC_7_544 b_7 NI_7 NS_544 0 1.8994901360482345e-06
GC_7_545 b_7 NI_7 NS_545 0 -9.0391646664637700e-05
GC_7_546 b_7 NI_7 NS_546 0 -5.8816387867082406e-05
GC_7_547 b_7 NI_7 NS_547 0 -1.2620480303474628e-03
GC_7_548 b_7 NI_7 NS_548 0 -3.0052300024630717e-04
GC_7_549 b_7 NI_7 NS_549 0 -1.6884323678572589e-03
GC_7_550 b_7 NI_7 NS_550 0 2.6375240576266483e-03
GC_7_551 b_7 NI_7 NS_551 0 4.9218035389979092e-04
GC_7_552 b_7 NI_7 NS_552 0 5.4232981927563786e-03
GC_7_553 b_7 NI_7 NS_553 0 7.0976984383705382e-03
GC_7_554 b_7 NI_7 NS_554 0 6.5580771321231473e-04
GC_7_555 b_7 NI_7 NS_555 0 6.4693545868062610e-04
GC_7_556 b_7 NI_7 NS_556 0 -6.5981442366279223e-04
GC_7_557 b_7 NI_7 NS_557 0 1.0491635822243541e-03
GC_7_558 b_7 NI_7 NS_558 0 1.5730867822218706e-03
GC_7_559 b_7 NI_7 NS_559 0 1.2639593617938720e-02
GC_7_560 b_7 NI_7 NS_560 0 1.3143543386492604e-02
GC_7_561 b_7 NI_7 NS_561 0 8.7648818817715676e-03
GC_7_562 b_7 NI_7 NS_562 0 -2.0356147047613904e-02
GC_7_563 b_7 NI_7 NS_563 0 8.3908943884454714e-03
GC_7_564 b_7 NI_7 NS_564 0 -2.8818702216267126e-03
GC_7_565 b_7 NI_7 NS_565 0 -1.2619354401647647e-02
GC_7_566 b_7 NI_7 NS_566 0 -3.8807125112067846e-02
GC_7_567 b_7 NI_7 NS_567 0 -7.2444869205233698e-03
GC_7_568 b_7 NI_7 NS_568 0 -2.1485688651118975e-03
GC_7_569 b_7 NI_7 NS_569 0 -5.2275000100849435e-02
GC_7_570 b_7 NI_7 NS_570 0 -1.8767871918635125e-03
GC_7_571 b_7 NI_7 NS_571 0 1.4892259625091711e-02
GC_7_572 b_7 NI_7 NS_572 0 8.6975590112820470e-03
GC_7_573 b_7 NI_7 NS_573 0 -5.9275337045537908e-03
GC_7_574 b_7 NI_7 NS_574 0 4.9905441768660543e-03
GC_7_575 b_7 NI_7 NS_575 0 8.3533718485947310e-03
GC_7_576 b_7 NI_7 NS_576 0 1.1690138962478914e-02
GC_7_577 b_7 NI_7 NS_577 0 4.5590097186728584e-03
GC_7_578 b_7 NI_7 NS_578 0 -2.9247916110241739e-03
GC_7_579 b_7 NI_7 NS_579 0 -7.8932468882798104e-03
GC_7_580 b_7 NI_7 NS_580 0 -8.1501572449078977e-03
GC_7_581 b_7 NI_7 NS_581 0 -5.6782670060520632e-03
GC_7_582 b_7 NI_7 NS_582 0 -6.1945380440555774e-04
GC_7_583 b_7 NI_7 NS_583 0 -1.8070910423911013e-02
GC_7_584 b_7 NI_7 NS_584 0 1.3562270005776356e-02
GC_7_585 b_7 NI_7 NS_585 0 4.7006670348608620e-03
GC_7_586 b_7 NI_7 NS_586 0 4.3832608868873595e-03
GC_7_587 b_7 NI_7 NS_587 0 6.4907980629585354e-04
GC_7_588 b_7 NI_7 NS_588 0 -1.1064122178835259e-04
GC_7_589 b_7 NI_7 NS_589 0 -3.7967884222323955e-03
GC_7_590 b_7 NI_7 NS_590 0 8.8034052782955802e-04
GC_7_591 b_7 NI_7 NS_591 0 -1.1248806869058599e-03
GC_7_592 b_7 NI_7 NS_592 0 1.6693625499625869e-02
GC_7_593 b_7 NI_7 NS_593 0 4.4443841504801691e-03
GC_7_594 b_7 NI_7 NS_594 0 7.1164003370832198e-04
GC_7_595 b_7 NI_7 NS_595 0 -5.2105034649928847e-04
GC_7_596 b_7 NI_7 NS_596 0 -2.2476782272340522e-03
GC_7_597 b_7 NI_7 NS_597 0 -4.9869185777709404e-03
GC_7_598 b_7 NI_7 NS_598 0 2.1058931895509008e-03
GC_7_599 b_7 NI_7 NS_599 0 7.3345854317744732e-03
GC_7_600 b_7 NI_7 NS_600 0 1.4346774374826956e-02
GC_7_601 b_7 NI_7 NS_601 0 4.1867521639659643e-03
GC_7_602 b_7 NI_7 NS_602 0 -1.6800211307715807e-03
GC_7_603 b_7 NI_7 NS_603 0 -3.3979285374385582e-03
GC_7_604 b_7 NI_7 NS_604 0 -2.1020210630134854e-03
GC_7_605 b_7 NI_7 NS_605 0 -5.4224785520090831e-03
GC_7_606 b_7 NI_7 NS_606 0 4.3763691520097266e-03
GC_7_607 b_7 NI_7 NS_607 0 1.3191411504853843e-02
GC_7_608 b_7 NI_7 NS_608 0 8.4408863589655204e-03
GC_7_609 b_7 NI_7 NS_609 0 2.8354700790539666e-03
GC_7_610 b_7 NI_7 NS_610 0 -4.1274251979498021e-03
GC_7_611 b_7 NI_7 NS_611 0 -5.3215591020414430e-03
GC_7_612 b_7 NI_7 NS_612 0 1.1333302092413056e-03
GC_7_613 b_7 NI_7 NS_613 0 -4.4370912591425215e-03
GC_7_614 b_7 NI_7 NS_614 0 8.3056987081650876e-03
GC_7_615 b_7 NI_7 NS_615 0 1.4614310659805320e-02
GC_7_616 b_7 NI_7 NS_616 0 -4.5696925851574413e-04
GC_7_617 b_7 NI_7 NS_617 0 -1.1788295653810254e-03
GC_7_618 b_7 NI_7 NS_618 0 -4.5487508157614669e-03
GC_7_619 b_7 NI_7 NS_619 0 -2.2870885734375471e-03
GC_7_620 b_7 NI_7 NS_620 0 4.3793440722958727e-03
GC_7_621 b_7 NI_7 NS_621 0 1.8255978652452984e-10
GC_7_622 b_7 NI_7 NS_622 0 -1.5799966821607916e-09
GC_7_623 b_7 NI_7 NS_623 0 1.4387717869203476e-03
GC_7_624 b_7 NI_7 NS_624 0 8.2177742587030405e-03
GC_7_625 b_7 NI_7 NS_625 0 -8.7491034336598778e-04
GC_7_626 b_7 NI_7 NS_626 0 -2.2094176141329532e-03
GC_7_627 b_7 NI_7 NS_627 0 -1.4716792739190912e-03
GC_7_628 b_7 NI_7 NS_628 0 2.7485700099440106e-03
GC_7_629 b_7 NI_7 NS_629 0 1.7223950886657998e-03
GC_7_630 b_7 NI_7 NS_630 0 7.6102898128641129e-03
GC_7_631 b_7 NI_7 NS_631 0 7.5930424150376097e-03
GC_7_632 b_7 NI_7 NS_632 0 -3.8216231342411799e-03
GC_7_633 b_7 NI_7 NS_633 0 -4.7008126272817050e-08
GC_7_634 b_7 NI_7 NS_634 0 -2.0170256389230800e-08
GC_7_635 b_7 NI_7 NS_635 0 1.1386078508430243e-02
GC_7_636 b_7 NI_7 NS_636 0 4.4716364368288537e-03
GC_7_637 b_7 NI_7 NS_637 0 -8.6429611557318608e-04
GC_7_638 b_7 NI_7 NS_638 0 6.4881769132780044e-03
GC_7_639 b_7 NI_7 NS_639 0 3.6256398046802148e-03
GC_7_640 b_7 NI_7 NS_640 0 4.0760137328029047e-04
GC_7_641 b_7 NI_7 NS_641 0 6.0652186025416457e-03
GC_7_642 b_7 NI_7 NS_642 0 -4.6566353957973846e-03
GC_7_643 b_7 NI_7 NS_643 0 -3.3846298142849603e-03
GC_7_644 b_7 NI_7 NS_644 0 -1.3607984889027435e-03
GC_7_645 b_7 NI_7 NS_645 0 1.0687130397943615e-04
GC_7_646 b_7 NI_7 NS_646 0 4.4902871994920287e-03
GC_7_647 b_7 NI_7 NS_647 0 7.2784000406350803e-03
GC_7_648 b_7 NI_7 NS_648 0 5.5303118943313360e-03
GC_7_649 b_7 NI_7 NS_649 0 -1.3590089392699114e-02
GC_7_650 b_7 NI_7 NS_650 0 5.7574152498781587e-09
GC_7_651 b_7 NI_7 NS_651 0 -1.0755252268142798e-06
GC_7_652 b_7 NI_7 NS_652 0 -2.3265199713856121e-05
GC_7_653 b_7 NI_7 NS_653 0 3.4981896186587222e-04
GC_7_654 b_7 NI_7 NS_654 0 -1.9740617794120256e-04
GC_7_655 b_7 NI_7 NS_655 0 -1.5437475694336465e-03
GC_7_656 b_7 NI_7 NS_656 0 -2.3356984989387521e-03
GC_7_657 b_7 NI_7 NS_657 0 -5.1338576158407424e-05
GC_7_658 b_7 NI_7 NS_658 0 4.3605105822488686e-03
GC_7_659 b_7 NI_7 NS_659 0 1.6175854247142774e-03
GC_7_660 b_7 NI_7 NS_660 0 -5.9520447551457941e-03
GC_7_661 b_7 NI_7 NS_661 0 -4.9853642799082267e-03
GC_7_662 b_7 NI_7 NS_662 0 6.4563496909199889e-03
GC_7_663 b_7 NI_7 NS_663 0 1.1341369443483389e-03
GC_7_664 b_7 NI_7 NS_664 0 -5.0676047520778109e-04
GC_7_665 b_7 NI_7 NS_665 0 2.7870925906266150e-03
GC_7_666 b_7 NI_7 NS_666 0 2.3388070901896596e-03
GC_7_667 b_7 NI_7 NS_667 0 -4.3321840737588517e-03
GC_7_668 b_7 NI_7 NS_668 0 -1.3583569026987050e-02
GC_7_669 b_7 NI_7 NS_669 0 1.5695054733302852e-03
GC_7_670 b_7 NI_7 NS_670 0 1.7683056108125223e-02
GC_7_671 b_7 NI_7 NS_671 0 9.8323100585864433e-03
GC_7_672 b_7 NI_7 NS_672 0 -2.3109433971130354e-03
GC_7_673 b_7 NI_7 NS_673 0 -1.3157076653895131e-02
GC_7_674 b_7 NI_7 NS_674 0 2.2142577719871078e-03
GC_7_675 b_7 NI_7 NS_675 0 9.1925801996316971e-03
GC_7_676 b_7 NI_7 NS_676 0 1.9425128055761706e-03
GC_7_677 b_7 NI_7 NS_677 0 -1.8069416737093048e-02
GC_7_678 b_7 NI_7 NS_678 0 -6.4922072793173963e-03
GC_7_679 b_7 NI_7 NS_679 0 1.5725031894717332e-02
GC_7_680 b_7 NI_7 NS_680 0 6.4951372716309857e-03
GC_7_681 b_7 NI_7 NS_681 0 8.1032021061081209e-03
GC_7_682 b_7 NI_7 NS_682 0 -4.2110865808055445e-03
GC_7_683 b_7 NI_7 NS_683 0 -7.5660733787598442e-03
GC_7_684 b_7 NI_7 NS_684 0 2.0432108254831364e-03
GC_7_685 b_7 NI_7 NS_685 0 6.6854403795751829e-03
GC_7_686 b_7 NI_7 NS_686 0 -2.7541191547744105e-03
GC_7_687 b_7 NI_7 NS_687 0 -6.6055143819589487e-03
GC_7_688 b_7 NI_7 NS_688 0 2.9142089168934042e-03
GC_7_689 b_7 NI_7 NS_689 0 7.6544550432042181e-03
GC_7_690 b_7 NI_7 NS_690 0 4.7731847373014589e-04
GC_7_691 b_7 NI_7 NS_691 0 -9.4088383419283876e-03
GC_7_692 b_7 NI_7 NS_692 0 -5.1695913268953253e-03
GC_7_693 b_7 NI_7 NS_693 0 6.8169860777995061e-03
GC_7_694 b_7 NI_7 NS_694 0 4.1131838889597316e-03
GC_7_695 b_7 NI_7 NS_695 0 -3.9575075777864267e-04
GC_7_696 b_7 NI_7 NS_696 0 -9.3603865378936611e-04
GC_7_697 b_7 NI_7 NS_697 0 5.6653330903600231e-03
GC_7_698 b_7 NI_7 NS_698 0 -1.3801763521175095e-03
GC_7_699 b_7 NI_7 NS_699 0 -9.2023055604558996e-03
GC_7_700 b_7 NI_7 NS_700 0 -1.2455924515792157e-03
GC_7_701 b_7 NI_7 NS_701 0 5.9915361490972992e-03
GC_7_702 b_7 NI_7 NS_702 0 7.3808288926772287e-04
GC_7_703 b_7 NI_7 NS_703 0 -2.6544499887793493e-03
GC_7_704 b_7 NI_7 NS_704 0 2.4842218286510217e-04
GC_7_705 b_7 NI_7 NS_705 0 6.6958869570911891e-03
GC_7_706 b_7 NI_7 NS_706 0 -2.2582332604381469e-03
GC_7_707 b_7 NI_7 NS_707 0 -9.3158034337999952e-03
GC_7_708 b_7 NI_7 NS_708 0 1.5268579780517778e-03
GC_7_709 b_7 NI_7 NS_709 0 5.7300528240279685e-03
GC_7_710 b_7 NI_7 NS_710 0 -1.5007464209294875e-03
GC_7_711 b_7 NI_7 NS_711 0 -3.3211786392641422e-03
GC_7_712 b_7 NI_7 NS_712 0 2.4082406838792899e-03
GC_7_713 b_7 NI_7 NS_713 0 7.2643748459257917e-03
GC_7_714 b_7 NI_7 NS_714 0 -4.0966020234659744e-03
GC_7_715 b_7 NI_7 NS_715 0 -8.5936626208300542e-03
GC_7_716 b_7 NI_7 NS_716 0 4.2025458057810602e-03
GC_7_717 b_7 NI_7 NS_717 0 4.8158718107756595e-03
GC_7_718 b_7 NI_7 NS_718 0 -3.8696534356426502e-03
GC_7_719 b_7 NI_7 NS_719 0 -2.4037832577575684e-03
GC_7_720 b_7 NI_7 NS_720 0 4.7598869813827134e-03
GC_7_721 b_7 NI_7 NS_721 0 7.0540650269529112e-03
GC_7_722 b_7 NI_7 NS_722 0 -7.3479411359844296e-03
GC_7_723 b_7 NI_7 NS_723 0 -7.1270973131398437e-03
GC_7_724 b_7 NI_7 NS_724 0 6.8936460130061836e-03
GC_7_725 b_7 NI_7 NS_725 0 1.6683535826806420e-03
GC_7_726 b_7 NI_7 NS_726 0 -5.2972271114586399e-03
GC_7_727 b_7 NI_7 NS_727 0 5.9423054445024959e-04
GC_7_728 b_7 NI_7 NS_728 0 5.4734750972633764e-03
GC_7_729 b_7 NI_7 NS_729 0 -4.1995963854246135e-09
GC_7_730 b_7 NI_7 NS_730 0 -1.3215418100235201e-08
GC_7_731 b_7 NI_7 NS_731 0 2.7118337317610826e-03
GC_7_732 b_7 NI_7 NS_732 0 -8.5806168970764384e-03
GC_7_733 b_7 NI_7 NS_733 0 8.7189177798857977e-04
GC_7_734 b_7 NI_7 NS_734 0 -3.4318677496628651e-03
GC_7_735 b_7 NI_7 NS_735 0 6.2897519477440303e-04
GC_7_736 b_7 NI_7 NS_736 0 4.0346891063129438e-03
GC_7_737 b_7 NI_7 NS_737 0 2.1766552368069174e-03
GC_7_738 b_7 NI_7 NS_738 0 -8.1586502032182876e-03
GC_7_739 b_7 NI_7 NS_739 0 -3.4870473344026519e-03
GC_7_740 b_7 NI_7 NS_740 0 7.0184761649911805e-03
GC_7_741 b_7 NI_7 NS_741 0 -9.0339788463068094e-08
GC_7_742 b_7 NI_7 NS_742 0 -3.0341137820754849e-07
GC_7_743 b_7 NI_7 NS_743 0 -8.0011228498603117e-03
GC_7_744 b_7 NI_7 NS_744 0 5.3809315920449498e-03
GC_7_745 b_7 NI_7 NS_745 0 4.1753805465283879e-03
GC_7_746 b_7 NI_7 NS_746 0 -6.8471567929904303e-03
GC_7_747 b_7 NI_7 NS_747 0 5.3267681360825271e-03
GC_7_748 b_7 NI_7 NS_748 0 7.4221548312965646e-04
GC_7_749 b_7 NI_7 NS_749 0 -2.3672741529545526e-03
GC_7_750 b_7 NI_7 NS_750 0 6.8575158556994590e-03
GC_7_751 b_7 NI_7 NS_751 0 -1.4866263327028761e-03
GC_7_752 b_7 NI_7 NS_752 0 -4.2154565571034574e-03
GC_7_753 b_7 NI_7 NS_753 0 2.3568559828399311e-03
GC_7_754 b_7 NI_7 NS_754 0 5.0372654950294731e-03
GC_7_755 b_7 NI_7 NS_755 0 -1.9997028978518201e-03
GC_7_756 b_7 NI_7 NS_756 0 -8.9736634094011031e-03
GC_7_757 b_7 NI_7 NS_757 0 -1.0963348981826430e-02
GC_7_758 b_7 NI_7 NS_758 0 8.3273459788010237e-09
GC_7_759 b_7 NI_7 NS_759 0 9.8608137541309655e-07
GC_7_760 b_7 NI_7 NS_760 0 3.6177580692637438e-05
GC_7_761 b_7 NI_7 NS_761 0 4.3739130100030089e-03
GC_7_762 b_7 NI_7 NS_762 0 -3.4750208144883866e-03
GC_7_763 b_7 NI_7 NS_763 0 -3.7382650588349020e-03
GC_7_764 b_7 NI_7 NS_764 0 6.2463706263140252e-03
GC_7_765 b_7 NI_7 NS_765 0 -8.7586408136103074e-03
GC_7_766 b_7 NI_7 NS_766 0 -5.9567967208995808e-03
GC_7_767 b_7 NI_7 NS_767 0 9.2115220543326926e-03
GC_7_768 b_7 NI_7 NS_768 0 -5.9461552367250049e-03
GC_7_769 b_7 NI_7 NS_769 0 7.1478496073212536e-03
GC_7_770 b_7 NI_7 NS_770 0 1.1907364851750354e-02
GC_7_771 b_7 NI_7 NS_771 0 -4.2314406862432805e-03
GC_7_772 b_7 NI_7 NS_772 0 -1.1324311754482670e-03
GC_7_773 b_7 NI_7 NS_773 0 -8.8598538031035897e-03
GC_7_774 b_7 NI_7 NS_774 0 -4.7416934372835739e-04
GC_7_775 b_7 NI_7 NS_775 0 1.4618428117404434e-02
GC_7_776 b_7 NI_7 NS_776 0 -1.0343814043206388e-02
GC_7_777 b_7 NI_7 NS_777 0 1.6441829610098921e-02
GC_7_778 b_7 NI_7 NS_778 0 4.0225220955532317e-03
GC_7_779 b_7 NI_7 NS_779 0 -1.1482359602821597e-02
GC_7_780 b_7 NI_7 NS_780 0 -2.4511076715170093e-04
GC_7_781 b_7 NI_7 NS_781 0 -1.6636907869808815e-02
GC_7_782 b_7 NI_7 NS_782 0 -4.4573833539531739e-02
GC_7_783 b_7 NI_7 NS_783 0 1.0652627781026205e-02
GC_7_784 b_7 NI_7 NS_784 0 1.1245836704824759e-03
GC_7_785 b_7 NI_7 NS_785 0 -4.8294133162753633e-02
GC_7_786 b_7 NI_7 NS_786 0 1.1061825357444450e-02
GC_7_787 b_7 NI_7 NS_787 0 -1.0433724890290598e-02
GC_7_788 b_7 NI_7 NS_788 0 4.8880722943306398e-04
GC_7_789 b_7 NI_7 NS_789 0 9.7769814577245238e-03
GC_7_790 b_7 NI_7 NS_790 0 -5.7678189360910387e-04
GC_7_791 b_7 NI_7 NS_791 0 4.6096264294178384e-03
GC_7_792 b_7 NI_7 NS_792 0 2.4174063328432173e-02
GC_7_793 b_7 NI_7 NS_793 0 -1.0735334757404506e-02
GC_7_794 b_7 NI_7 NS_794 0 1.9692205285333675e-03
GC_7_795 b_7 NI_7 NS_795 0 -8.4726763358986650e-03
GC_7_796 b_7 NI_7 NS_796 0 -1.3537888744257891e-02
GC_7_797 b_7 NI_7 NS_797 0 1.0150146799700815e-02
GC_7_798 b_7 NI_7 NS_798 0 9.8140578254577826e-04
GC_7_799 b_7 NI_7 NS_799 0 -1.9163081124141737e-02
GC_7_800 b_7 NI_7 NS_800 0 2.8679163645573689e-02
GC_7_801 b_7 NI_7 NS_801 0 -9.6128534059335673e-03
GC_7_802 b_7 NI_7 NS_802 0 -9.6555955252516381e-04
GC_7_803 b_7 NI_7 NS_803 0 1.8914255743890747e-03
GC_7_804 b_7 NI_7 NS_804 0 -1.3780579732376864e-03
GC_7_805 b_7 NI_7 NS_805 0 9.4683004623363556e-03
GC_7_806 b_7 NI_7 NS_806 0 -2.4742048931168523e-04
GC_7_807 b_7 NI_7 NS_807 0 -1.4944029195498548e-04
GC_7_808 b_7 NI_7 NS_808 0 3.0270110750136282e-02
GC_7_809 b_7 NI_7 NS_809 0 -8.5288571474533385e-03
GC_7_810 b_7 NI_7 NS_810 0 1.5479029107857520e-04
GC_7_811 b_7 NI_7 NS_811 0 2.1683696568205440e-04
GC_7_812 b_7 NI_7 NS_812 0 -5.4812504195694460e-03
GC_7_813 b_7 NI_7 NS_813 0 1.0036183359561534e-02
GC_7_814 b_7 NI_7 NS_814 0 -3.3857046458688161e-04
GC_7_815 b_7 NI_7 NS_815 0 8.9342197380139505e-03
GC_7_816 b_7 NI_7 NS_816 0 2.6365790566234219e-02
GC_7_817 b_7 NI_7 NS_817 0 -8.3555257129623705e-03
GC_7_818 b_7 NI_7 NS_818 0 1.3766353521306978e-03
GC_7_819 b_7 NI_7 NS_819 0 -2.5869003037965813e-03
GC_7_820 b_7 NI_7 NS_820 0 -7.3539855532168954e-03
GC_7_821 b_7 NI_7 NS_821 0 1.0553574481281474e-02
GC_7_822 b_7 NI_7 NS_822 0 -8.2350362934182318e-04
GC_7_823 b_7 NI_7 NS_823 0 1.4438990691573983e-02
GC_7_824 b_7 NI_7 NS_824 0 1.9950572998707252e-02
GC_7_825 b_7 NI_7 NS_825 0 -8.2760929479172261e-03
GC_7_826 b_7 NI_7 NS_826 0 2.9305026858324913e-03
GC_7_827 b_7 NI_7 NS_827 0 -5.5941981722551666e-03
GC_7_828 b_7 NI_7 NS_828 0 -6.9177081116038337e-03
GC_7_829 b_7 NI_7 NS_829 0 1.1244066907563639e-02
GC_7_830 b_7 NI_7 NS_830 0 -1.3754115571425990e-03
GC_7_831 b_7 NI_7 NS_831 0 1.5700535733520513e-02
GC_7_832 b_7 NI_7 NS_832 0 1.2945582787109602e-02
GC_7_833 b_7 NI_7 NS_833 0 -7.1893581632682642e-03
GC_7_834 b_7 NI_7 NS_834 0 5.1106031408532518e-03
GC_7_835 b_7 NI_7 NS_835 0 -6.8765855225411832e-03
GC_7_836 b_7 NI_7 NS_836 0 -4.8360476722872411e-03
GC_7_837 b_7 NI_7 NS_837 0 4.7733861887687582e-09
GC_7_838 b_7 NI_7 NS_838 0 4.4198788423842333e-08
GC_7_839 b_7 NI_7 NS_839 0 1.2004109539084519e-02
GC_7_840 b_7 NI_7 NS_840 0 -2.5766667985547792e-03
GC_7_841 b_7 NI_7 NS_841 0 -5.2510748822878059e-03
GC_7_842 b_7 NI_7 NS_842 0 4.7015434585164634e-03
GC_7_843 b_7 NI_7 NS_843 0 -6.1588977770092729e-03
GC_7_844 b_7 NI_7 NS_844 0 -4.3232047873268649e-03
GC_7_845 b_7 NI_7 NS_845 0 1.1774222757480588e-02
GC_7_846 b_7 NI_7 NS_846 0 -3.7297245581477466e-03
GC_7_847 b_7 NI_7 NS_847 0 1.2978425484962117e-02
GC_7_848 b_7 NI_7 NS_848 0 9.4653912116303748e-03
GC_7_849 b_7 NI_7 NS_849 0 3.9180865256078189e-06
GC_7_850 b_7 NI_7 NS_850 0 -9.4184499384502609e-07
GC_7_851 b_7 NI_7 NS_851 0 1.6087880668846286e-02
GC_7_852 b_7 NI_7 NS_852 0 1.6769944407268818e-02
GC_7_853 b_7 NI_7 NS_853 0 1.2047068907067899e-02
GC_7_854 b_7 NI_7 NS_854 0 -2.4806934766404940e-03
GC_7_855 b_7 NI_7 NS_855 0 -8.3607712443942439e-03
GC_7_856 b_7 NI_7 NS_856 0 7.9691115098588070e-05
GC_7_857 b_7 NI_7 NS_857 0 1.1309399053679902e-02
GC_7_858 b_7 NI_7 NS_858 0 7.3306425655571723e-03
GC_7_859 b_7 NI_7 NS_859 0 -4.6732532631951216e-03
GC_7_860 b_7 NI_7 NS_860 0 7.3569206939826208e-03
GC_7_861 b_7 NI_7 NS_861 0 -8.0809736139068524e-03
GC_7_862 b_7 NI_7 NS_862 0 -3.7224024938438639e-03
GC_7_863 b_7 NI_7 NS_863 0 1.5958294213797873e-02
GC_7_864 b_7 NI_7 NS_864 0 -7.7554800609770866e-03
GC_7_865 b_7 NI_7 NS_865 0 5.6902093423388727e-05
GC_7_866 b_7 NI_7 NS_866 0 -1.2101497968766654e-10
GC_7_867 b_7 NI_7 NS_867 0 -2.0303366611081539e-09
GC_7_868 b_7 NI_7 NS_868 0 3.4201182266648488e-08
GC_7_869 b_7 NI_7 NS_869 0 -5.1436491854061222e-07
GC_7_870 b_7 NI_7 NS_870 0 -3.8156305152981841e-07
GC_7_871 b_7 NI_7 NS_871 0 -8.7410298584905201e-07
GC_7_872 b_7 NI_7 NS_872 0 9.5756911806380033e-06
GC_7_873 b_7 NI_7 NS_873 0 1.2647595038002632e-05
GC_7_874 b_7 NI_7 NS_874 0 -1.2046156964301665e-05
GC_7_875 b_7 NI_7 NS_875 0 -1.7539276855345540e-05
GC_7_876 b_7 NI_7 NS_876 0 8.8319931092852381e-06
GC_7_877 b_7 NI_7 NS_877 0 2.8401356102728134e-05
GC_7_878 b_7 NI_7 NS_878 0 -6.5602080510244538e-06
GC_7_879 b_7 NI_7 NS_879 0 -3.2049432553514889e-06
GC_7_880 b_7 NI_7 NS_880 0 -3.0960968420523310e-06
GC_7_881 b_7 NI_7 NS_881 0 -2.8498746517432749e-06
GC_7_882 b_7 NI_7 NS_882 0 -1.4497135355042237e-05
GC_7_883 b_7 NI_7 NS_883 0 -2.4758797607658901e-05
GC_7_884 b_7 NI_7 NS_884 0 4.0215888953601763e-05
GC_7_885 b_7 NI_7 NS_885 0 3.7734251543373230e-05
GC_7_886 b_7 NI_7 NS_886 0 -4.7032653194256001e-05
GC_7_887 b_7 NI_7 NS_887 0 -3.0428739551672947e-05
GC_7_888 b_7 NI_7 NS_888 0 -2.0941082668923348e-05
GC_7_889 b_7 NI_7 NS_889 0 3.3065697995894667e-05
GC_7_890 b_7 NI_7 NS_890 0 2.6831766976384883e-05
GC_7_891 b_7 NI_7 NS_891 0 -1.8367588008954196e-05
GC_7_892 b_7 NI_7 NS_892 0 -2.8795047652233076e-05
GC_7_893 b_7 NI_7 NS_893 0 2.1463776587106759e-05
GC_7_894 b_7 NI_7 NS_894 0 6.0257593036310044e-05
GC_7_895 b_7 NI_7 NS_895 0 -2.1175885143587752e-05
GC_7_896 b_7 NI_7 NS_896 0 -5.5544466880166393e-05
GC_7_897 b_7 NI_7 NS_897 0 -3.1395988025785353e-05
GC_7_898 b_7 NI_7 NS_898 0 -1.1645823528632582e-05
GC_7_899 b_7 NI_7 NS_899 0 2.0313078482073281e-05
GC_7_900 b_7 NI_7 NS_900 0 1.3868917036846245e-05
GC_7_901 b_7 NI_7 NS_901 0 -2.4579282099446013e-05
GC_7_902 b_7 NI_7 NS_902 0 -1.0925906040923385e-05
GC_7_903 b_7 NI_7 NS_903 0 2.0765200319146652e-05
GC_7_904 b_7 NI_7 NS_904 0 1.0076894291539012e-05
GC_7_905 b_7 NI_7 NS_905 0 -1.8224310152157206e-05
GC_7_906 b_7 NI_7 NS_906 0 -2.0845754904284453e-05
GC_7_907 b_7 NI_7 NS_907 0 5.4971700006793713e-06
GC_7_908 b_7 NI_7 NS_908 0 3.2160028343369790e-05
GC_7_909 b_7 NI_7 NS_909 0 -8.2126411937722956e-06
GC_7_910 b_7 NI_7 NS_910 0 -2.6520248110671897e-05
GC_7_911 b_7 NI_7 NS_911 0 -1.8293638144835498e-06
GC_7_912 b_7 NI_7 NS_912 0 1.6901090469052797e-06
GC_7_913 b_7 NI_7 NS_913 0 -1.9229428525516533e-05
GC_7_914 b_7 NI_7 NS_914 0 -1.1940389295159550e-05
GC_7_915 b_7 NI_7 NS_915 0 6.9715891916813242e-06
GC_7_916 b_7 NI_7 NS_916 0 2.0939279618377833e-05
GC_7_917 b_7 NI_7 NS_917 0 -1.5976584568600856e-05
GC_7_918 b_7 NI_7 NS_918 0 -1.4813682394233148e-05
GC_7_919 b_7 NI_7 NS_919 0 1.3385310440314107e-06
GC_7_920 b_7 NI_7 NS_920 0 5.3014194841579197e-06
GC_7_921 b_7 NI_7 NS_921 0 -2.4841398268693000e-05
GC_7_922 b_7 NI_7 NS_922 0 -9.8244215834397053e-06
GC_7_923 b_7 NI_7 NS_923 0 8.5458021642558965e-06
GC_7_924 b_7 NI_7 NS_924 0 2.3051008505913615e-05
GC_7_925 b_7 NI_7 NS_925 0 -2.0672703839776976e-05
GC_7_926 b_7 NI_7 NS_926 0 -5.6252260129033698e-06
GC_7_927 b_7 NI_7 NS_927 0 6.2604061522386173e-06
GC_7_928 b_7 NI_7 NS_928 0 7.5159774017725214e-06
GC_7_929 b_7 NI_7 NS_929 0 -3.0565110074478262e-05
GC_7_930 b_7 NI_7 NS_930 0 -2.5578435869723339e-06
GC_7_931 b_7 NI_7 NS_931 0 1.8794275591178957e-05
GC_7_932 b_7 NI_7 NS_932 0 2.5290693985582271e-05
GC_7_933 b_7 NI_7 NS_933 0 -2.1787356163786520e-05
GC_7_934 b_7 NI_7 NS_934 0 6.9643264419352430e-06
GC_7_935 b_7 NI_7 NS_935 0 1.5266699242892035e-05
GC_7_936 b_7 NI_7 NS_936 0 3.9769083095713419e-06
GC_7_937 b_7 NI_7 NS_937 0 -3.4533195713567385e-05
GC_7_938 b_7 NI_7 NS_938 0 1.3723106986026460e-05
GC_7_939 b_7 NI_7 NS_939 0 3.7468926805963499e-05
GC_7_940 b_7 NI_7 NS_940 0 1.2337879234222103e-05
GC_7_941 b_7 NI_7 NS_941 0 -7.7468826747346917e-06
GC_7_942 b_7 NI_7 NS_942 0 1.8808846610432296e-05
GC_7_943 b_7 NI_7 NS_943 0 1.2774791679486795e-05
GC_7_944 b_7 NI_7 NS_944 0 -1.1287274821811191e-05
GC_7_945 b_7 NI_7 NS_945 0 1.0984712330284056e-10
GC_7_946 b_7 NI_7 NS_946 0 3.5338508198594203e-11
GC_7_947 b_7 NI_7 NS_947 0 -1.3692658994745888e-05
GC_7_948 b_7 NI_7 NS_948 0 2.5942031526095177e-05
GC_7_949 b_7 NI_7 NS_949 0 -2.0635045549449428e-06
GC_7_950 b_7 NI_7 NS_950 0 1.0503207275281666e-05
GC_7_951 b_7 NI_7 NS_951 0 6.1728472679227264e-06
GC_7_952 b_7 NI_7 NS_952 0 -8.5363569231054215e-06
GC_7_953 b_7 NI_7 NS_953 0 -8.1127304160819484e-06
GC_7_954 b_7 NI_7 NS_954 0 2.5390652982189230e-05
GC_7_955 b_7 NI_7 NS_955 0 2.4972769473836168e-05
GC_7_956 b_7 NI_7 NS_956 0 -1.0420768266848149e-05
GC_7_957 b_7 NI_7 NS_957 0 4.8846708363307946e-09
GC_7_958 b_7 NI_7 NS_958 0 -1.2244750555021914e-09
GC_7_959 b_7 NI_7 NS_959 0 2.6368527704139106e-05
GC_7_960 b_7 NI_7 NS_960 0 -1.2610361652808703e-05
GC_7_961 b_7 NI_7 NS_961 0 -8.2494856152927020e-06
GC_7_962 b_7 NI_7 NS_962 0 1.8114633529210649e-05
GC_7_963 b_7 NI_7 NS_963 0 -1.0378260542242953e-05
GC_7_964 b_7 NI_7 NS_964 0 -3.0219654485094672e-07
GC_7_965 b_7 NI_7 NS_965 0 1.9390177844513017e-05
GC_7_966 b_7 NI_7 NS_966 0 -1.4388822649680083e-05
GC_7_967 b_7 NI_7 NS_967 0 7.1948773173901266e-06
GC_7_968 b_7 NI_7 NS_968 0 1.1599588890965741e-05
GC_7_969 b_7 NI_7 NS_969 0 -2.2864918042583392e-07
GC_7_970 b_7 NI_7 NS_970 0 -1.4637611558960359e-05
GC_7_971 b_7 NI_7 NS_971 0 1.3160146689539436e-05
GC_7_972 b_7 NI_7 NS_972 0 2.7988798207563730e-05
GC_7_973 b_7 NI_7 NS_973 0 -6.3809589100370006e-04
GC_7_974 b_7 NI_7 NS_974 0 -9.7135985355233427e-11
GC_7_975 b_7 NI_7 NS_975 0 3.8809012817708924e-09
GC_7_976 b_7 NI_7 NS_976 0 -6.7422274949627611e-08
GC_7_977 b_7 NI_7 NS_977 0 -1.1286634338698946e-05
GC_7_978 b_7 NI_7 NS_978 0 -9.3365543637775104e-06
GC_7_979 b_7 NI_7 NS_979 0 -2.2471556609682971e-06
GC_7_980 b_7 NI_7 NS_980 0 2.3210495738364341e-07
GC_7_981 b_7 NI_7 NS_981 0 -3.0313696705542765e-05
GC_7_982 b_7 NI_7 NS_982 0 2.7072956297279158e-05
GC_7_983 b_7 NI_7 NS_983 0 -3.3247384458935047e-05
GC_7_984 b_7 NI_7 NS_984 0 8.1286562346541068e-06
GC_7_985 b_7 NI_7 NS_985 0 3.1755754034795042e-05
GC_7_986 b_7 NI_7 NS_986 0 2.7371065044610979e-05
GC_7_987 b_7 NI_7 NS_987 0 -9.0592365607737122e-06
GC_7_988 b_7 NI_7 NS_988 0 1.4745493117446728e-05
GC_7_989 b_7 NI_7 NS_989 0 1.2657458209755026e-05
GC_7_990 b_7 NI_7 NS_990 0 3.6938816717762177e-05
GC_7_991 b_7 NI_7 NS_991 0 -1.0625069484968271e-05
GC_7_992 b_7 NI_7 NS_992 0 6.8145131275435068e-05
GC_7_993 b_7 NI_7 NS_993 0 9.5462337680982353e-05
GC_7_994 b_7 NI_7 NS_994 0 -6.6200955206056067e-05
GC_7_995 b_7 NI_7 NS_995 0 2.7086627864076785e-05
GC_7_996 b_7 NI_7 NS_996 0 3.1697630810383419e-05
GC_7_997 b_7 NI_7 NS_997 0 -7.3750444451776447e-06
GC_7_998 b_7 NI_7 NS_998 0 -7.2639306672962544e-05
GC_7_999 b_7 NI_7 NS_999 0 -9.8543925208709574e-06
GC_7_1000 b_7 NI_7 NS_1000 0 -3.3996033600476389e-05
GC_7_1001 b_7 NI_7 NS_1001 0 -7.7016997498360152e-05
GC_7_1002 b_7 NI_7 NS_1002 0 1.9071607922172825e-05
GC_7_1003 b_7 NI_7 NS_1003 0 2.4929646163584060e-05
GC_7_1004 b_7 NI_7 NS_1004 0 5.0927035276202100e-05
GC_7_1005 b_7 NI_7 NS_1005 0 -2.3148587796001884e-05
GC_7_1006 b_7 NI_7 NS_1006 0 -3.5473797730263880e-06
GC_7_1007 b_7 NI_7 NS_1007 0 6.9848633035912860e-05
GC_7_1008 b_7 NI_7 NS_1008 0 4.4676895603441971e-05
GC_7_1009 b_7 NI_7 NS_1009 0 2.9208030456246231e-05
GC_7_1010 b_7 NI_7 NS_1010 0 1.9693885759761100e-05
GC_7_1011 b_7 NI_7 NS_1011 0 -7.3329286185316995e-06
GC_7_1012 b_7 NI_7 NS_1012 0 -2.5741690024422878e-05
GC_7_1013 b_7 NI_7 NS_1013 0 -7.5876248188038902e-06
GC_7_1014 b_7 NI_7 NS_1014 0 -2.5167217829747839e-05
GC_7_1015 b_7 NI_7 NS_1015 0 6.7364185748551757e-06
GC_7_1016 b_7 NI_7 NS_1016 0 4.9241814029544812e-05
GC_7_1017 b_7 NI_7 NS_1017 0 1.2922943614808559e-05
GC_7_1018 b_7 NI_7 NS_1018 0 2.7360377523625716e-05
GC_7_1019 b_7 NI_7 NS_1019 0 5.8665038648906798e-06
GC_7_1020 b_7 NI_7 NS_1020 0 2.1248438208371524e-06
GC_7_1021 b_7 NI_7 NS_1021 0 -6.3215456580183611e-07
GC_7_1022 b_7 NI_7 NS_1022 0 -1.5379666031993652e-05
GC_7_1023 b_7 NI_7 NS_1023 0 5.6145726161734163e-05
GC_7_1024 b_7 NI_7 NS_1024 0 3.8184732187509650e-05
GC_7_1025 b_7 NI_7 NS_1025 0 1.9943094176905348e-05
GC_7_1026 b_7 NI_7 NS_1026 0 1.4808803766565994e-05
GC_7_1027 b_7 NI_7 NS_1027 0 8.3810729239559633e-06
GC_7_1028 b_7 NI_7 NS_1028 0 -1.2844653484838514e-05
GC_7_1029 b_7 NI_7 NS_1029 0 -5.6561618513691115e-06
GC_7_1030 b_7 NI_7 NS_1030 0 -1.3981126542408287e-05
GC_7_1031 b_7 NI_7 NS_1031 0 6.6094138757294372e-05
GC_7_1032 b_7 NI_7 NS_1032 0 1.3028891582634993e-05
GC_7_1033 b_7 NI_7 NS_1033 0 2.2769668837713581e-05
GC_7_1034 b_7 NI_7 NS_1034 0 4.9311356817032155e-06
GC_7_1035 b_7 NI_7 NS_1035 0 -5.5540359488588195e-06
GC_7_1036 b_7 NI_7 NS_1036 0 -2.1975719204796177e-05
GC_7_1037 b_7 NI_7 NS_1037 0 -9.1463352557649051e-06
GC_7_1038 b_7 NI_7 NS_1038 0 -7.0651012264413655e-06
GC_7_1039 b_7 NI_7 NS_1039 0 6.0665964719695408e-05
GC_7_1040 b_7 NI_7 NS_1040 0 -9.4701623989225406e-06
GC_7_1041 b_7 NI_7 NS_1041 0 2.1425125660485143e-05
GC_7_1042 b_7 NI_7 NS_1042 0 -7.3811012174990269e-06
GC_7_1043 b_7 NI_7 NS_1043 0 -2.3068068868007783e-05
GC_7_1044 b_7 NI_7 NS_1044 0 -1.3110914697563906e-05
GC_7_1045 b_7 NI_7 NS_1045 0 -8.6671553808734461e-06
GC_7_1046 b_7 NI_7 NS_1046 0 4.4627804793682517e-06
GC_7_1047 b_7 NI_7 NS_1047 0 4.5473391861639589e-05
GC_7_1048 b_7 NI_7 NS_1048 0 -2.5661818385631497e-05
GC_7_1049 b_7 NI_7 NS_1049 0 6.0269477960900150e-06
GC_7_1050 b_7 NI_7 NS_1050 0 -1.6485832030230712e-05
GC_7_1051 b_7 NI_7 NS_1051 0 -1.8722678595157823e-05
GC_7_1052 b_7 NI_7 NS_1052 0 8.6301690229459830e-06
GC_7_1053 b_7 NI_7 NS_1053 0 -4.6983879414721009e-11
GC_7_1054 b_7 NI_7 NS_1054 0 -1.7787115840534583e-10
GC_7_1055 b_7 NI_7 NS_1055 0 1.7486976986880226e-06
GC_7_1056 b_7 NI_7 NS_1056 0 8.7729613863640251e-06
GC_7_1057 b_7 NI_7 NS_1057 0 2.2060668170288899e-06
GC_7_1058 b_7 NI_7 NS_1058 0 -7.0028082450527230e-06
GC_7_1059 b_7 NI_7 NS_1059 0 -9.0193539593989135e-06
GC_7_1060 b_7 NI_7 NS_1060 0 5.7725428025680062e-06
GC_7_1061 b_7 NI_7 NS_1061 0 4.7628863931968367e-06
GC_7_1062 b_7 NI_7 NS_1062 0 1.1522803286950406e-05
GC_7_1063 b_7 NI_7 NS_1063 0 2.4566772071145011e-05
GC_7_1064 b_7 NI_7 NS_1064 0 -2.1153857919134811e-05
GC_7_1065 b_7 NI_7 NS_1065 0 -5.7421782045878141e-09
GC_7_1066 b_7 NI_7 NS_1066 0 -5.6214288493594294e-09
GC_7_1067 b_7 NI_7 NS_1067 0 3.0633018313586341e-05
GC_7_1068 b_7 NI_7 NS_1068 0 7.5206529009410168e-06
GC_7_1069 b_7 NI_7 NS_1069 0 -2.6889442654711343e-06
GC_7_1070 b_7 NI_7 NS_1070 0 1.1036276927505903e-05
GC_7_1071 b_7 NI_7 NS_1071 0 8.0385273229214092e-06
GC_7_1072 b_7 NI_7 NS_1072 0 1.1983682472872218e-06
GC_7_1073 b_7 NI_7 NS_1073 0 1.9085223137004534e-05
GC_7_1074 b_7 NI_7 NS_1074 0 -2.1544589911361024e-05
GC_7_1075 b_7 NI_7 NS_1075 0 -6.5775870974882853e-06
GC_7_1076 b_7 NI_7 NS_1076 0 -7.4340050883479901e-06
GC_7_1077 b_7 NI_7 NS_1077 0 -5.4042926599403817e-06
GC_7_1078 b_7 NI_7 NS_1078 0 1.2516897398937941e-05
GC_7_1079 b_7 NI_7 NS_1079 0 1.6097136864025916e-05
GC_7_1080 b_7 NI_7 NS_1080 0 7.3672698972032669e-06
GC_7_1081 b_7 NI_7 NS_1081 0 -5.0477230321812300e-05
GC_7_1082 b_7 NI_7 NS_1082 0 -7.9794554981852371e-12
GC_7_1083 b_7 NI_7 NS_1083 0 -2.0628673241437072e-10
GC_7_1084 b_7 NI_7 NS_1084 0 9.8384590385688702e-09
GC_7_1085 b_7 NI_7 NS_1085 0 5.6375621180128711e-07
GC_7_1086 b_7 NI_7 NS_1086 0 4.4381074681424582e-08
GC_7_1087 b_7 NI_7 NS_1087 0 2.9366447355701418e-06
GC_7_1088 b_7 NI_7 NS_1088 0 -1.4886584018811337e-06
GC_7_1089 b_7 NI_7 NS_1089 0 -3.1321941535235076e-06
GC_7_1090 b_7 NI_7 NS_1090 0 -2.6552915144783717e-06
GC_7_1091 b_7 NI_7 NS_1091 0 4.5743593691778643e-06
GC_7_1092 b_7 NI_7 NS_1092 0 -4.2831838769972379e-07
GC_7_1093 b_7 NI_7 NS_1093 0 -7.3616119657349265e-06
GC_7_1094 b_7 NI_7 NS_1094 0 -7.5350577766040880e-06
GC_7_1095 b_7 NI_7 NS_1095 0 -2.4585706000201301e-07
GC_7_1096 b_7 NI_7 NS_1096 0 -1.3969578215031932e-06
GC_7_1097 b_7 NI_7 NS_1097 0 -5.8994749214835779e-06
GC_7_1098 b_7 NI_7 NS_1098 0 2.4069591611359547e-06
GC_7_1099 b_7 NI_7 NS_1099 0 5.0799358816161482e-06
GC_7_1100 b_7 NI_7 NS_1100 0 -5.0478327027837558e-06
GC_7_1101 b_7 NI_7 NS_1101 0 -1.6513908413215353e-05
GC_7_1102 b_7 NI_7 NS_1102 0 4.9731464227449840e-06
GC_7_1103 b_7 NI_7 NS_1103 0 -1.2104003908863980e-06
GC_7_1104 b_7 NI_7 NS_1104 0 7.3647401393215794e-06
GC_7_1105 b_7 NI_7 NS_1105 0 -6.6058683428436764e-06
GC_7_1106 b_7 NI_7 NS_1106 0 -3.9243501578819963e-06
GC_7_1107 b_7 NI_7 NS_1107 0 -3.2757672774511088e-06
GC_7_1108 b_7 NI_7 NS_1108 0 8.1805471506399537e-06
GC_7_1109 b_7 NI_7 NS_1109 0 -1.4123073940839566e-06
GC_7_1110 b_7 NI_7 NS_1110 0 -3.8938058231810697e-06
GC_7_1111 b_7 NI_7 NS_1111 0 -3.9336561432386659e-06
GC_7_1112 b_7 NI_7 NS_1112 0 1.1229367990804589e-05
GC_7_1113 b_7 NI_7 NS_1113 0 -1.1559740002342472e-07
GC_7_1114 b_7 NI_7 NS_1114 0 7.5148536290910078e-06
GC_7_1115 b_7 NI_7 NS_1115 0 -3.6231367223372806e-06
GC_7_1116 b_7 NI_7 NS_1116 0 1.5253185900289507e-06
GC_7_1117 b_7 NI_7 NS_1117 0 -4.3432149261770756e-07
GC_7_1118 b_7 NI_7 NS_1118 0 8.2698466722233608e-06
GC_7_1119 b_7 NI_7 NS_1119 0 -5.5569844576101104e-07
GC_7_1120 b_7 NI_7 NS_1120 0 2.2142469182767329e-06
GC_7_1121 b_7 NI_7 NS_1121 0 -2.3137636054259028e-06
GC_7_1122 b_7 NI_7 NS_1122 0 8.3308447343469453e-06
GC_7_1123 b_7 NI_7 NS_1123 0 6.0315795096390426e-07
GC_7_1124 b_7 NI_7 NS_1124 0 9.9619461899240410e-06
GC_7_1125 b_7 NI_7 NS_1125 0 -6.8797673852283587e-07
GC_7_1126 b_7 NI_7 NS_1126 0 8.8045970442275277e-06
GC_7_1127 b_7 NI_7 NS_1127 0 -1.2376794038065644e-06
GC_7_1128 b_7 NI_7 NS_1128 0 4.0443129561998239e-06
GC_7_1129 b_7 NI_7 NS_1129 0 1.2364271983300757e-06
GC_7_1130 b_7 NI_7 NS_1130 0 1.2169058445979296e-05
GC_7_1131 b_7 NI_7 NS_1131 0 1.8569135898999737e-05
GC_7_1132 b_7 NI_7 NS_1132 0 1.6970585799512243e-05
GC_7_1133 b_7 NI_7 NS_1133 0 4.9794873003784954e-06
GC_7_1134 b_7 NI_7 NS_1134 0 7.7555437561003196e-06
GC_7_1135 b_7 NI_7 NS_1135 0 1.0278856022417668e-05
GC_7_1136 b_7 NI_7 NS_1136 0 3.8769448248975357e-06
GC_7_1137 b_7 NI_7 NS_1137 0 6.7691301721138843e-06
GC_7_1138 b_7 NI_7 NS_1138 0 1.0908029076929664e-05
GC_7_1139 b_7 NI_7 NS_1139 0 3.3282822979810613e-05
GC_7_1140 b_7 NI_7 NS_1140 0 -6.0912170509587346e-06
GC_7_1141 b_7 NI_7 NS_1141 0 8.1276576973491634e-06
GC_7_1142 b_7 NI_7 NS_1142 0 3.4130678633804635e-06
GC_7_1143 b_7 NI_7 NS_1143 0 1.1915390989017211e-05
GC_7_1144 b_7 NI_7 NS_1144 0 -1.0252449304110118e-05
GC_7_1145 b_7 NI_7 NS_1145 0 1.0732664768642318e-05
GC_7_1146 b_7 NI_7 NS_1146 0 6.4703327354191275e-06
GC_7_1147 b_7 NI_7 NS_1147 0 1.6861236152848839e-05
GC_7_1148 b_7 NI_7 NS_1148 0 -3.0702836787832926e-05
GC_7_1149 b_7 NI_7 NS_1149 0 8.0800696456886783e-06
GC_7_1150 b_7 NI_7 NS_1150 0 -2.9184897481682489e-06
GC_7_1151 b_7 NI_7 NS_1151 0 -3.2230745204389401e-06
GC_7_1152 b_7 NI_7 NS_1152 0 -1.6215595630258714e-05
GC_7_1153 b_7 NI_7 NS_1153 0 1.1759403285943833e-05
GC_7_1154 b_7 NI_7 NS_1154 0 -1.5875024335789592e-06
GC_7_1155 b_7 NI_7 NS_1155 0 -1.2692758148261150e-05
GC_7_1156 b_7 NI_7 NS_1156 0 -2.5024419936263744e-05
GC_7_1157 b_7 NI_7 NS_1157 0 -1.5671325212595702e-07
GC_7_1158 b_7 NI_7 NS_1158 0 -6.5860906053057561e-06
GC_7_1159 b_7 NI_7 NS_1159 0 -9.5588616820519839e-06
GC_7_1160 b_7 NI_7 NS_1160 0 -2.6136598800748877e-06
GC_7_1161 b_7 NI_7 NS_1161 0 1.0214438537466626e-10
GC_7_1162 b_7 NI_7 NS_1162 0 4.7347223125480885e-11
GC_7_1163 b_7 NI_7 NS_1163 0 1.4916303707474074e-06
GC_7_1164 b_7 NI_7 NS_1164 0 -4.6685481578400495e-06
GC_7_1165 b_7 NI_7 NS_1165 0 -1.3624857473710703e-06
GC_7_1166 b_7 NI_7 NS_1166 0 -1.3366695079904711e-06
GC_7_1167 b_7 NI_7 NS_1167 0 -4.8492451210010704e-06
GC_7_1168 b_7 NI_7 NS_1168 0 -9.9200203491614105e-07
GC_7_1169 b_7 NI_7 NS_1169 0 -1.1407274613556098e-06
GC_7_1170 b_7 NI_7 NS_1170 0 -2.7064160585852566e-06
GC_7_1171 b_7 NI_7 NS_1171 0 -9.9964601441018025e-06
GC_7_1172 b_7 NI_7 NS_1172 0 -4.0330070143323939e-06
GC_7_1173 b_7 NI_7 NS_1173 0 6.6625988499472914e-09
GC_7_1174 b_7 NI_7 NS_1174 0 5.4065805071009712e-09
GC_7_1175 b_7 NI_7 NS_1175 0 1.7627794378037294e-06
GC_7_1176 b_7 NI_7 NS_1176 0 4.8652326875520583e-07
GC_7_1177 b_7 NI_7 NS_1177 0 -1.6104309019592795e-06
GC_7_1178 b_7 NI_7 NS_1178 0 3.2255924130736961e-06
GC_7_1179 b_7 NI_7 NS_1179 0 -8.2940680221948207e-07
GC_7_1180 b_7 NI_7 NS_1180 0 7.0026344314977093e-07
GC_7_1181 b_7 NI_7 NS_1181 0 -7.6527107816609632e-06
GC_7_1182 b_7 NI_7 NS_1182 0 5.4683776836790579e-07
GC_7_1183 b_7 NI_7 NS_1183 0 -2.2162358769792994e-06
GC_7_1184 b_7 NI_7 NS_1184 0 2.0035048378365251e-06
GC_7_1185 b_7 NI_7 NS_1185 0 -2.0640123859388496e-06
GC_7_1186 b_7 NI_7 NS_1186 0 1.9717473550805969e-06
GC_7_1187 b_7 NI_7 NS_1187 0 1.2832744836875838e-06
GC_7_1188 b_7 NI_7 NS_1188 0 2.8361931164707395e-06
GC_7_1189 b_7 NI_7 NS_1189 0 -1.5116974816513267e-04
GC_7_1190 b_7 NI_7 NS_1190 0 3.7546613985139118e-11
GC_7_1191 b_7 NI_7 NS_1191 0 1.7615049595068684e-11
GC_7_1192 b_7 NI_7 NS_1192 0 8.7388023639138293e-10
GC_7_1193 b_7 NI_7 NS_1193 0 -2.3302531617206880e-06
GC_7_1194 b_7 NI_7 NS_1194 0 -1.6501624994826903e-06
GC_7_1195 b_7 NI_7 NS_1195 0 1.4540859300646731e-06
GC_7_1196 b_7 NI_7 NS_1196 0 3.8965294260650798e-06
GC_7_1197 b_7 NI_7 NS_1197 0 2.9654313717934649e-06
GC_7_1198 b_7 NI_7 NS_1198 0 5.4214117431294718e-06
GC_7_1199 b_7 NI_7 NS_1199 0 5.3772066465548715e-06
GC_7_1200 b_7 NI_7 NS_1200 0 -8.4804855966351445e-06
GC_7_1201 b_7 NI_7 NS_1201 0 -2.2508555118987447e-06
GC_7_1202 b_7 NI_7 NS_1202 0 -1.2662152480601633e-05
GC_7_1203 b_7 NI_7 NS_1203 0 -3.7274336870485032e-06
GC_7_1204 b_7 NI_7 NS_1204 0 2.7451157872100370e-06
GC_7_1205 b_7 NI_7 NS_1205 0 4.4942029329419126e-06
GC_7_1206 b_7 NI_7 NS_1206 0 1.5804116041397220e-06
GC_7_1207 b_7 NI_7 NS_1207 0 8.5384649794823791e-06
GC_7_1208 b_7 NI_7 NS_1208 0 -3.8252125141911908e-05
GC_7_1209 b_7 NI_7 NS_1209 0 -4.2843638902332613e-05
GC_7_1210 b_7 NI_7 NS_1210 0 -1.4538419196101190e-06
GC_7_1211 b_7 NI_7 NS_1211 0 -1.4647394672845111e-05
GC_7_1212 b_7 NI_7 NS_1212 0 -8.2775789683787145e-06
GC_7_1213 b_7 NI_7 NS_1213 0 -7.0243590072052186e-05
GC_7_1214 b_7 NI_7 NS_1214 0 7.5186050112088342e-05
GC_7_1215 b_7 NI_7 NS_1215 0 4.8693965777547285e-06
GC_7_1216 b_7 NI_7 NS_1216 0 1.3024168574190676e-05
GC_7_1217 b_7 NI_7 NS_1217 0 6.5219907725124233e-05
GC_7_1218 b_7 NI_7 NS_1218 0 1.2202210589645455e-04
GC_7_1219 b_7 NI_7 NS_1219 0 -2.7571959546207018e-07
GC_7_1220 b_7 NI_7 NS_1220 0 -3.7368893097601352e-05
GC_7_1221 b_7 NI_7 NS_1221 0 1.6806415000677518e-05
GC_7_1222 b_7 NI_7 NS_1222 0 4.1840187991344472e-06
GC_7_1223 b_7 NI_7 NS_1223 0 2.5159053641993270e-05
GC_7_1224 b_7 NI_7 NS_1224 0 -3.0985798306936698e-05
GC_7_1225 b_7 NI_7 NS_1225 0 -8.5163888435333739e-06
GC_7_1226 b_7 NI_7 NS_1226 0 -2.5733018738001182e-06
GC_7_1227 b_7 NI_7 NS_1227 0 -8.0803339051272540e-06
GC_7_1228 b_7 NI_7 NS_1228 0 2.4256733965716711e-05
GC_7_1229 b_7 NI_7 NS_1229 0 6.0403015165832173e-06
GC_7_1230 b_7 NI_7 NS_1230 0 8.3879398679446879e-06
GC_7_1231 b_7 NI_7 NS_1231 0 5.7351158412203006e-05
GC_7_1232 b_7 NI_7 NS_1232 0 2.3736636305631379e-05
GC_7_1233 b_7 NI_7 NS_1233 0 3.5347113435515709e-06
GC_7_1234 b_7 NI_7 NS_1234 0 -1.2244131266048427e-05
GC_7_1235 b_7 NI_7 NS_1235 0 -7.4155436410681434e-08
GC_7_1236 b_7 NI_7 NS_1236 0 -1.3740072243584064e-06
GC_7_1237 b_7 NI_7 NS_1237 0 7.1802710929492608e-06
GC_7_1238 b_7 NI_7 NS_1238 0 2.7779090491769501e-06
GC_7_1239 b_7 NI_7 NS_1239 0 4.2417148439695124e-05
GC_7_1240 b_7 NI_7 NS_1240 0 -1.9012479449699167e-05
GC_7_1241 b_7 NI_7 NS_1241 0 -2.5057099833908493e-06
GC_7_1242 b_7 NI_7 NS_1242 0 -7.6313015071477028e-06
GC_7_1243 b_7 NI_7 NS_1243 0 -2.8031655036561363e-06
GC_7_1244 b_7 NI_7 NS_1244 0 1.0883302356709432e-06
GC_7_1245 b_7 NI_7 NS_1245 0 9.8314153433488927e-06
GC_7_1246 b_7 NI_7 NS_1246 0 2.5417452190593787e-06
GC_7_1247 b_7 NI_7 NS_1247 0 2.2416083247945541e-05
GC_7_1248 b_7 NI_7 NS_1248 0 -3.3139468859819468e-05
GC_7_1249 b_7 NI_7 NS_1249 0 -5.7255560835556010e-06
GC_7_1250 b_7 NI_7 NS_1250 0 -4.2016003516442760e-06
GC_7_1251 b_7 NI_7 NS_1251 0 -8.8988093342705095e-07
GC_7_1252 b_7 NI_7 NS_1252 0 4.2524272336476864e-06
GC_7_1253 b_7 NI_7 NS_1253 0 1.2480231037941978e-05
GC_7_1254 b_7 NI_7 NS_1254 0 -2.7947779116093408e-07
GC_7_1255 b_7 NI_7 NS_1255 0 4.7407457181550132e-07
GC_7_1256 b_7 NI_7 NS_1256 0 -3.2834917606565192e-05
GC_7_1257 b_7 NI_7 NS_1257 0 -6.9267934891142545e-06
GC_7_1258 b_7 NI_7 NS_1258 0 4.0680066469883679e-07
GC_7_1259 b_7 NI_7 NS_1259 0 3.8410670811787340e-06
GC_7_1260 b_7 NI_7 NS_1260 0 3.5676048903140439e-06
GC_7_1261 b_7 NI_7 NS_1261 0 1.4108535928568072e-05
GC_7_1262 b_7 NI_7 NS_1262 0 -6.6872350694861107e-06
GC_7_1263 b_7 NI_7 NS_1263 0 -1.5604809407279362e-05
GC_7_1264 b_7 NI_7 NS_1264 0 -1.9003792469655514e-05
GC_7_1265 b_7 NI_7 NS_1265 0 -2.9951985159487196e-06
GC_7_1266 b_7 NI_7 NS_1266 0 5.1042289840157399e-06
GC_7_1267 b_7 NI_7 NS_1267 0 4.2096659402540220e-06
GC_7_1268 b_7 NI_7 NS_1268 0 -1.8810295851789860e-06
GC_7_1269 b_7 NI_7 NS_1269 0 -2.7916694458960362e-11
GC_7_1270 b_7 NI_7 NS_1270 0 5.8150969482684282e-12
GC_7_1271 b_7 NI_7 NS_1271 0 4.8699137906540009e-06
GC_7_1272 b_7 NI_7 NS_1272 0 -1.1668169730033340e-05
GC_7_1273 b_7 NI_7 NS_1273 0 -5.0904552801596064e-07
GC_7_1274 b_7 NI_7 NS_1274 0 2.7992316332495055e-06
GC_7_1275 b_7 NI_7 NS_1275 0 2.3509281489058503e-06
GC_7_1276 b_7 NI_7 NS_1276 0 -1.5716763985951608e-06
GC_7_1277 b_7 NI_7 NS_1277 0 2.1314589935884512e-06
GC_7_1278 b_7 NI_7 NS_1278 0 -9.8974506031493253e-06
GC_7_1279 b_7 NI_7 NS_1279 0 -1.0613671233307990e-05
GC_7_1280 b_7 NI_7 NS_1280 0 -3.5263815370770148e-06
GC_7_1281 b_7 NI_7 NS_1281 0 -2.3906789558815852e-10
GC_7_1282 b_7 NI_7 NS_1282 0 4.4559234698778725e-10
GC_7_1283 b_7 NI_7 NS_1283 0 -9.1766890084382757e-06
GC_7_1284 b_7 NI_7 NS_1284 0 -5.6138461064269551e-06
GC_7_1285 b_7 NI_7 NS_1285 0 1.9952308960928147e-06
GC_7_1286 b_7 NI_7 NS_1286 0 -6.7132345849226938e-06
GC_7_1287 b_7 NI_7 NS_1287 0 -3.3605892940498525e-06
GC_7_1288 b_7 NI_7 NS_1288 0 -1.7941587249152314e-07
GC_7_1289 b_7 NI_7 NS_1289 0 -8.5928704864844082e-06
GC_7_1290 b_7 NI_7 NS_1290 0 5.9552771838913034e-07
GC_7_1291 b_7 NI_7 NS_1291 0 2.6078614450589012e-06
GC_7_1292 b_7 NI_7 NS_1292 0 2.8392946982038250e-06
GC_7_1293 b_7 NI_7 NS_1293 0 9.9242063428482553e-07
GC_7_1294 b_7 NI_7 NS_1294 0 -3.6889661768747719e-06
GC_7_1295 b_7 NI_7 NS_1295 0 -5.4153669596692585e-06
GC_7_1296 b_7 NI_7 NS_1296 0 -4.2328094175612535e-06
GD_7_1 b_7 NI_7 NA_1 0 -2.6035567090653045e-06
GD_7_2 b_7 NI_7 NA_2 0 1.1368429267067173e-05
GD_7_3 b_7 NI_7 NA_3 0 -6.7345348115469480e-07
GD_7_4 b_7 NI_7 NA_4 0 1.6002508354826357e-05
GD_7_5 b_7 NI_7 NA_5 0 1.0577033559931800e-02
GD_7_6 b_7 NI_7 NA_6 0 -1.1498023080688546e-03
GD_7_7 b_7 NI_7 NA_7 0 -1.1040267719203507e-02
GD_7_8 b_7 NI_7 NA_8 0 -4.9039720174917948e-03
GD_7_9 b_7 NI_7 NA_9 0 2.6301362904956894e-05
GD_7_10 b_7 NI_7 NA_10 0 1.0461289839228412e-04
GD_7_11 b_7 NI_7 NA_11 0 2.6760858875997496e-06
GD_7_12 b_7 NI_7 NA_12 0 1.9066309295319530e-05
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 -8.9827477565911261e-05
GC_8_2 b_8 NI_8 NS_2 0 3.3242005650471814e-12
GC_8_3 b_8 NI_8 NS_3 0 -4.3152827204773593e-11
GC_8_4 b_8 NI_8 NS_4 0 3.0281097488476864e-10
GC_8_5 b_8 NI_8 NS_5 0 -1.5652915128417047e-06
GC_8_6 b_8 NI_8 NS_6 0 -1.5563384536993090e-06
GC_8_7 b_8 NI_8 NS_7 0 9.4716797769954153e-07
GC_8_8 b_8 NI_8 NS_8 0 7.1437250210312804e-07
GC_8_9 b_8 NI_8 NS_9 0 -2.7263894436313070e-06
GC_8_10 b_8 NI_8 NS_10 0 3.0058194397671323e-06
GC_8_11 b_8 NI_8 NS_11 0 -3.0650239933520425e-06
GC_8_12 b_8 NI_8 NS_12 0 -2.5788292223348386e-06
GC_8_13 b_8 NI_8 NS_13 0 1.4936491761315348e-06
GC_8_14 b_8 NI_8 NS_14 0 1.1481036062095533e-07
GC_8_15 b_8 NI_8 NS_15 0 -1.6611509913478407e-06
GC_8_16 b_8 NI_8 NS_16 0 1.7822155953479825e-06
GC_8_17 b_8 NI_8 NS_17 0 8.5990611832396805e-07
GC_8_18 b_8 NI_8 NS_18 0 4.1352253866174127e-06
GC_8_19 b_8 NI_8 NS_19 0 -4.3810515542332666e-06
GC_8_20 b_8 NI_8 NS_20 0 -1.9846150037142261e-06
GC_8_21 b_8 NI_8 NS_21 0 2.4929788910399087e-06
GC_8_22 b_8 NI_8 NS_22 0 -1.8455358161143965e-06
GC_8_23 b_8 NI_8 NS_23 0 -1.1634615259156321e-06
GC_8_24 b_8 NI_8 NS_24 0 3.2977044769439517e-06
GC_8_25 b_8 NI_8 NS_25 0 -8.1357990646615057e-06
GC_8_26 b_8 NI_8 NS_26 0 1.1093579496551894e-05
GC_8_27 b_8 NI_8 NS_27 0 1.2697839722840948e-06
GC_8_28 b_8 NI_8 NS_28 0 -1.6862494691287143e-06
GC_8_29 b_8 NI_8 NS_29 0 9.8771721882999585e-06
GC_8_30 b_8 NI_8 NS_30 0 1.6972996785253655e-05
GC_8_31 b_8 NI_8 NS_31 0 -7.1199368208360647e-07
GC_8_32 b_8 NI_8 NS_32 0 -4.4201306239547393e-07
GC_8_33 b_8 NI_8 NS_33 0 4.0869273386203470e-07
GC_8_34 b_8 NI_8 NS_34 0 -1.4042432752672766e-06
GC_8_35 b_8 NI_8 NS_35 0 6.8711715976939374e-06
GC_8_36 b_8 NI_8 NS_36 0 -1.2535127521387594e-07
GC_8_37 b_8 NI_8 NS_37 0 7.0587983537688731e-07
GC_8_38 b_8 NI_8 NS_38 0 3.0247942221758663e-06
GC_8_39 b_8 NI_8 NS_39 0 5.1850942183359399e-07
GC_8_40 b_8 NI_8 NS_40 0 2.8703461043321816e-06
GC_8_41 b_8 NI_8 NS_41 0 1.1686954045464061e-06
GC_8_42 b_8 NI_8 NS_42 0 -1.4312838563183692e-06
GC_8_43 b_8 NI_8 NS_43 0 9.2306171473456087e-06
GC_8_44 b_8 NI_8 NS_44 0 5.0868160435306424e-06
GC_8_45 b_8 NI_8 NS_45 0 5.3876564637369625e-07
GC_8_46 b_8 NI_8 NS_46 0 1.1688122885922442e-06
GC_8_47 b_8 NI_8 NS_47 0 4.7182574069914724e-08
GC_8_48 b_8 NI_8 NS_48 0 4.6163602122646449e-07
GC_8_49 b_8 NI_8 NS_49 0 1.2781466762017103e-06
GC_8_50 b_8 NI_8 NS_50 0 -8.5245171853529547e-07
GC_8_51 b_8 NI_8 NS_51 0 9.0033505219645287e-06
GC_8_52 b_8 NI_8 NS_52 0 7.1340339607380236e-07
GC_8_53 b_8 NI_8 NS_53 0 8.3038630242768916e-07
GC_8_54 b_8 NI_8 NS_54 0 1.4741778667541672e-06
GC_8_55 b_8 NI_8 NS_55 0 1.0390717779819093e-06
GC_8_56 b_8 NI_8 NS_56 0 6.2172831354114025e-07
GC_8_57 b_8 NI_8 NS_57 0 1.3551398390147330e-06
GC_8_58 b_8 NI_8 NS_58 0 -9.5010374995671753e-07
GC_8_59 b_8 NI_8 NS_59 0 7.9167174348644161e-06
GC_8_60 b_8 NI_8 NS_60 0 -2.0394120708880360e-06
GC_8_61 b_8 NI_8 NS_61 0 1.1753942484714661e-06
GC_8_62 b_8 NI_8 NS_62 0 1.5633821695218288e-06
GC_8_63 b_8 NI_8 NS_63 0 1.6188837427560199e-06
GC_8_64 b_8 NI_8 NS_64 0 -2.2250595761041297e-07
GC_8_65 b_8 NI_8 NS_65 0 1.3149938865425409e-06
GC_8_66 b_8 NI_8 NS_66 0 -9.9060639467716218e-07
GC_8_67 b_8 NI_8 NS_67 0 5.7974590961176807e-06
GC_8_68 b_8 NI_8 NS_68 0 -3.8075830686117384e-06
GC_8_69 b_8 NI_8 NS_69 0 1.8131055595039410e-06
GC_8_70 b_8 NI_8 NS_70 0 1.4425427048956999e-06
GC_8_71 b_8 NI_8 NS_71 0 1.1283305302398639e-06
GC_8_72 b_8 NI_8 NS_72 0 -1.3977655145668385e-06
GC_8_73 b_8 NI_8 NS_73 0 1.4102950324081137e-06
GC_8_74 b_8 NI_8 NS_74 0 -1.1060954032069588e-06
GC_8_75 b_8 NI_8 NS_75 0 2.9944002848615209e-06
GC_8_76 b_8 NI_8 NS_76 0 -4.1483176038548089e-06
GC_8_77 b_8 NI_8 NS_77 0 2.2296545952858967e-06
GC_8_78 b_8 NI_8 NS_78 0 3.1298443969812815e-07
GC_8_79 b_8 NI_8 NS_79 0 -3.1154206363302453e-07
GC_8_80 b_8 NI_8 NS_80 0 -1.1925988681398563e-06
GC_8_81 b_8 NI_8 NS_81 0 2.5423220965464837e-11
GC_8_82 b_8 NI_8 NS_82 0 -4.1101297741697924e-11
GC_8_83 b_8 NI_8 NS_83 0 8.0347227619132519e-07
GC_8_84 b_8 NI_8 NS_84 0 -1.5695291248422986e-06
GC_8_85 b_8 NI_8 NS_85 0 1.2661365991387119e-06
GC_8_86 b_8 NI_8 NS_86 0 2.2070188455484463e-07
GC_8_87 b_8 NI_8 NS_87 0 1.6021636243117797e-07
GC_8_88 b_8 NI_8 NS_88 0 -5.5094468347318413e-07
GC_8_89 b_8 NI_8 NS_89 0 5.5034027897380227e-07
GC_8_90 b_8 NI_8 NS_90 0 -8.6165058478781618e-07
GC_8_91 b_8 NI_8 NS_91 0 1.3129411429602754e-06
GC_8_92 b_8 NI_8 NS_92 0 -2.0695644791391218e-06
GC_8_93 b_8 NI_8 NS_93 0 4.8975006972119856e-10
GC_8_94 b_8 NI_8 NS_94 0 -1.2287919683883264e-09
GC_8_95 b_8 NI_8 NS_95 0 5.5017491809434667e-07
GC_8_96 b_8 NI_8 NS_96 0 -8.6030143423961329e-07
GC_8_97 b_8 NI_8 NS_97 0 7.1448037661488829e-07
GC_8_98 b_8 NI_8 NS_98 0 -9.5257238633543859e-07
GC_8_99 b_8 NI_8 NS_99 0 9.1157337373000175e-08
GC_8_100 b_8 NI_8 NS_100 0 4.9897436910693628e-08
GC_8_101 b_8 NI_8 NS_101 0 1.3758223413260241e-06
GC_8_102 b_8 NI_8 NS_102 0 -1.2408283157489187e-06
GC_8_103 b_8 NI_8 NS_103 0 1.6631097294172730e-06
GC_8_104 b_8 NI_8 NS_104 0 -3.1895780974394368e-07
GC_8_105 b_8 NI_8 NS_105 0 -2.4124578416145467e-07
GC_8_106 b_8 NI_8 NS_106 0 -7.4502378872088228e-07
GC_8_107 b_8 NI_8 NS_107 0 7.3810168609135753e-07
GC_8_108 b_8 NI_8 NS_108 0 2.9282298880966152e-07
GC_8_109 b_8 NI_8 NS_109 0 4.7667632269475806e-05
GC_8_110 b_8 NI_8 NS_110 0 7.4777264111531709e-12
GC_8_111 b_8 NI_8 NS_111 0 -1.8812330297467647e-11
GC_8_112 b_8 NI_8 NS_112 0 9.9179817694731620e-10
GC_8_113 b_8 NI_8 NS_113 0 -6.5157772919276652e-08
GC_8_114 b_8 NI_8 NS_114 0 2.4828596924332408e-07
GC_8_115 b_8 NI_8 NS_115 0 2.2372325303152989e-07
GC_8_116 b_8 NI_8 NS_116 0 4.0478121261771895e-07
GC_8_117 b_8 NI_8 NS_117 0 -1.7409009899152110e-07
GC_8_118 b_8 NI_8 NS_118 0 2.7593237182474479e-07
GC_8_119 b_8 NI_8 NS_119 0 7.2779057256869352e-07
GC_8_120 b_8 NI_8 NS_120 0 1.4717946334717668e-06
GC_8_121 b_8 NI_8 NS_121 0 1.0335877202586945e-06
GC_8_122 b_8 NI_8 NS_122 0 -4.2692940603476937e-07
GC_8_123 b_8 NI_8 NS_123 0 3.0382895555919639e-07
GC_8_124 b_8 NI_8 NS_124 0 9.1841932931212856e-07
GC_8_125 b_8 NI_8 NS_125 0 7.7986183201780100e-07
GC_8_126 b_8 NI_8 NS_126 0 -3.1608309715519218e-07
GC_8_127 b_8 NI_8 NS_127 0 4.3388029694833279e-06
GC_8_128 b_8 NI_8 NS_128 0 1.5030456575535356e-06
GC_8_129 b_8 NI_8 NS_129 0 -1.5184038384996943e-06
GC_8_130 b_8 NI_8 NS_130 0 -3.5718099898283821e-06
GC_8_131 b_8 NI_8 NS_131 0 2.4364831101187593e-07
GC_8_132 b_8 NI_8 NS_132 0 1.5787640513570830e-06
GC_8_133 b_8 NI_8 NS_133 0 3.1022177059500977e-06
GC_8_134 b_8 NI_8 NS_134 0 -4.6733355551125369e-06
GC_8_135 b_8 NI_8 NS_135 0 -7.4687476663351928e-07
GC_8_136 b_8 NI_8 NS_136 0 5.6934744720914763e-07
GC_8_137 b_8 NI_8 NS_137 0 5.7285804037791956e-06
GC_8_138 b_8 NI_8 NS_138 0 -5.7347849558217713e-06
GC_8_139 b_8 NI_8 NS_139 0 -3.3214859844983585e-06
GC_8_140 b_8 NI_8 NS_140 0 1.7576635033084148e-06
GC_8_141 b_8 NI_8 NS_141 0 8.8321671233361232e-07
GC_8_142 b_8 NI_8 NS_142 0 1.2580676533736260e-06
GC_8_143 b_8 NI_8 NS_143 0 1.6925155551497138e-06
GC_8_144 b_8 NI_8 NS_144 0 -4.0851793568462532e-06
GC_8_145 b_8 NI_8 NS_145 0 6.1027160316104840e-07
GC_8_146 b_8 NI_8 NS_146 0 2.1452820216946979e-07
GC_8_147 b_8 NI_8 NS_147 0 2.5203328064130463e-07
GC_8_148 b_8 NI_8 NS_148 0 -4.0638362763948222e-06
GC_8_149 b_8 NI_8 NS_149 0 -1.5631460282022353e-07
GC_8_150 b_8 NI_8 NS_150 0 1.7770659249180450e-07
GC_8_151 b_8 NI_8 NS_151 0 4.7896805006934913e-06
GC_8_152 b_8 NI_8 NS_152 0 -6.3217697871400315e-06
GC_8_153 b_8 NI_8 NS_153 0 -1.7965573698903114e-06
GC_8_154 b_8 NI_8 NS_154 0 -1.3136931980465541e-06
GC_8_155 b_8 NI_8 NS_155 0 1.3999546101867824e-06
GC_8_156 b_8 NI_8 NS_156 0 -1.1893439469619954e-06
GC_8_157 b_8 NI_8 NS_157 0 4.3391054957203330e-07
GC_8_158 b_8 NI_8 NS_158 0 -2.1052475281099815e-06
GC_8_159 b_8 NI_8 NS_159 0 -1.3418247478405380e-06
GC_8_160 b_8 NI_8 NS_160 0 -1.1874133675675553e-05
GC_8_161 b_8 NI_8 NS_161 0 -2.2438006008028916e-06
GC_8_162 b_8 NI_8 NS_162 0 -1.7319021262954637e-06
GC_8_163 b_8 NI_8 NS_163 0 -2.3535062918731839e-06
GC_8_164 b_8 NI_8 NS_164 0 -4.0395592190843313e-06
GC_8_165 b_8 NI_8 NS_165 0 -1.4505101052171528e-06
GC_8_166 b_8 NI_8 NS_166 0 -2.4379032007769178e-06
GC_8_167 b_8 NI_8 NS_167 0 -1.0686776675526253e-05
GC_8_168 b_8 NI_8 NS_168 0 -7.2206318043142947e-06
GC_8_169 b_8 NI_8 NS_169 0 -3.1790011965332975e-06
GC_8_170 b_8 NI_8 NS_170 0 -8.7765646518000480e-07
GC_8_171 b_8 NI_8 NS_171 0 -5.7557871294543013e-06
GC_8_172 b_8 NI_8 NS_172 0 -4.1572902406081303e-07
GC_8_173 b_8 NI_8 NS_173 0 -3.1006023500652938e-06
GC_8_174 b_8 NI_8 NS_174 0 -1.7564430058366173e-06
GC_8_175 b_8 NI_8 NS_175 0 -1.0631076197779632e-05
GC_8_176 b_8 NI_8 NS_176 0 3.2969262070772249e-06
GC_8_177 b_8 NI_8 NS_177 0 -3.6194758798094701e-06
GC_8_178 b_8 NI_8 NS_178 0 8.1861918120580391e-07
GC_8_179 b_8 NI_8 NS_179 0 -2.8825397396461652e-06
GC_8_180 b_8 NI_8 NS_180 0 3.9154067911771946e-06
GC_8_181 b_8 NI_8 NS_181 0 -4.3323123751007068e-06
GC_8_182 b_8 NI_8 NS_182 0 1.7065232408438311e-07
GC_8_183 b_8 NI_8 NS_183 0 -1.8686334012278774e-06
GC_8_184 b_8 NI_8 NS_184 0 7.2154269506615735e-06
GC_8_185 b_8 NI_8 NS_185 0 -1.5642572413585173e-06
GC_8_186 b_8 NI_8 NS_186 0 2.7942571527040632e-06
GC_8_187 b_8 NI_8 NS_187 0 9.2411103741672378e-07
GC_8_188 b_8 NI_8 NS_188 0 1.8150574412506581e-06
GC_8_189 b_8 NI_8 NS_189 0 -3.0215514610862273e-11
GC_8_190 b_8 NI_8 NS_190 0 -3.9734410970963791e-12
GC_8_191 b_8 NI_8 NS_191 0 -1.7144583806931508e-06
GC_8_192 b_8 NI_8 NS_192 0 2.1408166427240492e-06
GC_8_193 b_8 NI_8 NS_193 0 -3.2467229274689556e-07
GC_8_194 b_8 NI_8 NS_194 0 1.0491055111534087e-06
GC_8_195 b_8 NI_8 NS_195 0 1.4393956449961329e-07
GC_8_196 b_8 NI_8 NS_196 0 6.2162088765516036e-07
GC_8_197 b_8 NI_8 NS_197 0 -1.0469793175834481e-06
GC_8_198 b_8 NI_8 NS_198 0 1.2713193869565789e-06
GC_8_199 b_8 NI_8 NS_199 0 9.7964309572781799e-07
GC_8_200 b_8 NI_8 NS_200 0 1.8202533537832965e-06
GC_8_201 b_8 NI_8 NS_201 0 -1.5166092414231499e-09
GC_8_202 b_8 NI_8 NS_202 0 -7.8069319230606050e-10
GC_8_203 b_8 NI_8 NS_203 0 -4.8493305091404293e-07
GC_8_204 b_8 NI_8 NS_204 0 -2.7294816345482374e-08
GC_8_205 b_8 NI_8 NS_205 0 -3.1063966726438798e-07
GC_8_206 b_8 NI_8 NS_206 0 1.7482712986492983e-07
GC_8_207 b_8 NI_8 NS_207 0 -5.5091838387353150e-07
GC_8_208 b_8 NI_8 NS_208 0 1.5193412401346080e-07
GC_8_209 b_8 NI_8 NS_209 0 6.6426780590835902e-07
GC_8_210 b_8 NI_8 NS_210 0 8.1167763052997333e-07
GC_8_211 b_8 NI_8 NS_211 0 2.1767294518340445e-07
GC_8_212 b_8 NI_8 NS_212 0 6.9613020287924208e-07
GC_8_213 b_8 NI_8 NS_213 0 1.1062253611695690e-08
GC_8_214 b_8 NI_8 NS_214 0 -1.3787271269862562e-07
GC_8_215 b_8 NI_8 NS_215 0 -3.4802846365162224e-07
GC_8_216 b_8 NI_8 NS_216 0 2.9432596662741921e-07
GC_8_217 b_8 NI_8 NS_217 0 -1.4436792034942754e-04
GC_8_218 b_8 NI_8 NS_218 0 3.3291263638535018e-11
GC_8_219 b_8 NI_8 NS_219 0 3.9883323515726886e-11
GC_8_220 b_8 NI_8 NS_220 0 9.0899662366808083e-10
GC_8_221 b_8 NI_8 NS_221 0 -2.1101234913528491e-06
GC_8_222 b_8 NI_8 NS_222 0 -1.6555661824002921e-06
GC_8_223 b_8 NI_8 NS_223 0 1.8946752501709343e-06
GC_8_224 b_8 NI_8 NS_224 0 3.8512532432831858e-06
GC_8_225 b_8 NI_8 NS_225 0 3.3113080539623584e-06
GC_8_226 b_8 NI_8 NS_226 0 4.9314976659244260e-06
GC_8_227 b_8 NI_8 NS_227 0 5.8707439286202048e-06
GC_8_228 b_8 NI_8 NS_228 0 -9.1115038491762851e-06
GC_8_229 b_8 NI_8 NS_229 0 -2.5610765229387163e-06
GC_8_230 b_8 NI_8 NS_230 0 -1.3919643302191962e-05
GC_8_231 b_8 NI_8 NS_231 0 -3.5429763029552249e-06
GC_8_232 b_8 NI_8 NS_232 0 2.1898513222213143e-06
GC_8_233 b_8 NI_8 NS_233 0 3.6503654141512055e-06
GC_8_234 b_8 NI_8 NS_234 0 1.2870366555765749e-06
GC_8_235 b_8 NI_8 NS_235 0 8.0002037603203853e-06
GC_8_236 b_8 NI_8 NS_236 0 -3.9897461343154713e-05
GC_8_237 b_8 NI_8 NS_237 0 -4.4314026475122865e-05
GC_8_238 b_8 NI_8 NS_238 0 -9.3723455087355680e-07
GC_8_239 b_8 NI_8 NS_239 0 -1.4827663582030518e-05
GC_8_240 b_8 NI_8 NS_240 0 -8.5762708433326660e-06
GC_8_241 b_8 NI_8 NS_241 0 -7.2940073275988389e-05
GC_8_242 b_8 NI_8 NS_242 0 7.5520857811787011e-05
GC_8_243 b_8 NI_8 NS_243 0 4.6287942721334772e-06
GC_8_244 b_8 NI_8 NS_244 0 1.3120197965391489e-05
GC_8_245 b_8 NI_8 NS_245 0 6.2840577430081738e-05
GC_8_246 b_8 NI_8 NS_246 0 1.2320096567797510e-04
GC_8_247 b_8 NI_8 NS_247 0 3.6368155448938129e-07
GC_8_248 b_8 NI_8 NS_248 0 -3.7020253081094690e-05
GC_8_249 b_8 NI_8 NS_249 0 1.6508675420718759e-05
GC_8_250 b_8 NI_8 NS_250 0 3.9674561201948944e-06
GC_8_251 b_8 NI_8 NS_251 0 2.4448290583456979e-05
GC_8_252 b_8 NI_8 NS_252 0 -3.0458303807775926e-05
GC_8_253 b_8 NI_8 NS_253 0 -8.8966496737748901e-06
GC_8_254 b_8 NI_8 NS_254 0 -2.3403611160863872e-06
GC_8_255 b_8 NI_8 NS_255 0 -8.8833970207453705e-06
GC_8_256 b_8 NI_8 NS_256 0 2.5237539293250701e-05
GC_8_257 b_8 NI_8 NS_257 0 5.8265839490299515e-06
GC_8_258 b_8 NI_8 NS_258 0 8.4672013698882566e-06
GC_8_259 b_8 NI_8 NS_259 0 5.6328874977444184e-05
GC_8_260 b_8 NI_8 NS_260 0 2.4970425089962572e-05
GC_8_261 b_8 NI_8 NS_261 0 3.5274172437146670e-06
GC_8_262 b_8 NI_8 NS_262 0 -1.1687206780677178e-05
GC_8_263 b_8 NI_8 NS_263 0 -4.0890973922978874e-07
GC_8_264 b_8 NI_8 NS_264 0 -1.3155488169292618e-06
GC_8_265 b_8 NI_8 NS_265 0 6.8059207769344937e-06
GC_8_266 b_8 NI_8 NS_266 0 3.0643937484580538e-06
GC_8_267 b_8 NI_8 NS_267 0 4.1947955595114279e-05
GC_8_268 b_8 NI_8 NS_268 0 -1.7198990320837099e-05
GC_8_269 b_8 NI_8 NS_269 0 -2.5585877680052339e-06
GC_8_270 b_8 NI_8 NS_270 0 -7.0970249139496231e-06
GC_8_271 b_8 NI_8 NS_271 0 -3.0311225837043117e-06
GC_8_272 b_8 NI_8 NS_272 0 1.7555037782321981e-06
GC_8_273 b_8 NI_8 NS_273 0 9.5694291041690855e-06
GC_8_274 b_8 NI_8 NS_274 0 2.9162043472269061e-06
GC_8_275 b_8 NI_8 NS_275 0 2.2976242444743221e-05
GC_8_276 b_8 NI_8 NS_276 0 -3.1187887378373403e-05
GC_8_277 b_8 NI_8 NS_277 0 -5.6936489462956411e-06
GC_8_278 b_8 NI_8 NS_278 0 -3.6758075589723143e-06
GC_8_279 b_8 NI_8 NS_279 0 -5.6141031777975998e-07
GC_8_280 b_8 NI_8 NS_280 0 5.0284082927310699e-06
GC_8_281 b_8 NI_8 NS_281 0 1.2292664335172909e-05
GC_8_282 b_8 NI_8 NS_282 0 2.0426180932153119e-07
GC_8_283 b_8 NI_8 NS_283 0 1.9186210978126755e-06
GC_8_284 b_8 NI_8 NS_284 0 -3.1503873427529073e-05
GC_8_285 b_8 NI_8 NS_285 0 -6.7230948547608340e-06
GC_8_286 b_8 NI_8 NS_286 0 9.4617212355398266e-07
GC_8_287 b_8 NI_8 NS_287 0 4.5912205527027724e-06
GC_8_288 b_8 NI_8 NS_288 0 3.8667655021111777e-06
GC_8_289 b_8 NI_8 NS_289 0 1.4096640076457054e-05
GC_8_290 b_8 NI_8 NS_290 0 -6.0051890717049046e-06
GC_8_291 b_8 NI_8 NS_291 0 -1.3991427910446774e-05
GC_8_292 b_8 NI_8 NS_292 0 -1.8834468892604709e-05
GC_8_293 b_8 NI_8 NS_293 0 -2.5005397984537574e-06
GC_8_294 b_8 NI_8 NS_294 0 5.3958763419262372e-06
GC_8_295 b_8 NI_8 NS_295 0 4.6402124658436853e-06
GC_8_296 b_8 NI_8 NS_296 0 -2.0953729759096263e-06
GC_8_297 b_8 NI_8 NS_297 0 -1.4467203819336474e-11
GC_8_298 b_8 NI_8 NS_298 0 3.9854440640962562e-12
GC_8_299 b_8 NI_8 NS_299 0 5.2050960028510581e-06
GC_8_300 b_8 NI_8 NS_300 0 -1.1255676100881105e-05
GC_8_301 b_8 NI_8 NS_301 0 -2.6207483451538596e-07
GC_8_302 b_8 NI_8 NS_302 0 2.9240504789927813e-06
GC_8_303 b_8 NI_8 NS_303 0 2.6491355159381732e-06
GC_8_304 b_8 NI_8 NS_304 0 -1.6106328041309598e-06
GC_8_305 b_8 NI_8 NS_305 0 2.4311685242360061e-06
GC_8_306 b_8 NI_8 NS_306 0 -9.4257315562704093e-06
GC_8_307 b_8 NI_8 NS_307 0 -9.9191354997037469e-06
GC_8_308 b_8 NI_8 NS_308 0 -3.6953382402418912e-06
GC_8_309 b_8 NI_8 NS_309 0 3.1959576745307867e-10
GC_8_310 b_8 NI_8 NS_310 0 2.6398845668252210e-10
GC_8_311 b_8 NI_8 NS_311 0 -8.5810764932905832e-06
GC_8_312 b_8 NI_8 NS_312 0 -5.7196784681706965e-06
GC_8_313 b_8 NI_8 NS_313 0 2.2759196056090958e-06
GC_8_314 b_8 NI_8 NS_314 0 -6.4442966917237831e-06
GC_8_315 b_8 NI_8 NS_315 0 -3.0692684469155330e-06
GC_8_316 b_8 NI_8 NS_316 0 -1.3767749195140599e-07
GC_8_317 b_8 NI_8 NS_317 0 -7.9176037216204242e-06
GC_8_318 b_8 NI_8 NS_318 0 4.8798269273138725e-07
GC_8_319 b_8 NI_8 NS_319 0 3.0157302746342652e-06
GC_8_320 b_8 NI_8 NS_320 0 2.8670037214396178e-06
GC_8_321 b_8 NI_8 NS_321 0 1.2342815438852571e-06
GC_8_322 b_8 NI_8 NS_322 0 -3.9109860546643406e-06
GC_8_323 b_8 NI_8 NS_323 0 -4.8692369627726337e-06
GC_8_324 b_8 NI_8 NS_324 0 -3.9053575391677449e-06
GC_8_325 b_8 NI_8 NS_325 0 -2.7355549187334252e-05
GC_8_326 b_8 NI_8 NS_326 0 -9.2004689892783815e-13
GC_8_327 b_8 NI_8 NS_327 0 -2.3520845443555046e-10
GC_8_328 b_8 NI_8 NS_328 0 1.0469206551463542e-08
GC_8_329 b_8 NI_8 NS_329 0 7.2942593018628223e-07
GC_8_330 b_8 NI_8 NS_330 0 1.1057570962313732e-07
GC_8_331 b_8 NI_8 NS_331 0 3.2329357931047078e-06
GC_8_332 b_8 NI_8 NS_332 0 -1.3955668494514933e-06
GC_8_333 b_8 NI_8 NS_333 0 -2.7334272365116766e-06
GC_8_334 b_8 NI_8 NS_334 0 -2.8887393023741341e-06
GC_8_335 b_8 NI_8 NS_335 0 5.0379778691549045e-06
GC_8_336 b_8 NI_8 NS_336 0 -5.9339284499749817e-07
GC_8_337 b_8 NI_8 NS_337 0 -7.0890005853333228e-06
GC_8_338 b_8 NI_8 NS_338 0 -8.3126032004067880e-06
GC_8_339 b_8 NI_8 NS_339 0 8.1233385608381881e-08
GC_8_340 b_8 NI_8 NS_340 0 -1.6105146417779089e-06
GC_8_341 b_8 NI_8 NS_341 0 -6.1810005306529682e-06
GC_8_342 b_8 NI_8 NS_342 0 1.8479514206333340e-06
GC_8_343 b_8 NI_8 NS_343 0 5.4033090185818387e-06
GC_8_344 b_8 NI_8 NS_344 0 -6.0039260941607976e-06
GC_8_345 b_8 NI_8 NS_345 0 -1.7425745602737103e-05
GC_8_346 b_8 NI_8 NS_346 0 4.6515788429650981e-06
GC_8_347 b_8 NI_8 NS_347 0 -1.1775864511319057e-06
GC_8_348 b_8 NI_8 NS_348 0 7.0644007101828345e-06
GC_8_349 b_8 NI_8 NS_349 0 -7.5195207804442351e-06
GC_8_350 b_8 NI_8 NS_350 0 -4.7823985853109301e-06
GC_8_351 b_8 NI_8 NS_351 0 -3.4396136863063548e-06
GC_8_352 b_8 NI_8 NS_352 0 8.0393797142925918e-06
GC_8_353 b_8 NI_8 NS_353 0 -2.5304455328029584e-06
GC_8_354 b_8 NI_8 NS_354 0 -4.9642132651771849e-06
GC_8_355 b_8 NI_8 NS_355 0 -3.8886553429736438e-06
GC_8_356 b_8 NI_8 NS_356 0 1.1491298781604422e-05
GC_8_357 b_8 NI_8 NS_357 0 -1.9009364602597598e-07
GC_8_358 b_8 NI_8 NS_358 0 7.1731154155505965e-06
GC_8_359 b_8 NI_8 NS_359 0 -4.3615428081983640e-06
GC_8_360 b_8 NI_8 NS_360 0 1.1394837868455241e-06
GC_8_361 b_8 NI_8 NS_361 0 -6.9161337388884301e-07
GC_8_362 b_8 NI_8 NS_362 0 7.9938193940055170e-06
GC_8_363 b_8 NI_8 NS_363 0 -1.2344329094977882e-06
GC_8_364 b_8 NI_8 NS_364 0 2.1996722749807628e-06
GC_8_365 b_8 NI_8 NS_365 0 -2.4841809839038011e-06
GC_8_366 b_8 NI_8 NS_366 0 8.1284199573628565e-06
GC_8_367 b_8 NI_8 NS_367 0 -4.1621089905891762e-07
GC_8_368 b_8 NI_8 NS_368 0 9.3187009804518404e-06
GC_8_369 b_8 NI_8 NS_369 0 -9.6408195955614881e-07
GC_8_370 b_8 NI_8 NS_370 0 8.8146488276622710e-06
GC_8_371 b_8 NI_8 NS_371 0 -1.3883421701659043e-06
GC_8_372 b_8 NI_8 NS_372 0 3.8439572113941904e-06
GC_8_373 b_8 NI_8 NS_373 0 8.6419623397476754e-07
GC_8_374 b_8 NI_8 NS_374 0 1.1901958933401049e-05
GC_8_375 b_8 NI_8 NS_375 0 1.7097639427919700e-05
GC_8_376 b_8 NI_8 NS_376 0 1.6762494472821039e-05
GC_8_377 b_8 NI_8 NS_377 0 4.6416751066790113e-06
GC_8_378 b_8 NI_8 NS_378 0 7.7284892974222504e-06
GC_8_379 b_8 NI_8 NS_379 0 9.7558219955344957e-06
GC_8_380 b_8 NI_8 NS_380 0 3.9053284851497372e-06
GC_8_381 b_8 NI_8 NS_381 0 6.3770738348050761e-06
GC_8_382 b_8 NI_8 NS_382 0 1.0690285848842254e-05
GC_8_383 b_8 NI_8 NS_383 0 3.1851231990195633e-05
GC_8_384 b_8 NI_8 NS_384 0 -5.6094600821076868e-06
GC_8_385 b_8 NI_8 NS_385 0 7.7676141374849534e-06
GC_8_386 b_8 NI_8 NS_386 0 3.4156077066310829e-06
GC_8_387 b_8 NI_8 NS_387 0 1.1409488058873613e-05
GC_8_388 b_8 NI_8 NS_388 0 -9.8749562238320672e-06
GC_8_389 b_8 NI_8 NS_389 0 1.0301967794167643e-05
GC_8_390 b_8 NI_8 NS_390 0 6.2888529873386936e-06
GC_8_391 b_8 NI_8 NS_391 0 1.5924363443576804e-05
GC_8_392 b_8 NI_8 NS_392 0 -2.9747673223493136e-05
GC_8_393 b_8 NI_8 NS_393 0 7.6974773749466651e-06
GC_8_394 b_8 NI_8 NS_394 0 -2.8352584169027767e-06
GC_8_395 b_8 NI_8 NS_395 0 -3.4077940023007342e-06
GC_8_396 b_8 NI_8 NS_396 0 -1.5676420752981393e-05
GC_8_397 b_8 NI_8 NS_397 0 1.1261364478014304e-05
GC_8_398 b_8 NI_8 NS_398 0 -1.6843780008378871e-06
GC_8_399 b_8 NI_8 NS_399 0 -1.2932101805171953e-05
GC_8_400 b_8 NI_8 NS_400 0 -2.4084155053322922e-05
GC_8_401 b_8 NI_8 NS_401 0 -4.1147736752860135e-07
GC_8_402 b_8 NI_8 NS_402 0 -6.3604263657400408e-06
GC_8_403 b_8 NI_8 NS_403 0 -9.4858826989094438e-06
GC_8_404 b_8 NI_8 NS_404 0 -2.3359066229229365e-06
GC_8_405 b_8 NI_8 NS_405 0 9.8167979746012557e-11
GC_8_406 b_8 NI_8 NS_406 0 5.4215173643891974e-11
GC_8_407 b_8 NI_8 NS_407 0 1.1810245428980056e-06
GC_8_408 b_8 NI_8 NS_408 0 -4.5943646829897436e-06
GC_8_409 b_8 NI_8 NS_409 0 -1.4778922544044982e-06
GC_8_410 b_8 NI_8 NS_410 0 -1.2797107614446277e-06
GC_8_411 b_8 NI_8 NS_411 0 -4.9247463389521385e-06
GC_8_412 b_8 NI_8 NS_412 0 -8.6882694000754574e-07
GC_8_413 b_8 NI_8 NS_413 0 -1.3801279406145654e-06
GC_8_414 b_8 NI_8 NS_414 0 -2.8355647841123515e-06
GC_8_415 b_8 NI_8 NS_415 0 -1.0039741470687459e-05
GC_8_416 b_8 NI_8 NS_416 0 -3.6814544966089865e-06
GC_8_417 b_8 NI_8 NS_417 0 6.6579466269269080e-09
GC_8_418 b_8 NI_8 NS_418 0 5.7676982302497143e-09
GC_8_419 b_8 NI_8 NS_419 0 1.3984241976860616e-06
GC_8_420 b_8 NI_8 NS_420 0 6.7801362874168227e-07
GC_8_421 b_8 NI_8 NS_421 0 -1.7284102075742273e-06
GC_8_422 b_8 NI_8 NS_422 0 3.1540251826678959e-06
GC_8_423 b_8 NI_8 NS_423 0 -9.2400629022111193e-07
GC_8_424 b_8 NI_8 NS_424 0 7.7572763327212417e-07
GC_8_425 b_8 NI_8 NS_425 0 -7.9033355777707110e-06
GC_8_426 b_8 NI_8 NS_426 0 8.3212689592286366e-07
GC_8_427 b_8 NI_8 NS_427 0 -2.4107258891567869e-06
GC_8_428 b_8 NI_8 NS_428 0 2.0829178382818444e-06
GC_8_429 b_8 NI_8 NS_429 0 -2.1271855950981551e-06
GC_8_430 b_8 NI_8 NS_430 0 2.1516735458049076e-06
GC_8_431 b_8 NI_8 NS_431 0 1.1284198567745169e-06
GC_8_432 b_8 NI_8 NS_432 0 2.8125734742807797e-06
GC_8_433 b_8 NI_8 NS_433 0 -3.3197615081752346e-03
GC_8_434 b_8 NI_8 NS_434 0 1.8243968468152608e-09
GC_8_435 b_8 NI_8 NS_435 0 5.5833686493084548e-08
GC_8_436 b_8 NI_8 NS_436 0 1.8994900695693906e-06
GC_8_437 b_8 NI_8 NS_437 0 -9.0391575330406562e-05
GC_8_438 b_8 NI_8 NS_438 0 -5.8816093923958042e-05
GC_8_439 b_8 NI_8 NS_439 0 -1.2620478087040008e-03
GC_8_440 b_8 NI_8 NS_440 0 -3.0052236560685572e-04
GC_8_441 b_8 NI_8 NS_441 0 -1.6884314959595308e-03
GC_8_442 b_8 NI_8 NS_442 0 2.6375243457810731e-03
GC_8_443 b_8 NI_8 NS_443 0 4.9218123319088865e-04
GC_8_444 b_8 NI_8 NS_444 0 5.4232987542233027e-03
GC_8_445 b_8 NI_8 NS_445 0 7.0977003071595445e-03
GC_8_446 b_8 NI_8 NS_446 0 6.5580733309815182e-04
GC_8_447 b_8 NI_8 NS_447 0 6.4693661373288881e-04
GC_8_448 b_8 NI_8 NS_448 0 -6.5981382851704174e-04
GC_8_449 b_8 NI_8 NS_449 0 1.0491643622350293e-03
GC_8_450 b_8 NI_8 NS_450 0 1.5730848825106787e-03
GC_8_451 b_8 NI_8 NS_451 0 1.2639596499595221e-02
GC_8_452 b_8 NI_8 NS_452 0 1.3143541779121158e-02
GC_8_453 b_8 NI_8 NS_453 0 8.7648802085989966e-03
GC_8_454 b_8 NI_8 NS_454 0 -2.0356149451767436e-02
GC_8_455 b_8 NI_8 NS_455 0 8.3908950576227857e-03
GC_8_456 b_8 NI_8 NS_456 0 -2.8818704505541629e-03
GC_8_457 b_8 NI_8 NS_457 0 -1.2619354463904752e-02
GC_8_458 b_8 NI_8 NS_458 0 -3.8807130047440914e-02
GC_8_459 b_8 NI_8 NS_459 0 -7.2444872566046229e-03
GC_8_460 b_8 NI_8 NS_460 0 -2.1485695287368129e-03
GC_8_461 b_8 NI_8 NS_461 0 -5.2275002091325899e-02
GC_8_462 b_8 NI_8 NS_462 0 -1.8767942545632823e-03
GC_8_463 b_8 NI_8 NS_463 0 1.4892258823874656e-02
GC_8_464 b_8 NI_8 NS_464 0 8.6975609016882380e-03
GC_8_465 b_8 NI_8 NS_465 0 -5.9275334219211990e-03
GC_8_466 b_8 NI_8 NS_466 0 4.9905430455247212e-03
GC_8_467 b_8 NI_8 NS_467 0 8.3533688017224487e-03
GC_8_468 b_8 NI_8 NS_468 0 1.1690136307649283e-02
GC_8_469 b_8 NI_8 NS_469 0 4.5590086452082148e-03
GC_8_470 b_8 NI_8 NS_470 0 -2.9247924675703751e-03
GC_8_471 b_8 NI_8 NS_471 0 -7.8932497668077316e-03
GC_8_472 b_8 NI_8 NS_472 0 -8.1501573079923451e-03
GC_8_473 b_8 NI_8 NS_473 0 -5.6782675818886586e-03
GC_8_474 b_8 NI_8 NS_474 0 -6.1945400958126414e-04
GC_8_475 b_8 NI_8 NS_475 0 -1.8070913512968582e-02
GC_8_476 b_8 NI_8 NS_476 0 1.3562267899832786e-02
GC_8_477 b_8 NI_8 NS_477 0 4.7006660092960848e-03
GC_8_478 b_8 NI_8 NS_478 0 4.3832612388715669e-03
GC_8_479 b_8 NI_8 NS_479 0 6.4907931480250123e-04
GC_8_480 b_8 NI_8 NS_480 0 -1.1064190397761466e-04
GC_8_481 b_8 NI_8 NS_481 0 -3.7967898148776251e-03
GC_8_482 b_8 NI_8 NS_482 0 8.8034002849976349e-04
GC_8_483 b_8 NI_8 NS_483 0 -1.1248852085648164e-03
GC_8_484 b_8 NI_8 NS_484 0 1.6693626561085681e-02
GC_8_485 b_8 NI_8 NS_485 0 4.4443837140707735e-03
GC_8_486 b_8 NI_8 NS_486 0 7.1164090460713511e-04
GC_8_487 b_8 NI_8 NS_487 0 -5.2105051449812662e-04
GC_8_488 b_8 NI_8 NS_488 0 -2.2476775714394236e-03
GC_8_489 b_8 NI_8 NS_489 0 -4.9869184166386228e-03
GC_8_490 b_8 NI_8 NS_490 0 2.1058932028184384e-03
GC_8_491 b_8 NI_8 NS_491 0 7.3345843722000415e-03
GC_8_492 b_8 NI_8 NS_492 0 1.4346772732982627e-02
GC_8_493 b_8 NI_8 NS_493 0 4.1867517343199233e-03
GC_8_494 b_8 NI_8 NS_494 0 -1.6800221464522598e-03
GC_8_495 b_8 NI_8 NS_495 0 -3.3979308304660097e-03
GC_8_496 b_8 NI_8 NS_496 0 -2.1020221579586941e-03
GC_8_497 b_8 NI_8 NS_497 0 -5.4224795889632124e-03
GC_8_498 b_8 NI_8 NS_498 0 4.3763674872056733e-03
GC_8_499 b_8 NI_8 NS_499 0 1.3191405138831415e-02
GC_8_500 b_8 NI_8 NS_500 0 8.4408875032396437e-03
GC_8_501 b_8 NI_8 NS_501 0 2.8354678435713620e-03
GC_8_502 b_8 NI_8 NS_502 0 -4.1274253349838736e-03
GC_8_503 b_8 NI_8 NS_503 0 -5.3215613230068199e-03
GC_8_504 b_8 NI_8 NS_504 0 1.1333329869068157e-03
GC_8_505 b_8 NI_8 NS_505 0 -4.4370944731322711e-03
GC_8_506 b_8 NI_8 NS_506 0 8.3056982999971472e-03
GC_8_507 b_8 NI_8 NS_507 0 1.4614309671755638e-02
GC_8_508 b_8 NI_8 NS_508 0 -4.5696282968979164e-04
GC_8_509 b_8 NI_8 NS_509 0 -1.1788303179443309e-03
GC_8_510 b_8 NI_8 NS_510 0 -4.5487487055275297e-03
GC_8_511 b_8 NI_8 NS_511 0 -2.2870873693187099e-03
GC_8_512 b_8 NI_8 NS_512 0 4.3793455117308502e-03
GC_8_513 b_8 NI_8 NS_513 0 1.8266346702042387e-10
GC_8_514 b_8 NI_8 NS_514 0 -1.5798165189790476e-09
GC_8_515 b_8 NI_8 NS_515 0 1.4387706854913055e-03
GC_8_516 b_8 NI_8 NS_516 0 8.2177758807079702e-03
GC_8_517 b_8 NI_8 NS_517 0 -8.7491003054830131e-04
GC_8_518 b_8 NI_8 NS_518 0 -2.2094167279764986e-03
GC_8_519 b_8 NI_8 NS_519 0 -1.4716785383793491e-03
GC_8_520 b_8 NI_8 NS_520 0 2.7485704243094028e-03
GC_8_521 b_8 NI_8 NS_521 0 1.7223951665609062e-03
GC_8_522 b_8 NI_8 NS_522 0 7.6102907946118004e-03
GC_8_523 b_8 NI_8 NS_523 0 7.5930439282453042e-03
GC_8_524 b_8 NI_8 NS_524 0 -3.8216212223364061e-03
GC_8_525 b_8 NI_8 NS_525 0 -4.7008113719748075e-08
GC_8_526 b_8 NI_8 NS_526 0 -2.0170175921527560e-08
GC_8_527 b_8 NI_8 NS_527 0 1.1386078511075155e-02
GC_8_528 b_8 NI_8 NS_528 0 4.4716365186009445e-03
GC_8_529 b_8 NI_8 NS_529 0 -8.6429611106076960e-04
GC_8_530 b_8 NI_8 NS_530 0 6.4881769365537556e-03
GC_8_531 b_8 NI_8 NS_531 0 3.6256397905615558e-03
GC_8_532 b_8 NI_8 NS_532 0 4.0760139183395434e-04
GC_8_533 b_8 NI_8 NS_533 0 6.0652196136451487e-03
GC_8_534 b_8 NI_8 NS_534 0 -4.6566352533665431e-03
GC_8_535 b_8 NI_8 NS_535 0 -3.3846294272645329e-03
GC_8_536 b_8 NI_8 NS_536 0 -1.3607984535558293e-03
GC_8_537 b_8 NI_8 NS_537 0 1.0687140882372673e-04
GC_8_538 b_8 NI_8 NS_538 0 4.4902870768095031e-03
GC_8_539 b_8 NI_8 NS_539 0 7.2783999813574004e-03
GC_8_540 b_8 NI_8 NS_540 0 5.5303118665791986e-03
GC_8_541 b_8 NI_8 NS_541 0 1.4425743160262673e-03
GC_8_542 b_8 NI_8 NS_542 0 -3.5904351902283599e-09
GC_8_543 b_8 NI_8 NS_543 0 -4.7342043005241280e-08
GC_8_544 b_8 NI_8 NS_544 0 -3.5032371879164385e-06
GC_8_545 b_8 NI_8 NS_545 0 -3.6675402894641808e-04
GC_8_546 b_8 NI_8 NS_546 0 1.3531650072534562e-04
GC_8_547 b_8 NI_8 NS_547 0 1.1270906275200328e-03
GC_8_548 b_8 NI_8 NS_548 0 1.9466317895270317e-03
GC_8_549 b_8 NI_8 NS_549 0 -5.2133196348722021e-05
GC_8_550 b_8 NI_8 NS_550 0 -3.4959654221104397e-03
GC_8_551 b_8 NI_8 NS_551 0 -1.5728294468906265e-03
GC_8_552 b_8 NI_8 NS_552 0 5.0835061312654610e-03
GC_8_553 b_8 NI_8 NS_553 0 4.2660497518821339e-03
GC_8_554 b_8 NI_8 NS_554 0 -4.9897929468884755e-03
GC_8_555 b_8 NI_8 NS_555 0 -1.0071498220759027e-03
GC_8_556 b_8 NI_8 NS_556 0 5.5941855889054973e-04
GC_8_557 b_8 NI_8 NS_557 0 -2.0791294208185309e-03
GC_8_558 b_8 NI_8 NS_558 0 -1.8719561555057042e-03
GC_8_559 b_8 NI_8 NS_559 0 3.6235023872610182e-03
GC_8_560 b_8 NI_8 NS_560 0 1.1644121608893448e-02
GC_8_561 b_8 NI_8 NS_561 0 -8.7672707288609787e-04
GC_8_562 b_8 NI_8 NS_562 0 -1.4855229397094554e-02
GC_8_563 b_8 NI_8 NS_563 0 -8.1250075395500349e-03
GC_8_564 b_8 NI_8 NS_564 0 1.9028461769213844e-03
GC_8_565 b_8 NI_8 NS_565 0 1.1255574772855069e-02
GC_8_566 b_8 NI_8 NS_566 0 -1.8013331580536425e-03
GC_8_567 b_8 NI_8 NS_567 0 -7.5649379527732855e-03
GC_8_568 b_8 NI_8 NS_568 0 -1.6931181123028608e-03
GC_8_569 b_8 NI_8 NS_569 0 1.5263484583700115e-02
GC_8_570 b_8 NI_8 NS_570 0 5.3089269192998752e-03
GC_8_571 b_8 NI_8 NS_571 0 -1.3074208595461044e-02
GC_8_572 b_8 NI_8 NS_572 0 -5.4740973546441984e-03
GC_8_573 b_8 NI_8 NS_573 0 -6.6401728312199546e-03
GC_8_574 b_8 NI_8 NS_574 0 3.4469264611769719e-03
GC_8_575 b_8 NI_8 NS_575 0 6.3571561981592157e-03
GC_8_576 b_8 NI_8 NS_576 0 -1.8769364689313543e-03
GC_8_577 b_8 NI_8 NS_577 0 -5.4767784277633697e-03
GC_8_578 b_8 NI_8 NS_578 0 2.1761635009273470e-03
GC_8_579 b_8 NI_8 NS_579 0 5.3904709118370977e-03
GC_8_580 b_8 NI_8 NS_580 0 -2.6291409473561582e-03
GC_8_581 b_8 NI_8 NS_581 0 -6.3068613159885214e-03
GC_8_582 b_8 NI_8 NS_582 0 -4.8944545977234772e-04
GC_8_583 b_8 NI_8 NS_583 0 7.6383029679271642e-03
GC_8_584 b_8 NI_8 NS_584 0 3.6283278652217924e-03
GC_8_585 b_8 NI_8 NS_585 0 -5.8333234857385497e-03
GC_8_586 b_8 NI_8 NS_586 0 -3.4684301852644598e-03
GC_8_587 b_8 NI_8 NS_587 0 2.9592189498357135e-04
GC_8_588 b_8 NI_8 NS_588 0 5.5702925731856414e-04
GC_8_589 b_8 NI_8 NS_589 0 -4.9284028648939751e-03
GC_8_590 b_8 NI_8 NS_590 0 8.8733927749224620e-04
GC_8_591 b_8 NI_8 NS_591 0 6.2016451885348513e-03
GC_8_592 b_8 NI_8 NS_592 0 6.8248095452391017e-04
GC_8_593 b_8 NI_8 NS_593 0 -5.3226827125025192e-03
GC_8_594 b_8 NI_8 NS_594 0 -4.8918923172083708e-04
GC_8_595 b_8 NI_8 NS_595 0 1.5482736461423169e-03
GC_8_596 b_8 NI_8 NS_596 0 -4.6609139365975398e-05
GC_8_597 b_8 NI_8 NS_597 0 -6.0242735099149194e-03
GC_8_598 b_8 NI_8 NS_598 0 1.9161515657498943e-03
GC_8_599 b_8 NI_8 NS_599 0 6.2494033097370630e-03
GC_8_600 b_8 NI_8 NS_600 0 2.0850478901609910e-04
GC_8_601 b_8 NI_8 NS_601 0 -5.0636589797220426e-03
GC_8_602 b_8 NI_8 NS_602 0 1.6954532442549862e-03
GC_8_603 b_8 NI_8 NS_603 0 2.4806587508527894e-03
GC_8_604 b_8 NI_8 NS_604 0 -9.6015729719453569e-04
GC_8_605 b_8 NI_8 NS_605 0 -6.5381321213502132e-03
GC_8_606 b_8 NI_8 NS_606 0 3.8750074616024205e-03
GC_8_607 b_8 NI_8 NS_607 0 7.4722546541910219e-03
GC_8_608 b_8 NI_8 NS_608 0 -1.0944729819687170e-03
GC_8_609 b_8 NI_8 NS_609 0 -3.9943218736882245e-03
GC_8_610 b_8 NI_8 NS_610 0 4.0357752344018557e-03
GC_8_611 b_8 NI_8 NS_611 0 2.8552013767557606e-03
GC_8_612 b_8 NI_8 NS_612 0 -3.0472624895248311e-03
GC_8_613 b_8 NI_8 NS_613 0 -6.0351388958250736e-03
GC_8_614 b_8 NI_8 NS_614 0 7.2276062148212226e-03
GC_8_615 b_8 NI_8 NS_615 0 7.9782887147300530e-03
GC_8_616 b_8 NI_8 NS_616 0 -4.7935801973903987e-03
GC_8_617 b_8 NI_8 NS_617 0 -5.4799474981498202e-04
GC_8_618 b_8 NI_8 NS_618 0 5.0230804901846803e-03
GC_8_619 b_8 NI_8 NS_619 0 2.5034134627312601e-04
GC_8_620 b_8 NI_8 NS_620 0 -4.7520661386947919e-03
GC_8_621 b_8 NI_8 NS_621 0 1.7366272814732665e-09
GC_8_622 b_8 NI_8 NS_622 0 3.2860222505096964e-09
GC_8_623 b_8 NI_8 NS_623 0 -1.4394125008006711e-03
GC_8_624 b_8 NI_8 NS_624 0 7.8706604761739751e-03
GC_8_625 b_8 NI_8 NS_625 0 -1.8574746928496201e-04
GC_8_626 b_8 NI_8 NS_626 0 3.0287972688730781e-03
GC_8_627 b_8 NI_8 NS_627 0 -1.2900533406371567e-04
GC_8_628 b_8 NI_8 NS_628 0 -3.3736684302623963e-03
GC_8_629 b_8 NI_8 NS_629 0 -8.9083181786642196e-04
GC_8_630 b_8 NI_8 NS_630 0 7.5293774121917194e-03
GC_8_631 b_8 NI_8 NS_631 0 3.7906243928354458e-03
GC_8_632 b_8 NI_8 NS_632 0 -6.1490577388281231e-03
GC_8_633 b_8 NI_8 NS_633 0 8.8448813607638299e-08
GC_8_634 b_8 NI_8 NS_634 0 -3.5531433518670525e-07
GC_8_635 b_8 NI_8 NS_635 0 6.7115065628059571e-03
GC_8_636 b_8 NI_8 NS_636 0 -5.3183245754123785e-03
GC_8_637 b_8 NI_8 NS_637 0 -2.6127433872478044e-03
GC_8_638 b_8 NI_8 NS_638 0 6.0487711501957470e-03
GC_8_639 b_8 NI_8 NS_639 0 -4.2945275038195592e-03
GC_8_640 b_8 NI_8 NS_640 0 1.3261562382252643e-05
GC_8_641 b_8 NI_8 NS_641 0 2.7224992724420517e-03
GC_8_642 b_8 NI_8 NS_642 0 -6.1956590818551156e-03
GC_8_643 b_8 NI_8 NS_643 0 2.0898364046733242e-03
GC_8_644 b_8 NI_8 NS_644 0 3.2611136183944987e-03
GC_8_645 b_8 NI_8 NS_645 0 -1.9638287424718730e-03
GC_8_646 b_8 NI_8 NS_646 0 -4.4203348237130550e-03
GC_8_647 b_8 NI_8 NS_647 0 2.8567435015331199e-03
GC_8_648 b_8 NI_8 NS_648 0 8.0017787545880788e-03
GC_8_649 b_8 NI_8 NS_649 0 -1.0963267163615556e-02
GC_8_650 b_8 NI_8 NS_650 0 8.3273558240227229e-09
GC_8_651 b_8 NI_8 NS_651 0 9.8608133417170609e-07
GC_8_652 b_8 NI_8 NS_652 0 3.6177581400220342e-05
GC_8_653 b_8 NI_8 NS_653 0 4.3739133121249206e-03
GC_8_654 b_8 NI_8 NS_654 0 -3.4750208858145815e-03
GC_8_655 b_8 NI_8 NS_655 0 -3.7382649263803117e-03
GC_8_656 b_8 NI_8 NS_656 0 6.2463704875684728e-03
GC_8_657 b_8 NI_8 NS_657 0 -8.7586408382760560e-03
GC_8_658 b_8 NI_8 NS_658 0 -5.9567965015504898e-03
GC_8_659 b_8 NI_8 NS_659 0 9.2115224594777664e-03
GC_8_660 b_8 NI_8 NS_660 0 -5.9461545218707492e-03
GC_8_661 b_8 NI_8 NS_661 0 7.1478506730971794e-03
GC_8_662 b_8 NI_8 NS_662 0 1.1907364828146454e-02
GC_8_663 b_8 NI_8 NS_663 0 -4.2314406094072299e-03
GC_8_664 b_8 NI_8 NS_664 0 -1.1324311967114867e-03
GC_8_665 b_8 NI_8 NS_665 0 -8.8598536418343730e-03
GC_8_666 b_8 NI_8 NS_666 0 -4.7416849389066552e-04
GC_8_667 b_8 NI_8 NS_667 0 1.4618431657846705e-02
GC_8_668 b_8 NI_8 NS_668 0 -1.0343807410178374e-02
GC_8_669 b_8 NI_8 NS_669 0 1.6441834998184746e-02
GC_8_670 b_8 NI_8 NS_670 0 4.0225150480326481e-03
GC_8_671 b_8 NI_8 NS_671 0 -1.1482356389915647e-02
GC_8_672 b_8 NI_8 NS_672 0 -2.4511055153151690e-04
GC_8_673 b_8 NI_8 NS_673 0 -1.6636905693249070e-02
GC_8_674 b_8 NI_8 NS_674 0 -4.4573847593434746e-02
GC_8_675 b_8 NI_8 NS_675 0 1.0652626364474773e-02
GC_8_676 b_8 NI_8 NS_676 0 1.1245824546634081e-03
GC_8_677 b_8 NI_8 NS_677 0 -4.8294136626157780e-02
GC_8_678 b_8 NI_8 NS_678 0 1.1061815040578954e-02
GC_8_679 b_8 NI_8 NS_679 0 -1.0433725392419936e-02
GC_8_680 b_8 NI_8 NS_680 0 4.8881006466942054e-04
GC_8_681 b_8 NI_8 NS_681 0 9.7769820990579199e-03
GC_8_682 b_8 NI_8 NS_682 0 -5.7678142352605999e-04
GC_8_683 b_8 NI_8 NS_683 0 4.6096297805843581e-03
GC_8_684 b_8 NI_8 NS_684 0 2.4174057785829706e-02
GC_8_685 b_8 NI_8 NS_685 0 -1.0735332678457969e-02
GC_8_686 b_8 NI_8 NS_686 0 1.9692174283492091e-03
GC_8_687 b_8 NI_8 NS_687 0 -8.4726796466467955e-03
GC_8_688 b_8 NI_8 NS_688 0 -1.3537898486971126e-02
GC_8_689 b_8 NI_8 NS_689 0 1.0150146142671455e-02
GC_8_690 b_8 NI_8 NS_690 0 9.8140263034084347e-04
GC_8_691 b_8 NI_8 NS_691 0 -1.9163084845158392e-02
GC_8_692 b_8 NI_8 NS_692 0 2.8679143996748226e-02
GC_8_693 b_8 NI_8 NS_693 0 -9.6128593052273101e-03
GC_8_694 b_8 NI_8 NS_694 0 -9.6556218531649641e-04
GC_8_695 b_8 NI_8 NS_695 0 1.8914256698378830e-03
GC_8_696 b_8 NI_8 NS_696 0 -1.3780642195261390e-03
GC_8_697 b_8 NI_8 NS_697 0 9.4682934906295483e-03
GC_8_698 b_8 NI_8 NS_698 0 -2.4742906784666765e-04
GC_8_699 b_8 NI_8 NS_699 0 -1.4947690032120667e-04
GC_8_700 b_8 NI_8 NS_700 0 3.0270099735804783e-02
GC_8_701 b_8 NI_8 NS_701 0 -8.5288666668267427e-03
GC_8_702 b_8 NI_8 NS_702 0 1.5479353290652112e-04
GC_8_703 b_8 NI_8 NS_703 0 2.1682367697665390e-04
GC_8_704 b_8 NI_8 NS_704 0 -5.4812459368185412e-03
GC_8_705 b_8 NI_8 NS_705 0 1.0036172398963972e-02
GC_8_706 b_8 NI_8 NS_706 0 -3.3856905311609712e-04
GC_8_707 b_8 NI_8 NS_707 0 8.9341986552970917e-03
GC_8_708 b_8 NI_8 NS_708 0 2.6365820649268686e-02
GC_8_709 b_8 NI_8 NS_709 0 -8.3555299518811906e-03
GC_8_710 b_8 NI_8 NS_710 0 1.3766425485373910e-03
GC_8_711 b_8 NI_8 NS_711 0 -2.5868995912225919e-03
GC_8_712 b_8 NI_8 NS_712 0 -7.3539695158887468e-03
GC_8_713 b_8 NI_8 NS_713 0 1.0553570375689646e-02
GC_8_714 b_8 NI_8 NS_714 0 -8.2349532403831098e-04
GC_8_715 b_8 NI_8 NS_715 0 1.4439005330395492e-02
GC_8_716 b_8 NI_8 NS_716 0 1.9950592749697335e-02
GC_8_717 b_8 NI_8 NS_717 0 -8.2760901444011124e-03
GC_8_718 b_8 NI_8 NS_718 0 2.9305080491009408e-03
GC_8_719 b_8 NI_8 NS_719 0 -5.5941898644445579e-03
GC_8_720 b_8 NI_8 NS_720 0 -6.9177066985703717e-03
GC_8_721 b_8 NI_8 NS_721 0 1.1244068786109772e-02
GC_8_722 b_8 NI_8 NS_722 0 -1.3754067091735658e-03
GC_8_723 b_8 NI_8 NS_723 0 1.5700544491828585e-02
GC_8_724 b_8 NI_8 NS_724 0 1.2945581178294334e-02
GC_8_725 b_8 NI_8 NS_725 0 -7.1893561392462873e-03
GC_8_726 b_8 NI_8 NS_726 0 5.1106036735557980e-03
GC_8_727 b_8 NI_8 NS_727 0 -6.8765841756682905e-03
GC_8_728 b_8 NI_8 NS_728 0 -4.8360484640687521e-03
GC_8_729 b_8 NI_8 NS_729 0 4.7735848894475902e-09
GC_8_730 b_8 NI_8 NS_730 0 4.4198496642633848e-08
GC_8_731 b_8 NI_8 NS_731 0 1.2004110238625411e-02
GC_8_732 b_8 NI_8 NS_732 0 -2.5766647096991985e-03
GC_8_733 b_8 NI_8 NS_733 0 -5.2510735941698160e-03
GC_8_734 b_8 NI_8 NS_734 0 4.7015438422580167e-03
GC_8_735 b_8 NI_8 NS_735 0 -6.1588966197801539e-03
GC_8_736 b_8 NI_8 NS_736 0 -4.3232052598594813e-03
GC_8_737 b_8 NI_8 NS_737 0 1.1774224067196677e-02
GC_8_738 b_8 NI_8 NS_738 0 -3.7297236083615195e-03
GC_8_739 b_8 NI_8 NS_739 0 1.2978428655534760e-02
GC_8_740 b_8 NI_8 NS_740 0 9.4653911577906157e-03
GC_8_741 b_8 NI_8 NS_741 0 3.9180865997499054e-06
GC_8_742 b_8 NI_8 NS_742 0 -9.4184571939958278e-07
GC_8_743 b_8 NI_8 NS_743 0 1.6087881053032115e-02
GC_8_744 b_8 NI_8 NS_744 0 1.6769943948052275e-02
GC_8_745 b_8 NI_8 NS_745 0 1.2047069299917234e-02
GC_8_746 b_8 NI_8 NS_746 0 -2.4806934562173252e-03
GC_8_747 b_8 NI_8 NS_747 0 -8.3607711567733368e-03
GC_8_748 b_8 NI_8 NS_748 0 7.9691057007696069e-05
GC_8_749 b_8 NI_8 NS_749 0 1.1309400430646627e-02
GC_8_750 b_8 NI_8 NS_750 0 7.3306414636073215e-03
GC_8_751 b_8 NI_8 NS_751 0 -4.6732525219133738e-03
GC_8_752 b_8 NI_8 NS_752 0 7.3569202905622282e-03
GC_8_753 b_8 NI_8 NS_753 0 -8.0809734698303569e-03
GC_8_754 b_8 NI_8 NS_754 0 -3.7224029866739436e-03
GC_8_755 b_8 NI_8 NS_755 0 1.5958294466899683e-02
GC_8_756 b_8 NI_8 NS_756 0 -7.7554798974917554e-03
GC_8_757 b_8 NI_8 NS_757 0 -1.3590089392699197e-02
GC_8_758 b_8 NI_8 NS_758 0 5.7574152498708389e-09
GC_8_759 b_8 NI_8 NS_759 0 -1.0755252268141780e-06
GC_8_760 b_8 NI_8 NS_760 0 -2.3265199713856362e-05
GC_8_761 b_8 NI_8 NS_761 0 3.4981896186587450e-04
GC_8_762 b_8 NI_8 NS_762 0 -1.9740617794120080e-04
GC_8_763 b_8 NI_8 NS_763 0 -1.5437475694336450e-03
GC_8_764 b_8 NI_8 NS_764 0 -2.3356984989387447e-03
GC_8_765 b_8 NI_8 NS_765 0 -5.1338576158386038e-05
GC_8_766 b_8 NI_8 NS_766 0 4.3605105822488738e-03
GC_8_767 b_8 NI_8 NS_767 0 1.6175854247143014e-03
GC_8_768 b_8 NI_8 NS_768 0 -5.9520447551457568e-03
GC_8_769 b_8 NI_8 NS_769 0 -4.9853642799081487e-03
GC_8_770 b_8 NI_8 NS_770 0 6.4563496909199637e-03
GC_8_771 b_8 NI_8 NS_771 0 1.1341369443484291e-03
GC_8_772 b_8 NI_8 NS_772 0 -5.0676047520777122e-04
GC_8_773 b_8 NI_8 NS_773 0 2.7870925906266081e-03
GC_8_774 b_8 NI_8 NS_774 0 2.3388070901895299e-03
GC_8_775 b_8 NI_8 NS_775 0 -4.3321840737588291e-03
GC_8_776 b_8 NI_8 NS_776 0 -1.3583569026987262e-02
GC_8_777 b_8 NI_8 NS_777 0 1.5695054733301118e-03
GC_8_778 b_8 NI_8 NS_778 0 1.7683056108125275e-02
GC_8_779 b_8 NI_8 NS_779 0 9.8323100585864381e-03
GC_8_780 b_8 NI_8 NS_780 0 -2.3109433971130354e-03
GC_8_781 b_8 NI_8 NS_781 0 -1.3157076653895183e-02
GC_8_782 b_8 NI_8 NS_782 0 2.2142577719870432e-03
GC_8_783 b_8 NI_8 NS_783 0 9.1925801996316798e-03
GC_8_784 b_8 NI_8 NS_784 0 1.9425128055761535e-03
GC_8_785 b_8 NI_8 NS_785 0 -1.8069416737093169e-02
GC_8_786 b_8 NI_8 NS_786 0 -6.4922072793175811e-03
GC_8_787 b_8 NI_8 NS_787 0 1.5725031894717315e-02
GC_8_788 b_8 NI_8 NS_788 0 6.4951372716310603e-03
GC_8_789 b_8 NI_8 NS_789 0 8.1032021061081139e-03
GC_8_790 b_8 NI_8 NS_790 0 -4.2110865808055722e-03
GC_8_791 b_8 NI_8 NS_791 0 -7.5660733787599700e-03
GC_8_792 b_8 NI_8 NS_792 0 2.0432108254830844e-03
GC_8_793 b_8 NI_8 NS_793 0 6.6854403795751473e-03
GC_8_794 b_8 NI_8 NS_794 0 -2.7541191547744469e-03
GC_8_795 b_8 NI_8 NS_795 0 -6.6055143819591091e-03
GC_8_796 b_8 NI_8 NS_796 0 2.9142089168934229e-03
GC_8_797 b_8 NI_8 NS_797 0 7.6544550432041565e-03
GC_8_798 b_8 NI_8 NS_798 0 4.7731847373014285e-04
GC_8_799 b_8 NI_8 NS_799 0 -9.4088383419286842e-03
GC_8_800 b_8 NI_8 NS_800 0 -5.1695913268952863e-03
GC_8_801 b_8 NI_8 NS_801 0 6.8169860777994714e-03
GC_8_802 b_8 NI_8 NS_802 0 4.1131838889598201e-03
GC_8_803 b_8 NI_8 NS_803 0 -3.9575075777870084e-04
GC_8_804 b_8 NI_8 NS_804 0 -9.3603865378935928e-04
GC_8_805 b_8 NI_8 NS_805 0 5.6653330903599433e-03
GC_8_806 b_8 NI_8 NS_806 0 -1.3801763521174536e-03
GC_8_807 b_8 NI_8 NS_807 0 -9.2023055604560974e-03
GC_8_808 b_8 NI_8 NS_808 0 -1.2455924515789119e-03
GC_8_809 b_8 NI_8 NS_809 0 5.9915361490972922e-03
GC_8_810 b_8 NI_8 NS_810 0 7.3808288926781632e-04
GC_8_811 b_8 NI_8 NS_811 0 -2.6544499887793606e-03
GC_8_812 b_8 NI_8 NS_812 0 2.4842218286524653e-04
GC_8_813 b_8 NI_8 NS_813 0 6.6958869570911692e-03
GC_8_814 b_8 NI_8 NS_814 0 -2.2582332604380384e-03
GC_8_815 b_8 NI_8 NS_815 0 -9.3158034337997974e-03
GC_8_816 b_8 NI_8 NS_816 0 1.5268579780520007e-03
GC_8_817 b_8 NI_8 NS_817 0 5.7300528240279962e-03
GC_8_818 b_8 NI_8 NS_818 0 -1.5007464209294873e-03
GC_8_819 b_8 NI_8 NS_819 0 -3.3211786392641491e-03
GC_8_820 b_8 NI_8 NS_820 0 2.4082406838792907e-03
GC_8_821 b_8 NI_8 NS_821 0 7.2643748459256989e-03
GC_8_822 b_8 NI_8 NS_822 0 -4.0966020234659865e-03
GC_8_823 b_8 NI_8 NS_823 0 -8.5936626208301184e-03
GC_8_824 b_8 NI_8 NS_824 0 4.2025458057814288e-03
GC_8_825 b_8 NI_8 NS_825 0 4.8158718107755970e-03
GC_8_826 b_8 NI_8 NS_826 0 -3.8696534356424837e-03
GC_8_827 b_8 NI_8 NS_827 0 -2.4037832577573606e-03
GC_8_828 b_8 NI_8 NS_828 0 4.7598869813829416e-03
GC_8_829 b_8 NI_8 NS_829 0 7.0540650269528297e-03
GC_8_830 b_8 NI_8 NS_830 0 -7.3479411359841200e-03
GC_8_831 b_8 NI_8 NS_831 0 -7.1270973131391472e-03
GC_8_832 b_8 NI_8 NS_832 0 6.8936460130063172e-03
GC_8_833 b_8 NI_8 NS_833 0 1.6683535826809515e-03
GC_8_834 b_8 NI_8 NS_834 0 -5.2972271114585471e-03
GC_8_835 b_8 NI_8 NS_835 0 5.9423054445045223e-04
GC_8_836 b_8 NI_8 NS_836 0 5.4734750972631214e-03
GC_8_837 b_8 NI_8 NS_837 0 -4.1995963853196410e-09
GC_8_838 b_8 NI_8 NS_838 0 -1.3215418100257055e-08
GC_8_839 b_8 NI_8 NS_839 0 2.7118337317614347e-03
GC_8_840 b_8 NI_8 NS_840 0 -8.5806168970764679e-03
GC_8_841 b_8 NI_8 NS_841 0 8.7189177798861761e-04
GC_8_842 b_8 NI_8 NS_842 0 -3.4318677496630173e-03
GC_8_843 b_8 NI_8 NS_843 0 6.2897519477433451e-04
GC_8_844 b_8 NI_8 NS_844 0 4.0346891063128120e-03
GC_8_845 b_8 NI_8 NS_845 0 2.1766552368069460e-03
GC_8_846 b_8 NI_8 NS_846 0 -8.1586502032184594e-03
GC_8_847 b_8 NI_8 NS_847 0 -3.4870473344026129e-03
GC_8_848 b_8 NI_8 NS_848 0 7.0184761649907702e-03
GC_8_849 b_8 NI_8 NS_849 0 -9.0339788463211348e-08
GC_8_850 b_8 NI_8 NS_850 0 -3.0341137820751456e-07
GC_8_851 b_8 NI_8 NS_851 0 -8.0011228498603499e-03
GC_8_852 b_8 NI_8 NS_852 0 5.3809315920449602e-03
GC_8_853 b_8 NI_8 NS_853 0 4.1753805465283697e-03
GC_8_854 b_8 NI_8 NS_854 0 -6.8471567929904512e-03
GC_8_855 b_8 NI_8 NS_855 0 5.3267681360825193e-03
GC_8_856 b_8 NI_8 NS_856 0 7.4221548312965950e-04
GC_8_857 b_8 NI_8 NS_857 0 -2.3672741529547139e-03
GC_8_858 b_8 NI_8 NS_858 0 6.8575158556994000e-03
GC_8_859 b_8 NI_8 NS_859 0 -1.4866263327029422e-03
GC_8_860 b_8 NI_8 NS_860 0 -4.2154565571034825e-03
GC_8_861 b_8 NI_8 NS_861 0 2.3568559828398964e-03
GC_8_862 b_8 NI_8 NS_862 0 5.0372654950294922e-03
GC_8_863 b_8 NI_8 NS_863 0 -1.9997028978518314e-03
GC_8_864 b_8 NI_8 NS_864 0 -8.9736634094011065e-03
GC_8_865 b_8 NI_8 NS_865 0 -6.3819045123490454e-04
GC_8_866 b_8 NI_8 NS_866 0 -9.7139014931444971e-11
GC_8_867 b_8 NI_8 NS_867 0 3.8809212179849958e-09
GC_8_868 b_8 NI_8 NS_868 0 -6.7423154828811638e-08
GC_8_869 b_8 NI_8 NS_869 0 -1.1292055994835782e-05
GC_8_870 b_8 NI_8 NS_870 0 -9.3317586031021132e-06
GC_8_871 b_8 NI_8 NS_871 0 -2.2441885173982082e-06
GC_8_872 b_8 NI_8 NS_872 0 2.2643068851606957e-07
GC_8_873 b_8 NI_8 NS_873 0 -3.0298269682759658e-05
GC_8_874 b_8 NI_8 NS_874 0 2.7085504736751332e-05
GC_8_875 b_8 NI_8 NS_875 0 -3.3245382921988061e-05
GC_8_876 b_8 NI_8 NS_876 0 8.1393427424868165e-06
GC_8_877 b_8 NI_8 NS_877 0 3.1754283744020495e-05
GC_8_878 b_8 NI_8 NS_878 0 2.7340888068444269e-05
GC_8_879 b_8 NI_8 NS_879 0 -9.0548909826326032e-06
GC_8_880 b_8 NI_8 NS_880 0 1.4743919436254082e-05
GC_8_881 b_8 NI_8 NS_881 0 1.2670953744548778e-05
GC_8_882 b_8 NI_8 NS_882 0 3.6937562957687217e-05
GC_8_883 b_8 NI_8 NS_883 0 -1.0602077981935941e-05
GC_8_884 b_8 NI_8 NS_884 0 6.8138223591564768e-05
GC_8_885 b_8 NI_8 NS_885 0 9.5404371417307429e-05
GC_8_886 b_8 NI_8 NS_886 0 -6.6240437925171972e-05
GC_8_887 b_8 NI_8 NS_887 0 2.7099114554271931e-05
GC_8_888 b_8 NI_8 NS_888 0 3.1676109559132145e-05
GC_8_889 b_8 NI_8 NS_889 0 -7.4559443761429928e-06
GC_8_890 b_8 NI_8 NS_890 0 -7.2595415389403950e-05
GC_8_891 b_8 NI_8 NS_891 0 -9.8760710242854638e-06
GC_8_892 b_8 NI_8 NS_892 0 -3.3982285223095123e-05
GC_8_893 b_8 NI_8 NS_893 0 -7.7016022905310823e-05
GC_8_894 b_8 NI_8 NS_894 0 1.9174780943685061e-05
GC_8_895 b_8 NI_8 NS_895 0 2.4970781923444521e-05
GC_8_896 b_8 NI_8 NS_896 0 5.0900352288878994e-05
GC_8_897 b_8 NI_8 NS_897 0 -2.3151129821017979e-05
GC_8_898 b_8 NI_8 NS_898 0 -3.5305283279587725e-06
GC_8_899 b_8 NI_8 NS_899 0 6.9874070756373283e-05
GC_8_900 b_8 NI_8 NS_900 0 4.4645040927349702e-05
GC_8_901 b_8 NI_8 NS_901 0 2.9213306598011200e-05
GC_8_902 b_8 NI_8 NS_902 0 1.9680256533082643e-05
GC_8_903 b_8 NI_8 NS_903 0 -7.3499986729041596e-06
GC_8_904 b_8 NI_8 NS_904 0 -2.5717486598762058e-05
GC_8_905 b_8 NI_8 NS_905 0 -7.6009666873922395e-06
GC_8_906 b_8 NI_8 NS_906 0 -2.5156205006081675e-05
GC_8_907 b_8 NI_8 NS_907 0 6.7666630937238335e-06
GC_8_908 b_8 NI_8 NS_908 0 4.9266774407680884e-05
GC_8_909 b_8 NI_8 NS_909 0 1.2941336945077549e-05
GC_8_910 b_8 NI_8 NS_910 0 2.7354614959747736e-05
GC_8_911 b_8 NI_8 NS_911 0 5.8648271665993535e-06
GC_8_912 b_8 NI_8 NS_912 0 2.1243225216481801e-06
GC_8_913 b_8 NI_8 NS_913 0 -6.3929727130516110e-07
GC_8_914 b_8 NI_8 NS_914 0 -1.5371386934314199e-05
GC_8_915 b_8 NI_8 NS_915 0 5.6176805751887757e-05
GC_8_916 b_8 NI_8 NS_916 0 3.8178320032679190e-05
GC_8_917 b_8 NI_8 NS_917 0 1.9951189550193791e-05
GC_8_918 b_8 NI_8 NS_918 0 1.4801252536911883e-05
GC_8_919 b_8 NI_8 NS_919 0 8.3758527716061313e-06
GC_8_920 b_8 NI_8 NS_920 0 -1.2841470841841403e-05
GC_8_921 b_8 NI_8 NS_921 0 -5.6602023716809923e-06
GC_8_922 b_8 NI_8 NS_922 0 -1.3971556509401184e-05
GC_8_923 b_8 NI_8 NS_923 0 6.6117296272822550e-05
GC_8_924 b_8 NI_8 NS_924 0 1.3011960662674814e-05
GC_8_925 b_8 NI_8 NS_925 0 2.2771804031875316e-05
GC_8_926 b_8 NI_8 NS_926 0 4.9238786207864425e-06
GC_8_927 b_8 NI_8 NS_927 0 -5.5579226572840975e-06
GC_8_928 b_8 NI_8 NS_928 0 -2.1967464621292030e-05
GC_8_929 b_8 NI_8 NS_929 0 -9.1458147383241964e-06
GC_8_930 b_8 NI_8 NS_930 0 -7.0555574392312071e-06
GC_8_931 b_8 NI_8 NS_931 0 6.0678791954734983e-05
GC_8_932 b_8 NI_8 NS_932 0 -9.4911797076412862e-06
GC_8_933 b_8 NI_8 NS_933 0 2.1422961709231469e-05
GC_8_934 b_8 NI_8 NS_934 0 -7.3860865759842646e-06
GC_8_935 b_8 NI_8 NS_935 0 -2.3066440526547223e-05
GC_8_936 b_8 NI_8 NS_936 0 -1.3101703004514835e-05
GC_8_937 b_8 NI_8 NS_937 0 -8.6613436903313765e-06
GC_8_938 b_8 NI_8 NS_938 0 4.4700965331380755e-06
GC_8_939 b_8 NI_8 NS_939 0 4.5474465807806720e-05
GC_8_940 b_8 NI_8 NS_940 0 -2.5680596822803277e-05
GC_8_941 b_8 NI_8 NS_941 0 6.0237990555890736e-06
GC_8_942 b_8 NI_8 NS_942 0 -1.6485892677598157e-05
GC_8_943 b_8 NI_8 NS_943 0 -1.8717568031343225e-05
GC_8_944 b_8 NI_8 NS_944 0 8.6339136430437180e-06
GC_8_945 b_8 NI_8 NS_945 0 -4.6974363672918852e-11
GC_8_946 b_8 NI_8 NS_946 0 -1.7787531847675571e-10
GC_8_947 b_8 NI_8 NS_947 0 1.7546083573935669e-06
GC_8_948 b_8 NI_8 NS_948 0 8.7733201070267524e-06
GC_8_949 b_8 NI_8 NS_949 0 2.2050701519323272e-06
GC_8_950 b_8 NI_8 NS_950 0 -7.0025601151918258e-06
GC_8_951 b_8 NI_8 NS_951 0 -9.0168694753762524e-06
GC_8_952 b_8 NI_8 NS_952 0 5.7743114823211253e-06
GC_8_953 b_8 NI_8 NS_953 0 4.7670671507719605e-06
GC_8_954 b_8 NI_8 NS_954 0 1.1522878135479672e-05
GC_8_955 b_8 NI_8 NS_955 0 2.4563930009413276e-05
GC_8_956 b_8 NI_8 NS_956 0 -2.1161930798522632e-05
GC_8_957 b_8 NI_8 NS_957 0 -5.7418254590187436e-09
GC_8_958 b_8 NI_8 NS_958 0 -5.6212347014438031e-09
GC_8_959 b_8 NI_8 NS_959 0 3.0635560115706536e-05
GC_8_960 b_8 NI_8 NS_960 0 7.5175044757363027e-06
GC_8_961 b_8 NI_8 NS_961 0 -2.6868652444067729e-06
GC_8_962 b_8 NI_8 NS_962 0 1.1037125073486176e-05
GC_8_963 b_8 NI_8 NS_963 0 8.0388604854908106e-06
GC_8_964 b_8 NI_8 NS_964 0 1.1978104481997498e-06
GC_8_965 b_8 NI_8 NS_965 0 1.9083139015007503e-05
GC_8_966 b_8 NI_8 NS_966 0 -2.1548979016799908e-05
GC_8_967 b_8 NI_8 NS_967 0 -6.5779392854920620e-06
GC_8_968 b_8 NI_8 NS_968 0 -7.4324860823958453e-06
GC_8_969 b_8 NI_8 NS_969 0 -5.4018424427721841e-06
GC_8_970 b_8 NI_8 NS_970 0 1.2517278037592277e-05
GC_8_971 b_8 NI_8 NS_971 0 1.6097893688849034e-05
GC_8_972 b_8 NI_8 NS_972 0 7.3673295068162372e-06
GC_8_973 b_8 NI_8 NS_973 0 5.6901722234699898e-05
GC_8_974 b_8 NI_8 NS_974 0 -1.2101213396680895e-10
GC_8_975 b_8 NI_8 NS_975 0 -2.0303491978908874e-09
GC_8_976 b_8 NI_8 NS_976 0 3.4201750446067413e-08
GC_8_977 b_8 NI_8 NS_977 0 -5.1436526914665222e-07
GC_8_978 b_8 NI_8 NS_978 0 -3.8174198707382499e-07
GC_8_979 b_8 NI_8 NS_979 0 -8.7414463221608958e-07
GC_8_980 b_8 NI_8 NS_980 0 9.5753742581416140e-06
GC_8_981 b_8 NI_8 NS_981 0 1.2647197505952552e-05
GC_8_982 b_8 NI_8 NS_982 0 -1.2046359910200124e-05
GC_8_983 b_8 NI_8 NS_983 0 -1.7539602579849068e-05
GC_8_984 b_8 NI_8 NS_984 0 8.8316937674471000e-06
GC_8_985 b_8 NI_8 NS_985 0 2.8400590124129947e-05
GC_8_986 b_8 NI_8 NS_986 0 -6.5599990940890361e-06
GC_8_987 b_8 NI_8 NS_987 0 -3.2052664594929021e-06
GC_8_988 b_8 NI_8 NS_988 0 -3.0961922312946044e-06
GC_8_989 b_8 NI_8 NS_989 0 -2.8500834762846448e-06
GC_8_990 b_8 NI_8 NS_990 0 -1.4496618354800996e-05
GC_8_991 b_8 NI_8 NS_991 0 -2.4759453261573380e-05
GC_8_992 b_8 NI_8 NS_992 0 4.0216184418300817e-05
GC_8_993 b_8 NI_8 NS_993 0 3.7734461680274470e-05
GC_8_994 b_8 NI_8 NS_994 0 -4.7031954550059869e-05
GC_8_995 b_8 NI_8 NS_995 0 -3.0428897926950825e-05
GC_8_996 b_8 NI_8 NS_996 0 -2.0940879554682338e-05
GC_8_997 b_8 NI_8 NS_997 0 3.3065735172139707e-05
GC_8_998 b_8 NI_8 NS_998 0 2.6832551784231428e-05
GC_8_999 b_8 NI_8 NS_999 0 -1.8367596890140374e-05
GC_8_1000 b_8 NI_8 NS_1000 0 -2.8794840952361264e-05
GC_8_1001 b_8 NI_8 NS_1001 0 2.1463962106819636e-05
GC_8_1002 b_8 NI_8 NS_1002 0 6.0258496476065369e-05
GC_8_1003 b_8 NI_8 NS_1003 0 -2.1175879363390152e-05
GC_8_1004 b_8 NI_8 NS_1004 0 -5.5544526407234130e-05
GC_8_1005 b_8 NI_8 NS_1005 0 -3.1396081116130613e-05
GC_8_1006 b_8 NI_8 NS_1006 0 -1.1645549923517444e-05
GC_8_1007 b_8 NI_8 NS_1007 0 2.0313321371094030e-05
GC_8_1008 b_8 NI_8 NS_1008 0 1.3869333990396011e-05
GC_8_1009 b_8 NI_8 NS_1009 0 -2.4579255791235662e-05
GC_8_1010 b_8 NI_8 NS_1010 0 -1.0925619124135592e-05
GC_8_1011 b_8 NI_8 NS_1011 0 2.0765547233160952e-05
GC_8_1012 b_8 NI_8 NS_1012 0 1.0077085389928579e-05
GC_8_1013 b_8 NI_8 NS_1013 0 -1.8224323567180912e-05
GC_8_1014 b_8 NI_8 NS_1014 0 -2.0845546888318154e-05
GC_8_1015 b_8 NI_8 NS_1015 0 5.4975824210943436e-06
GC_8_1016 b_8 NI_8 NS_1016 0 3.2160679415450316e-05
GC_8_1017 b_8 NI_8 NS_1017 0 -8.2125209333517789e-06
GC_8_1018 b_8 NI_8 NS_1018 0 -2.6520146916278293e-05
GC_8_1019 b_8 NI_8 NS_1019 0 -1.8293146455222130e-06
GC_8_1020 b_8 NI_8 NS_1020 0 1.6902885315817333e-06
GC_8_1021 b_8 NI_8 NS_1021 0 -1.9229254596406557e-05
GC_8_1022 b_8 NI_8 NS_1022 0 -1.1940103514307731e-05
GC_8_1023 b_8 NI_8 NS_1023 0 6.9725826746085411e-06
GC_8_1024 b_8 NI_8 NS_1024 0 2.0939545235772656e-05
GC_8_1025 b_8 NI_8 NS_1025 0 -1.5976405886999928e-05
GC_8_1026 b_8 NI_8 NS_1026 0 -1.4813667294286718e-05
GC_8_1027 b_8 NI_8 NS_1027 0 1.3388594832552253e-06
GC_8_1028 b_8 NI_8 NS_1028 0 5.3013248127220865e-06
GC_8_1029 b_8 NI_8 NS_1029 0 -2.4841218600445859e-05
GC_8_1030 b_8 NI_8 NS_1030 0 -9.8243626096656753e-06
GC_8_1031 b_8 NI_8 NS_1031 0 8.5462507277628255e-06
GC_8_1032 b_8 NI_8 NS_1032 0 2.3050513033619908e-05
GC_8_1033 b_8 NI_8 NS_1033 0 -2.0672693998101101e-05
GC_8_1034 b_8 NI_8 NS_1034 0 -5.6252742587896056e-06
GC_8_1035 b_8 NI_8 NS_1035 0 6.2603548142835307e-06
GC_8_1036 b_8 NI_8 NS_1036 0 7.5158350350047385e-06
GC_8_1037 b_8 NI_8 NS_1037 0 -3.0565168948302942e-05
GC_8_1038 b_8 NI_8 NS_1038 0 -2.5578178142494448e-06
GC_8_1039 b_8 NI_8 NS_1039 0 1.8794227644801613e-05
GC_8_1040 b_8 NI_8 NS_1040 0 2.5290847560590359e-05
GC_8_1041 b_8 NI_8 NS_1041 0 -2.1787413981820226e-05
GC_8_1042 b_8 NI_8 NS_1042 0 6.9645038757859913e-06
GC_8_1043 b_8 NI_8 NS_1043 0 1.5266871400115835e-05
GC_8_1044 b_8 NI_8 NS_1044 0 3.9771038840503643e-06
GC_8_1045 b_8 NI_8 NS_1045 0 -3.4533265730569028e-05
GC_8_1046 b_8 NI_8 NS_1046 0 1.3723474281250743e-05
GC_8_1047 b_8 NI_8 NS_1047 0 3.7469639958417893e-05
GC_8_1048 b_8 NI_8 NS_1048 0 1.2338009037062751e-05
GC_8_1049 b_8 NI_8 NS_1049 0 -7.7465657120511851e-06
GC_8_1050 b_8 NI_8 NS_1050 0 1.8808998254187964e-05
GC_8_1051 b_8 NI_8 NS_1051 0 1.2775019175621911e-05
GC_8_1052 b_8 NI_8 NS_1052 0 -1.1287479124834744e-05
GC_8_1053 b_8 NI_8 NS_1053 0 1.0985023350478586e-10
GC_8_1054 b_8 NI_8 NS_1054 0 3.5334379739597272e-11
GC_8_1055 b_8 NI_8 NS_1055 0 -1.3692325165810239e-05
GC_8_1056 b_8 NI_8 NS_1056 0 2.5942177910078325e-05
GC_8_1057 b_8 NI_8 NS_1057 0 -2.0633484136615916e-06
GC_8_1058 b_8 NI_8 NS_1058 0 1.0503161247881810e-05
GC_8_1059 b_8 NI_8 NS_1059 0 6.1729255244477641e-06
GC_8_1060 b_8 NI_8 NS_1060 0 -8.5364898035949855e-06
GC_8_1061 b_8 NI_8 NS_1061 0 -8.1124828689221351e-06
GC_8_1062 b_8 NI_8 NS_1062 0 2.5390671883901396e-05
GC_8_1063 b_8 NI_8 NS_1063 0 2.4973015112174624e-05
GC_8_1064 b_8 NI_8 NS_1064 0 -1.0421081391876841e-05
GC_8_1065 b_8 NI_8 NS_1065 0 4.8846452159104946e-09
GC_8_1066 b_8 NI_8 NS_1066 0 -1.2242819436785700e-09
GC_8_1067 b_8 NI_8 NS_1067 0 2.6368704308076974e-05
GC_8_1068 b_8 NI_8 NS_1068 0 -1.2610269208584276e-05
GC_8_1069 b_8 NI_8 NS_1069 0 -8.2495149921631671e-06
GC_8_1070 b_8 NI_8 NS_1070 0 1.8114668642208773e-05
GC_8_1071 b_8 NI_8 NS_1071 0 -1.0378170863178244e-05
GC_8_1072 b_8 NI_8 NS_1072 0 -3.0217641234753045e-07
GC_8_1073 b_8 NI_8 NS_1073 0 1.9390226143353015e-05
GC_8_1074 b_8 NI_8 NS_1074 0 -1.4389078693484807e-05
GC_8_1075 b_8 NI_8 NS_1075 0 7.1949278675940190e-06
GC_8_1076 b_8 NI_8 NS_1076 0 1.1599497490776776e-05
GC_8_1077 b_8 NI_8 NS_1077 0 -2.2868233619537970e-07
GC_8_1078 b_8 NI_8 NS_1078 0 -1.4637668239716117e-05
GC_8_1079 b_8 NI_8 NS_1079 0 1.3160347761058939e-05
GC_8_1080 b_8 NI_8 NS_1080 0 2.7988961085857271e-05
GC_8_1081 b_8 NI_8 NS_1081 0 -1.5116578292907588e-04
GC_8_1082 b_8 NI_8 NS_1082 0 3.7546773408545184e-11
GC_8_1083 b_8 NI_8 NS_1083 0 1.7613689229908914e-11
GC_8_1084 b_8 NI_8 NS_1084 0 8.7391547346102015e-10
GC_8_1085 b_8 NI_8 NS_1085 0 -2.3302368727450964e-06
GC_8_1086 b_8 NI_8 NS_1086 0 -1.6501405799907008e-06
GC_8_1087 b_8 NI_8 NS_1087 0 1.4541338000362102e-06
GC_8_1088 b_8 NI_8 NS_1088 0 3.8965286645506939e-06
GC_8_1089 b_8 NI_8 NS_1089 0 2.9654764339535484e-06
GC_8_1090 b_8 NI_8 NS_1090 0 5.4214068528188574e-06
GC_8_1091 b_8 NI_8 NS_1091 0 5.3772552094806114e-06
GC_8_1092 b_8 NI_8 NS_1092 0 -8.4804552529554119e-06
GC_8_1093 b_8 NI_8 NS_1093 0 -2.2507482155869561e-06
GC_8_1094 b_8 NI_8 NS_1094 0 -1.2662235754551318e-05
GC_8_1095 b_8 NI_8 NS_1095 0 -3.7273768695479633e-06
GC_8_1096 b_8 NI_8 NS_1096 0 2.7450756072030121e-06
GC_8_1097 b_8 NI_8 NS_1097 0 4.4941470889546057e-06
GC_8_1098 b_8 NI_8 NS_1098 0 1.5803601763117893e-06
GC_8_1099 b_8 NI_8 NS_1099 0 8.5385429008253462e-06
GC_8_1100 b_8 NI_8 NS_1100 0 -3.8252064403339113e-05
GC_8_1101 b_8 NI_8 NS_1101 0 -4.2843506330045589e-05
GC_8_1102 b_8 NI_8 NS_1102 0 -1.4539738280627441e-06
GC_8_1103 b_8 NI_8 NS_1103 0 -1.4647321671212984e-05
GC_8_1104 b_8 NI_8 NS_1104 0 -8.2775488446371938e-06
GC_8_1105 b_8 NI_8 NS_1105 0 -7.0243415011378261e-05
GC_8_1106 b_8 NI_8 NS_1106 0 7.5185373052606228e-05
GC_8_1107 b_8 NI_8 NS_1107 0 4.8693910332070745e-06
GC_8_1108 b_8 NI_8 NS_1108 0 1.3024069957438032e-05
GC_8_1109 b_8 NI_8 NS_1109 0 6.5219389258840249e-05
GC_8_1110 b_8 NI_8 NS_1110 0 1.2202119012709182e-04
GC_8_1111 b_8 NI_8 NS_1111 0 -2.7583336906281945e-07
GC_8_1112 b_8 NI_8 NS_1112 0 -3.7368601349371732e-05
GC_8_1113 b_8 NI_8 NS_1113 0 1.6806380366035555e-05
GC_8_1114 b_8 NI_8 NS_1114 0 4.1838901850126294e-06
GC_8_1115 b_8 NI_8 NS_1115 0 2.5158699200995393e-05
GC_8_1116 b_8 NI_8 NS_1116 0 -3.0985675094655683e-05
GC_8_1117 b_8 NI_8 NS_1117 0 -8.5164686258604183e-06
GC_8_1118 b_8 NI_8 NS_1118 0 -2.5732809379440692e-06
GC_8_1119 b_8 NI_8 NS_1119 0 -8.0804277344840986e-06
GC_8_1120 b_8 NI_8 NS_1120 0 2.4256609943807490e-05
GC_8_1121 b_8 NI_8 NS_1121 0 6.0403101074231962e-06
GC_8_1122 b_8 NI_8 NS_1122 0 8.3878806810714611e-06
GC_8_1123 b_8 NI_8 NS_1123 0 5.7350641695724164e-05
GC_8_1124 b_8 NI_8 NS_1124 0 2.3736431325358169e-05
GC_8_1125 b_8 NI_8 NS_1125 0 3.5345618442382057e-06
GC_8_1126 b_8 NI_8 NS_1126 0 -1.2244040689402119e-05
GC_8_1127 b_8 NI_8 NS_1127 0 -7.4192211421473117e-08
GC_8_1128 b_8 NI_8 NS_1128 0 -1.3740254268568609e-06
GC_8_1129 b_8 NI_8 NS_1129 0 7.1802180880760278e-06
GC_8_1130 b_8 NI_8 NS_1130 0 2.7778761625266769e-06
GC_8_1131 b_8 NI_8 NS_1131 0 4.2416637362733929e-05
GC_8_1132 b_8 NI_8 NS_1132 0 -1.9012301542805821e-05
GC_8_1133 b_8 NI_8 NS_1133 0 -2.5057990506521963e-06
GC_8_1134 b_8 NI_8 NS_1134 0 -7.6312045984306559e-06
GC_8_1135 b_8 NI_8 NS_1135 0 -2.8031960760784652e-06
GC_8_1136 b_8 NI_8 NS_1136 0 1.0883859983538483e-06
GC_8_1137 b_8 NI_8 NS_1137 0 9.8313754423913632e-06
GC_8_1138 b_8 NI_8 NS_1138 0 2.5417290751212789e-06
GC_8_1139 b_8 NI_8 NS_1139 0 2.2415809203385402e-05
GC_8_1140 b_8 NI_8 NS_1140 0 -3.3139167121608181e-05
GC_8_1141 b_8 NI_8 NS_1141 0 -5.7255922281304711e-06
GC_8_1142 b_8 NI_8 NS_1142 0 -4.2015261251419790e-06
GC_8_1143 b_8 NI_8 NS_1143 0 -8.8987750649266219e-07
GC_8_1144 b_8 NI_8 NS_1144 0 4.2524697463421603e-06
GC_8_1145 b_8 NI_8 NS_1145 0 1.2480177626981187e-05
GC_8_1146 b_8 NI_8 NS_1146 0 -2.7949776519837514e-07
GC_8_1147 b_8 NI_8 NS_1147 0 4.7396010513989109e-07
GC_8_1148 b_8 NI_8 NS_1148 0 -3.2834662825340429e-05
GC_8_1149 b_8 NI_8 NS_1149 0 -6.9268197909284865e-06
GC_8_1150 b_8 NI_8 NS_1150 0 4.0684788043564599e-07
GC_8_1151 b_8 NI_8 NS_1151 0 3.8410642257109424e-06
GC_8_1152 b_8 NI_8 NS_1152 0 3.5676544395288592e-06
GC_8_1153 b_8 NI_8 NS_1153 0 1.4108455476504448e-05
GC_8_1154 b_8 NI_8 NS_1154 0 -6.6872319521418035e-06
GC_8_1155 b_8 NI_8 NS_1155 0 -1.5604802671619446e-05
GC_8_1156 b_8 NI_8 NS_1156 0 -1.9003612100759633e-05
GC_8_1157 b_8 NI_8 NS_1157 0 -2.9952190864105451e-06
GC_8_1158 b_8 NI_8 NS_1158 0 5.1042659168480706e-06
GC_8_1159 b_8 NI_8 NS_1159 0 4.2096737234037257e-06
GC_8_1160 b_8 NI_8 NS_1160 0 -1.8809873155290637e-06
GC_8_1161 b_8 NI_8 NS_1161 0 -2.7916063629710387e-11
GC_8_1162 b_8 NI_8 NS_1162 0 5.8158869804658266e-12
GC_8_1163 b_8 NI_8 NS_1163 0 4.8698608293622767e-06
GC_8_1164 b_8 NI_8 NS_1164 0 -1.1668132756184000e-05
GC_8_1165 b_8 NI_8 NS_1165 0 -5.0905766263651410e-07
GC_8_1166 b_8 NI_8 NS_1166 0 2.7992517191271374e-06
GC_8_1167 b_8 NI_8 NS_1167 0 2.3509246519691581e-06
GC_8_1168 b_8 NI_8 NS_1168 0 -1.5716513757587633e-06
GC_8_1169 b_8 NI_8 NS_1169 0 2.1314065912552961e-06
GC_8_1170 b_8 NI_8 NS_1170 0 -9.8974346559377429e-06
GC_8_1171 b_8 NI_8 NS_1171 0 -1.0613651051088620e-05
GC_8_1172 b_8 NI_8 NS_1172 0 -3.5263093768165573e-06
GC_8_1173 b_8 NI_8 NS_1173 0 -2.3907019582353944e-10
GC_8_1174 b_8 NI_8 NS_1174 0 4.4566934989896017e-10
GC_8_1175 b_8 NI_8 NS_1175 0 -9.1766904785067173e-06
GC_8_1176 b_8 NI_8 NS_1176 0 -5.6138362671568484e-06
GC_8_1177 b_8 NI_8 NS_1177 0 1.9952213416829358e-06
GC_8_1178 b_8 NI_8 NS_1178 0 -6.7132233631998266e-06
GC_8_1179 b_8 NI_8 NS_1179 0 -3.3605963503343478e-06
GC_8_1180 b_8 NI_8 NS_1180 0 -1.7941019693921135e-07
GC_8_1181 b_8 NI_8 NS_1181 0 -8.5928669258722031e-06
GC_8_1182 b_8 NI_8 NS_1182 0 5.9560211267403282e-07
GC_8_1183 b_8 NI_8 NS_1183 0 2.6078670348732246e-06
GC_8_1184 b_8 NI_8 NS_1184 0 2.8393330926642202e-06
GC_8_1185 b_8 NI_8 NS_1185 0 9.9244062586401734e-07
GC_8_1186 b_8 NI_8 NS_1186 0 -3.6889586660117102e-06
GC_8_1187 b_8 NI_8 NS_1187 0 -5.4153742151816157e-06
GC_8_1188 b_8 NI_8 NS_1188 0 -4.2328073567166690e-06
GC_8_1189 b_8 NI_8 NS_1189 0 -5.1646794666512383e-05
GC_8_1190 b_8 NI_8 NS_1190 0 -7.9566915510117766e-12
GC_8_1191 b_8 NI_8 NS_1191 0 -2.0642359462071570e-10
GC_8_1192 b_8 NI_8 NS_1192 0 9.8399898188375934e-09
GC_8_1193 b_8 NI_8 NS_1193 0 5.5721844989526019e-07
GC_8_1194 b_8 NI_8 NS_1194 0 5.0159590713096275e-08
GC_8_1195 b_8 NI_8 NS_1195 0 2.9182992135186413e-06
GC_8_1196 b_8 NI_8 NS_1196 0 -1.4785625960902526e-06
GC_8_1197 b_8 NI_8 NS_1197 0 -3.1221351145168077e-06
GC_8_1198 b_8 NI_8 NS_1198 0 -2.6253129677475220e-06
GC_8_1199 b_8 NI_8 NS_1199 0 4.5600550910977048e-06
GC_8_1200 b_8 NI_8 NS_1200 0 -4.1953988439605065e-07
GC_8_1201 b_8 NI_8 NS_1201 0 -7.3317357999927205e-06
GC_8_1202 b_8 NI_8 NS_1202 0 -7.4847503068486345e-06
GC_8_1203 b_8 NI_8 NS_1203 0 -2.4481668723586044e-07
GC_8_1204 b_8 NI_8 NS_1204 0 -1.3835222177170756e-06
GC_8_1205 b_8 NI_8 NS_1205 0 -5.8631656126871328e-06
GC_8_1206 b_8 NI_8 NS_1206 0 2.4072495361923689e-06
GC_8_1207 b_8 NI_8 NS_1207 0 5.0674514058068607e-06
GC_8_1208 b_8 NI_8 NS_1208 0 -5.0233992403471512e-06
GC_8_1209 b_8 NI_8 NS_1209 0 -1.6437325917166785e-05
GC_8_1210 b_8 NI_8 NS_1210 0 4.9721643273290921e-06
GC_8_1211 b_8 NI_8 NS_1211 0 -1.1936072948299605e-06
GC_8_1212 b_8 NI_8 NS_1212 0 7.3470965646782847e-06
GC_8_1213 b_8 NI_8 NS_1213 0 -6.5660733378204233e-06
GC_8_1214 b_8 NI_8 NS_1214 0 -3.8974729409905644e-06
GC_8_1215 b_8 NI_8 NS_1215 0 -3.2508502593184511e-06
GC_8_1216 b_8 NI_8 NS_1216 0 8.1592787430836238e-06
GC_8_1217 b_8 NI_8 NS_1217 0 -1.3863279942670564e-06
GC_8_1218 b_8 NI_8 NS_1218 0 -3.8634309997736837e-06
GC_8_1219 b_8 NI_8 NS_1219 0 -3.9088390714711643e-06
GC_8_1220 b_8 NI_8 NS_1220 0 1.1192659993417064e-05
GC_8_1221 b_8 NI_8 NS_1221 0 -1.0533516797335881e-07
GC_8_1222 b_8 NI_8 NS_1222 0 7.4969856528519335e-06
GC_8_1223 b_8 NI_8 NS_1223 0 -3.5950146782043827e-06
GC_8_1224 b_8 NI_8 NS_1224 0 1.5343056865398140e-06
GC_8_1225 b_8 NI_8 NS_1225 0 -4.2006651583756872e-07
GC_8_1226 b_8 NI_8 NS_1226 0 8.2501959207116159e-06
GC_8_1227 b_8 NI_8 NS_1227 0 -5.3672290699967248e-07
GC_8_1228 b_8 NI_8 NS_1228 0 2.2139596231731688e-06
GC_8_1229 b_8 NI_8 NS_1229 0 -2.2958979911232970e-06
GC_8_1230 b_8 NI_8 NS_1230 0 8.3126793789984176e-06
GC_8_1231 b_8 NI_8 NS_1231 0 6.2644668820497287e-07
GC_8_1232 b_8 NI_8 NS_1232 0 9.9677224134399762e-06
GC_8_1233 b_8 NI_8 NS_1233 0 -6.6638651277909378e-07
GC_8_1234 b_8 NI_8 NS_1234 0 8.7834119953533695e-06
GC_8_1235 b_8 NI_8 NS_1235 0 -1.2310800098916309e-06
GC_8_1236 b_8 NI_8 NS_1236 0 4.0450381657636236e-06
GC_8_1237 b_8 NI_8 NS_1237 0 1.2531594277236880e-06
GC_8_1238 b_8 NI_8 NS_1238 0 1.2151059542659122e-05
GC_8_1239 b_8 NI_8 NS_1239 0 1.8598606547261168e-05
GC_8_1240 b_8 NI_8 NS_1240 0 1.6955555723717928e-05
GC_8_1241 b_8 NI_8 NS_1241 0 4.9927745967830079e-06
GC_8_1242 b_8 NI_8 NS_1242 0 7.7348606953901600e-06
GC_8_1243 b_8 NI_8 NS_1243 0 1.0287804914393564e-05
GC_8_1244 b_8 NI_8 NS_1244 0 3.8686392852920068e-06
GC_8_1245 b_8 NI_8 NS_1245 0 6.7815816057385929e-06
GC_8_1246 b_8 NI_8 NS_1246 0 1.0888476652163074e-05
GC_8_1247 b_8 NI_8 NS_1247 0 3.3297997022294209e-05
GC_8_1248 b_8 NI_8 NS_1248 0 -6.1160188985235537e-06
GC_8_1249 b_8 NI_8 NS_1249 0 8.1345733110466286e-06
GC_8_1250 b_8 NI_8 NS_1250 0 3.3940891790671715e-06
GC_8_1251 b_8 NI_8 NS_1251 0 1.1919583791541920e-05
GC_8_1252 b_8 NI_8 NS_1252 0 -1.0263713578753234e-05
GC_8_1253 b_8 NI_8 NS_1253 0 1.0740952396971787e-05
GC_8_1254 b_8 NI_8 NS_1254 0 6.4520281090498001e-06
GC_8_1255 b_8 NI_8 NS_1255 0 1.6864072825719078e-05
GC_8_1256 b_8 NI_8 NS_1256 0 -3.0725039335417161e-05
GC_8_1257 b_8 NI_8 NS_1257 0 8.0822544583331121e-06
GC_8_1258 b_8 NI_8 NS_1258 0 -2.9351848037081178e-06
GC_8_1259 b_8 NI_8 NS_1259 0 -3.2232094595058498e-06
GC_8_1260 b_8 NI_8 NS_1260 0 -1.6225074518073567e-05
GC_8_1261 b_8 NI_8 NS_1261 0 1.1764426946159312e-05
GC_8_1262 b_8 NI_8 NS_1262 0 -1.6046712888120811e-06
GC_8_1263 b_8 NI_8 NS_1263 0 -1.2697691027377807e-05
GC_8_1264 b_8 NI_8 NS_1264 0 -2.5038899722243241e-05
GC_8_1265 b_8 NI_8 NS_1265 0 -1.6043446731099470e-07
GC_8_1266 b_8 NI_8 NS_1266 0 -6.5987142141084813e-06
GC_8_1267 b_8 NI_8 NS_1267 0 -9.5600451210935713e-06
GC_8_1268 b_8 NI_8 NS_1268 0 -2.6183609173092354e-06
GC_8_1269 b_8 NI_8 NS_1269 0 1.0192258940955909e-10
GC_8_1270 b_8 NI_8 NS_1270 0 4.7260122097064714e-11
GC_8_1271 b_8 NI_8 NS_1271 0 1.4895145074962471e-06
GC_8_1272 b_8 NI_8 NS_1272 0 -4.6804883382696362e-06
GC_8_1273 b_8 NI_8 NS_1273 0 -1.3643762994802377e-06
GC_8_1274 b_8 NI_8 NS_1274 0 -1.3419853090316462e-06
GC_8_1275 b_8 NI_8 NS_1275 0 -4.8481160809990949e-06
GC_8_1276 b_8 NI_8 NS_1276 0 -9.9610102182957589e-07
GC_8_1277 b_8 NI_8 NS_1277 0 -1.1402781723946506e-06
GC_8_1278 b_8 NI_8 NS_1278 0 -2.7145520074131250e-06
GC_8_1279 b_8 NI_8 NS_1279 0 -9.9975793931318279e-06
GC_8_1280 b_8 NI_8 NS_1280 0 -4.0377359720169821e-06
GC_8_1281 b_8 NI_8 NS_1281 0 6.6624156040485003e-09
GC_8_1282 b_8 NI_8 NS_1282 0 5.4072848029121264e-09
GC_8_1283 b_8 NI_8 NS_1283 0 1.7619933875713316e-06
GC_8_1284 b_8 NI_8 NS_1284 0 4.8751331554877116e-07
GC_8_1285 b_8 NI_8 NS_1285 0 -1.6125718751221595e-06
GC_8_1286 b_8 NI_8 NS_1286 0 3.2218635699892687e-06
GC_8_1287 b_8 NI_8 NS_1287 0 -8.2907771843737805e-07
GC_8_1288 b_8 NI_8 NS_1288 0 6.9895330929204260e-07
GC_8_1289 b_8 NI_8 NS_1289 0 -7.6542254276610198e-06
GC_8_1290 b_8 NI_8 NS_1290 0 5.4120117675070776e-07
GC_8_1291 b_8 NI_8 NS_1291 0 -2.2205061720973162e-06
GC_8_1292 b_8 NI_8 NS_1292 0 1.9993208223077728e-06
GC_8_1293 b_8 NI_8 NS_1293 0 -2.0646061155641264e-06
GC_8_1294 b_8 NI_8 NS_1294 0 1.9702201981795651e-06
GC_8_1295 b_8 NI_8 NS_1295 0 1.2826138561459737e-06
GC_8_1296 b_8 NI_8 NS_1296 0 2.8349435182638205e-06
GD_8_1 b_8 NI_8 NA_1 0 1.1360095432780715e-05
GD_8_2 b_8 NI_8 NA_2 0 -2.6048127175717560e-06
GD_8_3 b_8 NI_8 NA_3 0 1.6003152016725775e-05
GD_8_4 b_8 NI_8 NA_4 0 -1.0996154956985477e-06
GD_8_5 b_8 NI_8 NA_5 0 -1.1498071994856763e-03
GD_8_6 b_8 NI_8 NA_6 0 1.0577033561008330e-02
GD_8_7 b_8 NI_8 NA_7 0 -4.9039857217504984e-03
GD_8_8 b_8 NI_8 NA_8 0 -1.1040267719203445e-02
GD_8_9 b_8 NI_8 NA_9 0 1.0462077715570234e-04
GD_8_10 b_8 NI_8 NA_10 0 2.6298651096735911e-05
GD_8_11 b_8 NI_8 NA_11 0 1.9065698154610354e-05
GD_8_12 b_8 NI_8 NA_12 0 3.1120404058041692e-06
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 8.6319383121689767e-06
GC_9_2 b_9 NI_9 NS_2 0 3.7625843103615139e-12
GC_9_3 b_9 NI_9 NS_3 0 -7.8512301742958723e-11
GC_9_4 b_9 NI_9 NS_4 0 2.5462458372855821e-09
GC_9_5 b_9 NI_9 NS_5 0 1.6079125231448565e-08
GC_9_6 b_9 NI_9 NS_6 0 -8.4902388654905115e-08
GC_9_7 b_9 NI_9 NS_7 0 -2.4705996890674441e-07
GC_9_8 b_9 NI_9 NS_8 0 2.7069013861410124e-07
GC_9_9 b_9 NI_9 NS_9 0 7.4260421400957415e-07
GC_9_10 b_9 NI_9 NS_10 0 -2.8637928135034012e-07
GC_9_11 b_9 NI_9 NS_11 0 -9.6682259458690681e-07
GC_9_12 b_9 NI_9 NS_12 0 -2.3726220472240319e-07
GC_9_13 b_9 NI_9 NS_13 0 1.0246333441339078e-06
GC_9_14 b_9 NI_9 NS_14 0 3.9650967292431843e-07
GC_9_15 b_9 NI_9 NS_15 0 -1.1998860899489725e-07
GC_9_16 b_9 NI_9 NS_16 0 -2.7403598517103499e-07
GC_9_17 b_9 NI_9 NS_17 0 1.0759569143078997e-07
GC_9_18 b_9 NI_9 NS_18 0 -5.1241337831432990e-07
GC_9_19 b_9 NI_9 NS_19 0 -2.0819725333068791e-06
GC_9_20 b_9 NI_9 NS_20 0 8.5957038177547223e-07
GC_9_21 b_9 NI_9 NS_21 0 2.4262765487128591e-06
GC_9_22 b_9 NI_9 NS_22 0 -6.0722347038911063e-07
GC_9_23 b_9 NI_9 NS_23 0 -6.6432077788056827e-07
GC_9_24 b_9 NI_9 NS_24 0 -1.3962518842334804e-06
GC_9_25 b_9 NI_9 NS_25 0 4.2621864689227025e-07
GC_9_26 b_9 NI_9 NS_26 0 1.8418687470235601e-06
GC_9_27 b_9 NI_9 NS_27 0 -3.2462319816030022e-08
GC_9_28 b_9 NI_9 NS_28 0 -1.3222091853483832e-06
GC_9_29 b_9 NI_9 NS_29 0 -6.3303759574963710e-07
GC_9_30 b_9 NI_9 NS_30 0 2.5875866080660242e-06
GC_9_31 b_9 NI_9 NS_31 0 4.5137908305712524e-07
GC_9_32 b_9 NI_9 NS_32 0 -2.2404784684585114e-06
GC_9_33 b_9 NI_9 NS_33 0 -7.9996213002072162e-07
GC_9_34 b_9 NI_9 NS_34 0 -9.3018072891235706e-07
GC_9_35 b_9 NI_9 NS_35 0 3.5769579923321463e-07
GC_9_36 b_9 NI_9 NS_36 0 9.1028071512740066e-07
GC_9_37 b_9 NI_9 NS_37 0 -5.5738544170847897e-07
GC_9_38 b_9 NI_9 NS_38 0 -7.2413000697183498e-07
GC_9_39 b_9 NI_9 NS_39 0 4.7554854534556854e-07
GC_9_40 b_9 NI_9 NS_40 0 7.3859799427512354e-07
GC_9_41 b_9 NI_9 NS_41 0 -1.7484853358379581e-07
GC_9_42 b_9 NI_9 NS_42 0 -8.7651973904873237e-07
GC_9_43 b_9 NI_9 NS_43 0 -3.3814271679472129e-07
GC_9_44 b_9 NI_9 NS_44 0 1.1560695411760450e-06
GC_9_45 b_9 NI_9 NS_45 0 2.5205996528335621e-07
GC_9_46 b_9 NI_9 NS_46 0 -8.4271728589964874e-07
GC_9_47 b_9 NI_9 NS_47 0 -6.4710168501798599e-08
GC_9_48 b_9 NI_9 NS_48 0 6.6992884094778063e-08
GC_9_49 b_9 NI_9 NS_49 0 -2.6027232955497463e-07
GC_9_50 b_9 NI_9 NS_50 0 -5.4871456024335597e-07
GC_9_51 b_9 NI_9 NS_51 0 1.8495540521298502e-07
GC_9_52 b_9 NI_9 NS_52 0 7.1500674871055694e-07
GC_9_53 b_9 NI_9 NS_53 0 -8.1315843557788796e-08
GC_9_54 b_9 NI_9 NS_54 0 -6.3403707616123697e-07
GC_9_55 b_9 NI_9 NS_55 0 1.0163401118575239e-07
GC_9_56 b_9 NI_9 NS_56 0 1.0359627899328417e-07
GC_9_57 b_9 NI_9 NS_57 0 -2.9116994154983760e-07
GC_9_58 b_9 NI_9 NS_58 0 -5.9231367966335099e-07
GC_9_59 b_9 NI_9 NS_59 0 1.5984484823034814e-07
GC_9_60 b_9 NI_9 NS_60 0 2.2926814995088421e-07
GC_9_61 b_9 NI_9 NS_61 0 -2.5752807416136031e-07
GC_9_62 b_9 NI_9 NS_62 0 -5.0661429277901950e-07
GC_9_63 b_9 NI_9 NS_63 0 4.7615638160106517e-08
GC_9_64 b_9 NI_9 NS_64 0 -4.9953157079493193e-08
GC_9_65 b_9 NI_9 NS_65 0 -3.6863297662543963e-07
GC_9_66 b_9 NI_9 NS_66 0 -5.5617336069143617e-07
GC_9_67 b_9 NI_9 NS_67 0 -2.3513418263433291e-07
GC_9_68 b_9 NI_9 NS_68 0 2.1282020402495668e-08
GC_9_69 b_9 NI_9 NS_69 0 -4.3378988076867097e-07
GC_9_70 b_9 NI_9 NS_70 0 -3.3905185406171975e-07
GC_9_71 b_9 NI_9 NS_71 0 -1.2438546651731397e-07
GC_9_72 b_9 NI_9 NS_72 0 1.6436434228457487e-08
GC_9_73 b_9 NI_9 NS_73 0 -5.6302292711778575e-07
GC_9_74 b_9 NI_9 NS_74 0 -4.3710345147345969e-07
GC_9_75 b_9 NI_9 NS_75 0 -3.1810786991683247e-07
GC_9_76 b_9 NI_9 NS_76 0 3.1491347693963997e-07
GC_9_77 b_9 NI_9 NS_77 0 -4.9916086103586235e-07
GC_9_78 b_9 NI_9 NS_78 0 3.8171571696855711e-08
GC_9_79 b_9 NI_9 NS_79 0 -1.1417710857837392e-08
GC_9_80 b_9 NI_9 NS_80 0 6.1722323163852206e-08
GC_9_81 b_9 NI_9 NS_81 0 -3.2599403648065630e-12
GC_9_82 b_9 NI_9 NS_82 0 3.2063248940036361e-12
GC_9_83 b_9 NI_9 NS_83 0 -5.7550737772572609e-07
GC_9_84 b_9 NI_9 NS_84 0 4.7702490060796627e-08
GC_9_85 b_9 NI_9 NS_85 0 -2.8964073366469688e-07
GC_9_86 b_9 NI_9 NS_86 0 1.1817130298957596e-07
GC_9_87 b_9 NI_9 NS_87 0 -6.6623357185682624e-09
GC_9_88 b_9 NI_9 NS_88 0 -6.8740889114615179e-08
GC_9_89 b_9 NI_9 NS_89 0 -6.6032151425136588e-07
GC_9_90 b_9 NI_9 NS_90 0 1.4099315115568838e-07
GC_9_91 b_9 NI_9 NS_91 0 2.8401491307966163e-08
GC_9_92 b_9 NI_9 NS_92 0 1.2370079224566411e-07
GC_9_93 b_9 NI_9 NS_93 0 -6.1319525985534601e-11
GC_9_94 b_9 NI_9 NS_94 0 1.2860118233849345e-10
GC_9_95 b_9 NI_9 NS_95 0 -3.4592661182126455e-08
GC_9_96 b_9 NI_9 NS_96 0 1.9617205390253256e-07
GC_9_97 b_9 NI_9 NS_97 0 -3.6672513582852600e-07
GC_9_98 b_9 NI_9 NS_98 0 -4.3542075340560152e-08
GC_9_99 b_9 NI_9 NS_99 0 -1.8660690712984150e-07
GC_9_100 b_9 NI_9 NS_100 0 -2.4842173628889380e-09
GC_9_101 b_9 NI_9 NS_101 0 1.9220309586561946e-07
GC_9_102 b_9 NI_9 NS_102 0 8.1574251924125913e-08
GC_9_103 b_9 NI_9 NS_103 0 -2.6531329610263406e-07
GC_9_104 b_9 NI_9 NS_104 0 3.1380266774050670e-07
GC_9_105 b_9 NI_9 NS_105 0 1.2493619038562761e-07
GC_9_106 b_9 NI_9 NS_106 0 -1.4405353252625135e-07
GC_9_107 b_9 NI_9 NS_107 0 -5.7943757793691350e-08
GC_9_108 b_9 NI_9 NS_108 0 2.3859204394691626e-07
GC_9_109 b_9 NI_9 NS_109 0 -6.4268973832438655e-05
GC_9_110 b_9 NI_9 NS_110 0 3.5608811733735932e-12
GC_9_111 b_9 NI_9 NS_111 0 5.0181470779815156e-11
GC_9_112 b_9 NI_9 NS_112 0 -1.5818286805183439e-09
GC_9_113 b_9 NI_9 NS_113 0 -1.0723767181122845e-06
GC_9_114 b_9 NI_9 NS_114 0 -1.0588516769913819e-06
GC_9_115 b_9 NI_9 NS_115 0 4.0966222370045114e-07
GC_9_116 b_9 NI_9 NS_116 0 3.5701268161210770e-07
GC_9_117 b_9 NI_9 NS_117 0 -2.2606175521006920e-06
GC_9_118 b_9 NI_9 NS_118 0 2.1080724541520204e-06
GC_9_119 b_9 NI_9 NS_119 0 -2.5321028272465404e-06
GC_9_120 b_9 NI_9 NS_120 0 -1.2387511500446026e-06
GC_9_121 b_9 NI_9 NS_121 0 1.3985074863733191e-06
GC_9_122 b_9 NI_9 NS_122 0 9.9855178263645300e-07
GC_9_123 b_9 NI_9 NS_123 0 -1.1234335140143336e-06
GC_9_124 b_9 NI_9 NS_124 0 1.3407169812091740e-06
GC_9_125 b_9 NI_9 NS_125 0 7.2718043307545175e-07
GC_9_126 b_9 NI_9 NS_126 0 3.0410638315810906e-06
GC_9_127 b_9 NI_9 NS_127 0 -2.8465210242471716e-06
GC_9_128 b_9 NI_9 NS_128 0 4.7256353817824603e-07
GC_9_129 b_9 NI_9 NS_129 0 3.6884673292179762e-06
GC_9_130 b_9 NI_9 NS_130 0 -2.0179825145791963e-06
GC_9_131 b_9 NI_9 NS_131 0 -1.8787035326470180e-07
GC_9_132 b_9 NI_9 NS_132 0 2.5631989928180776e-06
GC_9_133 b_9 NI_9 NS_133 0 -4.0642678676331408e-06
GC_9_134 b_9 NI_9 NS_134 0 4.8363275583174408e-06
GC_9_135 b_9 NI_9 NS_135 0 6.4243781730073412e-07
GC_9_136 b_9 NI_9 NS_136 0 -1.5864528594891733e-06
GC_9_137 b_9 NI_9 NS_137 0 4.6100754012492218e-06
GC_9_138 b_9 NI_9 NS_138 0 9.9431417688034680e-06
GC_9_139 b_9 NI_9 NS_139 0 -1.1102512738898258e-07
GC_9_140 b_9 NI_9 NS_140 0 5.2377553798849037e-07
GC_9_141 b_9 NI_9 NS_141 0 -6.3326477438059365e-09
GC_9_142 b_9 NI_9 NS_142 0 -7.8556209593878724e-07
GC_9_143 b_9 NI_9 NS_143 0 5.3518681477106396e-06
GC_9_144 b_9 NI_9 NS_144 0 4.9529420927014422e-07
GC_9_145 b_9 NI_9 NS_145 0 8.4638405682791566e-07
GC_9_146 b_9 NI_9 NS_146 0 1.9176013022286493e-06
GC_9_147 b_9 NI_9 NS_147 0 3.0812572357416208e-08
GC_9_148 b_9 NI_9 NS_148 0 1.1332187831024110e-06
GC_9_149 b_9 NI_9 NS_149 0 5.8507452051162455e-07
GC_9_150 b_9 NI_9 NS_150 0 -1.1108412052988983e-06
GC_9_151 b_9 NI_9 NS_151 0 5.8253731629484397e-06
GC_9_152 b_9 NI_9 NS_152 0 4.0748048078532346e-06
GC_9_153 b_9 NI_9 NS_153 0 6.0627424537070819e-07
GC_9_154 b_9 NI_9 NS_154 0 8.5952656432851220e-07
GC_9_155 b_9 NI_9 NS_155 0 1.9691787149379871e-07
GC_9_156 b_9 NI_9 NS_156 0 2.4098279403892837e-07
GC_9_157 b_9 NI_9 NS_157 0 8.4525406209373880e-07
GC_9_158 b_9 NI_9 NS_158 0 -6.7216232539348124e-07
GC_9_159 b_9 NI_9 NS_159 0 6.6650680022715593e-06
GC_9_160 b_9 NI_9 NS_160 0 7.5450001439376136e-07
GC_9_161 b_9 NI_9 NS_161 0 7.7455345781197034e-07
GC_9_162 b_9 NI_9 NS_162 0 7.4913763950816948e-07
GC_9_163 b_9 NI_9 NS_163 0 6.6483808111120954e-07
GC_9_164 b_9 NI_9 NS_164 0 -6.6192010960418920e-08
GC_9_165 b_9 NI_9 NS_165 0 8.7154930984792029e-07
GC_9_166 b_9 NI_9 NS_166 0 -6.4038523460401364e-07
GC_9_167 b_9 NI_9 NS_167 0 5.7752035409058771e-06
GC_9_168 b_9 NI_9 NS_168 0 -1.5909579004649881e-06
GC_9_169 b_9 NI_9 NS_169 0 8.2383268143557782e-07
GC_9_170 b_9 NI_9 NS_170 0 5.6703544276976561e-07
GC_9_171 b_9 NI_9 NS_171 0 6.2584752106258432e-07
GC_9_172 b_9 NI_9 NS_172 0 -5.5331126512951171e-07
GC_9_173 b_9 NI_9 NS_173 0 9.3777214075065234e-07
GC_9_174 b_9 NI_9 NS_174 0 -4.4580594499758347e-07
GC_9_175 b_9 NI_9 NS_175 0 3.9036527975080192e-06
GC_9_176 b_9 NI_9 NS_176 0 -2.9906976924276734e-06
GC_9_177 b_9 NI_9 NS_177 0 8.9571159853093252e-07
GC_9_178 b_9 NI_9 NS_178 0 3.2738015239698209e-07
GC_9_179 b_9 NI_9 NS_179 0 2.1611045769566047e-07
GC_9_180 b_9 NI_9 NS_180 0 -7.9556613937681483e-07
GC_9_181 b_9 NI_9 NS_181 0 1.1598922327421579e-06
GC_9_182 b_9 NI_9 NS_182 0 -3.2475017577326960e-07
GC_9_183 b_9 NI_9 NS_183 0 1.6774700532449030e-06
GC_9_184 b_9 NI_9 NS_184 0 -3.0902010840335071e-06
GC_9_185 b_9 NI_9 NS_185 0 7.9113464065757435e-07
GC_9_186 b_9 NI_9 NS_186 0 -1.0639022406434434e-07
GC_9_187 b_9 NI_9 NS_187 0 -1.9701920410353643e-07
GC_9_188 b_9 NI_9 NS_188 0 -4.0861220854972234e-07
GC_9_189 b_9 NI_9 NS_189 0 8.5880505021837861e-12
GC_9_190 b_9 NI_9 NS_190 0 -1.5730111163015284e-11
GC_9_191 b_9 NI_9 NS_191 0 8.3871732232196766e-07
GC_9_192 b_9 NI_9 NS_192 0 -5.9378072950965052e-07
GC_9_193 b_9 NI_9 NS_193 0 4.9464383582741553e-07
GC_9_194 b_9 NI_9 NS_194 0 -3.5991688488458075e-08
GC_9_195 b_9 NI_9 NS_195 0 1.7011370475271230e-08
GC_9_196 b_9 NI_9 NS_196 0 -8.9110360549662434e-08
GC_9_197 b_9 NI_9 NS_197 0 5.2142111292827032e-07
GC_9_198 b_9 NI_9 NS_198 0 -1.7665723239274968e-08
GC_9_199 b_9 NI_9 NS_199 0 7.0517832918479781e-07
GC_9_200 b_9 NI_9 NS_200 0 -1.5613966499217453e-06
GC_9_201 b_9 NI_9 NS_201 0 4.0969093044474210e-10
GC_9_202 b_9 NI_9 NS_202 0 -5.8070565674525218e-10
GC_9_203 b_9 NI_9 NS_203 0 1.0099571759541767e-06
GC_9_204 b_9 NI_9 NS_204 0 -2.7386426453291840e-07
GC_9_205 b_9 NI_9 NS_205 0 3.5400776289230581e-07
GC_9_206 b_9 NI_9 NS_206 0 -1.7369737280795063e-07
GC_9_207 b_9 NI_9 NS_207 0 2.5492753439939549e-07
GC_9_208 b_9 NI_9 NS_208 0 2.6554657336933125e-08
GC_9_209 b_9 NI_9 NS_209 0 1.0857954102463385e-06
GC_9_210 b_9 NI_9 NS_210 0 -1.1750248170863178e-06
GC_9_211 b_9 NI_9 NS_211 0 6.5375735792921663e-07
GC_9_212 b_9 NI_9 NS_212 0 -3.3455157774406295e-07
GC_9_213 b_9 NI_9 NS_213 0 -2.1221532316237273e-07
GC_9_214 b_9 NI_9 NS_214 0 -9.8558344386953799e-08
GC_9_215 b_9 NI_9 NS_215 0 7.5732163503027058e-07
GC_9_216 b_9 NI_9 NS_216 0 3.2283769143031115e-07
GC_9_217 b_9 NI_9 NS_217 0 3.7776793059158761e-05
GC_9_218 b_9 NI_9 NS_218 0 1.2388387498661432e-12
GC_9_219 b_9 NI_9 NS_219 0 -8.1189421476233326e-12
GC_9_220 b_9 NI_9 NS_220 0 3.0025156656481305e-09
GC_9_221 b_9 NI_9 NS_221 0 3.6864096140477088e-07
GC_9_222 b_9 NI_9 NS_222 0 9.8384375208727129e-08
GC_9_223 b_9 NI_9 NS_223 0 6.5834108424835108e-07
GC_9_224 b_9 NI_9 NS_224 0 3.5826323196178347e-07
GC_9_225 b_9 NI_9 NS_225 0 1.2346444828719008e-06
GC_9_226 b_9 NI_9 NS_226 0 -8.6742584047711034e-07
GC_9_227 b_9 NI_9 NS_227 0 7.8270821732259217e-07
GC_9_228 b_9 NI_9 NS_228 0 -5.3020285813964240e-07
GC_9_229 b_9 NI_9 NS_229 0 8.2388488451075353e-07
GC_9_230 b_9 NI_9 NS_230 0 -2.1816060755568735e-06
GC_9_231 b_9 NI_9 NS_231 0 6.7227948741547858e-07
GC_9_232 b_9 NI_9 NS_232 0 -8.4321342257758818e-07
GC_9_233 b_9 NI_9 NS_233 0 -1.1291327394520202e-06
GC_9_234 b_9 NI_9 NS_234 0 -1.5078929035092817e-06
GC_9_235 b_9 NI_9 NS_235 0 -4.8950885484672692e-07
GC_9_236 b_9 NI_9 NS_236 0 -2.1010055549630162e-06
GC_9_237 b_9 NI_9 NS_237 0 -1.7840769191436358e-06
GC_9_238 b_9 NI_9 NS_238 0 -6.5666044625133552e-07
GC_9_239 b_9 NI_9 NS_239 0 -5.8884157148688778e-07
GC_9_240 b_9 NI_9 NS_240 0 -1.1663525112834538e-06
GC_9_241 b_9 NI_9 NS_241 0 -2.5818289991119619e-06
GC_9_242 b_9 NI_9 NS_242 0 -7.0827744473402031e-07
GC_9_243 b_9 NI_9 NS_243 0 -7.1488910397717744e-07
GC_9_244 b_9 NI_9 NS_244 0 -6.2489467981221662e-07
GC_9_245 b_9 NI_9 NS_245 0 -3.5725257144444890e-06
GC_9_246 b_9 NI_9 NS_246 0 -4.6960489232952820e-07
GC_9_247 b_9 NI_9 NS_247 0 2.3206992262364214e-07
GC_9_248 b_9 NI_9 NS_248 0 -2.1170858963077545e-07
GC_9_249 b_9 NI_9 NS_249 0 -9.1740987651137415e-07
GC_9_250 b_9 NI_9 NS_250 0 -9.0468444035514671e-07
GC_9_251 b_9 NI_9 NS_251 0 -1.9019688796405151e-06
GC_9_252 b_9 NI_9 NS_252 0 1.9079338181215280e-07
GC_9_253 b_9 NI_9 NS_253 0 -1.1727251356695167e-06
GC_9_254 b_9 NI_9 NS_254 0 -4.8228536860679057e-07
GC_9_255 b_9 NI_9 NS_255 0 -1.3189947265032804e-06
GC_9_256 b_9 NI_9 NS_256 0 9.6811866978736451e-07
GC_9_257 b_9 NI_9 NS_257 0 -7.9967662495712040e-07
GC_9_258 b_9 NI_9 NS_258 0 -4.7983605372566410e-07
GC_9_259 b_9 NI_9 NS_259 0 -3.1176934116338781e-06
GC_9_260 b_9 NI_9 NS_260 0 3.9714448933535231e-07
GC_9_261 b_9 NI_9 NS_261 0 -6.0262007509222107e-07
GC_9_262 b_9 NI_9 NS_262 0 1.6123629798434410e-07
GC_9_263 b_9 NI_9 NS_263 0 -6.6728219895732326e-07
GC_9_264 b_9 NI_9 NS_264 0 -1.5681799310467037e-07
GC_9_265 b_9 NI_9 NS_265 0 -1.3447998348427451e-06
GC_9_266 b_9 NI_9 NS_266 0 -7.5295134716512393e-08
GC_9_267 b_9 NI_9 NS_267 0 -3.0787569088162543e-06
GC_9_268 b_9 NI_9 NS_268 0 2.3443937154252810e-06
GC_9_269 b_9 NI_9 NS_269 0 -7.5438808434588358e-07
GC_9_270 b_9 NI_9 NS_270 0 3.5807973517605594e-07
GC_9_271 b_9 NI_9 NS_271 0 -8.0000269046748477e-07
GC_9_272 b_9 NI_9 NS_272 0 1.0728589591953658e-06
GC_9_273 b_9 NI_9 NS_273 0 -1.2382200312892323e-06
GC_9_274 b_9 NI_9 NS_274 0 1.6928107977453573e-07
GC_9_275 b_9 NI_9 NS_275 0 -1.0795274282556417e-06
GC_9_276 b_9 NI_9 NS_276 0 3.5773163085495202e-06
GC_9_277 b_9 NI_9 NS_277 0 -6.8450354945262966e-07
GC_9_278 b_9 NI_9 NS_278 0 4.6096066426239952e-07
GC_9_279 b_9 NI_9 NS_279 0 1.7787792485276478e-07
GC_9_280 b_9 NI_9 NS_280 0 1.4971790750980267e-06
GC_9_281 b_9 NI_9 NS_281 0 -1.1956615221775686e-06
GC_9_282 b_9 NI_9 NS_282 0 3.1705710691171730e-07
GC_9_283 b_9 NI_9 NS_283 0 9.5833922079459183e-07
GC_9_284 b_9 NI_9 NS_284 0 3.0173142727059990e-06
GC_9_285 b_9 NI_9 NS_285 0 -5.5639873335740708e-07
GC_9_286 b_9 NI_9 NS_286 0 6.1271405495831585e-07
GC_9_287 b_9 NI_9 NS_287 0 1.0073495239800170e-06
GC_9_288 b_9 NI_9 NS_288 0 8.4909695380614445e-07
GC_9_289 b_9 NI_9 NS_289 0 -1.1354680794339095e-06
GC_9_290 b_9 NI_9 NS_290 0 5.7364291894271997e-07
GC_9_291 b_9 NI_9 NS_291 0 1.7677963202681086e-06
GC_9_292 b_9 NI_9 NS_292 0 1.3974325455662546e-06
GC_9_293 b_9 NI_9 NS_293 0 -1.4090581337468607e-07
GC_9_294 b_9 NI_9 NS_294 0 6.5189410162294185e-07
GC_9_295 b_9 NI_9 NS_295 0 6.9857723477036288e-07
GC_9_296 b_9 NI_9 NS_296 0 -1.8042707923041638e-08
GC_9_297 b_9 NI_9 NS_297 0 2.1846692109162719e-11
GC_9_298 b_9 NI_9 NS_298 0 1.4146797539594427e-11
GC_9_299 b_9 NI_9 NS_299 0 -5.3445526427249712e-07
GC_9_300 b_9 NI_9 NS_300 0 6.6480557333264759e-07
GC_9_301 b_9 NI_9 NS_301 0 -1.6746126984844937e-08
GC_9_302 b_9 NI_9 NS_302 0 3.0212499387548956e-07
GC_9_303 b_9 NI_9 NS_303 0 2.1121858407397158e-07
GC_9_304 b_9 NI_9 NS_304 0 1.5832844038768925e-07
GC_9_305 b_9 NI_9 NS_305 0 -1.8419973012270505e-07
GC_9_306 b_9 NI_9 NS_306 0 5.6372911611541835e-07
GC_9_307 b_9 NI_9 NS_307 0 8.6158165321880489e-07
GC_9_308 b_9 NI_9 NS_308 0 4.0477746253451237e-07
GC_9_309 b_9 NI_9 NS_309 0 7.9125258963766665e-10
GC_9_310 b_9 NI_9 NS_310 0 5.1026630458007299e-10
GC_9_311 b_9 NI_9 NS_311 0 1.2590894748485795e-06
GC_9_312 b_9 NI_9 NS_312 0 1.3277660919117045e-07
GC_9_313 b_9 NI_9 NS_313 0 -1.4104368055506146e-07
GC_9_314 b_9 NI_9 NS_314 0 8.3427642969274922e-07
GC_9_315 b_9 NI_9 NS_315 0 8.2109303768951596e-08
GC_9_316 b_9 NI_9 NS_316 0 4.1437494257948261e-08
GC_9_317 b_9 NI_9 NS_317 0 3.4449309783900058e-07
GC_9_318 b_9 NI_9 NS_318 0 3.3673996544483408e-07
GC_9_319 b_9 NI_9 NS_319 0 3.0905318599837565e-07
GC_9_320 b_9 NI_9 NS_320 0 4.0930286866619064e-07
GC_9_321 b_9 NI_9 NS_321 0 6.5356327505369636e-08
GC_9_322 b_9 NI_9 NS_322 0 5.9259656048406198e-08
GC_9_323 b_9 NI_9 NS_323 0 7.1106427730296290e-07
GC_9_324 b_9 NI_9 NS_324 0 8.9929471251213676e-07
GC_9_325 b_9 NI_9 NS_325 0 -7.7897755178497040e-06
GC_9_326 b_9 NI_9 NS_326 0 -1.0504384210231227e-11
GC_9_327 b_9 NI_9 NS_327 0 7.2834305343675158e-11
GC_9_328 b_9 NI_9 NS_328 0 -4.8050177105270724e-09
GC_9_329 b_9 NI_9 NS_329 0 -9.4013969298927402e-07
GC_9_330 b_9 NI_9 NS_330 0 -7.1654523912861288e-07
GC_9_331 b_9 NI_9 NS_331 0 6.8854958059456982e-07
GC_9_332 b_9 NI_9 NS_332 0 1.1986222021131561e-06
GC_9_333 b_9 NI_9 NS_333 0 -6.6100439596982664e-07
GC_9_334 b_9 NI_9 NS_334 0 2.7641652125432837e-06
GC_9_335 b_9 NI_9 NS_335 0 -1.7497665202282307e-07
GC_9_336 b_9 NI_9 NS_336 0 -8.3646259564527563e-07
GC_9_337 b_9 NI_9 NS_337 0 3.2529126099732215e-06
GC_9_338 b_9 NI_9 NS_338 0 -1.7247914410889513e-06
GC_9_339 b_9 NI_9 NS_339 0 -2.9874406605742488e-07
GC_9_340 b_9 NI_9 NS_340 0 1.3039956725208411e-06
GC_9_341 b_9 NI_9 NS_341 0 1.3767943682889687e-06
GC_9_342 b_9 NI_9 NS_342 0 1.3767902737600688e-06
GC_9_343 b_9 NI_9 NS_343 0 2.3876606493858103e-06
GC_9_344 b_9 NI_9 NS_344 0 -3.3965039474772125e-06
GC_9_345 b_9 NI_9 NS_345 0 -2.0837819973429387e-06
GC_9_346 b_9 NI_9 NS_346 0 -6.2972585089709747e-06
GC_9_347 b_9 NI_9 NS_347 0 -1.0480082429528079e-07
GC_9_348 b_9 NI_9 NS_348 0 5.0287915235959996e-07
GC_9_349 b_9 NI_9 NS_349 0 -1.2562664484121109e-05
GC_9_350 b_9 NI_9 NS_350 0 3.3121737456051184e-06
GC_9_351 b_9 NI_9 NS_351 0 -1.5084708261694680e-07
GC_9_352 b_9 NI_9 NS_352 0 -6.4681367911661098e-07
GC_9_353 b_9 NI_9 NS_353 0 3.1495034106914135e-06
GC_9_354 b_9 NI_9 NS_354 0 1.5214634523510912e-05
GC_9_355 b_9 NI_9 NS_355 0 1.0368191831909943e-06
GC_9_356 b_9 NI_9 NS_356 0 -1.0548175863696154e-06
GC_9_357 b_9 NI_9 NS_357 0 1.1266687922505035e-06
GC_9_358 b_9 NI_9 NS_358 0 -3.1887869867129060e-07
GC_9_359 b_9 NI_9 NS_359 0 6.6856639590401625e-06
GC_9_360 b_9 NI_9 NS_360 0 -3.1044276687575103e-06
GC_9_361 b_9 NI_9 NS_361 0 3.3083090263185698e-07
GC_9_362 b_9 NI_9 NS_362 0 3.9509260934992563e-07
GC_9_363 b_9 NI_9 NS_363 0 -2.9432285754885246e-06
GC_9_364 b_9 NI_9 NS_364 0 8.3275607248522578e-07
GC_9_365 b_9 NI_9 NS_365 0 1.7555516527109533e-07
GC_9_366 b_9 NI_9 NS_366 0 -8.8267505722861004e-07
GC_9_367 b_9 NI_9 NS_367 0 6.7910587929880289e-06
GC_9_368 b_9 NI_9 NS_368 0 3.5401068494706750e-06
GC_9_369 b_9 NI_9 NS_369 0 3.3550311684064455e-07
GC_9_370 b_9 NI_9 NS_370 0 8.9039137907046030e-09
GC_9_371 b_9 NI_9 NS_371 0 2.4547534064459883e-07
GC_9_372 b_9 NI_9 NS_372 0 -6.0588451713230681e-07
GC_9_373 b_9 NI_9 NS_373 0 4.0057199029230229e-07
GC_9_374 b_9 NI_9 NS_374 0 -1.3949656546656928e-06
GC_9_375 b_9 NI_9 NS_375 0 6.0103726151808368e-06
GC_9_376 b_9 NI_9 NS_376 0 -2.3488855263706700e-06
GC_9_377 b_9 NI_9 NS_377 0 2.3332536786187373e-08
GC_9_378 b_9 NI_9 NS_378 0 -2.5588299940332057e-07
GC_9_379 b_9 NI_9 NS_379 0 -9.3826688212882049e-07
GC_9_380 b_9 NI_9 NS_380 0 -1.1597849797356862e-06
GC_9_381 b_9 NI_9 NS_381 0 3.0914674513940292e-07
GC_9_382 b_9 NI_9 NS_382 0 -1.3347759895946143e-06
GC_9_383 b_9 NI_9 NS_383 0 3.0251029869675590e-06
GC_9_384 b_9 NI_9 NS_384 0 -4.1459970243136622e-06
GC_9_385 b_9 NI_9 NS_385 0 -1.7543382277815890e-07
GC_9_386 b_9 NI_9 NS_386 0 -3.4365978919129670e-07
GC_9_387 b_9 NI_9 NS_387 0 -1.9736555184533427e-06
GC_9_388 b_9 NI_9 NS_388 0 -6.6869931604301837e-07
GC_9_389 b_9 NI_9 NS_389 0 2.0799733237903739e-07
GC_9_390 b_9 NI_9 NS_390 0 -1.4276259202841291e-06
GC_9_391 b_9 NI_9 NS_391 0 9.0915890973965364e-08
GC_9_392 b_9 NI_9 NS_392 0 -3.5637762141807373e-06
GC_9_393 b_9 NI_9 NS_393 0 -4.5635455283404521e-07
GC_9_394 b_9 NI_9 NS_394 0 -3.7736039551604835e-07
GC_9_395 b_9 NI_9 NS_395 0 -2.1515974650472914e-06
GC_9_396 b_9 NI_9 NS_396 0 5.3436247650383030e-07
GC_9_397 b_9 NI_9 NS_397 0 -6.9689873553403656e-08
GC_9_398 b_9 NI_9 NS_398 0 -1.6164296626926941e-06
GC_9_399 b_9 NI_9 NS_399 0 -1.2654800281132049e-06
GC_9_400 b_9 NI_9 NS_400 0 -1.4050915176992110e-06
GC_9_401 b_9 NI_9 NS_401 0 -8.0777186361641247e-07
GC_9_402 b_9 NI_9 NS_402 0 9.5484858608632625e-08
GC_9_403 b_9 NI_9 NS_403 0 -9.4861233090604695e-07
GC_9_404 b_9 NI_9 NS_404 0 1.0889515254061357e-06
GC_9_405 b_9 NI_9 NS_405 0 -1.7801297954637844e-11
GC_9_406 b_9 NI_9 NS_406 0 1.0630471834665305e-11
GC_9_407 b_9 NI_9 NS_407 0 -5.7532575618422243e-07
GC_9_408 b_9 NI_9 NS_408 0 -1.1642953118212305e-06
GC_9_409 b_9 NI_9 NS_409 0 -3.7975205228178491e-07
GC_9_410 b_9 NI_9 NS_410 0 2.2310881886639307e-07
GC_9_411 b_9 NI_9 NS_411 0 -5.0948352272290323e-07
GC_9_412 b_9 NI_9 NS_412 0 3.9880774207621382e-07
GC_9_413 b_9 NI_9 NS_413 0 -1.9110851818781462e-07
GC_9_414 b_9 NI_9 NS_414 0 -1.0234486491294976e-06
GC_9_415 b_9 NI_9 NS_415 0 -4.4605791238369709e-07
GC_9_416 b_9 NI_9 NS_416 0 -2.0182535310980208e-07
GC_9_417 b_9 NI_9 NS_417 0 -9.1683370650581271e-10
GC_9_418 b_9 NI_9 NS_418 0 1.5474433498851082e-10
GC_9_419 b_9 NI_9 NS_419 0 -2.2824754562418505e-07
GC_9_420 b_9 NI_9 NS_420 0 -1.9835505380535849e-07
GC_9_421 b_9 NI_9 NS_421 0 -1.7951605212935118e-07
GC_9_422 b_9 NI_9 NS_422 0 -3.4653935248410290e-07
GC_9_423 b_9 NI_9 NS_423 0 -3.9555960468929039e-07
GC_9_424 b_9 NI_9 NS_424 0 -1.3726968866999598e-07
GC_9_425 b_9 NI_9 NS_425 0 -9.9082675076481331e-07
GC_9_426 b_9 NI_9 NS_426 0 5.0307644082112362e-08
GC_9_427 b_9 NI_9 NS_427 0 -5.8387934640009407e-07
GC_9_428 b_9 NI_9 NS_428 0 4.7571068636246209e-07
GC_9_429 b_9 NI_9 NS_429 0 -1.3188452292748047e-08
GC_9_430 b_9 NI_9 NS_430 0 4.1222541935232678e-07
GC_9_431 b_9 NI_9 NS_431 0 -8.6504626112622037e-07
GC_9_432 b_9 NI_9 NS_432 0 -9.7526959576591296e-07
GC_9_433 b_9 NI_9 NS_433 0 -3.0637390258745653e-05
GC_9_434 b_9 NI_9 NS_434 0 -1.9702128922295207e-12
GC_9_435 b_9 NI_9 NS_435 0 -2.2725987935251676e-10
GC_9_436 b_9 NI_9 NS_436 0 1.0440683091420875e-08
GC_9_437 b_9 NI_9 NS_437 0 6.9327075772895857e-07
GC_9_438 b_9 NI_9 NS_438 0 1.0332693965227134e-07
GC_9_439 b_9 NI_9 NS_439 0 3.1648136551990708e-06
GC_9_440 b_9 NI_9 NS_440 0 -1.3944687587093970e-06
GC_9_441 b_9 NI_9 NS_441 0 -2.7897599395051306e-06
GC_9_442 b_9 NI_9 NS_442 0 -2.8314313765396396e-06
GC_9_443 b_9 NI_9 NS_443 0 4.9208217412362675e-06
GC_9_444 b_9 NI_9 NS_444 0 -5.3538931394146047e-07
GC_9_445 b_9 NI_9 NS_445 0 -7.0691796697171877e-06
GC_9_446 b_9 NI_9 NS_446 0 -8.1237002977537784e-06
GC_9_447 b_9 NI_9 NS_447 0 1.8606051713759501e-08
GC_9_448 b_9 NI_9 NS_448 0 -1.5534374181940269e-06
GC_9_449 b_9 NI_9 NS_449 0 -6.0814386712905951e-06
GC_9_450 b_9 NI_9 NS_450 0 1.9319035635267397e-06
GC_9_451 b_9 NI_9 NS_451 0 5.3119888684153384e-06
GC_9_452 b_9 NI_9 NS_452 0 -5.7335802720794026e-06
GC_9_453 b_9 NI_9 NS_453 0 -1.7096906214453850e-05
GC_9_454 b_9 NI_9 NS_454 0 4.6242225024036597e-06
GC_9_455 b_9 NI_9 NS_455 0 -1.1944686810243358e-06
GC_9_456 b_9 NI_9 NS_456 0 7.0592835206899497e-06
GC_9_457 b_9 NI_9 NS_457 0 -7.2285774152580770e-06
GC_9_458 b_9 NI_9 NS_458 0 -4.5688871340496629e-06
GC_9_459 b_9 NI_9 NS_459 0 -3.3893053534737101e-06
GC_9_460 b_9 NI_9 NS_460 0 7.9766987742465969e-06
GC_9_461 b_9 NI_9 NS_461 0 -2.2427661929853413e-06
GC_9_462 b_9 NI_9 NS_462 0 -4.6665000747328514e-06
GC_9_463 b_9 NI_9 NS_463 0 -3.8807669557381958e-06
GC_9_464 b_9 NI_9 NS_464 0 1.1289712317303322e-05
GC_9_465 b_9 NI_9 NS_465 0 -1.9128086870098292e-07
GC_9_466 b_9 NI_9 NS_466 0 7.1636505475757842e-06
GC_9_467 b_9 NI_9 NS_467 0 -4.1441825791170350e-06
GC_9_468 b_9 NI_9 NS_468 0 1.2150895285208924e-06
GC_9_469 b_9 NI_9 NS_469 0 -6.4403629797339984e-07
GC_9_470 b_9 NI_9 NS_470 0 7.9591241556368631e-06
GC_9_471 b_9 NI_9 NS_471 0 -1.0603802441712649e-06
GC_9_472 b_9 NI_9 NS_472 0 2.1884900028547649e-06
GC_9_473 b_9 NI_9 NS_473 0 -2.4285512724725666e-06
GC_9_474 b_9 NI_9 NS_474 0 8.0706354233291110e-06
GC_9_475 b_9 NI_9 NS_475 0 -1.7503960537922478e-07
GC_9_476 b_9 NI_9 NS_476 0 9.4003712245883445e-06
GC_9_477 b_9 NI_9 NS_477 0 -8.8143827315388563e-07
GC_9_478 b_9 NI_9 NS_478 0 8.6988676273124995e-06
GC_9_479 b_9 NI_9 NS_479 0 -1.3355221743032494e-06
GC_9_480 b_9 NI_9 NS_480 0 3.8589146976407710e-06
GC_9_481 b_9 NI_9 NS_481 0 9.5135058797662191e-07
GC_9_482 b_9 NI_9 NS_482 0 1.1830488778823846e-05
GC_9_483 b_9 NI_9 NS_483 0 1.7339678797240731e-05
GC_9_484 b_9 NI_9 NS_484 0 1.6620957308255897e-05
GC_9_485 b_9 NI_9 NS_485 0 4.6876736494517663e-06
GC_9_486 b_9 NI_9 NS_486 0 7.6215653602616897e-06
GC_9_487 b_9 NI_9 NS_487 0 9.8092201296377697e-06
GC_9_488 b_9 NI_9 NS_488 0 3.8277640482981294e-06
GC_9_489 b_9 NI_9 NS_489 0 6.4308510021047979e-06
GC_9_490 b_9 NI_9 NS_490 0 1.0600263064961318e-05
GC_9_491 b_9 NI_9 NS_491 0 3.1894622300475022e-05
GC_9_492 b_9 NI_9 NS_492 0 -5.8207807636128487e-06
GC_9_493 b_9 NI_9 NS_493 0 7.7815650272817109e-06
GC_9_494 b_9 NI_9 NS_494 0 3.3341157194248052e-06
GC_9_495 b_9 NI_9 NS_495 0 1.1392291086949541e-05
GC_9_496 b_9 NI_9 NS_496 0 -9.9543852558921988e-06
GC_9_497 b_9 NI_9 NS_497 0 1.0335937958678393e-05
GC_9_498 b_9 NI_9 NS_498 0 6.2186470346401225e-06
GC_9_499 b_9 NI_9 NS_499 0 1.5858030035394574e-05
GC_9_500 b_9 NI_9 NS_500 0 -2.9884766570321333e-05
GC_9_501 b_9 NI_9 NS_501 0 7.7006040061302838e-06
GC_9_502 b_9 NI_9 NS_502 0 -2.8908265031752880e-06
GC_9_503 b_9 NI_9 NS_503 0 -3.4539416534743921e-06
GC_9_504 b_9 NI_9 NS_504 0 -1.5715634424896563e-05
GC_9_505 b_9 NI_9 NS_505 0 1.1293336772111315e-05
GC_9_506 b_9 NI_9 NS_506 0 -1.7359447748475528e-06
GC_9_507 b_9 NI_9 NS_507 0 -1.3020290219530934e-05
GC_9_508 b_9 NI_9 NS_508 0 -2.4148618105014092e-05
GC_9_509 b_9 NI_9 NS_509 0 -4.2214980552864209e-07
GC_9_510 b_9 NI_9 NS_510 0 -6.3952476250105969e-06
GC_9_511 b_9 NI_9 NS_511 0 -9.5214716047993739e-06
GC_9_512 b_9 NI_9 NS_512 0 -2.3393118156211000e-06
GC_9_513 b_9 NI_9 NS_513 0 9.7737450807189109e-11
GC_9_514 b_9 NI_9 NS_514 0 5.3682968097319237e-11
GC_9_515 b_9 NI_9 NS_515 0 1.1864487812216120e-06
GC_9_516 b_9 NI_9 NS_516 0 -4.6217718853373054e-06
GC_9_517 b_9 NI_9 NS_517 0 -1.4846153495081745e-06
GC_9_518 b_9 NI_9 NS_518 0 -1.2851850047218688e-06
GC_9_519 b_9 NI_9 NS_519 0 -4.9361112590830248e-06
GC_9_520 b_9 NI_9 NS_520 0 -8.7754697161409676e-07
GC_9_521 b_9 NI_9 NS_521 0 -1.3873432706784373e-06
GC_9_522 b_9 NI_9 NS_522 0 -2.8331814892647540e-06
GC_9_523 b_9 NI_9 NS_523 0 -1.0078501326314437e-05
GC_9_524 b_9 NI_9 NS_524 0 -3.6998808006242207e-06
GC_9_525 b_9 NI_9 NS_525 0 6.6046402380156052e-09
GC_9_526 b_9 NI_9 NS_526 0 5.7463000433130731e-09
GC_9_527 b_9 NI_9 NS_527 0 1.3894889417729582e-06
GC_9_528 b_9 NI_9 NS_528 0 6.7846017556909592e-07
GC_9_529 b_9 NI_9 NS_529 0 -1.7344558979559085e-06
GC_9_530 b_9 NI_9 NS_530 0 3.1417316171108086e-06
GC_9_531 b_9 NI_9 NS_531 0 -9.2518103183885618e-07
GC_9_532 b_9 NI_9 NS_532 0 7.7635647951149957e-07
GC_9_533 b_9 NI_9 NS_533 0 -7.9006817086351804e-06
GC_9_534 b_9 NI_9 NS_534 0 8.1641424483464110e-07
GC_9_535 b_9 NI_9 NS_535 0 -2.4105963279546957e-06
GC_9_536 b_9 NI_9 NS_536 0 2.0859203883758027e-06
GC_9_537 b_9 NI_9 NS_537 0 -2.1253694461879582e-06
GC_9_538 b_9 NI_9 NS_538 0 2.1337376796243204e-06
GC_9_539 b_9 NI_9 NS_539 0 1.1308767477586115e-06
GC_9_540 b_9 NI_9 NS_540 0 2.8161632054237241e-06
GC_9_541 b_9 NI_9 NS_541 0 -1.4324487330469199e-04
GC_9_542 b_9 NI_9 NS_542 0 3.4599467413052740e-11
GC_9_543 b_9 NI_9 NS_543 0 3.0173709435680436e-11
GC_9_544 b_9 NI_9 NS_544 0 9.4205983492422668e-10
GC_9_545 b_9 NI_9 NS_545 0 -2.1091114572365045e-06
GC_9_546 b_9 NI_9 NS_546 0 -1.6534016903911216e-06
GC_9_547 b_9 NI_9 NS_547 0 1.8892532615790832e-06
GC_9_548 b_9 NI_9 NS_548 0 3.8450042742583117e-06
GC_9_549 b_9 NI_9 NS_549 0 3.2880814857221841e-06
GC_9_550 b_9 NI_9 NS_550 0 4.9269039539685649e-06
GC_9_551 b_9 NI_9 NS_551 0 5.8303633159812734e-06
GC_9_552 b_9 NI_9 NS_552 0 -9.0831332799048900e-06
GC_9_553 b_9 NI_9 NS_553 0 -2.5401375317783300e-06
GC_9_554 b_9 NI_9 NS_554 0 -1.3836005451209194e-05
GC_9_555 b_9 NI_9 NS_555 0 -3.5342175278354143e-06
GC_9_556 b_9 NI_9 NS_556 0 2.1965935209234460e-06
GC_9_557 b_9 NI_9 NS_557 0 3.6390200670882789e-06
GC_9_558 b_9 NI_9 NS_558 0 1.2969560792705312e-06
GC_9_559 b_9 NI_9 NS_559 0 7.8997169570542283e-06
GC_9_560 b_9 NI_9 NS_560 0 -3.9683457076451259e-05
GC_9_561 b_9 NI_9 NS_561 0 -4.4005703656238965e-05
GC_9_562 b_9 NI_9 NS_562 0 -8.8268777709008879e-07
GC_9_563 b_9 NI_9 NS_563 0 -1.4766093497203224e-05
GC_9_564 b_9 NI_9 NS_564 0 -8.4725309764088267e-06
GC_9_565 b_9 NI_9 NS_565 0 -7.2348312401145337e-05
GC_9_566 b_9 NI_9 NS_566 0 7.5140007938084206e-05
GC_9_567 b_9 NI_9 NS_567 0 4.6496204966377330e-06
GC_9_568 b_9 NI_9 NS_568 0 1.3009890318642478e-05
GC_9_569 b_9 NI_9 NS_569 0 6.2664895123892416e-05
GC_9_570 b_9 NI_9 NS_570 0 1.2224105928877594e-04
GC_9_571 b_9 NI_9 NS_571 0 2.4432286803255246e-07
GC_9_572 b_9 NI_9 NS_572 0 -3.6753045522304275e-05
GC_9_573 b_9 NI_9 NS_573 0 1.6411266024218295e-05
GC_9_574 b_9 NI_9 NS_574 0 3.8870354784114661e-06
GC_9_575 b_9 NI_9 NS_575 0 2.4218752682674635e-05
GC_9_576 b_9 NI_9 NS_576 0 -3.0243867620374805e-05
GC_9_577 b_9 NI_9 NS_577 0 -8.8438580316228302e-06
GC_9_578 b_9 NI_9 NS_578 0 -2.2760875918115729e-06
GC_9_579 b_9 NI_9 NS_579 0 -8.7280266962045885e-06
GC_9_580 b_9 NI_9 NS_580 0 2.5050836428464080e-05
GC_9_581 b_9 NI_9 NS_581 0 5.8326436131262786e-06
GC_9_582 b_9 NI_9 NS_582 0 8.3787532165186872e-06
GC_9_583 b_9 NI_9 NS_583 0 5.5968998100025125e-05
GC_9_584 b_9 NI_9 NS_584 0 2.4647272650315577e-05
GC_9_585 b_9 NI_9 NS_585 0 3.4490056979279019e-06
GC_9_586 b_9 NI_9 NS_586 0 -1.1606188993900533e-05
GC_9_587 b_9 NI_9 NS_587 0 -4.0623963328018797e-07
GC_9_588 b_9 NI_9 NS_588 0 -1.2992062548705400e-06
GC_9_589 b_9 NI_9 NS_589 0 6.7879557742943439e-06
GC_9_590 b_9 NI_9 NS_590 0 3.0205339665738351e-06
GC_9_591 b_9 NI_9 NS_591 0 4.1591493957191341e-05
GC_9_592 b_9 NI_9 NS_592 0 -1.7165556407216300e-05
GC_9_593 b_9 NI_9 NS_593 0 -2.5739638972008553e-06
GC_9_594 b_9 NI_9 NS_594 0 -7.0282436432026678e-06
GC_9_595 b_9 NI_9 NS_595 0 -2.9900961912380127e-06
GC_9_596 b_9 NI_9 NS_596 0 1.7603693193363226e-06
GC_9_597 b_9 NI_9 NS_597 0 9.5385224671499211e-06
GC_9_598 b_9 NI_9 NS_598 0 2.8682580273595621e-06
GC_9_599 b_9 NI_9 NS_599 0 2.2731242079705236e-05
GC_9_600 b_9 NI_9 NS_600 0 -3.1037334052771686e-05
GC_9_601 b_9 NI_9 NS_601 0 -5.6872056827168597e-06
GC_9_602 b_9 NI_9 NS_602 0 -3.6245387664927025e-06
GC_9_603 b_9 NI_9 NS_603 0 -5.2396148009239352e-07
GC_9_604 b_9 NI_9 NS_604 0 5.0176564252489972e-06
GC_9_605 b_9 NI_9 NS_605 0 1.2253621314045922e-05
GC_9_606 b_9 NI_9 NS_606 0 1.7526947027216957e-07
GC_9_607 b_9 NI_9 NS_607 0 1.8081448188586922e-06
GC_9_608 b_9 NI_9 NS_608 0 -3.1349624740910630e-05
GC_9_609 b_9 NI_9 NS_609 0 -6.7180800695120862e-06
GC_9_610 b_9 NI_9 NS_610 0 9.7556963357286584e-07
GC_9_611 b_9 NI_9 NS_611 0 4.6118407332583356e-06
GC_9_612 b_9 NI_9 NS_612 0 3.8655555583483718e-06
GC_9_613 b_9 NI_9 NS_613 0 1.4061772046009059e-05
GC_9_614 b_9 NI_9 NS_614 0 -6.0101884678337119e-06
GC_9_615 b_9 NI_9 NS_615 0 -1.4015860688176883e-05
GC_9_616 b_9 NI_9 NS_616 0 -1.8746801196373944e-05
GC_9_617 b_9 NI_9 NS_617 0 -2.5061575703374167e-06
GC_9_618 b_9 NI_9 NS_618 0 5.4162640386069681e-06
GC_9_619 b_9 NI_9 NS_619 0 4.6576662901954450e-06
GC_9_620 b_9 NI_9 NS_620 0 -2.0834543373339985e-06
GC_9_621 b_9 NI_9 NS_621 0 -1.4565910006074132e-11
GC_9_622 b_9 NI_9 NS_622 0 4.2060440282703927e-12
GC_9_623 b_9 NI_9 NS_623 0 5.1979353402652667e-06
GC_9_624 b_9 NI_9 NS_624 0 -1.1242576754087001e-05
GC_9_625 b_9 NI_9 NS_625 0 -2.6677167481414741e-07
GC_9_626 b_9 NI_9 NS_626 0 2.9264747688262533e-06
GC_9_627 b_9 NI_9 NS_627 0 2.6445008217943786e-06
GC_9_628 b_9 NI_9 NS_628 0 -1.5935795607822244e-06
GC_9_629 b_9 NI_9 NS_629 0 2.4075831164431022e-06
GC_9_630 b_9 NI_9 NS_630 0 -9.4307995867632093e-06
GC_9_631 b_9 NI_9 NS_631 0 -9.9265724179344562e-06
GC_9_632 b_9 NI_9 NS_632 0 -3.6883835363550907e-06
GC_9_633 b_9 NI_9 NS_633 0 3.1234678021024361e-10
GC_9_634 b_9 NI_9 NS_634 0 2.7704243155543102e-10
GC_9_635 b_9 NI_9 NS_635 0 -8.5916119905036413e-06
GC_9_636 b_9 NI_9 NS_636 0 -5.6864935232245213e-06
GC_9_637 b_9 NI_9 NS_637 0 2.2662276392309312e-06
GC_9_638 b_9 NI_9 NS_638 0 -6.4520067025861817e-06
GC_9_639 b_9 NI_9 NS_639 0 -3.0674012774411139e-06
GC_9_640 b_9 NI_9 NS_640 0 -1.3540167405187163e-07
GC_9_641 b_9 NI_9 NS_641 0 -7.9220186819051894e-06
GC_9_642 b_9 NI_9 NS_642 0 4.8459928122780466e-07
GC_9_643 b_9 NI_9 NS_643 0 3.0018513797385119e-06
GC_9_644 b_9 NI_9 NS_644 0 2.8730924786954239e-06
GC_9_645 b_9 NI_9 NS_645 0 1.2172140123650646e-06
GC_9_646 b_9 NI_9 NS_646 0 -3.8814878695881873e-06
GC_9_647 b_9 NI_9 NS_647 0 -4.8738055419244665e-06
GC_9_648 b_9 NI_9 NS_648 0 -3.9067779273018356e-06
GC_9_649 b_9 NI_9 NS_649 0 5.6901722858630906e-05
GC_9_650 b_9 NI_9 NS_650 0 -1.2101214696902654e-10
GC_9_651 b_9 NI_9 NS_651 0 -2.0303492180511211e-09
GC_9_652 b_9 NI_9 NS_652 0 3.4201751865296745e-08
GC_9_653 b_9 NI_9 NS_653 0 -5.1436525338421706e-07
GC_9_654 b_9 NI_9 NS_654 0 -3.8174198074055462e-07
GC_9_655 b_9 NI_9 NS_655 0 -8.7414460132438866e-07
GC_9_656 b_9 NI_9 NS_656 0 9.5753742718516656e-06
GC_9_657 b_9 NI_9 NS_657 0 1.2647197559549357e-05
GC_9_658 b_9 NI_9 NS_658 0 -1.2046359928505865e-05
GC_9_659 b_9 NI_9 NS_659 0 -1.7539602496435053e-05
GC_9_660 b_9 NI_9 NS_660 0 8.8316937569634122e-06
GC_9_661 b_9 NI_9 NS_661 0 2.8400590187642023e-05
GC_9_662 b_9 NI_9 NS_662 0 -6.5599992345446662e-06
GC_9_663 b_9 NI_9 NS_663 0 -3.2052663771441450e-06
GC_9_664 b_9 NI_9 NS_664 0 -3.0961922735083450e-06
GC_9_665 b_9 NI_9 NS_665 0 -2.8500835465075323e-06
GC_9_666 b_9 NI_9 NS_666 0 -1.4496618491843491e-05
GC_9_667 b_9 NI_9 NS_667 0 -2.4759453236327353e-05
GC_9_668 b_9 NI_9 NS_668 0 4.0216184098678795e-05
GC_9_669 b_9 NI_9 NS_669 0 3.7734461362250143e-05
GC_9_670 b_9 NI_9 NS_670 0 -4.7031954491313228e-05
GC_9_671 b_9 NI_9 NS_671 0 -3.0428897985625818e-05
GC_9_672 b_9 NI_9 NS_672 0 -2.0940879609513644e-05
GC_9_673 b_9 NI_9 NS_673 0 3.3065734946937343e-05
GC_9_674 b_9 NI_9 NS_674 0 2.6832551869096672e-05
GC_9_675 b_9 NI_9 NS_675 0 -1.8367596889521854e-05
GC_9_676 b_9 NI_9 NS_676 0 -2.8794840948235055e-05
GC_9_677 b_9 NI_9 NS_677 0 2.1463961944456878e-05
GC_9_678 b_9 NI_9 NS_678 0 6.0258496213280377e-05
GC_9_679 b_9 NI_9 NS_679 0 -2.1175879407106407e-05
GC_9_680 b_9 NI_9 NS_680 0 -5.5544526317301132e-05
GC_9_681 b_9 NI_9 NS_681 0 -3.1396081126751017e-05
GC_9_682 b_9 NI_9 NS_682 0 -1.1645550077974733e-05
GC_9_683 b_9 NI_9 NS_683 0 2.0313320790889322e-05
GC_9_684 b_9 NI_9 NS_684 0 1.3869333986479771e-05
GC_9_685 b_9 NI_9 NS_685 0 -2.4579256005700782e-05
GC_9_686 b_9 NI_9 NS_686 0 -1.0925619028646579e-05
GC_9_687 b_9 NI_9 NS_687 0 2.0765547116127809e-05
GC_9_688 b_9 NI_9 NS_688 0 1.0077085812366526e-05
GC_9_689 b_9 NI_9 NS_689 0 -1.8224323606800499e-05
GC_9_690 b_9 NI_9 NS_690 0 -2.0845546805780225e-05
GC_9_691 b_9 NI_9 NS_691 0 5.4975821143041202e-06
GC_9_692 b_9 NI_9 NS_692 0 3.2160679956752230e-05
GC_9_693 b_9 NI_9 NS_693 0 -8.2125207951843117e-06
GC_9_694 b_9 NI_9 NS_694 0 -2.6520146726066688e-05
GC_9_695 b_9 NI_9 NS_695 0 -1.8293146698927648e-06
GC_9_696 b_9 NI_9 NS_696 0 1.6902887215291423e-06
GC_9_697 b_9 NI_9 NS_697 0 -1.9229254423503023e-05
GC_9_698 b_9 NI_9 NS_698 0 -1.1940103298075982e-05
GC_9_699 b_9 NI_9 NS_699 0 6.9725833410388860e-06
GC_9_700 b_9 NI_9 NS_700 0 2.0939545459448216e-05
GC_9_701 b_9 NI_9 NS_701 0 -1.5976405731800880e-05
GC_9_702 b_9 NI_9 NS_702 0 -1.4813667358462449e-05
GC_9_703 b_9 NI_9 NS_703 0 1.3388596766199003e-06
GC_9_704 b_9 NI_9 NS_704 0 5.3013247072635318e-06
GC_9_705 b_9 NI_9 NS_705 0 -2.4841218466113813e-05
GC_9_706 b_9 NI_9 NS_706 0 -9.8243626611648414e-06
GC_9_707 b_9 NI_9 NS_707 0 8.5462509717283991e-06
GC_9_708 b_9 NI_9 NS_708 0 2.3050512592887988e-05
GC_9_709 b_9 NI_9 NS_709 0 -2.0672693912653576e-05
GC_9_710 b_9 NI_9 NS_710 0 -5.6252743822772404e-06
GC_9_711 b_9 NI_9 NS_711 0 6.2603548248657980e-06
GC_9_712 b_9 NI_9 NS_712 0 7.5158346809360109e-06
GC_9_713 b_9 NI_9 NS_713 0 -3.0565168717394374e-05
GC_9_714 b_9 NI_9 NS_714 0 -2.5578181338808562e-06
GC_9_715 b_9 NI_9 NS_715 0 1.8794226505983732e-05
GC_9_716 b_9 NI_9 NS_716 0 2.5290846671332918e-05
GC_9_717 b_9 NI_9 NS_717 0 -2.1787414660029742e-05
GC_9_718 b_9 NI_9 NS_718 0 6.9645035808395984e-06
GC_9_719 b_9 NI_9 NS_719 0 1.5266870746895403e-05
GC_9_720 b_9 NI_9 NS_720 0 3.9771046859446234e-06
GC_9_721 b_9 NI_9 NS_721 0 -3.4533266394194799e-05
GC_9_722 b_9 NI_9 NS_722 0 1.3723474401827054e-05
GC_9_723 b_9 NI_9 NS_723 0 3.7469640110972260e-05
GC_9_724 b_9 NI_9 NS_724 0 1.2338010272661636e-05
GC_9_725 b_9 NI_9 NS_725 0 -7.7465657423676141e-06
GC_9_726 b_9 NI_9 NS_726 0 1.8808998669165939e-05
GC_9_727 b_9 NI_9 NS_727 0 1.2775019477040576e-05
GC_9_728 b_9 NI_9 NS_728 0 -1.1287478919010131e-05
GC_9_729 b_9 NI_9 NS_729 0 1.0985023700363512e-10
GC_9_730 b_9 NI_9 NS_730 0 3.5334384136850538e-11
GC_9_731 b_9 NI_9 NS_731 0 -1.3692325264420816e-05
GC_9_732 b_9 NI_9 NS_732 0 2.5942178261406131e-05
GC_9_733 b_9 NI_9 NS_733 0 -2.0633483795435707e-06
GC_9_734 b_9 NI_9 NS_734 0 1.0503161437866458e-05
GC_9_735 b_9 NI_9 NS_735 0 6.1729256970711120e-06
GC_9_736 b_9 NI_9 NS_736 0 -8.5364896176953737e-06
GC_9_737 b_9 NI_9 NS_737 0 -8.1124828757664882e-06
GC_9_738 b_9 NI_9 NS_738 0 2.5390672393033168e-05
GC_9_739 b_9 NI_9 NS_739 0 2.4973015458427218e-05
GC_9_740 b_9 NI_9 NS_740 0 -1.0421081112522697e-05
GC_9_741 b_9 NI_9 NS_741 0 4.8846458436102481e-09
GC_9_742 b_9 NI_9 NS_742 0 -1.2242819030942906e-09
GC_9_743 b_9 NI_9 NS_743 0 2.6368704707249266e-05
GC_9_744 b_9 NI_9 NS_744 0 -1.2610269330606921e-05
GC_9_745 b_9 NI_9 NS_745 0 -8.2495148329796757e-06
GC_9_746 b_9 NI_9 NS_746 0 1.8114668802010426e-05
GC_9_747 b_9 NI_9 NS_747 0 -1.0378170770127183e-05
GC_9_748 b_9 NI_9 NS_748 0 -3.0217642067771631e-07
GC_9_749 b_9 NI_9 NS_749 0 1.9390226743584523e-05
GC_9_750 b_9 NI_9 NS_750 0 -1.4389078589537210e-05
GC_9_751 b_9 NI_9 NS_751 0 7.1949281939545464e-06
GC_9_752 b_9 NI_9 NS_752 0 1.1599497571888150e-05
GC_9_753 b_9 NI_9 NS_753 0 -2.2868214949040899e-07
GC_9_754 b_9 NI_9 NS_754 0 -1.4637668358797035e-05
GC_9_755 b_9 NI_9 NS_755 0 1.3160348027878964e-05
GC_9_756 b_9 NI_9 NS_756 0 2.7988961318822774e-05
GC_9_757 b_9 NI_9 NS_757 0 -6.3809595178207306e-04
GC_9_758 b_9 NI_9 NS_758 0 -9.7135980855898662e-11
GC_9_759 b_9 NI_9 NS_759 0 3.8809011749551905e-09
GC_9_760 b_9 NI_9 NS_760 0 -6.7422274741723916e-08
GC_9_761 b_9 NI_9 NS_761 0 -1.1286635238526398e-05
GC_9_762 b_9 NI_9 NS_762 0 -9.3365547946119337e-06
GC_9_763 b_9 NI_9 NS_763 0 -2.2471565876233769e-06
GC_9_764 b_9 NI_9 NS_764 0 2.3210492418880009e-07
GC_9_765 b_9 NI_9 NS_765 0 -3.0313696629227993e-05
GC_9_766 b_9 NI_9 NS_766 0 2.7072955824765312e-05
GC_9_767 b_9 NI_9 NS_767 0 -3.3247384051705323e-05
GC_9_768 b_9 NI_9 NS_768 0 8.1286507295039923e-06
GC_9_769 b_9 NI_9 NS_769 0 3.1755740671884641e-05
GC_9_770 b_9 NI_9 NS_770 0 2.7371062582158002e-05
GC_9_771 b_9 NI_9 NS_771 0 -9.0592455326207185e-06
GC_9_772 b_9 NI_9 NS_772 0 1.4745488688867908e-05
GC_9_773 b_9 NI_9 NS_773 0 1.2657452693869481e-05
GC_9_774 b_9 NI_9 NS_774 0 3.6938831232147876e-05
GC_9_775 b_9 NI_9 NS_775 0 -1.0625090512655731e-05
GC_9_776 b_9 NI_9 NS_776 0 6.8145150523449586e-05
GC_9_777 b_9 NI_9 NS_777 0 9.5462361546343010e-05
GC_9_778 b_9 NI_9 NS_778 0 -6.6200939362170009e-05
GC_9_779 b_9 NI_9 NS_779 0 2.7086625673307029e-05
GC_9_780 b_9 NI_9 NS_780 0 3.1697639280339858e-05
GC_9_781 b_9 NI_9 NS_781 0 -7.3750072361536536e-06
GC_9_782 b_9 NI_9 NS_782 0 -7.2639290827336111e-05
GC_9_783 b_9 NI_9 NS_783 0 -9.8543873519437713e-06
GC_9_784 b_9 NI_9 NS_784 0 -3.3996036020446728e-05
GC_9_785 b_9 NI_9 NS_785 0 -7.7016952071555595e-05
GC_9_786 b_9 NI_9 NS_786 0 1.9071595377477670e-05
GC_9_787 b_9 NI_9 NS_787 0 2.4929631884834399e-05
GC_9_788 b_9 NI_9 NS_788 0 5.0927030183106003e-05
GC_9_789 b_9 NI_9 NS_789 0 -2.3148581531051638e-05
GC_9_790 b_9 NI_9 NS_790 0 -3.5473839802586377e-06
GC_9_791 b_9 NI_9 NS_791 0 6.9848628601674876e-05
GC_9_792 b_9 NI_9 NS_792 0 4.4676877423808920e-05
GC_9_793 b_9 NI_9 NS_793 0 2.9208026797332296e-05
GC_9_794 b_9 NI_9 NS_794 0 1.9693880966242524e-05
GC_9_795 b_9 NI_9 NS_795 0 -7.3329400660922800e-06
GC_9_796 b_9 NI_9 NS_796 0 -2.5741687239305675e-05
GC_9_797 b_9 NI_9 NS_797 0 -7.5876273770167362e-06
GC_9_798 b_9 NI_9 NS_798 0 -2.5167214221424882e-05
GC_9_799 b_9 NI_9 NS_799 0 6.7364215277651590e-06
GC_9_800 b_9 NI_9 NS_800 0 4.9241831237592936e-05
GC_9_801 b_9 NI_9 NS_801 0 1.2922949907309970e-05
GC_9_802 b_9 NI_9 NS_802 0 2.7360377784838086e-05
GC_9_803 b_9 NI_9 NS_803 0 5.8665065587317712e-06
GC_9_804 b_9 NI_9 NS_804 0 2.1248473506562489e-06
GC_9_805 b_9 NI_9 NS_805 0 -6.3214814524509036e-07
GC_9_806 b_9 NI_9 NS_806 0 -1.5379664158684778e-05
GC_9_807 b_9 NI_9 NS_807 0 5.6145747998505798e-05
GC_9_808 b_9 NI_9 NS_808 0 3.8184728937167638e-05
GC_9_809 b_9 NI_9 NS_809 0 1.9943098803950866e-05
GC_9_810 b_9 NI_9 NS_810 0 1.4808800471371668e-05
GC_9_811 b_9 NI_9 NS_811 0 8.3810801999019918e-06
GC_9_812 b_9 NI_9 NS_812 0 -1.2844658496124913e-05
GC_9_813 b_9 NI_9 NS_813 0 -5.6561555814100697e-06
GC_9_814 b_9 NI_9 NS_814 0 -1.3981129443443264e-05
GC_9_815 b_9 NI_9 NS_815 0 6.6094147513344389e-05
GC_9_816 b_9 NI_9 NS_816 0 1.3028870095685336e-05
GC_9_817 b_9 NI_9 NS_817 0 2.2769670615442580e-05
GC_9_818 b_9 NI_9 NS_818 0 4.9311308052096838e-06
GC_9_819 b_9 NI_9 NS_819 0 -5.5540365311244962e-06
GC_9_820 b_9 NI_9 NS_820 0 -2.1975728530530918e-05
GC_9_821 b_9 NI_9 NS_821 0 -9.1463308359853417e-06
GC_9_822 b_9 NI_9 NS_822 0 -7.0651058045965897e-06
GC_9_823 b_9 NI_9 NS_823 0 6.0665957290699438e-05
GC_9_824 b_9 NI_9 NS_824 0 -9.4701819154580705e-06
GC_9_825 b_9 NI_9 NS_825 0 2.1425124861513092e-05
GC_9_826 b_9 NI_9 NS_826 0 -7.3811074379501653e-06
GC_9_827 b_9 NI_9 NS_827 0 -2.3068076918328013e-05
GC_9_828 b_9 NI_9 NS_828 0 -1.3110919461531548e-05
GC_9_829 b_9 NI_9 NS_829 0 -8.6671540266394147e-06
GC_9_830 b_9 NI_9 NS_830 0 4.4627732214031369e-06
GC_9_831 b_9 NI_9 NS_831 0 4.5473376943922713e-05
GC_9_832 b_9 NI_9 NS_832 0 -2.5661823167711394e-05
GC_9_833 b_9 NI_9 NS_833 0 6.0269434172810541e-06
GC_9_834 b_9 NI_9 NS_834 0 -1.6485835936117598e-05
GC_9_835 b_9 NI_9 NS_835 0 -1.8722684202156870e-05
GC_9_836 b_9 NI_9 NS_836 0 8.6301705064291936e-06
GC_9_837 b_9 NI_9 NS_837 0 -4.6983778657638287e-11
GC_9_838 b_9 NI_9 NS_838 0 -1.7787081282066339e-10
GC_9_839 b_9 NI_9 NS_839 0 1.7486926917940410e-06
GC_9_840 b_9 NI_9 NS_840 0 8.7729554932131744e-06
GC_9_841 b_9 NI_9 NS_841 0 2.2060636794003548e-06
GC_9_842 b_9 NI_9 NS_842 0 -7.0028074670855852e-06
GC_9_843 b_9 NI_9 NS_843 0 -9.0193558926148486e-06
GC_9_844 b_9 NI_9 NS_844 0 5.7725449241821562e-06
GC_9_845 b_9 NI_9 NS_845 0 4.7628827956065172e-06
GC_9_846 b_9 NI_9 NS_846 0 1.1522802080245294e-05
GC_9_847 b_9 NI_9 NS_847 0 2.4566763680301080e-05
GC_9_848 b_9 NI_9 NS_848 0 -2.1153853200860300e-05
GC_9_849 b_9 NI_9 NS_849 0 -5.7421773142849572e-09
GC_9_850 b_9 NI_9 NS_850 0 -5.6214187853346790e-09
GC_9_851 b_9 NI_9 NS_851 0 3.0633017830220606e-05
GC_9_852 b_9 NI_9 NS_852 0 7.5206554419129426e-06
GC_9_853 b_9 NI_9 NS_853 0 -2.6889461084653131e-06
GC_9_854 b_9 NI_9 NS_854 0 1.1036277354993729e-05
GC_9_855 b_9 NI_9 NS_855 0 8.0385272225943326e-06
GC_9_856 b_9 NI_9 NS_856 0 1.1983685410935221e-06
GC_9_857 b_9 NI_9 NS_857 0 1.9085220456489907e-05
GC_9_858 b_9 NI_9 NS_858 0 -2.1544586533416968e-05
GC_9_859 b_9 NI_9 NS_859 0 -6.5775891761729278e-06
GC_9_860 b_9 NI_9 NS_860 0 -7.4340037716176146e-06
GC_9_861 b_9 NI_9 NS_861 0 -5.4042930956811705e-06
GC_9_862 b_9 NI_9 NS_862 0 1.2516899148487792e-05
GC_9_863 b_9 NI_9 NS_863 0 1.6097136293338694e-05
GC_9_864 b_9 NI_9 NS_864 0 7.3672696961396570e-06
GC_9_865 b_9 NI_9 NS_865 0 -1.4246400256028493e-02
GC_9_866 b_9 NI_9 NS_866 0 6.2293160768327371e-09
GC_9_867 b_9 NI_9 NS_867 0 -1.0771399406067467e-06
GC_9_868 b_9 NI_9 NS_868 0 -2.3238215206440901e-05
GC_9_869 b_9 NI_9 NS_869 0 3.4199266343491519e-04
GC_9_870 b_9 NI_9 NS_870 0 -1.9835114711510228e-04
GC_9_871 b_9 NI_9 NS_871 0 -1.5573869762491889e-03
GC_9_872 b_9 NI_9 NS_872 0 -2.3367645319626756e-03
GC_9_873 b_9 NI_9 NS_873 0 -6.7656858961289294e-05
GC_9_874 b_9 NI_9 NS_874 0 4.3764648565271158e-03
GC_9_875 b_9 NI_9 NS_875 0 1.6012909917152746e-03
GC_9_876 b_9 NI_9 NS_876 0 -5.9363791255958153e-03
GC_9_877 b_9 NI_9 NS_877 0 -4.9862942191484993e-03
GC_9_878 b_9 NI_9 NS_878 0 6.4938569038296510e-03
GC_9_879 b_9 NI_9 NS_879 0 1.1242574208519920e-03
GC_9_880 b_9 NI_9 NS_880 0 -4.9042309876351563e-04
GC_9_881 b_9 NI_9 NS_881 0 2.8092071387608572e-03
GC_9_882 b_9 NI_9 NS_882 0 2.3585353006908027e-03
GC_9_883 b_9 NI_9 NS_883 0 -4.3182735494993350e-03
GC_9_884 b_9 NI_9 NS_884 0 -1.3539567903205919e-02
GC_9_885 b_9 NI_9 NS_885 0 1.6031707990065366e-03
GC_9_886 b_9 NI_9 NS_886 0 1.7677776973712638e-02
GC_9_887 b_9 NI_9 NS_887 0 9.8386853699242906e-03
GC_9_888 b_9 NI_9 NS_888 0 -2.2919452674643819e-03
GC_9_889 b_9 NI_9 NS_889 0 -1.3104487520470351e-02
GC_9_890 b_9 NI_9 NS_890 0 2.2186351324758216e-03
GC_9_891 b_9 NI_9 NS_891 0 9.2001458916820874e-03
GC_9_892 b_9 NI_9 NS_892 0 1.9506148644372902e-03
GC_9_893 b_9 NI_9 NS_893 0 -1.7998043609793842e-02
GC_9_894 b_9 NI_9 NS_894 0 -6.4920163427329746e-03
GC_9_895 b_9 NI_9 NS_895 0 1.5711166851321900e-02
GC_9_896 b_9 NI_9 NS_896 0 6.4981549055296720e-03
GC_9_897 b_9 NI_9 NS_897 0 8.1166025771046337e-03
GC_9_898 b_9 NI_9 NS_898 0 -4.1938599544669268e-03
GC_9_899 b_9 NI_9 NS_899 0 -7.5320604141213780e-03
GC_9_900 b_9 NI_9 NS_900 0 2.0324522546205071e-03
GC_9_901 b_9 NI_9 NS_901 0 6.7023914700824524e-03
GC_9_902 b_9 NI_9 NS_902 0 -2.7451417078800987e-03
GC_9_903 b_9 NI_9 NS_903 0 -6.5840314599313133e-03
GC_9_904 b_9 NI_9 NS_904 0 2.8920091767600364e-03
GC_9_905 b_9 NI_9 NS_905 0 7.6634824591408929e-03
GC_9_906 b_9 NI_9 NS_906 0 4.8601602431004305e-04
GC_9_907 b_9 NI_9 NS_907 0 -9.3542684002521567e-03
GC_9_908 b_9 NI_9 NS_908 0 -5.1821823155192110e-03
GC_9_909 b_9 NI_9 NS_909 0 6.8205079141039114e-03
GC_9_910 b_9 NI_9 NS_910 0 4.1105978305452512e-03
GC_9_911 b_9 NI_9 NS_911 0 -3.8505593707250909e-04
GC_9_912 b_9 NI_9 NS_912 0 -9.3423498820469476e-04
GC_9_913 b_9 NI_9 NS_913 0 5.6830560567739464e-03
GC_9_914 b_9 NI_9 NS_914 0 -1.3773210671378590e-03
GC_9_915 b_9 NI_9 NS_915 0 -9.1525589686269043e-03
GC_9_916 b_9 NI_9 NS_916 0 -1.2845549510713376e-03
GC_9_917 b_9 NI_9 NS_917 0 5.9995912358443539e-03
GC_9_918 b_9 NI_9 NS_918 0 7.3474949662837952e-04
GC_9_919 b_9 NI_9 NS_919 0 -2.6407532414300930e-03
GC_9_920 b_9 NI_9 NS_920 0 2.3246011121313796e-04
GC_9_921 b_9 NI_9 NS_921 0 6.7119817333128676e-03
GC_9_922 b_9 NI_9 NS_922 0 -2.2566059982605906e-03
GC_9_923 b_9 NI_9 NS_923 0 -9.2876748456727273e-03
GC_9_924 b_9 NI_9 NS_924 0 1.4716659449829088e-03
GC_9_925 b_9 NI_9 NS_925 0 5.7396120360619389e-03
GC_9_926 b_9 NI_9 NS_926 0 -1.5055499470721973e-03
GC_9_927 b_9 NI_9 NS_927 0 -3.3169903661786643e-03
GC_9_928 b_9 NI_9 NS_928 0 2.3821024421813923e-03
GC_9_929 b_9 NI_9 NS_929 0 7.2818936807726659e-03
GC_9_930 b_9 NI_9 NS_930 0 -4.0976796271507878e-03
GC_9_931 b_9 NI_9 NS_931 0 -8.5931345432160473e-03
GC_9_932 b_9 NI_9 NS_932 0 4.1427763954092669e-03
GC_9_933 b_9 NI_9 NS_933 0 4.8244396283538835e-03
GC_9_934 b_9 NI_9 NS_934 0 -3.8807312376370512e-03
GC_9_935 b_9 NI_9 NS_935 0 -2.4175655609639567e-03
GC_9_936 b_9 NI_9 NS_936 0 4.7355196559177833e-03
GC_9_937 b_9 NI_9 NS_937 0 7.0698660120572911e-03
GC_9_938 b_9 NI_9 NS_938 0 -7.3594026153951083e-03
GC_9_939 b_9 NI_9 NS_939 0 -7.1573588934082484e-03
GC_9_940 b_9 NI_9 NS_940 0 6.8575791856932047e-03
GC_9_941 b_9 NI_9 NS_941 0 1.6629097338057275e-03
GC_9_942 b_9 NI_9 NS_942 0 -5.3099127673498113e-03
GC_9_943 b_9 NI_9 NS_943 0 5.8005351314567761e-04
GC_9_944 b_9 NI_9 NS_944 0 5.4707649844615647e-03
GC_9_945 b_9 NI_9 NS_945 0 -4.5818073807837382e-09
GC_9_946 b_9 NI_9 NS_946 0 -1.3467649890965799e-08
GC_9_947 b_9 NI_9 NS_947 0 2.7089365488078628e-03
GC_9_948 b_9 NI_9 NS_948 0 -8.5910067713740618e-03
GC_9_949 b_9 NI_9 NS_949 0 8.6608706430432497e-04
GC_9_950 b_9 NI_9 NS_950 0 -3.4347604172176439e-03
GC_9_951 b_9 NI_9 NS_951 0 6.2756551860495289e-04
GC_9_952 b_9 NI_9 NS_952 0 4.0313415341298323e-03
GC_9_953 b_9 NI_9 NS_953 0 2.1670484566328990e-03
GC_9_954 b_9 NI_9 NS_954 0 -8.1665277093597027e-03
GC_9_955 b_9 NI_9 NS_955 0 -3.4991635045163627e-03
GC_9_956 b_9 NI_9 NS_956 0 7.0126788784464064e-03
GC_9_957 b_9 NI_9 NS_957 0 -1.0829860079749097e-07
GC_9_958 b_9 NI_9 NS_958 0 -3.0048166007698173e-07
GC_9_959 b_9 NI_9 NS_959 0 -8.0240632959310849e-03
GC_9_960 b_9 NI_9 NS_960 0 5.3776059369875229e-03
GC_9_961 b_9 NI_9 NS_961 0 4.1768102857436809e-03
GC_9_962 b_9 NI_9 NS_962 0 -6.8620734780150093e-03
GC_9_963 b_9 NI_9 NS_963 0 5.3214177374611288e-03
GC_9_964 b_9 NI_9 NS_964 0 7.4369283070834912e-04
GC_9_965 b_9 NI_9 NS_965 0 -2.3651597210068696e-03
GC_9_966 b_9 NI_9 NS_966 0 6.8561897696883820e-03
GC_9_967 b_9 NI_9 NS_967 0 -1.4960016228829085e-03
GC_9_968 b_9 NI_9 NS_968 0 -4.2193424589338719e-03
GC_9_969 b_9 NI_9 NS_969 0 2.3601153783920506e-03
GC_9_970 b_9 NI_9 NS_970 0 5.0361467955909447e-03
GC_9_971 b_9 NI_9 NS_971 0 -2.0068772397933586e-03
GC_9_972 b_9 NI_9 NS_972 0 -8.9761631515452665e-03
GC_9_973 b_9 NI_9 NS_973 0 -1.0575774344971856e-02
GC_9_974 b_9 NI_9 NS_974 0 9.5594887915491672e-09
GC_9_975 b_9 NI_9 NS_975 0 9.8516036529254084e-07
GC_9_976 b_9 NI_9 NS_976 0 3.6184052898170068e-05
GC_9_977 b_9 NI_9 NS_977 0 4.3796872631612811e-03
GC_9_978 b_9 NI_9 NS_978 0 -3.4738145892704068e-03
GC_9_979 b_9 NI_9 NS_979 0 -3.7302937390053903e-03
GC_9_980 b_9 NI_9 NS_980 0 6.2452078499370643e-03
GC_9_981 b_9 NI_9 NS_981 0 -8.7505776398336364e-03
GC_9_982 b_9 NI_9 NS_982 0 -5.9709534917151514e-03
GC_9_983 b_9 NI_9 NS_983 0 9.2221604719982132e-03
GC_9_984 b_9 NI_9 NS_984 0 -5.9539857747886241e-03
GC_9_985 b_9 NI_9 NS_985 0 7.1415969970234743e-03
GC_9_986 b_9 NI_9 NS_986 0 1.1891209555263446e-02
GC_9_987 b_9 NI_9 NS_987 0 -4.2237323549645881e-03
GC_9_988 b_9 NI_9 NS_988 0 -1.1434325744962479e-03
GC_9_989 b_9 NI_9 NS_989 0 -8.8759714399074627e-03
GC_9_990 b_9 NI_9 NS_990 0 -4.8953589312983998e-04
GC_9_991 b_9 NI_9 NS_991 0 1.4613659188457721e-02
GC_9_992 b_9 NI_9 NS_992 0 -1.0366887955436634e-02
GC_9_993 b_9 NI_9 NS_993 0 1.6417972793514500e-02
GC_9_994 b_9 NI_9 NS_994 0 4.0448629043991352e-03
GC_9_995 b_9 NI_9 NS_995 0 -1.1484874502364639e-02
GC_9_996 b_9 NI_9 NS_996 0 -2.5535024427150173e-04
GC_9_997 b_9 NI_9 NS_997 0 -1.6636070051176451e-02
GC_9_998 b_9 NI_9 NS_998 0 -4.4594455804944838e-02
GC_9_999 b_9 NI_9 NS_999 0 1.0649429618427063e-02
GC_9_1000 b_9 NI_9 NS_1000 0 1.1313046844154578e-03
GC_9_1001 b_9 NI_9 NS_1001 0 -4.8338823264733016e-02
GC_9_1002 b_9 NI_9 NS_1002 0 1.1008374278087492e-02
GC_9_1003 b_9 NI_9 NS_1003 0 -1.0431880825344686e-02
GC_9_1004 b_9 NI_9 NS_1004 0 4.9175332268411266e-04
GC_9_1005 b_9 NI_9 NS_1005 0 9.7750184355797978e-03
GC_9_1006 b_9 NI_9 NS_1006 0 -5.7660630482914295e-04
GC_9_1007 b_9 NI_9 NS_1007 0 4.5630906760372241e-03
GC_9_1008 b_9 NI_9 NS_1008 0 2.4175324745685945e-02
GC_9_1009 b_9 NI_9 NS_1009 0 -1.0747431121523959e-02
GC_9_1010 b_9 NI_9 NS_1010 0 1.9593872761877597e-03
GC_9_1011 b_9 NI_9 NS_1011 0 -8.4817642342787727e-03
GC_9_1012 b_9 NI_9 NS_1012 0 -1.3531506014886409e-02
GC_9_1013 b_9 NI_9 NS_1013 0 1.0144375276298858e-02
GC_9_1014 b_9 NI_9 NS_1014 0 9.9163999690206252e-04
GC_9_1015 b_9 NI_9 NS_1015 0 -1.9215613754864649e-02
GC_9_1016 b_9 NI_9 NS_1016 0 2.8664616511138288e-02
GC_9_1017 b_9 NI_9 NS_1017 0 -9.6176083690540648e-03
GC_9_1018 b_9 NI_9 NS_1018 0 -9.6671756683572752e-04
GC_9_1019 b_9 NI_9 NS_1019 0 1.8850217211049773e-03
GC_9_1020 b_9 NI_9 NS_1020 0 -1.3790988094074545e-03
GC_9_1021 b_9 NI_9 NS_1021 0 9.4567904444767814e-03
GC_9_1022 b_9 NI_9 NS_1022 0 -2.3685211886363632e-04
GC_9_1023 b_9 NI_9 NS_1023 0 -2.0769122372691598e-04
GC_9_1024 b_9 NI_9 NS_1024 0 3.0287226914972033e-02
GC_9_1025 b_9 NI_9 NS_1025 0 -8.5365006859136651e-03
GC_9_1026 b_9 NI_9 NS_1026 0 1.5565108158540613e-04
GC_9_1027 b_9 NI_9 NS_1027 0 2.0685614831006629e-04
GC_9_1028 b_9 NI_9 NS_1028 0 -5.4692331968237851e-03
GC_9_1029 b_9 NI_9 NS_1029 0 1.0024590641568933e-02
GC_9_1030 b_9 NI_9 NS_1030 0 -3.2645329195833683e-04
GC_9_1031 b_9 NI_9 NS_1031 0 8.8940609144675976e-03
GC_9_1032 b_9 NI_9 NS_1032 0 2.6408655915439106e-02
GC_9_1033 b_9 NI_9 NS_1033 0 -8.3634759220739888e-03
GC_9_1034 b_9 NI_9 NS_1034 0 1.3809659287109966e-03
GC_9_1035 b_9 NI_9 NS_1035 0 -2.5879996554086611e-03
GC_9_1036 b_9 NI_9 NS_1036 0 -7.3315703572979611e-03
GC_9_1037 b_9 NI_9 NS_1037 0 1.0540527218066437e-02
GC_9_1038 b_9 NI_9 NS_1038 0 -8.1039258793280742e-04
GC_9_1039 b_9 NI_9 NS_1039 0 1.4431148071945628e-02
GC_9_1040 b_9 NI_9 NS_1040 0 2.0002722624435816e-02
GC_9_1041 b_9 NI_9 NS_1041 0 -8.2822084206109394e-03
GC_9_1042 b_9 NI_9 NS_1042 0 2.9406883298634754e-03
GC_9_1043 b_9 NI_9 NS_1043 0 -5.5808165852560283e-03
GC_9_1044 b_9 NI_9 NS_1044 0 -6.8969412193629195e-03
GC_9_1045 b_9 NI_9 NS_1045 0 1.1228146951872402e-02
GC_9_1046 b_9 NI_9 NS_1046 0 -1.3571951651239430e-03
GC_9_1047 b_9 NI_9 NS_1047 0 1.5726414818171070e-02
GC_9_1048 b_9 NI_9 NS_1048 0 1.2982437375539932e-02
GC_9_1049 b_9 NI_9 NS_1049 0 -7.1842600170538336e-03
GC_9_1050 b_9 NI_9 NS_1050 0 5.1249171225878484e-03
GC_9_1051 b_9 NI_9 NS_1051 0 -6.8612401525741983e-03
GC_9_1052 b_9 NI_9 NS_1052 0 -4.8303580716637902e-03
GC_9_1053 b_9 NI_9 NS_1053 0 5.1293978529190900e-09
GC_9_1054 b_9 NI_9 NS_1054 0 4.4375939771903200e-08
GC_9_1055 b_9 NI_9 NS_1055 0 1.2002066621692222e-02
GC_9_1056 b_9 NI_9 NS_1056 0 -2.5554187856198793e-03
GC_9_1057 b_9 NI_9 NS_1057 0 -5.2431712474782398e-03
GC_9_1058 b_9 NI_9 NS_1058 0 4.7077251126198027e-03
GC_9_1059 b_9 NI_9 NS_1059 0 -6.1541426639683938e-03
GC_9_1060 b_9 NI_9 NS_1060 0 -4.3159714527651622e-03
GC_9_1061 b_9 NI_9 NS_1061 0 1.1759644470661005e-02
GC_9_1062 b_9 NI_9 NS_1062 0 -3.7148810384935028e-03
GC_9_1063 b_9 NI_9 NS_1063 0 1.3000692755248818e-02
GC_9_1064 b_9 NI_9 NS_1064 0 9.4708304140755789e-03
GC_9_1065 b_9 NI_9 NS_1065 0 3.9444980155269995e-06
GC_9_1066 b_9 NI_9 NS_1066 0 -9.3341884547428572e-07
GC_9_1067 b_9 NI_9 NS_1067 0 1.6111759272943997e-02
GC_9_1068 b_9 NI_9 NS_1068 0 1.6784783951932173e-02
GC_9_1069 b_9 NI_9 NS_1069 0 1.2052346388523776e-02
GC_9_1070 b_9 NI_9 NS_1070 0 -2.4747670936221479e-03
GC_9_1071 b_9 NI_9 NS_1071 0 -8.3473624943100917e-03
GC_9_1072 b_9 NI_9 NS_1072 0 8.3965843540299053e-05
GC_9_1073 b_9 NI_9 NS_1073 0 1.1340547357927900e-02
GC_9_1074 b_9 NI_9 NS_1074 0 7.3400065017338685e-03
GC_9_1075 b_9 NI_9 NS_1075 0 -4.6549262453052364e-03
GC_9_1076 b_9 NI_9 NS_1076 0 7.3654590976730836e-03
GC_9_1077 b_9 NI_9 NS_1077 0 -8.0793072060614569e-03
GC_9_1078 b_9 NI_9 NS_1078 0 -3.7190022515168407e-03
GC_9_1079 b_9 NI_9 NS_1079 0 1.5982962397912484e-02
GC_9_1080 b_9 NI_9 NS_1080 0 -7.7384993131403533e-03
GC_9_1081 b_9 NI_9 NS_1081 0 1.1808601739345403e-03
GC_9_1082 b_9 NI_9 NS_1082 0 -3.5561504517818890e-09
GC_9_1083 b_9 NI_9 NS_1083 0 -4.8002201619295907e-08
GC_9_1084 b_9 NI_9 NS_1084 0 -3.4752337930980621e-06
GC_9_1085 b_9 NI_9 NS_1085 0 -3.6811894665245419e-04
GC_9_1086 b_9 NI_9 NS_1086 0 1.3598159843515576e-04
GC_9_1087 b_9 NI_9 NS_1087 0 1.1297148004086330e-03
GC_9_1088 b_9 NI_9 NS_1088 0 1.9432455940075811e-03
GC_9_1089 b_9 NI_9 NS_1089 0 -6.5025362219099531e-05
GC_9_1090 b_9 NI_9 NS_1090 0 -3.4937339203136770e-03
GC_9_1091 b_9 NI_9 NS_1091 0 -1.5644030835218136e-03
GC_9_1092 b_9 NI_9 NS_1092 0 5.0905614508097042e-03
GC_9_1093 b_9 NI_9 NS_1093 0 4.2534104358233323e-03
GC_9_1094 b_9 NI_9 NS_1094 0 -4.9937797865619929e-03
GC_9_1095 b_9 NI_9 NS_1095 0 -1.0085420667727239e-03
GC_9_1096 b_9 NI_9 NS_1096 0 5.6396308343254994e-04
GC_9_1097 b_9 NI_9 NS_1097 0 -2.0807418986295637e-03
GC_9_1098 b_9 NI_9 NS_1098 0 -1.8633296175920790e-03
GC_9_1099 b_9 NI_9 NS_1099 0 3.6453743243149588e-03
GC_9_1100 b_9 NI_9 NS_1100 0 1.1647299721461420e-02
GC_9_1101 b_9 NI_9 NS_1101 0 -8.9809376412818530e-04
GC_9_1102 b_9 NI_9 NS_1102 0 -1.4854264015549987e-02
GC_9_1103 b_9 NI_9 NS_1103 0 -8.1235082744215009e-03
GC_9_1104 b_9 NI_9 NS_1104 0 1.9195541370244941e-03
GC_9_1105 b_9 NI_9 NS_1105 0 1.1262993899966392e-02
GC_9_1106 b_9 NI_9 NS_1106 0 -1.8122030646776197e-03
GC_9_1107 b_9 NI_9 NS_1107 0 -7.5672396693017199e-03
GC_9_1108 b_9 NI_9 NS_1108 0 -1.6812110656908249e-03
GC_9_1109 b_9 NI_9 NS_1109 0 1.5281607338987563e-02
GC_9_1110 b_9 NI_9 NS_1110 0 5.3008467150268612e-03
GC_9_1111 b_9 NI_9 NS_1111 0 -1.3082790601246279e-02
GC_9_1112 b_9 NI_9 NS_1112 0 -5.4613195741109099e-03
GC_9_1113 b_9 NI_9 NS_1113 0 -6.6370644341743265e-03
GC_9_1114 b_9 NI_9 NS_1114 0 3.4566491501496041e-03
GC_9_1115 b_9 NI_9 NS_1115 0 6.3615686418213102e-03
GC_9_1116 b_9 NI_9 NS_1116 0 -1.8793111909258396e-03
GC_9_1117 b_9 NI_9 NS_1117 0 -5.4737174823897769e-03
GC_9_1118 b_9 NI_9 NS_1118 0 2.1829945210677278e-03
GC_9_1119 b_9 NI_9 NS_1119 0 5.3937402484606749e-03
GC_9_1120 b_9 NI_9 NS_1120 0 -2.6324139397167837e-03
GC_9_1121 b_9 NI_9 NS_1121 0 -6.3064434681043766e-03
GC_9_1122 b_9 NI_9 NS_1122 0 -4.8383766170783808e-04
GC_9_1123 b_9 NI_9 NS_1123 0 7.6452212090595273e-03
GC_9_1124 b_9 NI_9 NS_1124 0 3.6298699377661880e-03
GC_9_1125 b_9 NI_9 NS_1125 0 -5.8336100716466794e-03
GC_9_1126 b_9 NI_9 NS_1126 0 -3.4646020589867849e-03
GC_9_1127 b_9 NI_9 NS_1127 0 2.9619270154026872e-04
GC_9_1128 b_9 NI_9 NS_1128 0 5.5809921323421332e-04
GC_9_1129 b_9 NI_9 NS_1129 0 -4.9270674088371085e-03
GC_9_1130 b_9 NI_9 NS_1130 0 8.9217933472828372e-04
GC_9_1131 b_9 NI_9 NS_1131 0 6.2062906001026730e-03
GC_9_1132 b_9 NI_9 NS_1132 0 6.8829116828021078e-04
GC_9_1133 b_9 NI_9 NS_1133 0 -5.3209606423650089e-03
GC_9_1134 b_9 NI_9 NS_1134 0 -4.8420041089506559e-04
GC_9_1135 b_9 NI_9 NS_1135 0 1.5503170145523498e-03
GC_9_1136 b_9 NI_9 NS_1136 0 -4.3200389211300233e-05
GC_9_1137 b_9 NI_9 NS_1137 0 -6.0223399978072689e-03
GC_9_1138 b_9 NI_9 NS_1138 0 1.9232230871372869e-03
GC_9_1139 b_9 NI_9 NS_1139 0 6.2616320411048544e-03
GC_9_1140 b_9 NI_9 NS_1140 0 2.1740092674760932e-04
GC_9_1141 b_9 NI_9 NS_1141 0 -5.0592004869657948e-03
GC_9_1142 b_9 NI_9 NS_1142 0 1.7016082211229375e-03
GC_9_1143 b_9 NI_9 NS_1143 0 2.4884719812637217e-03
GC_9_1144 b_9 NI_9 NS_1144 0 -9.5763486206161780e-04
GC_9_1145 b_9 NI_9 NS_1145 0 -6.5329668169025823e-03
GC_9_1146 b_9 NI_9 NS_1146 0 3.8846211805320103e-03
GC_9_1147 b_9 NI_9 NS_1147 0 7.4932612544989499e-03
GC_9_1148 b_9 NI_9 NS_1148 0 -1.0960049926959493e-03
GC_9_1149 b_9 NI_9 NS_1149 0 -3.9851227910626614e-03
GC_9_1150 b_9 NI_9 NS_1150 0 4.0409663137630381e-03
GC_9_1151 b_9 NI_9 NS_1151 0 2.8633248923082711e-03
GC_9_1152 b_9 NI_9 NS_1152 0 -3.0534840298028073e-03
GC_9_1153 b_9 NI_9 NS_1153 0 -6.0227358976724862e-03
GC_9_1154 b_9 NI_9 NS_1154 0 7.2373634148455044e-03
GC_9_1155 b_9 NI_9 NS_1155 0 7.9896911475281929e-03
GC_9_1156 b_9 NI_9 NS_1156 0 -4.8114454952552215e-03
GC_9_1157 b_9 NI_9 NS_1157 0 -5.3743564158331258e-04
GC_9_1158 b_9 NI_9 NS_1158 0 5.0204611318347839e-03
GC_9_1159 b_9 NI_9 NS_1159 0 2.4825046595649999e-04
GC_9_1160 b_9 NI_9 NS_1160 0 -4.7581887208284872e-03
GC_9_1161 b_9 NI_9 NS_1161 0 1.8107928900694784e-09
GC_9_1162 b_9 NI_9 NS_1162 0 3.2741501040610477e-09
GC_9_1163 b_9 NI_9 NS_1163 0 -1.4272198943202567e-03
GC_9_1164 b_9 NI_9 NS_1164 0 7.8707210220527197e-03
GC_9_1165 b_9 NI_9 NS_1165 0 -1.7999304571094510e-04
GC_9_1166 b_9 NI_9 NS_1166 0 3.0272429820567058e-03
GC_9_1167 b_9 NI_9 NS_1167 0 -1.3039321363534197e-04
GC_9_1168 b_9 NI_9 NS_1168 0 -3.3752920552105122e-03
GC_9_1169 b_9 NI_9 NS_1169 0 -8.7633793226019714e-04
GC_9_1170 b_9 NI_9 NS_1170 0 7.5304798544569215e-03
GC_9_1171 b_9 NI_9 NS_1171 0 3.7887923511289970e-03
GC_9_1172 b_9 NI_9 NS_1172 0 -6.1573981675861842e-03
GC_9_1173 b_9 NI_9 NS_1173 0 8.6224200991830757e-08
GC_9_1174 b_9 NI_9 NS_1174 0 -3.5295605187739513e-07
GC_9_1175 b_9 NI_9 NS_1175 0 6.7186821084001848e-03
GC_9_1176 b_9 NI_9 NS_1176 0 -5.3194058456995531e-03
GC_9_1177 b_9 NI_9 NS_1177 0 -2.6111750021722232e-03
GC_9_1178 b_9 NI_9 NS_1178 0 6.0542434733270884e-03
GC_9_1179 b_9 NI_9 NS_1179 0 -4.2922721003970940e-03
GC_9_1180 b_9 NI_9 NS_1180 0 1.4428546680433891e-05
GC_9_1181 b_9 NI_9 NS_1181 0 2.7173858195240013e-03
GC_9_1182 b_9 NI_9 NS_1182 0 -6.2039927976012725e-03
GC_9_1183 b_9 NI_9 NS_1183 0 2.0957202069937977e-03
GC_9_1184 b_9 NI_9 NS_1184 0 3.2562858946082549e-03
GC_9_1185 b_9 NI_9 NS_1185 0 -1.9700288888946996e-03
GC_9_1186 b_9 NI_9 NS_1186 0 -4.4205336936084961e-03
GC_9_1187 b_9 NI_9 NS_1187 0 2.8640819012434363e-03
GC_9_1188 b_9 NI_9 NS_1188 0 8.0083594488233913e-03
GC_9_1189 b_9 NI_9 NS_1189 0 -3.3036440496388309e-03
GC_9_1190 b_9 NI_9 NS_1190 0 1.8493852990039438e-09
GC_9_1191 b_9 NI_9 NS_1191 0 5.6032181727570970e-08
GC_9_1192 b_9 NI_9 NS_1192 0 1.8929694726481910e-06
GC_9_1193 b_9 NI_9 NS_1193 0 -9.1167730377775055e-05
GC_9_1194 b_9 NI_9 NS_1194 0 -5.7737930953436403e-05
GC_9_1195 b_9 NI_9 NS_1195 0 -1.2657732650326302e-03
GC_9_1196 b_9 NI_9 NS_1196 0 -2.9559391213972711e-04
GC_9_1197 b_9 NI_9 NS_1197 0 -1.6792135009617308e-03
GC_9_1198 b_9 NI_9 NS_1198 0 2.6464975853239003e-03
GC_9_1199 b_9 NI_9 NS_1199 0 5.1121163694870734e-04
GC_9_1200 b_9 NI_9 NS_1200 0 5.4276087233707882e-03
GC_9_1201 b_9 NI_9 NS_1201 0 7.1034879093775892e-03
GC_9_1202 b_9 NI_9 NS_1202 0 6.3629218728458053e-04
GC_9_1203 b_9 NI_9 NS_1203 0 6.4432949284838224e-04
GC_9_1204 b_9 NI_9 NS_1204 0 -6.6091956934284733e-04
GC_9_1205 b_9 NI_9 NS_1205 0 1.0576978538098197e-03
GC_9_1206 b_9 NI_9 NS_1206 0 1.5711412082406503e-03
GC_9_1207 b_9 NI_9 NS_1207 0 1.2687514000960961e-02
GC_9_1208 b_9 NI_9 NS_1208 0 1.3123213842793620e-02
GC_9_1209 b_9 NI_9 NS_1209 0 8.7187980280740620e-03
GC_9_1210 b_9 NI_9 NS_1210 0 -2.0392080770404941e-02
GC_9_1211 b_9 NI_9 NS_1211 0 8.3891007675096149e-03
GC_9_1212 b_9 NI_9 NS_1212 0 -2.9045258231576486e-03
GC_9_1213 b_9 NI_9 NS_1213 0 -1.2701289616757108e-02
GC_9_1214 b_9 NI_9 NS_1214 0 -3.8806698559281830e-02
GC_9_1215 b_9 NI_9 NS_1215 0 -7.2523391607987623e-03
GC_9_1216 b_9 NI_9 NS_1216 0 -2.1332749486277251e-03
GC_9_1217 b_9 NI_9 NS_1217 0 -5.2307199518102629e-02
GC_9_1218 b_9 NI_9 NS_1218 0 -1.7936156154075005e-03
GC_9_1219 b_9 NI_9 NS_1219 0 1.4914415704611370e-02
GC_9_1220 b_9 NI_9 NS_1220 0 8.6735766433999103e-03
GC_9_1221 b_9 NI_9 NS_1221 0 -5.9233530129432872e-03
GC_9_1222 b_9 NI_9 NS_1222 0 5.0044974747570099e-03
GC_9_1223 b_9 NI_9 NS_1223 0 8.3724199730542733e-03
GC_9_1224 b_9 NI_9 NS_1224 0 1.1688363041629256e-02
GC_9_1225 b_9 NI_9 NS_1225 0 4.5592638427856668e-03
GC_9_1226 b_9 NI_9 NS_1226 0 -2.9327411502679656e-03
GC_9_1227 b_9 NI_9 NS_1227 0 -7.8986738210523374e-03
GC_9_1228 b_9 NI_9 NS_1228 0 -8.1490651708686825e-03
GC_9_1229 b_9 NI_9 NS_1229 0 -5.6808140380008344e-03
GC_9_1230 b_9 NI_9 NS_1230 0 -6.1281001254625373e-04
GC_9_1231 b_9 NI_9 NS_1231 0 -1.8070850582016330e-02
GC_9_1232 b_9 NI_9 NS_1232 0 1.3578965336294211e-02
GC_9_1233 b_9 NI_9 NS_1233 0 4.7069865927157669e-03
GC_9_1234 b_9 NI_9 NS_1234 0 4.3794388494791834e-03
GC_9_1235 b_9 NI_9 NS_1235 0 6.5015827899565564e-04
GC_9_1236 b_9 NI_9 NS_1236 0 -1.0995438866251910e-04
GC_9_1237 b_9 NI_9 NS_1237 0 -3.7964000712596988e-03
GC_9_1238 b_9 NI_9 NS_1238 0 8.8498888791788762e-04
GC_9_1239 b_9 NI_9 NS_1239 0 -1.1178276217446753e-03
GC_9_1240 b_9 NI_9 NS_1240 0 1.6699689447770082e-02
GC_9_1241 b_9 NI_9 NS_1241 0 4.4472808489183537e-03
GC_9_1242 b_9 NI_9 NS_1242 0 7.0796446279316474e-04
GC_9_1243 b_9 NI_9 NS_1243 0 -5.1995804564576825e-04
GC_9_1244 b_9 NI_9 NS_1244 0 -2.2477509841922040e-03
GC_9_1245 b_9 NI_9 NS_1245 0 -4.9864557315705835e-03
GC_9_1246 b_9 NI_9 NS_1246 0 2.1108879594370889e-03
GC_9_1247 b_9 NI_9 NS_1247 0 7.3425285253475572e-03
GC_9_1248 b_9 NI_9 NS_1248 0 1.4345855671288942e-02
GC_9_1249 b_9 NI_9 NS_1249 0 4.1872276218322896e-03
GC_9_1250 b_9 NI_9 NS_1250 0 -1.6838583578748683e-03
GC_9_1251 b_9 NI_9 NS_1251 0 -3.3981244613817841e-03
GC_9_1252 b_9 NI_9 NS_1252 0 -2.1006228483129922e-03
GC_9_1253 b_9 NI_9 NS_1253 0 -5.4204253675511349e-03
GC_9_1254 b_9 NI_9 NS_1254 0 4.3817251608101399e-03
GC_9_1255 b_9 NI_9 NS_1255 0 1.3196874516908940e-02
GC_9_1256 b_9 NI_9 NS_1256 0 8.4333068839489850e-03
GC_9_1257 b_9 NI_9 NS_1257 0 2.8324343455928464e-03
GC_9_1258 b_9 NI_9 NS_1258 0 -4.1306062545731345e-03
GC_9_1259 b_9 NI_9 NS_1259 0 -5.3207859139795480e-03
GC_9_1260 b_9 NI_9 NS_1260 0 1.1381580917244102e-03
GC_9_1261 b_9 NI_9 NS_1261 0 -4.4310202375813850e-03
GC_9_1262 b_9 NI_9 NS_1262 0 8.3104314799015838e-03
GC_9_1263 b_9 NI_9 NS_1263 0 1.4612787176392996e-02
GC_9_1264 b_9 NI_9 NS_1264 0 -4.6824808428590583e-04
GC_9_1265 b_9 NI_9 NS_1265 0 -1.1845312544063750e-03
GC_9_1266 b_9 NI_9 NS_1266 0 -4.5473900694159236e-03
GC_9_1267 b_9 NI_9 NS_1267 0 -2.2825675268084238e-03
GC_9_1268 b_9 NI_9 NS_1268 0 4.3832539464182209e-03
GC_9_1269 b_9 NI_9 NS_1269 0 1.3571801834910809e-10
GC_9_1270 b_9 NI_9 NS_1270 0 -1.5466404332868415e-09
GC_9_1271 b_9 NI_9 NS_1271 0 1.4460267395114291e-03
GC_9_1272 b_9 NI_9 NS_1272 0 8.2165466488516581e-03
GC_9_1273 b_9 NI_9 NS_1273 0 -8.7895013781721801e-04
GC_9_1274 b_9 NI_9 NS_1274 0 -2.2072129621422006e-03
GC_9_1275 b_9 NI_9 NS_1275 0 -1.4679136924828696e-03
GC_9_1276 b_9 NI_9 NS_1276 0 2.7519856011815826e-03
GC_9_1277 b_9 NI_9 NS_1277 0 1.7320146128120993e-03
GC_9_1278 b_9 NI_9 NS_1278 0 7.6059319906844336e-03
GC_9_1279 b_9 NI_9 NS_1279 0 7.5874087584804116e-03
GC_9_1280 b_9 NI_9 NS_1280 0 -3.8276835723259242e-03
GC_9_1281 b_9 NI_9 NS_1281 0 -5.2101127048442273e-08
GC_9_1282 b_9 NI_9 NS_1282 0 -2.0817452725125374e-08
GC_9_1283 b_9 NI_9 NS_1283 0 1.1391243353869363e-02
GC_9_1284 b_9 NI_9 NS_1284 0 4.4700328609421853e-03
GC_9_1285 b_9 NI_9 NS_1285 0 -8.6185040455332145e-04
GC_9_1286 b_9 NI_9 NS_1286 0 6.4916224558386739e-03
GC_9_1287 b_9 NI_9 NS_1287 0 3.6263738639324100e-03
GC_9_1288 b_9 NI_9 NS_1288 0 4.0710465875459486e-04
GC_9_1289 b_9 NI_9 NS_1289 0 6.0525104336892430e-03
GC_9_1290 b_9 NI_9 NS_1290 0 -4.6635404939705033e-03
GC_9_1291 b_9 NI_9 NS_1291 0 -3.3929752774385460e-03
GC_9_1292 b_9 NI_9 NS_1292 0 -1.3533960148467020e-03
GC_9_1293 b_9 NI_9 NS_1293 0 1.1237968653240769e-04
GC_9_1294 b_9 NI_9 NS_1294 0 4.4958002104339007e-03
GC_9_1295 b_9 NI_9 NS_1295 0 7.2795569588585815e-03
GC_9_1296 b_9 NI_9 NS_1296 0 5.5305048407844008e-03
GD_9_1 b_9 NI_9 NA_1 0 -1.1809815270069599e-06
GD_9_2 b_9 NI_9 NA_2 0 8.8077022209712270e-06
GD_9_3 b_9 NI_9 NA_3 0 -7.3787539613406628e-06
GD_9_4 b_9 NI_9 NA_4 0 2.0978275349305061e-06
GD_9_5 b_9 NI_9 NA_5 0 -3.7841747996511557e-07
GD_9_6 b_9 NI_9 NA_6 0 1.5903935805109086e-05
GD_9_7 b_9 NI_9 NA_7 0 2.6298650779412850e-05
GD_9_8 b_9 NI_9 NA_8 0 1.0461291060168750e-04
GD_9_9 b_9 NI_9 NA_9 0 -1.0894630938571586e-02
GD_9_10 b_9 NI_9 NA_10 0 -5.0003173062905405e-03
GD_9_11 b_9 NI_9 NA_11 0 1.0616351945255143e-02
GD_9_12 b_9 NI_9 NA_12 0 -1.1524162700684187e-03
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 -6.4269108890426031e-05
GC_10_2 b_10 NI_10 NS_2 0 3.5608758750194558e-12
GC_10_3 b_10 NI_10 NS_3 0 5.0181455014832888e-11
GC_10_4 b_10 NI_10 NS_4 0 -1.5818258186118837e-09
GC_10_5 b_10 NI_10 NS_5 0 -1.0723785347193048e-06
GC_10_6 b_10 NI_10 NS_6 0 -1.0588572002217353e-06
GC_10_7 b_10 NI_10 NS_7 0 4.0966300862679092e-07
GC_10_8 b_10 NI_10 NS_8 0 3.5700924166291026e-07
GC_10_9 b_10 NI_10 NS_9 0 -2.2606370969952933e-06
GC_10_10 b_10 NI_10 NS_10 0 2.1080754795648527e-06
GC_10_11 b_10 NI_10 NS_11 0 -2.5321226812747143e-06
GC_10_12 b_10 NI_10 NS_12 0 -1.2387507638221284e-06
GC_10_13 b_10 NI_10 NS_13 0 1.3985171664019561e-06
GC_10_14 b_10 NI_10 NS_14 0 9.9857056756006000e-07
GC_10_15 b_10 NI_10 NS_15 0 -1.1234361617478999e-06
GC_10_16 b_10 NI_10 NS_16 0 1.3407171178731672e-06
GC_10_17 b_10 NI_10 NS_17 0 7.2717033380081709e-07
GC_10_18 b_10 NI_10 NS_18 0 3.0410821437297618e-06
GC_10_19 b_10 NI_10 NS_19 0 -2.8465566244158362e-06
GC_10_20 b_10 NI_10 NS_20 0 4.7261396987540701e-07
GC_10_21 b_10 NI_10 NS_21 0 3.6885481355640843e-06
GC_10_22 b_10 NI_10 NS_22 0 -2.0179897534361182e-06
GC_10_23 b_10 NI_10 NS_23 0 -1.8785477894481499e-07
GC_10_24 b_10 NI_10 NS_24 0 2.5632237281484920e-06
GC_10_25 b_10 NI_10 NS_25 0 -4.0642271614605739e-06
GC_10_26 b_10 NI_10 NS_26 0 4.8362651360148793e-06
GC_10_27 b_10 NI_10 NS_27 0 6.4243497804642389e-07
GC_10_28 b_10 NI_10 NS_28 0 -1.5864771096893328e-06
GC_10_29 b_10 NI_10 NS_29 0 4.6099988334889110e-06
GC_10_30 b_10 NI_10 NS_30 0 9.9431005821945181e-06
GC_10_31 b_10 NI_10 NS_31 0 -1.1101182983381940e-07
GC_10_32 b_10 NI_10 NS_32 0 5.2381959014459952e-07
GC_10_33 b_10 NI_10 NS_33 0 -6.3534472844856835e-09
GC_10_34 b_10 NI_10 NS_34 0 -7.8556148182460921e-07
GC_10_35 b_10 NI_10 NS_35 0 5.3519045022033963e-06
GC_10_36 b_10 NI_10 NS_36 0 4.9534794708461480e-07
GC_10_37 b_10 NI_10 NS_37 0 8.4640691220787019e-07
GC_10_38 b_10 NI_10 NS_38 0 1.9176163953696913e-06
GC_10_39 b_10 NI_10 NS_39 0 3.0829094526442717e-08
GC_10_40 b_10 NI_10 NS_40 0 1.1331876659154334e-06
GC_10_41 b_10 NI_10 NS_41 0 5.8507489929243412e-07
GC_10_42 b_10 NI_10 NS_42 0 -1.1108574654615857e-06
GC_10_43 b_10 NI_10 NS_43 0 5.8253754159859358e-06
GC_10_44 b_10 NI_10 NS_44 0 4.0748102815353696e-06
GC_10_45 b_10 NI_10 NS_45 0 6.0627770353371994e-07
GC_10_46 b_10 NI_10 NS_46 0 8.5953268538909556e-07
GC_10_47 b_10 NI_10 NS_47 0 1.9692641404286799e-07
GC_10_48 b_10 NI_10 NS_48 0 2.4097902082097051e-07
GC_10_49 b_10 NI_10 NS_49 0 8.4525379212601115e-07
GC_10_50 b_10 NI_10 NS_50 0 -6.7217933148134213e-07
GC_10_51 b_10 NI_10 NS_51 0 6.6650675856957109e-06
GC_10_52 b_10 NI_10 NS_52 0 7.5450089134820570e-07
GC_10_53 b_10 NI_10 NS_53 0 7.7455830846526781e-07
GC_10_54 b_10 NI_10 NS_54 0 7.4914083012606946e-07
GC_10_55 b_10 NI_10 NS_55 0 6.6483861121411665e-07
GC_10_56 b_10 NI_10 NS_56 0 -6.6207048315799222e-08
GC_10_57 b_10 NI_10 NS_57 0 8.7154214197483277e-07
GC_10_58 b_10 NI_10 NS_58 0 -6.4039890914913032e-07
GC_10_59 b_10 NI_10 NS_59 0 5.7751873474465618e-06
GC_10_60 b_10 NI_10 NS_60 0 -1.5909440827247247e-06
GC_10_61 b_10 NI_10 NS_61 0 8.2383230968136076e-07
GC_10_62 b_10 NI_10 NS_62 0 5.6704141614970717e-07
GC_10_63 b_10 NI_10 NS_63 0 6.2584342657758000e-07
GC_10_64 b_10 NI_10 NS_64 0 -5.5330724255698057e-07
GC_10_65 b_10 NI_10 NS_65 0 9.3776534406016582e-07
GC_10_66 b_10 NI_10 NS_66 0 -4.4580075140251181e-07
GC_10_67 b_10 NI_10 NS_67 0 3.9036809076630920e-06
GC_10_68 b_10 NI_10 NS_68 0 -2.9906803793788682e-06
GC_10_69 b_10 NI_10 NS_69 0 8.9572364625214876e-07
GC_10_70 b_10 NI_10 NS_70 0 3.2737991597797378e-07
GC_10_71 b_10 NI_10 NS_71 0 2.1610865723822126e-07
GC_10_72 b_10 NI_10 NS_72 0 -7.9557875152650822e-07
GC_10_73 b_10 NI_10 NS_73 0 1.1598906744963746e-06
GC_10_74 b_10 NI_10 NS_74 0 -3.2475047855096002e-07
GC_10_75 b_10 NI_10 NS_75 0 1.6774796610394616e-06
GC_10_76 b_10 NI_10 NS_76 0 -3.0902024037437805e-06
GC_10_77 b_10 NI_10 NS_77 0 7.9113858640234788e-07
GC_10_78 b_10 NI_10 NS_78 0 -1.0639300978828699e-07
GC_10_79 b_10 NI_10 NS_79 0 -1.9702131690300841e-07
GC_10_80 b_10 NI_10 NS_80 0 -4.0861489060034292e-07
GC_10_81 b_10 NI_10 NS_81 0 8.5881251995136321e-12
GC_10_82 b_10 NI_10 NS_82 0 -1.5730105129151757e-11
GC_10_83 b_10 NI_10 NS_83 0 8.3872041058784440e-07
GC_10_84 b_10 NI_10 NS_84 0 -5.9377995317625628e-07
GC_10_85 b_10 NI_10 NS_85 0 4.9464521979581797e-07
GC_10_86 b_10 NI_10 NS_86 0 -3.5993780553851340e-08
GC_10_87 b_10 NI_10 NS_87 0 1.7010424530273983e-08
GC_10_88 b_10 NI_10 NS_88 0 -8.9112330998567741e-08
GC_10_89 b_10 NI_10 NS_89 0 5.2142270375326500e-07
GC_10_90 b_10 NI_10 NS_90 0 -1.7666132512227204e-08
GC_10_91 b_10 NI_10 NS_91 0 7.0518168166708437e-07
GC_10_92 b_10 NI_10 NS_92 0 -1.5614012758353395e-06
GC_10_93 b_10 NI_10 NS_93 0 4.0969092083715271e-10
GC_10_94 b_10 NI_10 NS_94 0 -5.8070917541870383e-10
GC_10_95 b_10 NI_10 NS_95 0 1.0099580941119874e-06
GC_10_96 b_10 NI_10 NS_96 0 -2.7386510703689203e-07
GC_10_97 b_10 NI_10 NS_97 0 3.5400836409920230e-07
GC_10_98 b_10 NI_10 NS_98 0 -1.7369728097408382e-07
GC_10_99 b_10 NI_10 NS_99 0 2.5492786403301221e-07
GC_10_100 b_10 NI_10 NS_100 0 2.6554572000272137e-08
GC_10_101 b_10 NI_10 NS_101 0 1.0857963314011963e-06
GC_10_102 b_10 NI_10 NS_102 0 -1.1750272418524408e-06
GC_10_103 b_10 NI_10 NS_103 0 6.5375759781831876e-07
GC_10_104 b_10 NI_10 NS_104 0 -3.3455320129086688e-07
GC_10_105 b_10 NI_10 NS_105 0 -2.1221596652350446e-07
GC_10_106 b_10 NI_10 NS_106 0 -9.8558852101661869e-08
GC_10_107 b_10 NI_10 NS_107 0 7.5732270626047558e-07
GC_10_108 b_10 NI_10 NS_108 0 3.2283849815584856e-07
GC_10_109 b_10 NI_10 NS_109 0 8.5353700624147858e-06
GC_10_110 b_10 NI_10 NS_110 0 3.7657768617705082e-12
GC_10_111 b_10 NI_10 NS_111 0 -7.8556130961095725e-11
GC_10_112 b_10 NI_10 NS_112 0 2.5472496702927444e-09
GC_10_113 b_10 NI_10 NS_113 0 1.5491020765872179e-08
GC_10_114 b_10 NI_10 NS_114 0 -8.4748458881662903e-08
GC_10_115 b_10 NI_10 NS_115 0 -2.4892835619274395e-07
GC_10_116 b_10 NI_10 NS_116 0 2.7099899152356496e-07
GC_10_117 b_10 NI_10 NS_117 0 7.4290255262160684e-07
GC_10_118 b_10 NI_10 NS_118 0 -2.8388539126079625e-07
GC_10_119 b_10 NI_10 NS_119 0 -9.6871922496031026e-07
GC_10_120 b_10 NI_10 NS_120 0 -2.3710765523206016e-07
GC_10_121 b_10 NI_10 NS_121 0 1.0260921059904393e-06
GC_10_122 b_10 NI_10 NS_122 0 4.0158025825205399e-07
GC_10_123 b_10 NI_10 NS_123 0 -1.2037277634538657e-07
GC_10_124 b_10 NI_10 NS_124 0 -2.7297926830364584e-07
GC_10_125 b_10 NI_10 NS_125 0 1.1063191900759817e-07
GC_10_126 b_10 NI_10 NS_126 0 -5.1161012849712046e-07
GC_10_127 b_10 NI_10 NS_127 0 -2.0841508442339258e-06
GC_10_128 b_10 NI_10 NS_128 0 8.6187339057261830e-07
GC_10_129 b_10 NI_10 NS_129 0 2.4334043652988738e-06
GC_10_130 b_10 NI_10 NS_130 0 -6.0600247408563596e-07
GC_10_131 b_10 NI_10 NS_131 0 -6.6287068478942835e-07
GC_10_132 b_10 NI_10 NS_132 0 -1.3976073131859868e-06
GC_10_133 b_10 NI_10 NS_133 0 4.2935248193319887e-07
GC_10_134 b_10 NI_10 NS_134 0 1.8452587732663383e-06
GC_10_135 b_10 NI_10 NS_135 0 -3.0162674146901214e-08
GC_10_136 b_10 NI_10 NS_136 0 -1.3237442430671560e-06
GC_10_137 b_10 NI_10 NS_137 0 -6.3111983789746830e-07
GC_10_138 b_10 NI_10 NS_138 0 2.5911451686118873e-06
GC_10_139 b_10 NI_10 NS_139 0 4.5382333845921617e-07
GC_10_140 b_10 NI_10 NS_140 0 -2.2434946956157334e-06
GC_10_141 b_10 NI_10 NS_141 0 -7.9908829542931484e-07
GC_10_142 b_10 NI_10 NS_142 0 -9.3142308863414328e-07
GC_10_143 b_10 NI_10 NS_143 0 3.6009684176601221e-07
GC_10_144 b_10 NI_10 NS_144 0 9.1166072207042383e-07
GC_10_145 b_10 NI_10 NS_145 0 -5.5608516347296237e-07
GC_10_146 b_10 NI_10 NS_146 0 -7.2540367862801529e-07
GC_10_147 b_10 NI_10 NS_147 0 4.7741247347118549e-07
GC_10_148 b_10 NI_10 NS_148 0 7.3899263488888040e-07
GC_10_149 b_10 NI_10 NS_149 0 -1.7328934405028428e-07
GC_10_150 b_10 NI_10 NS_150 0 -8.7767189638710877e-07
GC_10_151 b_10 NI_10 NS_151 0 -3.3590723320584951e-07
GC_10_152 b_10 NI_10 NS_152 0 1.1576102654953951e-06
GC_10_153 b_10 NI_10 NS_153 0 2.5415469249157632e-07
GC_10_154 b_10 NI_10 NS_154 0 -8.4414324156421600e-07
GC_10_155 b_10 NI_10 NS_155 0 -6.4136896819129982e-08
GC_10_156 b_10 NI_10 NS_156 0 6.7381110760600436e-08
GC_10_157 b_10 NI_10 NS_157 0 -2.5853724782441283e-07
GC_10_158 b_10 NI_10 NS_158 0 -5.4962212254448558e-07
GC_10_159 b_10 NI_10 NS_159 0 1.8909308094272547e-07
GC_10_160 b_10 NI_10 NS_160 0 7.1454065646060009e-07
GC_10_161 b_10 NI_10 NS_161 0 -7.9752782808398507e-08
GC_10_162 b_10 NI_10 NS_162 0 -6.3559736895309935e-07
GC_10_163 b_10 NI_10 NS_163 0 1.0309127192158649e-07
GC_10_164 b_10 NI_10 NS_164 0 1.0288960112750457e-07
GC_10_165 b_10 NI_10 NS_165 0 -2.8962091301816065e-07
GC_10_166 b_10 NI_10 NS_166 0 -5.9366746260631026e-07
GC_10_167 b_10 NI_10 NS_167 0 1.6267859619129108e-07
GC_10_168 b_10 NI_10 NS_168 0 2.2629219517892758e-07
GC_10_169 b_10 NI_10 NS_169 0 -2.5661136063185844e-07
GC_10_170 b_10 NI_10 NS_170 0 -5.0830136335299795e-07
GC_10_171 b_10 NI_10 NS_171 0 4.8280469242091466e-08
GC_10_172 b_10 NI_10 NS_172 0 -5.1510934363974057e-08
GC_10_173 b_10 NI_10 NS_173 0 -3.6755823972693761e-07
GC_10_174 b_10 NI_10 NS_174 0 -5.5772119588974828e-07
GC_10_175 b_10 NI_10 NS_175 0 -2.3473064752707004e-07
GC_10_176 b_10 NI_10 NS_176 0 1.8282672799804991e-08
GC_10_177 b_10 NI_10 NS_177 0 -4.3348900929002551e-07
GC_10_178 b_10 NI_10 NS_178 0 -3.4064050988712810e-07
GC_10_179 b_10 NI_10 NS_179 0 -1.2461967823361119e-07
GC_10_180 b_10 NI_10 NS_180 0 1.5315385421594747e-08
GC_10_181 b_10 NI_10 NS_181 0 -5.6246373021391801e-07
GC_10_182 b_10 NI_10 NS_182 0 -4.3868127399372494e-07
GC_10_183 b_10 NI_10 NS_183 0 -3.1884387224145043e-07
GC_10_184 b_10 NI_10 NS_184 0 3.1347573808402908e-07
GC_10_185 b_10 NI_10 NS_185 0 -4.9949272723744761e-07
GC_10_186 b_10 NI_10 NS_186 0 3.7092806758786055e-08
GC_10_187 b_10 NI_10 NS_187 0 -1.1552577779069757e-08
GC_10_188 b_10 NI_10 NS_188 0 6.1370299990161728e-08
GC_10_189 b_10 NI_10 NS_189 0 -3.2703261597867943e-12
GC_10_190 b_10 NI_10 NS_190 0 3.1967999152808639e-12
GC_10_191 b_10 NI_10 NS_191 0 -5.7559168562679915e-07
GC_10_192 b_10 NI_10 NS_192 0 4.6740601092655766e-08
GC_10_193 b_10 NI_10 NS_193 0 -2.8964972465063667e-07
GC_10_194 b_10 NI_10 NS_194 0 1.1772129605619192e-07
GC_10_195 b_10 NI_10 NS_195 0 -6.5539810391817466e-09
GC_10_196 b_10 NI_10 NS_196 0 -6.9121965074688752e-08
GC_10_197 b_10 NI_10 NS_197 0 -6.5992747763213768e-07
GC_10_198 b_10 NI_10 NS_198 0 1.4030089581685533e-07
GC_10_199 b_10 NI_10 NS_199 0 2.8354547143241159e-08
GC_10_200 b_10 NI_10 NS_200 0 1.2330380072297451e-07
GC_10_201 b_10 NI_10 NS_201 0 -6.1637907142462932e-11
GC_10_202 b_10 NI_10 NS_202 0 1.2851412777033574e-10
GC_10_203 b_10 NI_10 NS_203 0 -3.4587920567088551e-08
GC_10_204 b_10 NI_10 NS_204 0 1.9625711966471574e-07
GC_10_205 b_10 NI_10 NS_205 0 -3.6686783410728681e-07
GC_10_206 b_10 NI_10 NS_206 0 -4.3787001940233118e-08
GC_10_207 b_10 NI_10 NS_207 0 -1.8653370863054718e-07
GC_10_208 b_10 NI_10 NS_208 0 -2.5483454371866319e-09
GC_10_209 b_10 NI_10 NS_209 0 1.9191377815368131e-07
GC_10_210 b_10 NI_10 NS_210 0 8.0894788954571862e-08
GC_10_211 b_10 NI_10 NS_211 0 -2.6556159497573972e-07
GC_10_212 b_10 NI_10 NS_212 0 3.1336803394772729e-07
GC_10_213 b_10 NI_10 NS_213 0 1.2476995782362210e-07
GC_10_214 b_10 NI_10 NS_214 0 -1.4419545217123531e-07
GC_10_215 b_10 NI_10 NS_215 0 -5.7833727547586693e-08
GC_10_216 b_10 NI_10 NS_216 0 2.3865277845550552e-07
GC_10_217 b_10 NI_10 NS_217 0 -7.7926469607543148e-06
GC_10_218 b_10 NI_10 NS_218 0 -1.0504553293629061e-11
GC_10_219 b_10 NI_10 NS_219 0 7.2835290804815884e-11
GC_10_220 b_10 NI_10 NS_220 0 -4.8050685243348332e-09
GC_10_221 b_10 NI_10 NS_221 0 -9.4069119524022573e-07
GC_10_222 b_10 NI_10 NS_222 0 -7.1603752389800015e-07
GC_10_223 b_10 NI_10 NS_223 0 6.8892042719230800e-07
GC_10_224 b_10 NI_10 NS_224 0 1.1980952793237308e-06
GC_10_225 b_10 NI_10 NS_225 0 -6.5943776501471717e-07
GC_10_226 b_10 NI_10 NS_226 0 2.7654897297284690e-06
GC_10_227 b_10 NI_10 NS_227 0 -1.7473377694920539e-07
GC_10_228 b_10 NI_10 NS_228 0 -8.3537114387099478e-07
GC_10_229 b_10 NI_10 NS_229 0 3.2530593163678559e-06
GC_10_230 b_10 NI_10 NS_230 0 -1.7278300353205874e-06
GC_10_231 b_10 NI_10 NS_231 0 -2.9824403640242300e-07
GC_10_232 b_10 NI_10 NS_232 0 1.3038484784149684e-06
GC_10_233 b_10 NI_10 NS_233 0 1.3780609789381852e-06
GC_10_234 b_10 NI_10 NS_234 0 1.3766269098435844e-06
GC_10_235 b_10 NI_10 NS_235 0 2.3900049070998119e-06
GC_10_236 b_10 NI_10 NS_236 0 -3.3970808950463025e-06
GC_10_237 b_10 NI_10 NS_237 0 -2.0889460886765649e-06
GC_10_238 b_10 NI_10 NS_238 0 -6.3013853352959738e-06
GC_10_239 b_10 NI_10 NS_239 0 -1.0350518090256880e-07
GC_10_240 b_10 NI_10 NS_240 0 5.0098788942861864e-07
GC_10_241 b_10 NI_10 NS_241 0 -1.2570134044292774e-05
GC_10_242 b_10 NI_10 NS_242 0 3.3150828196484912e-06
GC_10_243 b_10 NI_10 NS_243 0 -1.5284618345830464e-07
GC_10_244 b_10 NI_10 NS_244 0 -6.4577807174638044e-07
GC_10_245 b_10 NI_10 NS_245 0 3.1485764027509264e-06
GC_10_246 b_10 NI_10 NS_246 0 1.5222934856195736e-05
GC_10_247 b_10 NI_10 NS_247 0 1.0404517162987888e-06
GC_10_248 b_10 NI_10 NS_248 0 -1.0566921706036249e-06
GC_10_249 b_10 NI_10 NS_249 0 1.1263352593330820e-06
GC_10_250 b_10 NI_10 NS_250 0 -3.1753828186526807e-07
GC_10_251 b_10 NI_10 NS_251 0 6.6877885662652865e-06
GC_10_252 b_10 NI_10 NS_252 0 -3.1068831068007271e-06
GC_10_253 b_10 NI_10 NS_253 0 3.3131394989124637e-07
GC_10_254 b_10 NI_10 NS_254 0 3.9399052531726174e-07
GC_10_255 b_10 NI_10 NS_255 0 -2.9448234408004386e-06
GC_10_256 b_10 NI_10 NS_256 0 8.3452676817408689e-07
GC_10_257 b_10 NI_10 NS_257 0 1.7440957487127260e-07
GC_10_258 b_10 NI_10 NS_258 0 -8.8189554307727281e-07
GC_10_259 b_10 NI_10 NS_259 0 6.7930818267240482e-06
GC_10_260 b_10 NI_10 NS_260 0 3.5421113432710583e-06
GC_10_261 b_10 NI_10 NS_261 0 3.3692415667420224e-07
GC_10_262 b_10 NI_10 NS_262 0 8.5653881910932970e-09
GC_10_263 b_10 NI_10 NS_263 0 2.4534233342955936e-07
GC_10_264 b_10 NI_10 NS_264 0 -6.0596655946302403e-07
GC_10_265 b_10 NI_10 NS_265 0 3.9992767100009707e-07
GC_10_266 b_10 NI_10 NS_266 0 -1.3944037017423760e-06
GC_10_267 b_10 NI_10 NS_267 0 6.0125195412989688e-06
GC_10_268 b_10 NI_10 NS_268 0 -2.3492484787712385e-06
GC_10_269 b_10 NI_10 NS_269 0 2.3933334004750826e-08
GC_10_270 b_10 NI_10 NS_270 0 -2.5641284093242423e-07
GC_10_271 b_10 NI_10 NS_271 0 -9.3874302861935655e-07
GC_10_272 b_10 NI_10 NS_272 0 -1.1595572122175209e-06
GC_10_273 b_10 NI_10 NS_273 0 3.0875209505423561e-07
GC_10_274 b_10 NI_10 NS_274 0 -1.3340650849100446e-06
GC_10_275 b_10 NI_10 NS_275 0 3.0267272818930983e-06
GC_10_276 b_10 NI_10 NS_276 0 -4.1471411109643444e-06
GC_10_277 b_10 NI_10 NS_277 0 -1.7529087202029956e-07
GC_10_278 b_10 NI_10 NS_278 0 -3.4421370556055743e-07
GC_10_279 b_10 NI_10 NS_279 0 -1.9740574017742036e-06
GC_10_280 b_10 NI_10 NS_280 0 -6.6802220718808026e-07
GC_10_281 b_10 NI_10 NS_281 0 2.0794851779546463e-07
GC_10_282 b_10 NI_10 NS_282 0 -1.4268871932576599e-06
GC_10_283 b_10 NI_10 NS_283 0 9.1799280787580999e-08
GC_10_284 b_10 NI_10 NS_284 0 -3.5652594358236103e-06
GC_10_285 b_10 NI_10 NS_285 0 -4.5658007187586009e-07
GC_10_286 b_10 NI_10 NS_286 0 -3.7774953588670830e-07
GC_10_287 b_10 NI_10 NS_287 0 -2.1515200859010554e-06
GC_10_288 b_10 NI_10 NS_288 0 5.3520821159976911e-07
GC_10_289 b_10 NI_10 NS_289 0 -6.9311927034650297e-08
GC_10_290 b_10 NI_10 NS_290 0 -1.6158303001597354e-06
GC_10_291 b_10 NI_10 NS_291 0 -1.2654301419610086e-06
GC_10_292 b_10 NI_10 NS_292 0 -1.4064598264882507e-06
GC_10_293 b_10 NI_10 NS_293 0 -8.0808678323128601e-07
GC_10_294 b_10 NI_10 NS_294 0 9.5515364185191276e-08
GC_10_295 b_10 NI_10 NS_295 0 -9.4819678469836846e-07
GC_10_296 b_10 NI_10 NS_296 0 1.0893409298813272e-06
GC_10_297 b_10 NI_10 NS_297 0 -1.7801084933251503e-11
GC_10_298 b_10 NI_10 NS_298 0 1.0630881941786959e-11
GC_10_299 b_10 NI_10 NS_299 0 -5.7491593033083039e-07
GC_10_300 b_10 NI_10 NS_300 0 -1.1642144528816073e-06
GC_10_301 b_10 NI_10 NS_301 0 -3.7984360502503945e-07
GC_10_302 b_10 NI_10 NS_302 0 2.2312045096140264e-07
GC_10_303 b_10 NI_10 NS_303 0 -5.0935911900977284e-07
GC_10_304 b_10 NI_10 NS_304 0 3.9895588553582338e-07
GC_10_305 b_10 NI_10 NS_305 0 -1.9090380692939389e-07
GC_10_306 b_10 NI_10 NS_306 0 -1.0234021995173510e-06
GC_10_307 b_10 NI_10 NS_307 0 -4.4623632876906560e-07
GC_10_308 b_10 NI_10 NS_308 0 -2.0242009810913807e-07
GC_10_309 b_10 NI_10 NS_309 0 -9.1682601589671989e-10
GC_10_310 b_10 NI_10 NS_310 0 1.5482536263965887e-10
GC_10_311 b_10 NI_10 NS_311 0 -2.2810807387781322e-07
GC_10_312 b_10 NI_10 NS_312 0 -1.9852561689200079e-07
GC_10_313 b_10 NI_10 NS_313 0 -1.7941654170894384e-07
GC_10_314 b_10 NI_10 NS_314 0 -3.4649156197352538e-07
GC_10_315 b_10 NI_10 NS_315 0 -3.9554559669743568e-07
GC_10_316 b_10 NI_10 NS_316 0 -1.3729807141218006e-07
GC_10_317 b_10 NI_10 NS_317 0 -9.9086725840121255e-07
GC_10_318 b_10 NI_10 NS_318 0 5.0093181013171943e-08
GC_10_319 b_10 NI_10 NS_319 0 -5.8386536116222042e-07
GC_10_320 b_10 NI_10 NS_320 0 4.7577279814751663e-07
GC_10_321 b_10 NI_10 NS_321 0 -1.3073757578218945e-08
GC_10_322 b_10 NI_10 NS_322 0 4.1221575381817186e-07
GC_10_323 b_10 NI_10 NS_323 0 -8.6500719903064591e-07
GC_10_324 b_10 NI_10 NS_324 0 -9.7526660286567506e-07
GC_10_325 b_10 NI_10 NS_325 0 3.7776220288571054e-05
GC_10_326 b_10 NI_10 NS_326 0 1.2388381391945491e-12
GC_10_327 b_10 NI_10 NS_327 0 -8.1190515026193420e-12
GC_10_328 b_10 NI_10 NS_328 0 3.0025196696692842e-09
GC_10_329 b_10 NI_10 NS_329 0 3.6863546891018801e-07
GC_10_330 b_10 NI_10 NS_330 0 9.8381714634245627e-08
GC_10_331 b_10 NI_10 NS_331 0 6.5833302869581074e-07
GC_10_332 b_10 NI_10 NS_332 0 3.5826078665336387e-07
GC_10_333 b_10 NI_10 NS_333 0 1.2346307675952701e-06
GC_10_334 b_10 NI_10 NS_334 0 -8.6742347459837909e-07
GC_10_335 b_10 NI_10 NS_335 0 7.8269091312090369e-07
GC_10_336 b_10 NI_10 NS_336 0 -5.3019534862595744e-07
GC_10_337 b_10 NI_10 NS_337 0 8.2387679916956559e-07
GC_10_338 b_10 NI_10 NS_338 0 -2.1815865999775592e-06
GC_10_339 b_10 NI_10 NS_339 0 6.7226779323324467e-07
GC_10_340 b_10 NI_10 NS_340 0 -8.4320819074894875e-07
GC_10_341 b_10 NI_10 NS_341 0 -1.1291288530828683e-06
GC_10_342 b_10 NI_10 NS_342 0 -1.5078759248046793e-06
GC_10_343 b_10 NI_10 NS_343 0 -4.8952429874035813e-07
GC_10_344 b_10 NI_10 NS_344 0 -2.1009697356980355e-06
GC_10_345 b_10 NI_10 NS_345 0 -1.7840493133516331e-06
GC_10_346 b_10 NI_10 NS_346 0 -6.5665271082569585e-07
GC_10_347 b_10 NI_10 NS_347 0 -5.8884957757418207e-07
GC_10_348 b_10 NI_10 NS_348 0 -1.1663417961726428e-06
GC_10_349 b_10 NI_10 NS_349 0 -2.5817961508666801e-06
GC_10_350 b_10 NI_10 NS_350 0 -7.0824160467612382e-07
GC_10_351 b_10 NI_10 NS_351 0 -7.1488744477433752e-07
GC_10_352 b_10 NI_10 NS_352 0 -6.2488995502938180e-07
GC_10_353 b_10 NI_10 NS_353 0 -3.5724825518431680e-06
GC_10_354 b_10 NI_10 NS_354 0 -4.6955674528674794e-07
GC_10_355 b_10 NI_10 NS_355 0 2.3206436357994382e-07
GC_10_356 b_10 NI_10 NS_356 0 -2.1172247072664742e-07
GC_10_357 b_10 NI_10 NS_357 0 -9.1741053745162611e-07
GC_10_358 b_10 NI_10 NS_358 0 -9.0467130342698208e-07
GC_10_359 b_10 NI_10 NS_359 0 -1.9019401387906308e-06
GC_10_360 b_10 NI_10 NS_360 0 1.9080907685598609e-07
GC_10_361 b_10 NI_10 NS_361 0 -1.1727179916730466e-06
GC_10_362 b_10 NI_10 NS_362 0 -4.8227499348525284e-07
GC_10_363 b_10 NI_10 NS_363 0 -1.3189678772717401e-06
GC_10_364 b_10 NI_10 NS_364 0 9.6812045173159703e-07
GC_10_365 b_10 NI_10 NS_365 0 -7.9967172811173072e-07
GC_10_366 b_10 NI_10 NS_366 0 -4.7982924578834642e-07
GC_10_367 b_10 NI_10 NS_367 0 -3.1176524076938382e-06
GC_10_368 b_10 NI_10 NS_368 0 3.9717227154412511e-07
GC_10_369 b_10 NI_10 NS_369 0 -6.0260883747479366e-07
GC_10_370 b_10 NI_10 NS_370 0 1.6123364825767504e-07
GC_10_371 b_10 NI_10 NS_371 0 -6.6727476242582864e-07
GC_10_372 b_10 NI_10 NS_372 0 -1.5680981752757446e-07
GC_10_373 b_10 NI_10 NS_373 0 -1.3447837412931022e-06
GC_10_374 b_10 NI_10 NS_374 0 -7.5287492266704022e-08
GC_10_375 b_10 NI_10 NS_375 0 -3.0786962646614466e-06
GC_10_376 b_10 NI_10 NS_376 0 2.3443902796002714e-06
GC_10_377 b_10 NI_10 NS_377 0 -7.5437663486093877e-07
GC_10_378 b_10 NI_10 NS_378 0 3.5807594785992426e-07
GC_10_379 b_10 NI_10 NS_379 0 -7.9998421411423021e-07
GC_10_380 b_10 NI_10 NS_380 0 1.0728520704217732e-06
GC_10_381 b_10 NI_10 NS_381 0 -1.2382060995612915e-06
GC_10_382 b_10 NI_10 NS_382 0 1.6928405711473574e-07
GC_10_383 b_10 NI_10 NS_383 0 -1.0794847885291676e-06
GC_10_384 b_10 NI_10 NS_384 0 3.5772850913182289e-06
GC_10_385 b_10 NI_10 NS_385 0 -6.8449390394910728e-07
GC_10_386 b_10 NI_10 NS_386 0 4.6095705576317645e-07
GC_10_387 b_10 NI_10 NS_387 0 1.7789017254130538e-07
GC_10_388 b_10 NI_10 NS_388 0 1.4971618211381142e-06
GC_10_389 b_10 NI_10 NS_389 0 -1.1956477428327266e-06
GC_10_390 b_10 NI_10 NS_390 0 3.1705872454518263e-07
GC_10_391 b_10 NI_10 NS_391 0 9.5835695191399473e-07
GC_10_392 b_10 NI_10 NS_392 0 3.0172741976837468e-06
GC_10_393 b_10 NI_10 NS_393 0 -5.5639036577292685e-07
GC_10_394 b_10 NI_10 NS_394 0 6.1270799907344599e-07
GC_10_395 b_10 NI_10 NS_395 0 1.0073478009264724e-06
GC_10_396 b_10 NI_10 NS_396 0 8.4907995384515472e-07
GC_10_397 b_10 NI_10 NS_397 0 -1.1354557625817660e-06
GC_10_398 b_10 NI_10 NS_398 0 5.7364219270568629e-07
GC_10_399 b_10 NI_10 NS_399 0 1.7677940966898031e-06
GC_10_400 b_10 NI_10 NS_400 0 1.3974058717223382e-06
GC_10_401 b_10 NI_10 NS_401 0 -1.4090126802628557e-07
GC_10_402 b_10 NI_10 NS_402 0 6.5188738321420302e-07
GC_10_403 b_10 NI_10 NS_403 0 6.9857278681583115e-07
GC_10_404 b_10 NI_10 NS_404 0 -1.8049620643413311e-08
GC_10_405 b_10 NI_10 NS_405 0 2.1846618922526439e-11
GC_10_406 b_10 NI_10 NS_406 0 1.4146775444213368e-11
GC_10_407 b_10 NI_10 NS_407 0 -5.3444744493007062e-07
GC_10_408 b_10 NI_10 NS_408 0 6.6480197274624728e-07
GC_10_409 b_10 NI_10 NS_409 0 -1.6743644148556701e-08
GC_10_410 b_10 NI_10 NS_410 0 3.0212225897502640e-07
GC_10_411 b_10 NI_10 NS_411 0 2.1121851933243082e-07
GC_10_412 b_10 NI_10 NS_412 0 1.5832440911237055e-07
GC_10_413 b_10 NI_10 NS_413 0 -1.8419242889331875e-07
GC_10_414 b_10 NI_10 NS_414 0 5.6372780530729515e-07
GC_10_415 b_10 NI_10 NS_415 0 8.6157926743891893e-07
GC_10_416 b_10 NI_10 NS_416 0 4.0476703737225424e-07
GC_10_417 b_10 NI_10 NS_417 0 7.9125327667396772e-10
GC_10_418 b_10 NI_10 NS_418 0 5.1026214141207431e-10
GC_10_419 b_10 NI_10 NS_419 0 1.2590913603713589e-06
GC_10_420 b_10 NI_10 NS_420 0 1.3277194062368242e-07
GC_10_421 b_10 NI_10 NS_421 0 -1.4104094816982340e-07
GC_10_422 b_10 NI_10 NS_422 0 8.3427619881604144e-07
GC_10_423 b_10 NI_10 NS_423 0 8.2109864346122023e-08
GC_10_424 b_10 NI_10 NS_424 0 4.1437008052444817e-08
GC_10_425 b_10 NI_10 NS_425 0 3.4449283246839274e-07
GC_10_426 b_10 NI_10 NS_426 0 3.3673142443173587e-07
GC_10_427 b_10 NI_10 NS_427 0 3.0905483530998112e-07
GC_10_428 b_10 NI_10 NS_428 0 4.0929891905796637e-07
GC_10_429 b_10 NI_10 NS_429 0 6.5355083477062854e-08
GC_10_430 b_10 NI_10 NS_430 0 5.9257338447030123e-08
GC_10_431 b_10 NI_10 NS_431 0 7.1106666759108083e-07
GC_10_432 b_10 NI_10 NS_432 0 8.9929616146302544e-07
GC_10_433 b_10 NI_10 NS_433 0 -1.4324861025282032e-04
GC_10_434 b_10 NI_10 NS_434 0 3.4599429970999890e-11
GC_10_435 b_10 NI_10 NS_435 0 3.0174888969782112e-11
GC_10_436 b_10 NI_10 NS_436 0 9.4201772421956121e-10
GC_10_437 b_10 NI_10 NS_437 0 -2.1091459556580796e-06
GC_10_438 b_10 NI_10 NS_438 0 -1.6534093682869667e-06
GC_10_439 b_10 NI_10 NS_439 0 1.8892050314652076e-06
GC_10_440 b_10 NI_10 NS_440 0 3.8449862697588235e-06
GC_10_441 b_10 NI_10 NS_441 0 3.2880590142055589e-06
GC_10_442 b_10 NI_10 NS_442 0 4.9269648232951067e-06
GC_10_443 b_10 NI_10 NS_443 0 5.8303024830013329e-06
GC_10_444 b_10 NI_10 NS_444 0 -9.0830949276066732e-06
GC_10_445 b_10 NI_10 NS_445 0 -2.5402010752916004e-06
GC_10_446 b_10 NI_10 NS_446 0 -1.3835967334667506e-05
GC_10_447 b_10 NI_10 NS_447 0 -3.5342725890626069e-06
GC_10_448 b_10 NI_10 NS_448 0 2.1966305697923715e-06
GC_10_449 b_10 NI_10 NS_449 0 3.6391266962433783e-06
GC_10_450 b_10 NI_10 NS_450 0 1.2970505518935621e-06
GC_10_451 b_10 NI_10 NS_451 0 7.8997684288469275e-06
GC_10_452 b_10 NI_10 NS_452 0 -3.9683339445140398e-05
GC_10_453 b_10 NI_10 NS_453 0 -4.4005795955361242e-05
GC_10_454 b_10 NI_10 NS_454 0 -8.8281784842177422e-07
GC_10_455 b_10 NI_10 NS_455 0 -1.4766052554575199e-05
GC_10_456 b_10 NI_10 NS_456 0 -8.4725927149341770e-06
GC_10_457 b_10 NI_10 NS_457 0 -7.2348592304007049e-05
GC_10_458 b_10 NI_10 NS_458 0 7.5140404776053606e-05
GC_10_459 b_10 NI_10 NS_459 0 4.6495324875952608e-06
GC_10_460 b_10 NI_10 NS_460 0 1.3009968469448146e-05
GC_10_461 b_10 NI_10 NS_461 0 6.2665099035800784e-05
GC_10_462 b_10 NI_10 NS_462 0 1.2224195416918459e-04
GC_10_463 b_10 NI_10 NS_463 0 2.4457542937450760e-07
GC_10_464 b_10 NI_10 NS_464 0 -3.6753280535911733e-05
GC_10_465 b_10 NI_10 NS_465 0 1.6411258195954708e-05
GC_10_466 b_10 NI_10 NS_466 0 3.8871954755495198e-06
GC_10_467 b_10 NI_10 NS_467 0 2.4219140037085866e-05
GC_10_468 b_10 NI_10 NS_468 0 -3.0244013755743459e-05
GC_10_469 b_10 NI_10 NS_469 0 -8.8437586386077631e-06
GC_10_470 b_10 NI_10 NS_470 0 -2.2761550027210164e-06
GC_10_471 b_10 NI_10 NS_471 0 -8.7280421249731384e-06
GC_10_472 b_10 NI_10 NS_472 0 2.5050968735191944e-05
GC_10_473 b_10 NI_10 NS_473 0 5.8325759078355851e-06
GC_10_474 b_10 NI_10 NS_474 0 8.3788302600318986e-06
GC_10_475 b_10 NI_10 NS_475 0 5.5969459801675242e-05
GC_10_476 b_10 NI_10 NS_476 0 2.4647582918710520e-05
GC_10_477 b_10 NI_10 NS_477 0 3.4492064062358255e-06
GC_10_478 b_10 NI_10 NS_478 0 -1.1606267738731554e-05
GC_10_479 b_10 NI_10 NS_479 0 -4.0620242380424786e-07
GC_10_480 b_10 NI_10 NS_480 0 -1.2991964397779393e-06
GC_10_481 b_10 NI_10 NS_481 0 6.7879704850620033e-06
GC_10_482 b_10 NI_10 NS_482 0 3.0205762289126828e-06
GC_10_483 b_10 NI_10 NS_483 0 4.1592015178744659e-05
GC_10_484 b_10 NI_10 NS_484 0 -1.7165665374976642e-05
GC_10_485 b_10 NI_10 NS_485 0 -2.5738436211535086e-06
GC_10_486 b_10 NI_10 NS_486 0 -7.0283376819833933e-06
GC_10_487 b_10 NI_10 NS_487 0 -2.9900644604569711e-06
GC_10_488 b_10 NI_10 NS_488 0 1.7603140982600878e-06
GC_10_489 b_10 NI_10 NS_489 0 9.5385432945228708e-06
GC_10_490 b_10 NI_10 NS_490 0 2.8682894334566471e-06
GC_10_491 b_10 NI_10 NS_491 0 2.2731564147989544e-05
GC_10_492 b_10 NI_10 NS_492 0 -3.1037617216230302e-05
GC_10_493 b_10 NI_10 NS_493 0 -5.6871501661912806e-06
GC_10_494 b_10 NI_10 NS_494 0 -3.6246204899398187e-06
GC_10_495 b_10 NI_10 NS_495 0 -5.2395997617335954e-07
GC_10_496 b_10 NI_10 NS_496 0 5.0176151610032377e-06
GC_10_497 b_10 NI_10 NS_497 0 1.2253681360214231e-05
GC_10_498 b_10 NI_10 NS_498 0 1.7530807766327591e-07
GC_10_499 b_10 NI_10 NS_499 0 1.8082954301829058e-06
GC_10_500 b_10 NI_10 NS_500 0 -3.1349948134845213e-05
GC_10_501 b_10 NI_10 NS_501 0 -6.7180534664305465e-06
GC_10_502 b_10 NI_10 NS_502 0 9.7548869986989034e-07
GC_10_503 b_10 NI_10 NS_503 0 4.6118094289440338e-06
GC_10_504 b_10 NI_10 NS_504 0 3.8655086263491989e-06
GC_10_505 b_10 NI_10 NS_505 0 1.4061847912579118e-05
GC_10_506 b_10 NI_10 NS_506 0 -6.0101960554777506e-06
GC_10_507 b_10 NI_10 NS_507 0 -1.4015900567442822e-05
GC_10_508 b_10 NI_10 NS_508 0 -1.8747000510165503e-05
GC_10_509 b_10 NI_10 NS_509 0 -2.5061634712958622e-06
GC_10_510 b_10 NI_10 NS_510 0 5.4162195799283912e-06
GC_10_511 b_10 NI_10 NS_511 0 4.6576523315815172e-06
GC_10_512 b_10 NI_10 NS_512 0 -2.0834692084549581e-06
GC_10_513 b_10 NI_10 NS_513 0 -1.4565941753593980e-11
GC_10_514 b_10 NI_10 NS_514 0 4.2048034221586431e-12
GC_10_515 b_10 NI_10 NS_515 0 5.1979769047532318e-06
GC_10_516 b_10 NI_10 NS_516 0 -1.1242606771714254e-05
GC_10_517 b_10 NI_10 NS_517 0 -2.6676768855521398e-07
GC_10_518 b_10 NI_10 NS_518 0 2.9264576171131015e-06
GC_10_519 b_10 NI_10 NS_519 0 2.6445018548753416e-06
GC_10_520 b_10 NI_10 NS_520 0 -1.5935934397612758e-06
GC_10_521 b_10 NI_10 NS_521 0 2.4076253787231408e-06
GC_10_522 b_10 NI_10 NS_522 0 -9.4308085524272477e-06
GC_10_523 b_10 NI_10 NS_523 0 -9.9265974818690249e-06
GC_10_524 b_10 NI_10 NS_524 0 -3.6884498915998644e-06
GC_10_525 b_10 NI_10 NS_525 0 3.1234724315884732e-10
GC_10_526 b_10 NI_10 NS_526 0 2.7697521026485995e-10
GC_10_527 b_10 NI_10 NS_527 0 -8.5916103485670579e-06
GC_10_528 b_10 NI_10 NS_528 0 -5.6865019292539686e-06
GC_10_529 b_10 NI_10 NS_529 0 2.2662364467159663e-06
GC_10_530 b_10 NI_10 NS_530 0 -6.4520167911088495e-06
GC_10_531 b_10 NI_10 NS_531 0 -3.0673944715153044e-06
GC_10_532 b_10 NI_10 NS_532 0 -1.3540710017181032e-07
GC_10_533 b_10 NI_10 NS_533 0 -7.9220167818713533e-06
GC_10_534 b_10 NI_10 NS_534 0 4.8453636854019418e-07
GC_10_535 b_10 NI_10 NS_535 0 3.0018484457339994e-06
GC_10_536 b_10 NI_10 NS_536 0 2.8730592517579312e-06
GC_10_537 b_10 NI_10 NS_537 0 1.2171965514011818e-06
GC_10_538 b_10 NI_10 NS_538 0 -3.8814953245347687e-06
GC_10_539 b_10 NI_10 NS_539 0 -4.8737996294447932e-06
GC_10_540 b_10 NI_10 NS_540 0 -3.9067810931837210e-06
GC_10_541 b_10 NI_10 NS_541 0 -3.1809059305217014e-05
GC_10_542 b_10 NI_10 NS_542 0 -1.9490474490220272e-12
GC_10_543 b_10 NI_10 NS_543 0 -2.2738568820249117e-10
GC_10_544 b_10 NI_10 NS_544 0 1.0441852117161765e-08
GC_10_545 b_10 NI_10 NS_545 0 6.8674751577302558e-07
GC_10_546 b_10 NI_10 NS_546 0 1.0912847713052050e-07
GC_10_547 b_10 NI_10 NS_547 0 3.1464725415515685e-06
GC_10_548 b_10 NI_10 NS_548 0 -1.3843757487774440e-06
GC_10_549 b_10 NI_10 NS_549 0 -2.7797116550689788e-06
GC_10_550 b_10 NI_10 NS_550 0 -2.8013711396961683e-06
GC_10_551 b_10 NI_10 NS_551 0 4.9066013164336570e-06
GC_10_552 b_10 NI_10 NS_552 0 -5.2641007260491574e-07
GC_10_553 b_10 NI_10 NS_553 0 -7.0388981145675631e-06
GC_10_554 b_10 NI_10 NS_554 0 -8.0734842770294906e-06
GC_10_555 b_10 NI_10 NS_555 0 1.9913894512022442e-08
GC_10_556 b_10 NI_10 NS_556 0 -1.5400079805498521e-06
GC_10_557 b_10 NI_10 NS_557 0 -6.0451837816403998e-06
GC_10_558 b_10 NI_10 NS_558 0 1.9318159384310007e-06
GC_10_559 b_10 NI_10 NS_559 0 5.2997093070917221e-06
GC_10_560 b_10 NI_10 NS_560 0 -5.7096591667012671e-06
GC_10_561 b_10 NI_10 NS_561 0 -1.7020825153362027e-05
GC_10_562 b_10 NI_10 NS_562 0 4.6231741982044338e-06
GC_10_563 b_10 NI_10 NS_563 0 -1.1776750505142961e-06
GC_10_564 b_10 NI_10 NS_564 0 7.0415494908454863e-06
GC_10_565 b_10 NI_10 NS_565 0 -7.1892211809480762e-06
GC_10_566 b_10 NI_10 NS_566 0 -4.5422170885806932e-06
GC_10_567 b_10 NI_10 NS_567 0 -3.3644348592024712e-06
GC_10_568 b_10 NI_10 NS_568 0 7.9554426755881966e-06
GC_10_569 b_10 NI_10 NS_569 0 -2.2172645287555157e-06
GC_10_570 b_10 NI_10 NS_570 0 -4.6363868500174537e-06
GC_10_571 b_10 NI_10 NS_571 0 -3.8558756938154314e-06
GC_10_572 b_10 NI_10 NS_572 0 1.1253137040755168e-05
GC_10_573 b_10 NI_10 NS_573 0 -1.8103187258957947e-07
GC_10_574 b_10 NI_10 NS_574 0 7.1456890390772864e-06
GC_10_575 b_10 NI_10 NS_575 0 -4.1163604896343898e-06
GC_10_576 b_10 NI_10 NS_576 0 1.2239893681119820e-06
GC_10_577 b_10 NI_10 NS_577 0 -6.2986810241564363e-07
GC_10_578 b_10 NI_10 NS_578 0 7.9394007743742448e-06
GC_10_579 b_10 NI_10 NS_579 0 -1.0416948870203981e-06
GC_10_580 b_10 NI_10 NS_580 0 2.1882199758278305e-06
GC_10_581 b_10 NI_10 NS_581 0 -2.4107594689369288e-06
GC_10_582 b_10 NI_10 NS_582 0 8.0524125220147169e-06
GC_10_583 b_10 NI_10 NS_583 0 -1.5236741075705701e-07
GC_10_584 b_10 NI_10 NS_584 0 9.4057521429355657e-06
GC_10_585 b_10 NI_10 NS_585 0 -8.6008091589355045e-07
GC_10_586 b_10 NI_10 NS_586 0 8.6777426423436119e-06
GC_10_587 b_10 NI_10 NS_587 0 -1.3290770475566425e-06
GC_10_588 b_10 NI_10 NS_588 0 3.8594417535181758e-06
GC_10_589 b_10 NI_10 NS_589 0 9.6762987328082351e-07
GC_10_590 b_10 NI_10 NS_590 0 1.1812355727470389e-05
GC_10_591 b_10 NI_10 NS_591 0 1.7367412035362374e-05
GC_10_592 b_10 NI_10 NS_592 0 1.6606440226795979e-05
GC_10_593 b_10 NI_10 NS_593 0 4.7005655512145674e-06
GC_10_594 b_10 NI_10 NS_594 0 7.6012305507460194e-06
GC_10_595 b_10 NI_10 NS_595 0 9.8175728001247055e-06
GC_10_596 b_10 NI_10 NS_596 0 3.8200676069308745e-06
GC_10_597 b_10 NI_10 NS_597 0 6.4427117978240272e-06
GC_10_598 b_10 NI_10 NS_598 0 1.0581087037468506e-05
GC_10_599 b_10 NI_10 NS_599 0 3.1909374859771068e-05
GC_10_600 b_10 NI_10 NS_600 0 -5.8429960836848804e-06
GC_10_601 b_10 NI_10 NS_601 0 7.7884074519920703e-06
GC_10_602 b_10 NI_10 NS_602 0 3.3158522216387464e-06
GC_10_603 b_10 NI_10 NS_603 0 1.1397117433050147e-05
GC_10_604 b_10 NI_10 NS_604 0 -9.9644756070637809e-06
GC_10_605 b_10 NI_10 NS_605 0 1.0344054312339736e-05
GC_10_606 b_10 NI_10 NS_606 0 6.2012170356266368e-06
GC_10_607 b_10 NI_10 NS_607 0 1.5863182284504304e-05
GC_10_608 b_10 NI_10 NS_608 0 -2.9905472199473169e-05
GC_10_609 b_10 NI_10 NS_609 0 7.7033687547793302e-06
GC_10_610 b_10 NI_10 NS_610 0 -2.9069263356953416e-06
GC_10_611 b_10 NI_10 NS_611 0 -3.4527977877439299e-06
GC_10_612 b_10 NI_10 NS_612 0 -1.5725352436016351e-05
GC_10_613 b_10 NI_10 NS_613 0 1.1298999549599578e-05
GC_10_614 b_10 NI_10 NS_614 0 -1.7523095027189883e-06
GC_10_615 b_10 NI_10 NS_615 0 -1.3023507330545018e-05
GC_10_616 b_10 NI_10 NS_616 0 -2.4164324100995707e-05
GC_10_617 b_10 NI_10 NS_617 0 -4.2518743728947021e-07
GC_10_618 b_10 NI_10 NS_618 0 -6.4081584911353400e-06
GC_10_619 b_10 NI_10 NS_619 0 -9.5225951954455687e-06
GC_10_620 b_10 NI_10 NS_620 0 -2.3446773851749633e-06
GC_10_621 b_10 NI_10 NS_621 0 9.7513649365775545e-11
GC_10_622 b_10 NI_10 NS_622 0 5.3586370485095460e-11
GC_10_623 b_10 NI_10 NS_623 0 1.1849083321267018e-06
GC_10_624 b_10 NI_10 NS_624 0 -4.6339014347782502e-06
GC_10_625 b_10 NI_10 NS_625 0 -1.4863760834301179e-06
GC_10_626 b_10 NI_10 NS_626 0 -1.2907053856757696e-06
GC_10_627 b_10 NI_10 NS_627 0 -4.9349922383034489e-06
GC_10_628 b_10 NI_10 NS_628 0 -8.8189376248682531e-07
GC_10_629 b_10 NI_10 NS_629 0 -1.3866100145644722e-06
GC_10_630 b_10 NI_10 NS_630 0 -2.8415046695241759e-06
GC_10_631 b_10 NI_10 NS_631 0 -1.0079602400428095e-05
GC_10_632 b_10 NI_10 NS_632 0 -3.7053046144993288e-06
GC_10_633 b_10 NI_10 NS_633 0 6.6047306059905226e-09
GC_10_634 b_10 NI_10 NS_634 0 5.7466231183883366e-09
GC_10_635 b_10 NI_10 NS_635 0 1.3885989502789948e-06
GC_10_636 b_10 NI_10 NS_636 0 6.7923793261236252e-07
GC_10_637 b_10 NI_10 NS_637 0 -1.7365100311679089e-06
GC_10_638 b_10 NI_10 NS_638 0 3.1379192391406338e-06
GC_10_639 b_10 NI_10 NS_639 0 -9.2489876556871306e-07
GC_10_640 b_10 NI_10 NS_640 0 7.7500973470929590e-07
GC_10_641 b_10 NI_10 NS_641 0 -7.9023120372615401e-06
GC_10_642 b_10 NI_10 NS_642 0 8.1042209666848402e-07
GC_10_643 b_10 NI_10 NS_643 0 -2.4148796965930569e-06
GC_10_644 b_10 NI_10 NS_644 0 2.0815635738673444e-06
GC_10_645 b_10 NI_10 NS_645 0 -2.1260357816936824e-06
GC_10_646 b_10 NI_10 NS_646 0 2.1321343939036211e-06
GC_10_647 b_10 NI_10 NS_647 0 1.1301419684912100e-06
GC_10_648 b_10 NI_10 NS_648 0 2.8148322384276432e-06
GC_10_649 b_10 NI_10 NS_649 0 -6.3819075348518371e-04
GC_10_650 b_10 NI_10 NS_650 0 -9.7138989804644198e-11
GC_10_651 b_10 NI_10 NS_651 0 3.8809213020749568e-09
GC_10_652 b_10 NI_10 NS_652 0 -6.7423153233845858e-08
GC_10_653 b_10 NI_10 NS_653 0 -1.1292057263862952e-05
GC_10_654 b_10 NI_10 NS_654 0 -9.3317597843433109e-06
GC_10_655 b_10 NI_10 NS_655 0 -2.2441912347374106e-06
GC_10_656 b_10 NI_10 NS_656 0 2.2642845401922535e-07
GC_10_657 b_10 NI_10 NS_657 0 -3.0298275459908922e-05
GC_10_658 b_10 NI_10 NS_658 0 2.7085505761474644e-05
GC_10_659 b_10 NI_10 NS_659 0 -3.3245391103317109e-05
GC_10_660 b_10 NI_10 NS_660 0 8.1393442525026905e-06
GC_10_661 b_10 NI_10 NS_661 0 3.1754280894125608e-05
GC_10_662 b_10 NI_10 NS_662 0 2.7340902019778223e-05
GC_10_663 b_10 NI_10 NS_663 0 -9.0548942961053751e-06
GC_10_664 b_10 NI_10 NS_664 0 1.4743928034458728e-05
GC_10_665 b_10 NI_10 NS_665 0 1.2670966010821840e-05
GC_10_666 b_10 NI_10 NS_666 0 3.6937564506495431e-05
GC_10_667 b_10 NI_10 NS_667 0 -1.0602068792454595e-05
GC_10_668 b_10 NI_10 NS_668 0 6.8138225566499619e-05
GC_10_669 b_10 NI_10 NS_669 0 9.5404370048703536e-05
GC_10_670 b_10 NI_10 NS_670 0 -6.6240443610732339e-05
GC_10_671 b_10 NI_10 NS_671 0 2.7099114329721589e-05
GC_10_672 b_10 NI_10 NS_672 0 3.1676108772077702e-05
GC_10_673 b_10 NI_10 NS_673 0 -7.4559479509472426e-06
GC_10_674 b_10 NI_10 NS_674 0 -7.2595413655826923e-05
GC_10_675 b_10 NI_10 NS_675 0 -9.8760715363145121e-06
GC_10_676 b_10 NI_10 NS_676 0 -3.3982284762719834e-05
GC_10_677 b_10 NI_10 NS_677 0 -7.7016034283787556e-05
GC_10_678 b_10 NI_10 NS_678 0 1.9174785957544022e-05
GC_10_679 b_10 NI_10 NS_679 0 2.4970785313462398e-05
GC_10_680 b_10 NI_10 NS_680 0 5.0900353670911029e-05
GC_10_681 b_10 NI_10 NS_681 0 -2.3151132545363912e-05
GC_10_682 b_10 NI_10 NS_682 0 -3.5305291180768160e-06
GC_10_683 b_10 NI_10 NS_683 0 6.9874061901191166e-05
GC_10_684 b_10 NI_10 NS_684 0 4.4645049537920434e-05
GC_10_685 b_10 NI_10 NS_685 0 2.9213302282090411e-05
GC_10_686 b_10 NI_10 NS_686 0 1.9680259923162727e-05
GC_10_687 b_10 NI_10 NS_687 0 -7.3500006149360051e-06
GC_10_688 b_10 NI_10 NS_688 0 -2.5717472693599477e-05
GC_10_689 b_10 NI_10 NS_689 0 -7.6009688242860110e-06
GC_10_690 b_10 NI_10 NS_690 0 -2.5156201215140217e-05
GC_10_691 b_10 NI_10 NS_691 0 6.7666484894973792e-06
GC_10_692 b_10 NI_10 NS_692 0 4.9266801949898238e-05
GC_10_693 b_10 NI_10 NS_693 0 1.2941341998740592e-05
GC_10_694 b_10 NI_10 NS_694 0 2.7354623773780945e-05
GC_10_695 b_10 NI_10 NS_695 0 5.8648218328080022e-06
GC_10_696 b_10 NI_10 NS_696 0 2.1243290417799161e-06
GC_10_697 b_10 NI_10 NS_697 0 -6.3929902258455820e-07
GC_10_698 b_10 NI_10 NS_698 0 -1.5371371862528264e-05
GC_10_699 b_10 NI_10 NS_699 0 5.6176831116005674e-05
GC_10_700 b_10 NI_10 NS_700 0 3.8178374829275704e-05
GC_10_701 b_10 NI_10 NS_701 0 1.9951205817163743e-05
GC_10_702 b_10 NI_10 NS_702 0 1.4801261902046074e-05
GC_10_703 b_10 NI_10 NS_703 0 8.3758764118362653e-06
GC_10_704 b_10 NI_10 NS_704 0 -1.2841463339293246e-05
GC_10_705 b_10 NI_10 NS_705 0 -5.6601888607229929e-06
GC_10_706 b_10 NI_10 NS_706 0 -1.3971550281960084e-05
GC_10_707 b_10 NI_10 NS_707 0 6.6117341609201339e-05
GC_10_708 b_10 NI_10 NS_708 0 1.3011952468918226e-05
GC_10_709 b_10 NI_10 NS_709 0 2.2771813794868498e-05
GC_10_710 b_10 NI_10 NS_710 0 4.9238765321780340e-06
GC_10_711 b_10 NI_10 NS_711 0 -5.5579099041640297e-06
GC_10_712 b_10 NI_10 NS_712 0 -2.1967476154490458e-05
GC_10_713 b_10 NI_10 NS_713 0 -9.1458067398642935e-06
GC_10_714 b_10 NI_10 NS_714 0 -7.0555601935873620e-06
GC_10_715 b_10 NI_10 NS_715 0 6.0678797961071843e-05
GC_10_716 b_10 NI_10 NS_716 0 -9.4911920514481574e-06
GC_10_717 b_10 NI_10 NS_717 0 2.1422964198437373e-05
GC_10_718 b_10 NI_10 NS_718 0 -7.3860835424353691e-06
GC_10_719 b_10 NI_10 NS_719 0 -2.3066431539390616e-05
GC_10_720 b_10 NI_10 NS_720 0 -1.3101705800712700e-05
GC_10_721 b_10 NI_10 NS_721 0 -8.6613366296168401e-06
GC_10_722 b_10 NI_10 NS_722 0 4.4701005309192796e-06
GC_10_723 b_10 NI_10 NS_723 0 4.5474475054313533e-05
GC_10_724 b_10 NI_10 NS_724 0 -2.5680606140023232e-05
GC_10_725 b_10 NI_10 NS_725 0 6.0238032383227525e-06
GC_10_726 b_10 NI_10 NS_726 0 -1.6485890145525831e-05
GC_10_727 b_10 NI_10 NS_727 0 -1.8717561847273327e-05
GC_10_728 b_10 NI_10 NS_728 0 8.6339108299133775e-06
GC_10_729 b_10 NI_10 NS_729 0 -4.6974532798100974e-11
GC_10_730 b_10 NI_10 NS_730 0 -1.7787557025782317e-10
GC_10_731 b_10 NI_10 NS_731 0 1.7546174895183273e-06
GC_10_732 b_10 NI_10 NS_732 0 8.7733268922510683e-06
GC_10_733 b_10 NI_10 NS_733 0 2.2050753387209847e-06
GC_10_734 b_10 NI_10 NS_734 0 -7.0025610832562191e-06
GC_10_735 b_10 NI_10 NS_735 0 -9.0168649745741640e-06
GC_10_736 b_10 NI_10 NS_736 0 5.7743082187514469e-06
GC_10_737 b_10 NI_10 NS_737 0 4.7670771916913970e-06
GC_10_738 b_10 NI_10 NS_738 0 1.1522884158036962e-05
GC_10_739 b_10 NI_10 NS_739 0 2.4563941346424643e-05
GC_10_740 b_10 NI_10 NS_740 0 -2.1161940120509821e-05
GC_10_741 b_10 NI_10 NS_741 0 -5.7418291353622801e-09
GC_10_742 b_10 NI_10 NS_742 0 -5.6212436215613893e-09
GC_10_743 b_10 NI_10 NS_743 0 3.0635563018055335e-05
GC_10_744 b_10 NI_10 NS_744 0 7.5174978425780822e-06
GC_10_745 b_10 NI_10 NS_745 0 -2.6868608061414452e-06
GC_10_746 b_10 NI_10 NS_746 0 1.1037124025663339e-05
GC_10_747 b_10 NI_10 NS_747 0 8.0388613665932933e-06
GC_10_748 b_10 NI_10 NS_748 0 1.1978095465852395e-06
GC_10_749 b_10 NI_10 NS_749 0 1.9083149471787286e-05
GC_10_750 b_10 NI_10 NS_750 0 -2.1548990614303349e-05
GC_10_751 b_10 NI_10 NS_751 0 -6.5779333799964184e-06
GC_10_752 b_10 NI_10 NS_752 0 -7.4324925366168556e-06
GC_10_753 b_10 NI_10 NS_753 0 -5.4018427610227658e-06
GC_10_754 b_10 NI_10 NS_754 0 1.2517272787458623e-05
GC_10_755 b_10 NI_10 NS_755 0 1.6097896779396038e-05
GC_10_756 b_10 NI_10 NS_756 0 7.3673312014929661e-06
GC_10_757 b_10 NI_10 NS_757 0 5.6902099855732724e-05
GC_10_758 b_10 NI_10 NS_758 0 -1.2101498766994265e-10
GC_10_759 b_10 NI_10 NS_759 0 -2.0303367219419840e-09
GC_10_760 b_10 NI_10 NS_760 0 3.4201184995939939e-08
GC_10_761 b_10 NI_10 NS_761 0 -5.1436485214084864e-07
GC_10_762 b_10 NI_10 NS_762 0 -3.8156302401383707e-07
GC_10_763 b_10 NI_10 NS_763 0 -8.7410285883448629e-07
GC_10_764 b_10 NI_10 NS_764 0 9.5756912232101723e-06
GC_10_765 b_10 NI_10 NS_765 0 1.2647595220759946e-05
GC_10_766 b_10 NI_10 NS_766 0 -1.2046157061810514e-05
GC_10_767 b_10 NI_10 NS_767 0 -1.7539276613558484e-05
GC_10_768 b_10 NI_10 NS_768 0 8.8319930232214526e-06
GC_10_769 b_10 NI_10 NS_769 0 2.8401356213346886e-05
GC_10_770 b_10 NI_10 NS_770 0 -6.5602084527167915e-06
GC_10_771 b_10 NI_10 NS_771 0 -3.2049430771493157e-06
GC_10_772 b_10 NI_10 NS_772 0 -3.0960969545231509e-06
GC_10_773 b_10 NI_10 NS_773 0 -2.8498748128382108e-06
GC_10_774 b_10 NI_10 NS_774 0 -1.4497135655540664e-05
GC_10_775 b_10 NI_10 NS_775 0 -2.4758797407387007e-05
GC_10_776 b_10 NI_10 NS_776 0 4.0215888297837489e-05
GC_10_777 b_10 NI_10 NS_777 0 3.7734250856548128e-05
GC_10_778 b_10 NI_10 NS_778 0 -4.7032653301687406e-05
GC_10_779 b_10 NI_10 NS_779 0 -3.0428739525600077e-05
GC_10_780 b_10 NI_10 NS_780 0 -2.0941082872033737e-05
GC_10_781 b_10 NI_10 NS_781 0 3.3065696919686832e-05
GC_10_782 b_10 NI_10 NS_782 0 2.6831766541901966e-05
GC_10_783 b_10 NI_10 NS_783 0 -1.8367588206145855e-05
GC_10_784 b_10 NI_10 NS_784 0 -2.8795047602126811e-05
GC_10_785 b_10 NI_10 NS_785 0 2.1463775174355082e-05
GC_10_786 b_10 NI_10 NS_786 0 6.0257593486086972e-05
GC_10_787 b_10 NI_10 NS_787 0 -2.1175884728206162e-05
GC_10_788 b_10 NI_10 NS_788 0 -5.5544466812222329e-05
GC_10_789 b_10 NI_10 NS_789 0 -3.1395988182654391e-05
GC_10_790 b_10 NI_10 NS_790 0 -1.1645823525445775e-05
GC_10_791 b_10 NI_10 NS_791 0 2.0313078232214476e-05
GC_10_792 b_10 NI_10 NS_792 0 1.3868917454410403e-05
GC_10_793 b_10 NI_10 NS_793 0 -2.4579282162969858e-05
GC_10_794 b_10 NI_10 NS_794 0 -1.0925905923322242e-05
GC_10_795 b_10 NI_10 NS_795 0 2.0765200347204598e-05
GC_10_796 b_10 NI_10 NS_796 0 1.0076894553900300e-05
GC_10_797 b_10 NI_10 NS_797 0 -1.8224310162295529e-05
GC_10_798 b_10 NI_10 NS_798 0 -2.0845754851241956e-05
GC_10_799 b_10 NI_10 NS_799 0 5.4971698738230652e-06
GC_10_800 b_10 NI_10 NS_800 0 3.2160028561156462e-05
GC_10_801 b_10 NI_10 NS_801 0 -8.2126411720176096e-06
GC_10_802 b_10 NI_10 NS_802 0 -2.6520248056848506e-05
GC_10_803 b_10 NI_10 NS_803 0 -1.8293638559269190e-06
GC_10_804 b_10 NI_10 NS_804 0 1.6901090709431998e-06
GC_10_805 b_10 NI_10 NS_805 0 -1.9229428560270311e-05
GC_10_806 b_10 NI_10 NS_806 0 -1.1940389222481743e-05
GC_10_807 b_10 NI_10 NS_807 0 6.9715891744153352e-06
GC_10_808 b_10 NI_10 NS_808 0 2.0939279883679893e-05
GC_10_809 b_10 NI_10 NS_809 0 -1.5976584542618341e-05
GC_10_810 b_10 NI_10 NS_810 0 -1.4813682333410816e-05
GC_10_811 b_10 NI_10 NS_811 0 1.3385310824420153e-06
GC_10_812 b_10 NI_10 NS_812 0 5.3014195794720317e-06
GC_10_813 b_10 NI_10 NS_813 0 -2.4841398253689556e-05
GC_10_814 b_10 NI_10 NS_814 0 -9.8244214895820123e-06
GC_10_815 b_10 NI_10 NS_815 0 8.5458025481600612e-06
GC_10_816 b_10 NI_10 NS_816 0 2.3051008654151455e-05
GC_10_817 b_10 NI_10 NS_817 0 -2.0672703662660086e-05
GC_10_818 b_10 NI_10 NS_818 0 -5.6252259885954029e-06
GC_10_819 b_10 NI_10 NS_819 0 6.2604064349023286e-06
GC_10_820 b_10 NI_10 NS_820 0 7.5159771654689443e-06
GC_10_821 b_10 NI_10 NS_821 0 -3.0565109760336192e-05
GC_10_822 b_10 NI_10 NS_822 0 -2.5578436695823663e-06
GC_10_823 b_10 NI_10 NS_823 0 1.8794275522848392e-05
GC_10_824 b_10 NI_10 NS_824 0 2.5290692919552269e-05
GC_10_825 b_10 NI_10 NS_825 0 -2.1787356141423068e-05
GC_10_826 b_10 NI_10 NS_826 0 6.9643260207717837e-06
GC_10_827 b_10 NI_10 NS_827 0 1.5266698662096949e-05
GC_10_828 b_10 NI_10 NS_828 0 3.9769079034624973e-06
GC_10_829 b_10 NI_10 NS_829 0 -3.4533195634599371e-05
GC_10_830 b_10 NI_10 NS_830 0 1.3723106174819480e-05
GC_10_831 b_10 NI_10 NS_831 0 3.7468924874153128e-05
GC_10_832 b_10 NI_10 NS_832 0 1.2337879215372577e-05
GC_10_833 b_10 NI_10 NS_833 0 -7.7468836914250586e-06
GC_10_834 b_10 NI_10 NS_834 0 1.8808846597873264e-05
GC_10_835 b_10 NI_10 NS_835 0 1.2774791343100730e-05
GC_10_836 b_10 NI_10 NS_836 0 -1.1287273921854961e-05
GC_10_837 b_10 NI_10 NS_837 0 1.0984716475357858e-10
GC_10_838 b_10 NI_10 NS_838 0 3.5338539478619712e-11
GC_10_839 b_10 NI_10 NS_839 0 -1.3692660051997675e-05
GC_10_840 b_10 NI_10 NS_840 0 2.5942031887171665e-05
GC_10_841 b_10 NI_10 NS_841 0 -2.0635045906463176e-06
GC_10_842 b_10 NI_10 NS_842 0 1.0503207742127529e-05
GC_10_843 b_10 NI_10 NS_843 0 6.1728475113391711e-06
GC_10_844 b_10 NI_10 NS_844 0 -8.5363565454743320e-06
GC_10_845 b_10 NI_10 NS_845 0 -8.1127306808112489e-06
GC_10_846 b_10 NI_10 NS_846 0 2.5390653583851210e-05
GC_10_847 b_10 NI_10 NS_847 0 2.4972769712954158e-05
GC_10_848 b_10 NI_10 NS_848 0 -1.0420766964574563e-05
GC_10_849 b_10 NI_10 NS_849 0 4.8846717358321208e-09
GC_10_850 b_10 NI_10 NS_850 0 -1.2244751306513728e-09
GC_10_851 b_10 NI_10 NS_851 0 2.6368528279490749e-05
GC_10_852 b_10 NI_10 NS_852 0 -1.2610361711836045e-05
GC_10_853 b_10 NI_10 NS_853 0 -8.2494854478138578e-06
GC_10_854 b_10 NI_10 NS_854 0 1.8114633830733751e-05
GC_10_855 b_10 NI_10 NS_855 0 -1.0378260422578782e-05
GC_10_856 b_10 NI_10 NS_856 0 -3.0219655162394557e-07
GC_10_857 b_10 NI_10 NS_857 0 1.9390178463993602e-05
GC_10_858 b_10 NI_10 NS_858 0 -1.4388822167994765e-05
GC_10_859 b_10 NI_10 NS_859 0 7.1948776390833339e-06
GC_10_860 b_10 NI_10 NS_860 0 1.1599589215816354e-05
GC_10_861 b_10 NI_10 NS_861 0 -2.2864885374817782e-07
GC_10_862 b_10 NI_10 NS_862 0 -1.4637611571913038e-05
GC_10_863 b_10 NI_10 NS_863 0 1.3160147010652816e-05
GC_10_864 b_10 NI_10 NS_864 0 2.7988798519227731e-05
GC_10_865 b_10 NI_10 NS_865 0 -1.0575813844565891e-02
GC_10_866 b_10 NI_10 NS_866 0 9.5595000797322291e-09
GC_10_867 b_10 NI_10 NS_867 0 9.8516030515516014e-07
GC_10_868 b_10 NI_10 NS_868 0 3.6184053568500416e-05
GC_10_869 b_10 NI_10 NS_869 0 4.3796987846204559e-03
GC_10_870 b_10 NI_10 NS_870 0 -3.4738273572151824e-03
GC_10_871 b_10 NI_10 NS_871 0 -3.7303087976085403e-03
GC_10_872 b_10 NI_10 NS_872 0 6.2452162897856517e-03
GC_10_873 b_10 NI_10 NS_873 0 -8.7506213698409635e-03
GC_10_874 b_10 NI_10 NS_874 0 -5.9709770293565629e-03
GC_10_875 b_10 NI_10 NS_875 0 9.2221481921875431e-03
GC_10_876 b_10 NI_10 NS_876 0 -5.9539987463148175e-03
GC_10_877 b_10 NI_10 NS_877 0 7.1415984118355759e-03
GC_10_878 b_10 NI_10 NS_878 0 1.1891295224266912e-02
GC_10_879 b_10 NI_10 NS_879 0 -4.2237505398800773e-03
GC_10_880 b_10 NI_10 NS_880 0 -1.1434212369576592e-03
GC_10_881 b_10 NI_10 NS_881 0 -8.8759814640091885e-03
GC_10_882 b_10 NI_10 NS_882 0 -4.8952057962337882e-04
GC_10_883 b_10 NI_10 NS_883 0 1.4613641196968881e-02
GC_10_884 b_10 NI_10 NS_884 0 -1.0366832197774839e-02
GC_10_885 b_10 NI_10 NS_885 0 1.6418114294333323e-02
GC_10_886 b_10 NI_10 NS_886 0 4.0449085602744872e-03
GC_10_887 b_10 NI_10 NS_887 0 -1.1484885642233411e-02
GC_10_888 b_10 NI_10 NS_888 0 -2.5531138660868504e-04
GC_10_889 b_10 NI_10 NS_889 0 -1.6635893694787171e-02
GC_10_890 b_10 NI_10 NS_890 0 -4.4594583733408251e-02
GC_10_891 b_10 NI_10 NS_891 0 1.0649465421879303e-02
GC_10_892 b_10 NI_10 NS_892 0 1.1312751632682825e-03
GC_10_893 b_10 NI_10 NS_893 0 -4.8338843232507325e-02
GC_10_894 b_10 NI_10 NS_894 0 1.1008114488516817e-02
GC_10_895 b_10 NI_10 NS_895 0 -1.0431960656455979e-02
GC_10_896 b_10 NI_10 NS_896 0 4.9182029671494072e-04
GC_10_897 b_10 NI_10 NS_897 0 9.7750129390908169e-03
GC_10_898 b_10 NI_10 NS_898 0 -5.7664994236781327e-04
GC_10_899 b_10 NI_10 NS_899 0 4.5629913452846990e-03
GC_10_900 b_10 NI_10 NS_900 0 2.4175388649885516e-02
GC_10_901 b_10 NI_10 NS_901 0 -1.0747452316886941e-02
GC_10_902 b_10 NI_10 NS_902 0 1.9594185762073658e-03
GC_10_903 b_10 NI_10 NS_903 0 -8.4817403504705863e-03
GC_10_904 b_10 NI_10 NS_904 0 -1.3531511683060460e-02
GC_10_905 b_10 NI_10 NS_905 0 1.0144391659537816e-02
GC_10_906 b_10 NI_10 NS_906 0 9.9163190992940589e-04
GC_10_907 b_10 NI_10 NS_907 0 -1.9215667499628625e-02
GC_10_908 b_10 NI_10 NS_908 0 2.8664614532787437e-02
GC_10_909 b_10 NI_10 NS_909 0 -9.6176245686748138e-03
GC_10_910 b_10 NI_10 NS_910 0 -9.6670243660712963e-04
GC_10_911 b_10 NI_10 NS_911 0 1.8850236376783587e-03
GC_10_912 b_10 NI_10 NS_912 0 -1.3790869189776265e-03
GC_10_913 b_10 NI_10 NS_913 0 9.4568126307968299e-03
GC_10_914 b_10 NI_10 NS_914 0 -2.3685228806114676e-04
GC_10_915 b_10 NI_10 NS_915 0 -2.0769913891800906e-04
GC_10_916 b_10 NI_10 NS_916 0 3.0287225815225197e-02
GC_10_917 b_10 NI_10 NS_917 0 -8.5365121254759573e-03
GC_10_918 b_10 NI_10 NS_918 0 1.5564869014196255e-04
GC_10_919 b_10 NI_10 NS_919 0 2.0684949366814382e-04
GC_10_920 b_10 NI_10 NS_920 0 -5.4692454922850124e-03
GC_10_921 b_10 NI_10 NS_921 0 1.0024581951580147e-02
GC_10_922 b_10 NI_10 NS_922 0 -3.2646578442430601e-04
GC_10_923 b_10 NI_10 NS_923 0 8.8940172499950860e-03
GC_10_924 b_10 NI_10 NS_924 0 2.6408722584590510e-02
GC_10_925 b_10 NI_10 NS_925 0 -8.3634730202592957e-03
GC_10_926 b_10 NI_10 NS_926 0 1.3809941229067442e-03
GC_10_927 b_10 NI_10 NS_927 0 -2.5879657944743555e-03
GC_10_928 b_10 NI_10 NS_928 0 -7.3315733123782900e-03
GC_10_929 b_10 NI_10 NS_929 0 1.0540538790800401e-02
GC_10_930 b_10 NI_10 NS_930 0 -8.1039972133489780e-04
GC_10_931 b_10 NI_10 NS_931 0 1.4431150419409948e-02
GC_10_932 b_10 NI_10 NS_932 0 2.0002733939750019e-02
GC_10_933 b_10 NI_10 NS_933 0 -8.2822059246821476e-03
GC_10_934 b_10 NI_10 NS_934 0 2.9406926195107977e-03
GC_10_935 b_10 NI_10 NS_935 0 -5.5808175597408293e-03
GC_10_936 b_10 NI_10 NS_936 0 -6.8969498956083083e-03
GC_10_937 b_10 NI_10 NS_937 0 1.1228136753316209e-02
GC_10_938 b_10 NI_10 NS_938 0 -1.3571923626691865e-03
GC_10_939 b_10 NI_10 NS_939 0 1.5726443230910735e-02
GC_10_940 b_10 NI_10 NS_940 0 1.2982464199572649e-02
GC_10_941 b_10 NI_10 NS_941 0 -7.1842400666946122e-03
GC_10_942 b_10 NI_10 NS_942 0 5.1249192588046126e-03
GC_10_943 b_10 NI_10 NS_943 0 -6.8612398462710132e-03
GC_10_944 b_10 NI_10 NS_944 0 -4.8303770995999423e-03
GC_10_945 b_10 NI_10 NS_945 0 5.1316152633800971e-09
GC_10_946 b_10 NI_10 NS_946 0 4.4376001550661304e-08
GC_10_947 b_10 NI_10 NS_947 0 1.2002073526814452e-02
GC_10_948 b_10 NI_10 NS_948 0 -2.5554187167626599e-03
GC_10_949 b_10 NI_10 NS_949 0 -5.2431605617128752e-03
GC_10_950 b_10 NI_10 NS_950 0 4.7077149664145829e-03
GC_10_951 b_10 NI_10 NS_951 0 -6.1541485641369974e-03
GC_10_952 b_10 NI_10 NS_952 0 -4.3159890494544537e-03
GC_10_953 b_10 NI_10 NS_953 0 1.1759641943645191e-02
GC_10_954 b_10 NI_10 NS_954 0 -3.7149034963143640e-03
GC_10_955 b_10 NI_10 NS_955 0 1.3000704445995869e-02
GC_10_956 b_10 NI_10 NS_956 0 9.4708226650160824e-03
GC_10_957 b_10 NI_10 NS_957 0 3.9444991209087498e-06
GC_10_958 b_10 NI_10 NS_958 0 -9.3342609517765419e-07
GC_10_959 b_10 NI_10 NS_959 0 1.6111759045012913e-02
GC_10_960 b_10 NI_10 NS_960 0 1.6784786458934973e-02
GC_10_961 b_10 NI_10 NS_961 0 1.2052345234300699e-02
GC_10_962 b_10 NI_10 NS_962 0 -2.4747655897065105e-03
GC_10_963 b_10 NI_10 NS_963 0 -8.3473626535816251e-03
GC_10_964 b_10 NI_10 NS_964 0 8.3966091170478043e-05
GC_10_965 b_10 NI_10 NS_965 0 1.1340524046310684e-02
GC_10_966 b_10 NI_10 NS_966 0 7.3400096830970865e-03
GC_10_967 b_10 NI_10 NS_967 0 -4.6549366351306192e-03
GC_10_968 b_10 NI_10 NS_968 0 7.3654636451295817e-03
GC_10_969 b_10 NI_10 NS_969 0 -8.0793067210239780e-03
GC_10_970 b_10 NI_10 NS_970 0 -3.7189954644689768e-03
GC_10_971 b_10 NI_10 NS_971 0 1.5982961900398968e-02
GC_10_972 b_10 NI_10 NS_972 0 -7.7384993754638200e-03
GC_10_973 b_10 NI_10 NS_973 0 -1.4246400256030944e-02
GC_10_974 b_10 NI_10 NS_974 0 6.2293160768216438e-09
GC_10_975 b_10 NI_10 NS_975 0 -1.0771399406067461e-06
GC_10_976 b_10 NI_10 NS_976 0 -2.3238215206440735e-05
GC_10_977 b_10 NI_10 NS_977 0 3.4199266343494576e-04
GC_10_978 b_10 NI_10 NS_978 0 -1.9835114711510098e-04
GC_10_979 b_10 NI_10 NS_979 0 -1.5573869762491497e-03
GC_10_980 b_10 NI_10 NS_980 0 -2.3367645319626856e-03
GC_10_981 b_10 NI_10 NS_981 0 -6.7656858961235585e-05
GC_10_982 b_10 NI_10 NS_982 0 4.3764648565270282e-03
GC_10_983 b_10 NI_10 NS_983 0 1.6012909917152984e-03
GC_10_984 b_10 NI_10 NS_984 0 -5.9363791255959263e-03
GC_10_985 b_10 NI_10 NS_985 0 -4.9862942191486164e-03
GC_10_986 b_10 NI_10 NS_986 0 6.4938569038295382e-03
GC_10_987 b_10 NI_10 NS_987 0 1.1242574208519831e-03
GC_10_988 b_10 NI_10 NS_988 0 -4.9042309876357471e-04
GC_10_989 b_10 NI_10 NS_989 0 2.8092071387607631e-03
GC_10_990 b_10 NI_10 NS_990 0 2.3585353006908101e-03
GC_10_991 b_10 NI_10 NS_991 0 -4.3182735494993983e-03
GC_10_992 b_10 NI_10 NS_992 0 -1.3539567903206089e-02
GC_10_993 b_10 NI_10 NS_993 0 1.6031707990063538e-03
GC_10_994 b_10 NI_10 NS_994 0 1.7677776973712766e-02
GC_10_995 b_10 NI_10 NS_995 0 9.8386853699242542e-03
GC_10_996 b_10 NI_10 NS_996 0 -2.2919452674644183e-03
GC_10_997 b_10 NI_10 NS_997 0 -1.3104487520470600e-02
GC_10_998 b_10 NI_10 NS_998 0 2.2186351324758997e-03
GC_10_999 b_10 NI_10 NS_999 0 9.2001458916820510e-03
GC_10_1000 b_10 NI_10 NS_1000 0 1.9506148644373145e-03
GC_10_1001 b_10 NI_10 NS_1001 0 -1.7998043609794144e-02
GC_10_1002 b_10 NI_10 NS_1002 0 -6.4920163427329095e-03
GC_10_1003 b_10 NI_10 NS_1003 0 1.5711166851321963e-02
GC_10_1004 b_10 NI_10 NS_1004 0 6.4981549055297162e-03
GC_10_1005 b_10 NI_10 NS_1005 0 8.1166025771045869e-03
GC_10_1006 b_10 NI_10 NS_1006 0 -4.1938599544669572e-03
GC_10_1007 b_10 NI_10 NS_1007 0 -7.5320604141215740e-03
GC_10_1008 b_10 NI_10 NS_1008 0 2.0324522546205787e-03
GC_10_1009 b_10 NI_10 NS_1009 0 6.7023914700823873e-03
GC_10_1010 b_10 NI_10 NS_1010 0 -2.7451417078800961e-03
GC_10_1011 b_10 NI_10 NS_1011 0 -6.5840314599315058e-03
GC_10_1012 b_10 NI_10 NS_1012 0 2.8920091767601699e-03
GC_10_1013 b_10 NI_10 NS_1013 0 7.6634824591408452e-03
GC_10_1014 b_10 NI_10 NS_1014 0 4.8601602431006213e-04
GC_10_1015 b_10 NI_10 NS_1015 0 -9.3542684002526928e-03
GC_10_1016 b_10 NI_10 NS_1016 0 -5.1821823155190445e-03
GC_10_1017 b_10 NI_10 NS_1017 0 6.8205079141039088e-03
GC_10_1018 b_10 NI_10 NS_1018 0 4.1105978305454073e-03
GC_10_1019 b_10 NI_10 NS_1019 0 -3.8505593707261957e-04
GC_10_1020 b_10 NI_10 NS_1020 0 -9.3423498820468078e-04
GC_10_1021 b_10 NI_10 NS_1021 0 5.6830560567737954e-03
GC_10_1022 b_10 NI_10 NS_1022 0 -1.3773210671377595e-03
GC_10_1023 b_10 NI_10 NS_1023 0 -9.1525589686274039e-03
GC_10_1024 b_10 NI_10 NS_1024 0 -1.2845549510707109e-03
GC_10_1025 b_10 NI_10 NS_1025 0 5.9995912358442897e-03
GC_10_1026 b_10 NI_10 NS_1026 0 7.3474949662859093e-04
GC_10_1027 b_10 NI_10 NS_1027 0 -2.6407532414302183e-03
GC_10_1028 b_10 NI_10 NS_1028 0 2.3246011121348884e-04
GC_10_1029 b_10 NI_10 NS_1029 0 6.7119817333126932e-03
GC_10_1030 b_10 NI_10 NS_1030 0 -2.2566059982603408e-03
GC_10_1031 b_10 NI_10 NS_1031 0 -9.2876748456725538e-03
GC_10_1032 b_10 NI_10 NS_1032 0 1.4716659449841003e-03
GC_10_1033 b_10 NI_10 NS_1033 0 5.7396120360619753e-03
GC_10_1034 b_10 NI_10 NS_1034 0 -1.5055499470718679e-03
GC_10_1035 b_10 NI_10 NS_1035 0 -3.3169903661782523e-03
GC_10_1036 b_10 NI_10 NS_1036 0 2.3821024421819010e-03
GC_10_1037 b_10 NI_10 NS_1037 0 7.2818936807726520e-03
GC_10_1038 b_10 NI_10 NS_1038 0 -4.0976796271503333e-03
GC_10_1039 b_10 NI_10 NS_1039 0 -8.5931345432147463e-03
GC_10_1040 b_10 NI_10 NS_1040 0 4.1427763954098445e-03
GC_10_1041 b_10 NI_10 NS_1041 0 4.8244396283542140e-03
GC_10_1042 b_10 NI_10 NS_1042 0 -3.8807312376367910e-03
GC_10_1043 b_10 NI_10 NS_1043 0 -2.4175655609633214e-03
GC_10_1044 b_10 NI_10 NS_1044 0 4.7355196559176020e-03
GC_10_1045 b_10 NI_10 NS_1045 0 7.0698660120576337e-03
GC_10_1046 b_10 NI_10 NS_1046 0 -7.3594026153947249e-03
GC_10_1047 b_10 NI_10 NS_1047 0 -7.1573588934073845e-03
GC_10_1048 b_10 NI_10 NS_1048 0 6.8575791856925836e-03
GC_10_1049 b_10 NI_10 NS_1049 0 1.6629097338060801e-03
GC_10_1050 b_10 NI_10 NS_1050 0 -5.3099127673499292e-03
GC_10_1051 b_10 NI_10 NS_1051 0 5.8005351314575763e-04
GC_10_1052 b_10 NI_10 NS_1052 0 5.4707649844612386e-03
GC_10_1053 b_10 NI_10 NS_1053 0 -4.5818073808091558e-09
GC_10_1054 b_10 NI_10 NS_1054 0 -1.3467649890979608e-08
GC_10_1055 b_10 NI_10 NS_1055 0 2.7089365488081898e-03
GC_10_1056 b_10 NI_10 NS_1056 0 -8.5910067713740774e-03
GC_10_1057 b_10 NI_10 NS_1057 0 8.6608706430445236e-04
GC_10_1058 b_10 NI_10 NS_1058 0 -3.4347604172177463e-03
GC_10_1059 b_10 NI_10 NS_1059 0 6.2756551860500102e-04
GC_10_1060 b_10 NI_10 NS_1060 0 4.0313415341296684e-03
GC_10_1061 b_10 NI_10 NS_1061 0 2.1670484566331375e-03
GC_10_1062 b_10 NI_10 NS_1062 0 -8.1665277093597704e-03
GC_10_1063 b_10 NI_10 NS_1063 0 -3.4991635045162226e-03
GC_10_1064 b_10 NI_10 NS_1064 0 7.0126788784460221e-03
GC_10_1065 b_10 NI_10 NS_1065 0 -1.0829860079787106e-07
GC_10_1066 b_10 NI_10 NS_1066 0 -3.0048166007703716e-07
GC_10_1067 b_10 NI_10 NS_1067 0 -8.0240632959311144e-03
GC_10_1068 b_10 NI_10 NS_1068 0 5.3776059369874257e-03
GC_10_1069 b_10 NI_10 NS_1069 0 4.1768102857437277e-03
GC_10_1070 b_10 NI_10 NS_1070 0 -6.8620734780150657e-03
GC_10_1071 b_10 NI_10 NS_1071 0 5.3214177374611279e-03
GC_10_1072 b_10 NI_10 NS_1072 0 7.4369283070833503e-04
GC_10_1073 b_10 NI_10 NS_1073 0 -2.3651597210068713e-03
GC_10_1074 b_10 NI_10 NS_1074 0 6.8561897696881010e-03
GC_10_1075 b_10 NI_10 NS_1075 0 -1.4960016228828792e-03
GC_10_1076 b_10 NI_10 NS_1076 0 -4.2193424589340115e-03
GC_10_1077 b_10 NI_10 NS_1077 0 2.3601153783920003e-03
GC_10_1078 b_10 NI_10 NS_1078 0 5.0361467955908666e-03
GC_10_1079 b_10 NI_10 NS_1079 0 -2.0068772397933460e-03
GC_10_1080 b_10 NI_10 NS_1080 0 -8.9761631515452682e-03
GC_10_1081 b_10 NI_10 NS_1081 0 -3.3036468467205803e-03
GC_10_1082 b_10 NI_10 NS_1082 0 1.8493852371142535e-09
GC_10_1083 b_10 NI_10 NS_1083 0 5.6032182830583812e-08
GC_10_1084 b_10 NI_10 NS_1084 0 1.8929694312798604e-06
GC_10_1085 b_10 NI_10 NS_1085 0 -9.1167743590498356e-05
GC_10_1086 b_10 NI_10 NS_1086 0 -5.7737884515204474e-05
GC_10_1087 b_10 NI_10 NS_1087 0 -1.2657732808128239e-03
GC_10_1088 b_10 NI_10 NS_1088 0 -2.9559373658780375e-04
GC_10_1089 b_10 NI_10 NS_1089 0 -1.6792131979911642e-03
GC_10_1090 b_10 NI_10 NS_1090 0 2.6464978146337535e-03
GC_10_1091 b_10 NI_10 NS_1091 0 5.1121228689390071e-04
GC_10_1092 b_10 NI_10 NS_1092 0 5.4276090903376730e-03
GC_10_1093 b_10 NI_10 NS_1093 0 7.1034889642706900e-03
GC_10_1094 b_10 NI_10 NS_1094 0 6.3629114794539951e-04
GC_10_1095 b_10 NI_10 NS_1095 0 6.4433017886676833e-04
GC_10_1096 b_10 NI_10 NS_1096 0 -6.6092009615995690e-04
GC_10_1097 b_10 NI_10 NS_1097 0 1.0576971634783552e-03
GC_10_1098 b_10 NI_10 NS_1098 0 1.5711403288683505e-03
GC_10_1099 b_10 NI_10 NS_1099 0 1.2687514716068831e-02
GC_10_1100 b_10 NI_10 NS_1100 0 1.3123212006357486e-02
GC_10_1101 b_10 NI_10 NS_1101 0 8.7187958059280687e-03
GC_10_1102 b_10 NI_10 NS_1102 0 -2.0392081307234116e-02
GC_10_1103 b_10 NI_10 NS_1103 0 8.3891006126972680e-03
GC_10_1104 b_10 NI_10 NS_1104 0 -2.9045267726896017e-03
GC_10_1105 b_10 NI_10 NS_1105 0 -1.2701294118210162e-02
GC_10_1106 b_10 NI_10 NS_1106 0 -3.8806698399796571e-02
GC_10_1107 b_10 NI_10 NS_1107 0 -7.2523396004929219e-03
GC_10_1108 b_10 NI_10 NS_1108 0 -2.1332744415701291e-03
GC_10_1109 b_10 NI_10 NS_1109 0 -5.2307204283657115e-02
GC_10_1110 b_10 NI_10 NS_1110 0 -1.7936126773729002e-03
GC_10_1111 b_10 NI_10 NS_1111 0 1.4914417235231995e-02
GC_10_1112 b_10 NI_10 NS_1112 0 8.6735768571818590e-03
GC_10_1113 b_10 NI_10 NS_1113 0 -5.9233541230436833e-03
GC_10_1114 b_10 NI_10 NS_1114 0 5.0044976616262140e-03
GC_10_1115 b_10 NI_10 NS_1115 0 8.3724192684992670e-03
GC_10_1116 b_10 NI_10 NS_1116 0 1.1688366973152635e-02
GC_10_1117 b_10 NI_10 NS_1117 0 4.5592638701915360e-03
GC_10_1118 b_10 NI_10 NS_1118 0 -2.9327397535174665e-03
GC_10_1119 b_10 NI_10 NS_1119 0 -7.8986718119426810e-03
GC_10_1120 b_10 NI_10 NS_1120 0 -8.1490630682327838e-03
GC_10_1121 b_10 NI_10 NS_1121 0 -5.6808135799187552e-03
GC_10_1122 b_10 NI_10 NS_1122 0 -6.1280929029166274e-04
GC_10_1123 b_10 NI_10 NS_1123 0 -1.8070847597754076e-02
GC_10_1124 b_10 NI_10 NS_1124 0 1.3578968444085435e-02
GC_10_1125 b_10 NI_10 NS_1125 0 4.7069876812876436e-03
GC_10_1126 b_10 NI_10 NS_1126 0 4.3794382429170383e-03
GC_10_1127 b_10 NI_10 NS_1127 0 6.5015895965032044e-04
GC_10_1128 b_10 NI_10 NS_1128 0 -1.0995412894793043e-04
GC_10_1129 b_10 NI_10 NS_1129 0 -3.7963992693998325e-03
GC_10_1130 b_10 NI_10 NS_1130 0 8.8498856452297011e-04
GC_10_1131 b_10 NI_10 NS_1131 0 -1.1178265542558536e-03
GC_10_1132 b_10 NI_10 NS_1132 0 1.6699689321745956e-02
GC_10_1133 b_10 NI_10 NS_1133 0 4.4472810558010599e-03
GC_10_1134 b_10 NI_10 NS_1134 0 7.0796491261417580e-04
GC_10_1135 b_10 NI_10 NS_1135 0 -5.1995706764918642e-04
GC_10_1136 b_10 NI_10 NS_1136 0 -2.2477503300167520e-03
GC_10_1137 b_10 NI_10 NS_1137 0 -4.9864550057338117e-03
GC_10_1138 b_10 NI_10 NS_1138 0 2.1108885148027647e-03
GC_10_1139 b_10 NI_10 NS_1139 0 7.3425321211990687e-03
GC_10_1140 b_10 NI_10 NS_1140 0 1.4345855450848603e-02
GC_10_1141 b_10 NI_10 NS_1141 0 4.1872288154565923e-03
GC_10_1142 b_10 NI_10 NS_1142 0 -1.6838584141340828e-03
GC_10_1143 b_10 NI_10 NS_1143 0 -3.3981227807577306e-03
GC_10_1144 b_10 NI_10 NS_1144 0 -2.1006244639393316e-03
GC_10_1145 b_10 NI_10 NS_1145 0 -5.4204239050152500e-03
GC_10_1146 b_10 NI_10 NS_1146 0 4.3817247946772789e-03
GC_10_1147 b_10 NI_10 NS_1147 0 1.3196875164562106e-02
GC_10_1148 b_10 NI_10 NS_1148 0 8.4333025960762215e-03
GC_10_1149 b_10 NI_10 NS_1149 0 2.8324347581599055e-03
GC_10_1150 b_10 NI_10 NS_1150 0 -4.1306074025395396e-03
GC_10_1151 b_10 NI_10 NS_1151 0 -5.3207869859125435e-03
GC_10_1152 b_10 NI_10 NS_1152 0 1.1381564650091301e-03
GC_10_1153 b_10 NI_10 NS_1153 0 -4.4310195627860777e-03
GC_10_1154 b_10 NI_10 NS_1154 0 8.3104298969830619e-03
GC_10_1155 b_10 NI_10 NS_1155 0 1.4612784030967715e-02
GC_10_1156 b_10 NI_10 NS_1156 0 -4.6824941615916286e-04
GC_10_1157 b_10 NI_10 NS_1157 0 -1.1845324017182325e-03
GC_10_1158 b_10 NI_10 NS_1158 0 -4.5473906517052905e-03
GC_10_1159 b_10 NI_10 NS_1159 0 -2.2825683634711859e-03
GC_10_1160 b_10 NI_10 NS_1160 0 4.3832546916945684e-03
GC_10_1161 b_10 NI_10 NS_1161 0 1.3572125749263832e-10
GC_10_1162 b_10 NI_10 NS_1162 0 -1.5466291439467210e-09
GC_10_1163 b_10 NI_10 NS_1163 0 1.4460258772959408e-03
GC_10_1164 b_10 NI_10 NS_1164 0 8.2165464976339253e-03
GC_10_1165 b_10 NI_10 NS_1165 0 -8.7895028612762450e-04
GC_10_1166 b_10 NI_10 NS_1166 0 -2.2072127801078967e-03
GC_10_1167 b_10 NI_10 NS_1167 0 -1.4679137055256259e-03
GC_10_1168 b_10 NI_10 NS_1168 0 2.7519857583777397e-03
GC_10_1169 b_10 NI_10 NS_1169 0 1.7320144525156832e-03
GC_10_1170 b_10 NI_10 NS_1170 0 7.6059319534155833e-03
GC_10_1171 b_10 NI_10 NS_1171 0 7.5874083955443442e-03
GC_10_1172 b_10 NI_10 NS_1172 0 -3.8276827721217786e-03
GC_10_1173 b_10 NI_10 NS_1173 0 -5.2101119458921127e-08
GC_10_1174 b_10 NI_10 NS_1174 0 -2.0817341836911985e-08
GC_10_1175 b_10 NI_10 NS_1175 0 1.1391243302973078e-02
GC_10_1176 b_10 NI_10 NS_1176 0 4.4700329649389140e-03
GC_10_1177 b_10 NI_10 NS_1177 0 -8.6185047828051496e-04
GC_10_1178 b_10 NI_10 NS_1178 0 6.4916224698060038e-03
GC_10_1179 b_10 NI_10 NS_1179 0 3.6263738522131434e-03
GC_10_1180 b_10 NI_10 NS_1180 0 4.0710467479625927e-04
GC_10_1181 b_10 NI_10 NS_1181 0 6.0525103069943628e-03
GC_10_1182 b_10 NI_10 NS_1182 0 -4.6635403232154074e-03
GC_10_1183 b_10 NI_10 NS_1183 0 -3.3929753833683639e-03
GC_10_1184 b_10 NI_10 NS_1184 0 -1.3533959440472391e-03
GC_10_1185 b_10 NI_10 NS_1185 0 1.1237967035868938e-04
GC_10_1186 b_10 NI_10 NS_1186 0 4.4958002999552216e-03
GC_10_1187 b_10 NI_10 NS_1187 0 7.2795569203941155e-03
GC_10_1188 b_10 NI_10 NS_1188 0 5.5305048222505033e-03
GC_10_1189 b_10 NI_10 NS_1189 0 1.1804777683495674e-03
GC_10_1190 b_10 NI_10 NS_1190 0 -3.5559914947529153e-09
GC_10_1191 b_10 NI_10 NS_1191 0 -4.8002576919061797e-08
GC_10_1192 b_10 NI_10 NS_1192 0 -3.4752161331347059e-06
GC_10_1193 b_10 NI_10 NS_1193 0 -3.6812591732166266e-04
GC_10_1194 b_10 NI_10 NS_1194 0 1.3598228422269945e-04
GC_10_1195 b_10 NI_10 NS_1195 0 1.1297229504253134e-03
GC_10_1196 b_10 NI_10 NS_1196 0 1.9432474187168031e-03
GC_10_1197 b_10 NI_10 NS_1197 0 -6.5058703572615884e-05
GC_10_1198 b_10 NI_10 NS_1198 0 -3.4937467840565101e-03
GC_10_1199 b_10 NI_10 NS_1199 0 -1.5644000874450823e-03
GC_10_1200 b_10 NI_10 NS_1200 0 5.0906047862238008e-03
GC_10_1201 b_10 NI_10 NS_1201 0 4.2534009791018301e-03
GC_10_1202 b_10 NI_10 NS_1202 0 -4.9938043723831991e-03
GC_10_1203 b_10 NI_10 NS_1203 0 -1.0085534104761970e-03
GC_10_1204 b_10 NI_10 NS_1204 0 5.6397848515128777e-04
GC_10_1205 b_10 NI_10 NS_1205 0 -2.0807522902705649e-03
GC_10_1206 b_10 NI_10 NS_1206 0 -1.8633136559348135e-03
GC_10_1207 b_10 NI_10 NS_1207 0 3.6454404149434895e-03
GC_10_1208 b_10 NI_10 NS_1208 0 1.1647363854914146e-02
GC_10_1209 b_10 NI_10 NS_1209 0 -8.9814490637171675e-04
GC_10_1210 b_10 NI_10 NS_1210 0 -1.4854322467497029e-02
GC_10_1211 b_10 NI_10 NS_1211 0 -8.1235366917756808e-03
GC_10_1212 b_10 NI_10 NS_1212 0 1.9196054013951708e-03
GC_10_1213 b_10 NI_10 NS_1213 0 1.1263052262444591e-02
GC_10_1214 b_10 NI_10 NS_1214 0 -1.8122303811994749e-03
GC_10_1215 b_10 NI_10 NS_1215 0 -7.5672721671333817e-03
GC_10_1216 b_10 NI_10 NS_1216 0 -1.6811809006930733e-03
GC_10_1217 b_10 NI_10 NS_1217 0 1.5281711704014636e-02
GC_10_1218 b_10 NI_10 NS_1218 0 5.3008478715180418e-03
GC_10_1219 b_10 NI_10 NS_1219 0 -1.3082857193876057e-02
GC_10_1220 b_10 NI_10 NS_1220 0 -5.4612980857567245e-03
GC_10_1221 b_10 NI_10 NS_1221 0 -6.6370720068815829e-03
GC_10_1222 b_10 NI_10 NS_1222 0 3.4566941278901492e-03
GC_10_1223 b_10 NI_10 NS_1223 0 6.3616038437344993e-03
GC_10_1224 b_10 NI_10 NS_1224 0 -1.8793238139981541e-03
GC_10_1225 b_10 NI_10 NS_1225 0 -5.4737178432874376e-03
GC_10_1226 b_10 NI_10 NS_1226 0 2.1830275702705280e-03
GC_10_1227 b_10 NI_10 NS_1227 0 5.3937685500656061e-03
GC_10_1228 b_10 NI_10 NS_1228 0 -2.6324368439134926e-03
GC_10_1229 b_10 NI_10 NS_1229 0 -6.3064548530876591e-03
GC_10_1230 b_10 NI_10 NS_1230 0 -4.8381422322162359e-04
GC_10_1231 b_10 NI_10 NS_1231 0 7.6452813373800721e-03
GC_10_1232 b_10 NI_10 NS_1232 0 3.6298748801943332e-03
GC_10_1233 b_10 NI_10 NS_1233 0 -5.8336237575828086e-03
GC_10_1234 b_10 NI_10 NS_1234 0 -3.4645950540191598e-03
GC_10_1235 b_10 NI_10 NS_1235 0 2.9620064699019242e-04
GC_10_1236 b_10 NI_10 NS_1236 0 5.5810490949433750e-04
GC_10_1237 b_10 NI_10 NS_1237 0 -4.9270622018716464e-03
GC_10_1238 b_10 NI_10 NS_1238 0 8.9219844387952805e-04
GC_10_1239 b_10 NI_10 NS_1239 0 6.2063433395615712e-03
GC_10_1240 b_10 NI_10 NS_1240 0 6.8827280037042496e-04
GC_10_1241 b_10 NI_10 NS_1241 0 -5.3209627948279659e-03
GC_10_1242 b_10 NI_10 NS_1242 0 -4.8419034240273438e-04
GC_10_1243 b_10 NI_10 NS_1243 0 1.5503311578845796e-03
GC_10_1244 b_10 NI_10 NS_1244 0 -4.3208426471623007e-05
GC_10_1245 b_10 NI_10 NS_1245 0 -6.0223341909894116e-03
GC_10_1246 b_10 NI_10 NS_1246 0 1.9232416158412493e-03
GC_10_1247 b_10 NI_10 NS_1247 0 6.2616668284918480e-03
GC_10_1248 b_10 NI_10 NS_1248 0 2.1736512536766315e-04
GC_10_1249 b_10 NI_10 NS_1249 0 -5.0591977956352735e-03
GC_10_1250 b_10 NI_10 NS_1250 0 1.7016169638886087e-03
GC_10_1251 b_10 NI_10 NS_1251 0 2.4884743734153018e-03
GC_10_1252 b_10 NI_10 NS_1252 0 -9.5765186686207996e-04
GC_10_1253 b_10 NI_10 NS_1253 0 -6.5329624741575377e-03
GC_10_1254 b_10 NI_10 NS_1254 0 3.8846374153698937e-03
GC_10_1255 b_10 NI_10 NS_1255 0 7.4932671045403118e-03
GC_10_1256 b_10 NI_10 NS_1256 0 -1.0960284059476624e-03
GC_10_1257 b_10 NI_10 NS_1257 0 -3.9851195992951565e-03
GC_10_1258 b_10 NI_10 NS_1258 0 4.0409800184820245e-03
GC_10_1259 b_10 NI_10 NS_1259 0 2.8633259784483058e-03
GC_10_1260 b_10 NI_10 NS_1260 0 -3.0534881857052169e-03
GC_10_1261 b_10 NI_10 NS_1261 0 -6.0227294634723587e-03
GC_10_1262 b_10 NI_10 NS_1262 0 7.2373898824168881e-03
GC_10_1263 b_10 NI_10 NS_1263 0 7.9897123603499300e-03
GC_10_1264 b_10 NI_10 NS_1264 0 -4.8114592221877809e-03
GC_10_1265 b_10 NI_10 NS_1265 0 -5.3741854794194053e-04
GC_10_1266 b_10 NI_10 NS_1266 0 5.0204729911852795e-03
GC_10_1267 b_10 NI_10 NS_1267 0 2.4825585937046733e-04
GC_10_1268 b_10 NI_10 NS_1268 0 -4.7581979868240613e-03
GC_10_1269 b_10 NI_10 NS_1269 0 1.8109009045382304e-09
GC_10_1270 b_10 NI_10 NS_1270 0 3.2745350759694328e-09
GC_10_1271 b_10 NI_10 NS_1271 0 -1.4271956704142406e-03
GC_10_1272 b_10 NI_10 NS_1272 0 7.8707399222079037e-03
GC_10_1273 b_10 NI_10 NS_1273 0 -1.7997912138199582e-04
GC_10_1274 b_10 NI_10 NS_1274 0 3.0272438861498278e-03
GC_10_1275 b_10 NI_10 NS_1275 0 -1.3038560981470660e-04
GC_10_1276 b_10 NI_10 NS_1276 0 -3.3753040658697246e-03
GC_10_1277 b_10 NI_10 NS_1277 0 -8.7631227784927372e-04
GC_10_1278 b_10 NI_10 NS_1278 0 7.5304822482262154e-03
GC_10_1279 b_10 NI_10 NS_1279 0 3.7888078988001267e-03
GC_10_1280 b_10 NI_10 NS_1280 0 -6.1574217064608271e-03
GC_10_1281 b_10 NI_10 NS_1281 0 8.6236192411829841e-08
GC_10_1282 b_10 NI_10 NS_1282 0 -3.5294023117688274e-07
GC_10_1283 b_10 NI_10 NS_1283 0 6.7186800340163838e-03
GC_10_1284 b_10 NI_10 NS_1284 0 -5.3194114838276199e-03
GC_10_1285 b_10 NI_10 NS_1285 0 -2.6111717720343763e-03
GC_10_1286 b_10 NI_10 NS_1286 0 6.0542407261782779e-03
GC_10_1287 b_10 NI_10 NS_1287 0 -4.2922715109812576e-03
GC_10_1288 b_10 NI_10 NS_1288 0 1.4429442712238376e-05
GC_10_1289 b_10 NI_10 NS_1289 0 2.7173883569819096e-03
GC_10_1290 b_10 NI_10 NS_1290 0 -6.2040232047717902e-03
GC_10_1291 b_10 NI_10 NS_1291 0 2.0957197437900294e-03
GC_10_1292 b_10 NI_10 NS_1292 0 3.2562724655940943e-03
GC_10_1293 b_10 NI_10 NS_1293 0 -1.9700345763534240e-03
GC_10_1294 b_10 NI_10 NS_1294 0 -4.4205367865173158e-03
GC_10_1295 b_10 NI_10 NS_1295 0 2.8640861259799835e-03
GC_10_1296 b_10 NI_10 NS_1296 0 8.0083630266011199e-03
GD_10_1 b_10 NI_10 NA_1 0 8.8077194058505180e-06
GD_10_2 b_10 NI_10 NA_2 0 -1.1492069396679217e-06
GD_10_3 b_10 NI_10 NA_3 0 2.0977618624591634e-06
GD_10_4 b_10 NI_10 NA_4 0 -7.3787014107040665e-06
GD_10_5 b_10 NI_10 NA_5 0 1.5904539956893246e-05
GD_10_6 b_10 NI_10 NA_6 0 5.7657636627220263e-08
GD_10_7 b_10 NI_10 NA_7 0 1.0462081506731580e-04
GD_10_8 b_10 NI_10 NA_8 0 2.6301361602033636e-05
GD_10_9 b_10 NI_10 NA_9 0 -5.0002986467510601e-03
GD_10_10 b_10 NI_10 NA_10 0 -1.0894630938571620e-02
GD_10_11 b_10 NI_10 NA_11 0 -1.1524164237483915e-03
GD_10_12 b_10 NI_10 NA_12 0 1.0616252270114096e-02
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 1.0244822794525164e-05
GC_11_2 b_11 NI_11 NS_2 0 -4.7957776193668679e-12
GC_11_3 b_11 NI_11 NS_3 0 1.0352126557291859e-11
GC_11_4 b_11 NI_11 NS_4 0 3.7845747542673630e-10
GC_11_5 b_11 NI_11 NS_5 0 1.3512318958511033e-07
GC_11_6 b_11 NI_11 NS_6 0 1.0761649168650469e-07
GC_11_7 b_11 NI_11 NS_7 0 7.2007398076211541e-07
GC_11_8 b_11 NI_11 NS_8 0 -1.8726838982061212e-07
GC_11_9 b_11 NI_11 NS_9 0 -5.9814074734497369e-07
GC_11_10 b_11 NI_11 NS_10 0 -3.6306362198031499e-07
GC_11_11 b_11 NI_11 NS_11 0 1.3989865035106945e-06
GC_11_12 b_11 NI_11 NS_12 0 3.2532219320448145e-07
GC_11_13 b_11 NI_11 NS_13 0 -9.9970701765863596e-07
GC_11_14 b_11 NI_11 NS_14 0 -1.7789572862708579e-06
GC_11_15 b_11 NI_11 NS_15 0 2.5545132789392265e-07
GC_11_16 b_11 NI_11 NS_16 0 -5.4830032526922591e-09
GC_11_17 b_11 NI_11 NS_17 0 -8.7354411997277704e-07
GC_11_18 b_11 NI_11 NS_18 0 9.7910845687819833e-08
GC_11_19 b_11 NI_11 NS_19 0 2.5713356278347616e-06
GC_11_20 b_11 NI_11 NS_20 0 -1.1143656760289906e-06
GC_11_21 b_11 NI_11 NS_21 0 -3.9892768220408415e-06
GC_11_22 b_11 NI_11 NS_22 0 -2.3994165281216005e-07
GC_11_23 b_11 NI_11 NS_23 0 1.2120544439697012e-08
GC_11_24 b_11 NI_11 NS_24 0 1.6053768102518516e-06
GC_11_25 b_11 NI_11 NS_25 0 -8.3045108079706851e-07
GC_11_26 b_11 NI_11 NS_26 0 -2.6088618446164441e-06
GC_11_27 b_11 NI_11 NS_27 0 -7.8261801358233647e-07
GC_11_28 b_11 NI_11 NS_28 0 1.4932820164380928e-06
GC_11_29 b_11 NI_11 NS_29 0 5.8174617884686882e-07
GC_11_30 b_11 NI_11 NS_30 0 -3.0275241142011333e-06
GC_11_31 b_11 NI_11 NS_31 0 -1.4471017856049872e-06
GC_11_32 b_11 NI_11 NS_32 0 2.5662003663756112e-06
GC_11_33 b_11 NI_11 NS_33 0 2.3925611709944086e-07
GC_11_34 b_11 NI_11 NS_34 0 1.2705123408307748e-06
GC_11_35 b_11 NI_11 NS_35 0 -6.9731593333334682e-07
GC_11_36 b_11 NI_11 NS_36 0 -1.1692999891687036e-06
GC_11_37 b_11 NI_11 NS_37 0 -5.8078326393000885e-08
GC_11_38 b_11 NI_11 NS_38 0 1.0861778267997847e-06
GC_11_39 b_11 NI_11 NS_39 0 -6.5276876328535746e-07
GC_11_40 b_11 NI_11 NS_40 0 -7.6713718649202940e-07
GC_11_41 b_11 NI_11 NS_41 0 -5.1252565493483295e-07
GC_11_42 b_11 NI_11 NS_42 0 1.1060716118469100e-06
GC_11_43 b_11 NI_11 NS_43 0 4.5034309802113077e-08
GC_11_44 b_11 NI_11 NS_44 0 -8.8826750259659145e-07
GC_11_45 b_11 NI_11 NS_45 0 -9.1170815607599308e-07
GC_11_46 b_11 NI_11 NS_46 0 1.0678781262246857e-06
GC_11_47 b_11 NI_11 NS_47 0 -1.1157805952305604e-07
GC_11_48 b_11 NI_11 NS_48 0 7.9119417002203291e-09
GC_11_49 b_11 NI_11 NS_49 0 -3.3924071482295499e-07
GC_11_50 b_11 NI_11 NS_50 0 1.0187664903525483e-06
GC_11_51 b_11 NI_11 NS_51 0 -9.8123095564665937e-08
GC_11_52 b_11 NI_11 NS_52 0 1.1222916177946031e-07
GC_11_53 b_11 NI_11 NS_53 0 -3.0038773289993305e-07
GC_11_54 b_11 NI_11 NS_54 0 1.0059083840470873e-06
GC_11_55 b_11 NI_11 NS_55 0 8.0898406716459302e-08
GC_11_56 b_11 NI_11 NS_56 0 1.6439248668201994e-07
GC_11_57 b_11 NI_11 NS_57 0 -7.9032990225881168e-08
GC_11_58 b_11 NI_11 NS_58 0 1.1304512681921052e-06
GC_11_59 b_11 NI_11 NS_59 0 7.8465118504263872e-07
GC_11_60 b_11 NI_11 NS_60 0 -9.7827390756301675e-09
GC_11_61 b_11 NI_11 NS_61 0 8.4849744427490190e-08
GC_11_62 b_11 NI_11 NS_62 0 8.2101101485749210e-07
GC_11_63 b_11 NI_11 NS_63 0 3.1725538645840096e-07
GC_11_64 b_11 NI_11 NS_64 0 -1.9311000217618422e-07
GC_11_65 b_11 NI_11 NS_65 0 1.9073676037172115e-07
GC_11_66 b_11 NI_11 NS_66 0 1.0069326472031314e-06
GC_11_67 b_11 NI_11 NS_67 0 7.9531979620802171e-07
GC_11_68 b_11 NI_11 NS_68 0 -8.1781879092168482e-07
GC_11_69 b_11 NI_11 NS_69 0 3.2999049945324142e-07
GC_11_70 b_11 NI_11 NS_70 0 5.3261479983676193e-07
GC_11_71 b_11 NI_11 NS_71 0 -5.5976464117050801e-09
GC_11_72 b_11 NI_11 NS_72 0 -5.5297834270144518e-07
GC_11_73 b_11 NI_11 NS_73 0 4.5646401315401706e-07
GC_11_74 b_11 NI_11 NS_74 0 7.5300361161787274e-07
GC_11_75 b_11 NI_11 NS_75 0 -9.7909721140035763e-09
GC_11_76 b_11 NI_11 NS_76 0 -1.1014051657417054e-06
GC_11_77 b_11 NI_11 NS_77 0 3.1840348298026744e-07
GC_11_78 b_11 NI_11 NS_78 0 1.0304780535832043e-07
GC_11_79 b_11 NI_11 NS_79 0 -3.9308689112672871e-07
GC_11_80 b_11 NI_11 NS_80 0 -2.5353730158931633e-07
GC_11_81 b_11 NI_11 NS_81 0 1.4515571478538346e-12
GC_11_82 b_11 NI_11 NS_82 0 3.4002188453955795e-12
GC_11_83 b_11 NI_11 NS_83 0 3.9032029330323289e-07
GC_11_84 b_11 NI_11 NS_84 0 2.2951833192143829e-07
GC_11_85 b_11 NI_11 NS_85 0 1.1980287161845008e-07
GC_11_86 b_11 NI_11 NS_86 0 3.5450126356735658e-08
GC_11_87 b_11 NI_11 NS_87 0 -2.7884548114104126e-07
GC_11_88 b_11 NI_11 NS_88 0 -1.0897739543940669e-07
GC_11_89 b_11 NI_11 NS_89 0 3.2156248411830503e-07
GC_11_90 b_11 NI_11 NS_90 0 6.8215246434227190e-08
GC_11_91 b_11 NI_11 NS_91 0 -3.5585231482699392e-07
GC_11_92 b_11 NI_11 NS_92 0 -4.5136759852891159e-07
GC_11_93 b_11 NI_11 NS_93 0 -1.0584805229259524e-11
GC_11_94 b_11 NI_11 NS_94 0 3.2224294609399470e-10
GC_11_95 b_11 NI_11 NS_95 0 1.8885858120686278e-07
GC_11_96 b_11 NI_11 NS_96 0 -1.9034151001852519e-07
GC_11_97 b_11 NI_11 NS_97 0 -7.7178512974942449e-08
GC_11_98 b_11 NI_11 NS_98 0 3.9129207523996657e-07
GC_11_99 b_11 NI_11 NS_99 0 -1.7579593363189687e-07
GC_11_100 b_11 NI_11 NS_100 0 6.2408030812996823e-08
GC_11_101 b_11 NI_11 NS_101 0 -5.3348876240287201e-07
GC_11_102 b_11 NI_11 NS_102 0 -2.6042869717021598e-07
GC_11_103 b_11 NI_11 NS_103 0 5.9194248093414513e-08
GC_11_104 b_11 NI_11 NS_104 0 2.3071610751678615e-08
GC_11_105 b_11 NI_11 NS_105 0 -3.6617554794634466e-07
GC_11_106 b_11 NI_11 NS_106 0 6.6093642204292523e-08
GC_11_107 b_11 NI_11 NS_107 0 1.0697471657171372e-07
GC_11_108 b_11 NI_11 NS_108 0 3.2656969951425695e-07
GC_11_109 b_11 NI_11 NS_109 0 -2.9911161707579539e-05
GC_11_110 b_11 NI_11 NS_110 0 1.1048132847921431e-11
GC_11_111 b_11 NI_11 NS_111 0 -3.3938051292743052e-11
GC_11_112 b_11 NI_11 NS_112 0 2.1481719843878497e-10
GC_11_113 b_11 NI_11 NS_113 0 -4.0868881292063674e-07
GC_11_114 b_11 NI_11 NS_114 0 -2.7774303279418284e-07
GC_11_115 b_11 NI_11 NS_115 0 -1.0550552681507772e-07
GC_11_116 b_11 NI_11 NS_116 0 5.6498379471847883e-07
GC_11_117 b_11 NI_11 NS_117 0 2.3968440168894882e-07
GC_11_118 b_11 NI_11 NS_118 0 1.4051825293880747e-06
GC_11_119 b_11 NI_11 NS_119 0 1.1112320351204262e-06
GC_11_120 b_11 NI_11 NS_120 0 -3.7354234343081379e-07
GC_11_121 b_11 NI_11 NS_121 0 6.7789966394659304e-07
GC_11_122 b_11 NI_11 NS_122 0 -2.0311523095445120e-06
GC_11_123 b_11 NI_11 NS_123 0 -6.4633558429412740e-07
GC_11_124 b_11 NI_11 NS_124 0 2.8079859852993205e-07
GC_11_125 b_11 NI_11 NS_125 0 1.0005711183277326e-06
GC_11_126 b_11 NI_11 NS_126 0 6.6400923777408325e-07
GC_11_127 b_11 NI_11 NS_127 0 3.8996124028758335e-06
GC_11_128 b_11 NI_11 NS_128 0 -3.7318011745422440e-06
GC_11_129 b_11 NI_11 NS_129 0 -5.6020141045821143e-06
GC_11_130 b_11 NI_11 NS_130 0 -3.8667583425199053e-06
GC_11_131 b_11 NI_11 NS_131 0 -9.1897809855672476e-07
GC_11_132 b_11 NI_11 NS_132 0 -2.0469360699519703e-06
GC_11_133 b_11 NI_11 NS_133 0 -1.3607680613791318e-05
GC_11_134 b_11 NI_11 NS_134 0 5.3832281349953715e-06
GC_11_135 b_11 NI_11 NS_135 0 -5.4034744042827497e-07
GC_11_136 b_11 NI_11 NS_136 0 1.8948094118119446e-06
GC_11_137 b_11 NI_11 NS_137 0 7.8102753208278756e-07
GC_11_138 b_11 NI_11 NS_138 0 1.9317332309021315e-05
GC_11_139 b_11 NI_11 NS_139 0 2.7701905865921138e-06
GC_11_140 b_11 NI_11 NS_140 0 -4.5964446365456098e-06
GC_11_141 b_11 NI_11 NS_141 0 1.4650389818155038e-06
GC_11_142 b_11 NI_11 NS_142 0 1.7125870602984472e-06
GC_11_143 b_11 NI_11 NS_143 0 5.3187248233344471e-06
GC_11_144 b_11 NI_11 NS_144 0 -2.2434174196270743e-06
GC_11_145 b_11 NI_11 NS_145 0 -4.1230615283114677e-07
GC_11_146 b_11 NI_11 NS_146 0 -8.1329353195240517e-07
GC_11_147 b_11 NI_11 NS_147 0 -2.0580558829392029e-06
GC_11_148 b_11 NI_11 NS_148 0 2.3269565748775576e-06
GC_11_149 b_11 NI_11 NS_149 0 -3.1364385036869037e-08
GC_11_150 b_11 NI_11 NS_150 0 1.2404834449775856e-06
GC_11_151 b_11 NI_11 NS_151 0 5.2823841922837669e-06
GC_11_152 b_11 NI_11 NS_152 0 5.9487379870582142e-06
GC_11_153 b_11 NI_11 NS_153 0 1.4530423712733087e-06
GC_11_154 b_11 NI_11 NS_154 0 -1.0228754146655851e-06
GC_11_155 b_11 NI_11 NS_155 0 1.1373660218386645e-07
GC_11_156 b_11 NI_11 NS_156 0 -4.7317199345628651e-08
GC_11_157 b_11 NI_11 NS_157 0 5.0717122606256377e-07
GC_11_158 b_11 NI_11 NS_158 0 7.4710285770137483e-07
GC_11_159 b_11 NI_11 NS_159 0 6.0612402040997282e-06
GC_11_160 b_11 NI_11 NS_160 0 4.9609741574904484e-07
GC_11_161 b_11 NI_11 NS_161 0 5.5847017534204021e-07
GC_11_162 b_11 NI_11 NS_162 0 -8.6793655509620613e-07
GC_11_163 b_11 NI_11 NS_163 0 -1.2621092861774065e-07
GC_11_164 b_11 NI_11 NS_164 0 -3.6192940669965447e-08
GC_11_165 b_11 NI_11 NS_165 0 6.7933528785878531e-07
GC_11_166 b_11 NI_11 NS_166 0 8.5069551298371271e-07
GC_11_167 b_11 NI_11 NS_167 0 4.7901342638046292e-06
GC_11_168 b_11 NI_11 NS_168 0 -1.9393531690170409e-06
GC_11_169 b_11 NI_11 NS_169 0 1.3625248623455341e-07
GC_11_170 b_11 NI_11 NS_170 0 -7.2246165135831387e-07
GC_11_171 b_11 NI_11 NS_171 0 -1.2136585834153347e-07
GC_11_172 b_11 NI_11 NS_172 0 1.4889792786772936e-07
GC_11_173 b_11 NI_11 NS_173 0 9.4361092978349277e-07
GC_11_174 b_11 NI_11 NS_174 0 7.7801140462892744e-07
GC_11_175 b_11 NI_11 NS_175 0 2.7633780059955155e-06
GC_11_176 b_11 NI_11 NS_176 0 -3.0197947455419984e-06
GC_11_177 b_11 NI_11 NS_177 0 -1.0372376210307649e-07
GC_11_178 b_11 NI_11 NS_178 0 -4.8471641262753846e-07
GC_11_179 b_11 NI_11 NS_179 0 8.9036105170688641e-08
GC_11_180 b_11 NI_11 NS_180 0 2.0200935518005624e-07
GC_11_181 b_11 NI_11 NS_181 0 1.3142787194827381e-06
GC_11_182 b_11 NI_11 NS_182 0 5.1190872831500703e-07
GC_11_183 b_11 NI_11 NS_183 0 6.6544904428229781e-07
GC_11_184 b_11 NI_11 NS_184 0 -2.7719655368978234e-06
GC_11_185 b_11 NI_11 NS_185 0 -1.6530791850499001e-07
GC_11_186 b_11 NI_11 NS_186 0 -1.3965379194367027e-07
GC_11_187 b_11 NI_11 NS_187 0 2.2791458354158658e-07
GC_11_188 b_11 NI_11 NS_188 0 2.3001717342262494e-08
GC_11_189 b_11 NI_11 NS_189 0 1.6157030185664873e-12
GC_11_190 b_11 NI_11 NS_190 0 -6.1868750422431226e-12
GC_11_191 b_11 NI_11 NS_191 0 9.8141713910577309e-07
GC_11_192 b_11 NI_11 NS_192 0 -2.6421990134292143e-07
GC_11_193 b_11 NI_11 NS_193 0 -2.6951743036423674e-08
GC_11_194 b_11 NI_11 NS_194 0 4.9063424516103392e-08
GC_11_195 b_11 NI_11 NS_195 0 2.6324977286028493e-07
GC_11_196 b_11 NI_11 NS_196 0 1.1274488173899972e-08
GC_11_197 b_11 NI_11 NS_197 0 8.3346104132126590e-07
GC_11_198 b_11 NI_11 NS_198 0 -1.5917973842263620e-07
GC_11_199 b_11 NI_11 NS_199 0 -6.3279065483576143e-08
GC_11_200 b_11 NI_11 NS_200 0 -1.0953395636559647e-06
GC_11_201 b_11 NI_11 NS_201 0 7.6569695851814386e-11
GC_11_202 b_11 NI_11 NS_202 0 -1.9331167472843489e-10
GC_11_203 b_11 NI_11 NS_203 0 6.8054874625314998e-07
GC_11_204 b_11 NI_11 NS_204 0 -4.3046093325857497e-07
GC_11_205 b_11 NI_11 NS_205 0 4.2750322639586565e-07
GC_11_206 b_11 NI_11 NS_206 0 1.6125226812403118e-07
GC_11_207 b_11 NI_11 NS_207 0 1.4001449673412343e-07
GC_11_208 b_11 NI_11 NS_208 0 -8.2569532692617981e-08
GC_11_209 b_11 NI_11 NS_209 0 -1.4342614803327999e-07
GC_11_210 b_11 NI_11 NS_210 0 -6.7675424117174636e-07
GC_11_211 b_11 NI_11 NS_211 0 2.4259828028390458e-08
GC_11_212 b_11 NI_11 NS_212 0 2.3629852973774312e-07
GC_11_213 b_11 NI_11 NS_213 0 3.3308573555303354e-07
GC_11_214 b_11 NI_11 NS_214 0 -5.5341486546891648e-08
GC_11_215 b_11 NI_11 NS_215 0 4.0226658212475853e-07
GC_11_216 b_11 NI_11 NS_216 0 2.2651269420919065e-07
GC_11_217 b_11 NI_11 NS_217 0 8.5535290096952099e-06
GC_11_218 b_11 NI_11 NS_218 0 3.7642528564441888e-12
GC_11_219 b_11 NI_11 NS_219 0 -7.8551930225641939e-11
GC_11_220 b_11 NI_11 NS_220 0 2.5470418010871218e-09
GC_11_221 b_11 NI_11 NS_221 0 1.5926580938613825e-08
GC_11_222 b_11 NI_11 NS_222 0 -8.5340732147958964e-08
GC_11_223 b_11 NI_11 NS_223 0 -2.5044501709378650e-07
GC_11_224 b_11 NI_11 NS_224 0 2.6988972840210725e-07
GC_11_225 b_11 NI_11 NS_225 0 7.4472050542182155e-07
GC_11_226 b_11 NI_11 NS_226 0 -2.8257742894721542e-07
GC_11_227 b_11 NI_11 NS_227 0 -9.7076232541472544e-07
GC_11_228 b_11 NI_11 NS_228 0 -2.4180541782182976e-07
GC_11_229 b_11 NI_11 NS_229 0 1.0253001983157930e-06
GC_11_230 b_11 NI_11 NS_230 0 4.0598744125163420e-07
GC_11_231 b_11 NI_11 NS_231 0 -1.2043552275546844e-07
GC_11_232 b_11 NI_11 NS_232 0 -2.7435486875136957e-07
GC_11_233 b_11 NI_11 NS_233 0 1.1179341566766751e-07
GC_11_234 b_11 NI_11 NS_234 0 -5.1154224541160299e-07
GC_11_235 b_11 NI_11 NS_235 0 -2.0930620661740532e-06
GC_11_236 b_11 NI_11 NS_236 0 8.5810262738141871e-07
GC_11_237 b_11 NI_11 NS_237 0 2.4408884888672626e-06
GC_11_238 b_11 NI_11 NS_238 0 -5.9923565079909285e-07
GC_11_239 b_11 NI_11 NS_239 0 -6.6143701309654581e-07
GC_11_240 b_11 NI_11 NS_240 0 -1.4026138040464731e-06
GC_11_241 b_11 NI_11 NS_241 0 4.2548592073409683e-07
GC_11_242 b_11 NI_11 NS_242 0 1.8523050649482303e-06
GC_11_243 b_11 NI_11 NS_243 0 -2.7461886132083222e-08
GC_11_244 b_11 NI_11 NS_244 0 -1.3270320331054105e-06
GC_11_245 b_11 NI_11 NS_245 0 -6.3828699998797494e-07
GC_11_246 b_11 NI_11 NS_246 0 2.5986442701086958e-06
GC_11_247 b_11 NI_11 NS_247 0 4.5949664081860429e-07
GC_11_248 b_11 NI_11 NS_248 0 -2.2490726539231804e-06
GC_11_249 b_11 NI_11 NS_249 0 -8.0030288893925862e-07
GC_11_250 b_11 NI_11 NS_250 0 -9.3521757893781803e-07
GC_11_251 b_11 NI_11 NS_251 0 3.5980072295991904e-07
GC_11_252 b_11 NI_11 NS_252 0 9.1582444886938376e-07
GC_11_253 b_11 NI_11 NS_253 0 -5.5704123332014562e-07
GC_11_254 b_11 NI_11 NS_254 0 -7.2806117483588784e-07
GC_11_255 b_11 NI_11 NS_255 0 4.7834203379101458e-07
GC_11_256 b_11 NI_11 NS_256 0 7.4258403393576302e-07
GC_11_257 b_11 NI_11 NS_257 0 -1.7303768964479531e-07
GC_11_258 b_11 NI_11 NS_258 0 -8.8058544293929973e-07
GC_11_259 b_11 NI_11 NS_259 0 -3.3837669292391448e-07
GC_11_260 b_11 NI_11 NS_260 0 1.1624991298721742e-06
GC_11_261 b_11 NI_11 NS_261 0 2.5595323510458913e-07
GC_11_262 b_11 NI_11 NS_262 0 -8.4667910868411739e-07
GC_11_263 b_11 NI_11 NS_263 0 -6.4574675279116858e-08
GC_11_264 b_11 NI_11 NS_264 0 6.7761705799691267e-08
GC_11_265 b_11 NI_11 NS_265 0 -2.5919670559911154e-07
GC_11_266 b_11 NI_11 NS_266 0 -5.5152744201854817e-07
GC_11_267 b_11 NI_11 NS_267 0 1.8905464347314762e-07
GC_11_268 b_11 NI_11 NS_268 0 7.1901969727640559e-07
GC_11_269 b_11 NI_11 NS_269 0 -7.9602560116447396e-08
GC_11_270 b_11 NI_11 NS_270 0 -6.3772380536086283e-07
GC_11_271 b_11 NI_11 NS_271 0 1.0329800214060183e-07
GC_11_272 b_11 NI_11 NS_272 0 1.0426218353444898e-07
GC_11_273 b_11 NI_11 NS_273 0 -2.9062616904547379e-07
GC_11_274 b_11 NI_11 NS_274 0 -5.9569102184132385e-07
GC_11_275 b_11 NI_11 NS_275 0 1.6437653502605574e-07
GC_11_276 b_11 NI_11 NS_276 0 2.3048497085709613e-07
GC_11_277 b_11 NI_11 NS_277 0 -2.5683232151565874e-07
GC_11_278 b_11 NI_11 NS_278 0 -5.1013987481336541e-07
GC_11_279 b_11 NI_11 NS_279 0 4.9680094279147830e-08
GC_11_280 b_11 NI_11 NS_280 0 -5.0623943625274384e-08
GC_11_281 b_11 NI_11 NS_281 0 -3.6842312906923460e-07
GC_11_282 b_11 NI_11 NS_282 0 -5.6019329737697475e-07
GC_11_283 b_11 NI_11 NS_283 0 -2.3359358698825428e-07
GC_11_284 b_11 NI_11 NS_284 0 2.0119413778834568e-08
GC_11_285 b_11 NI_11 NS_285 0 -4.3463044515080601e-07
GC_11_286 b_11 NI_11 NS_286 0 -3.4260327162895406e-07
GC_11_287 b_11 NI_11 NS_287 0 -1.2394298039170350e-07
GC_11_288 b_11 NI_11 NS_288 0 1.6157722068219209e-08
GC_11_289 b_11 NI_11 NS_289 0 -5.6455860657062528e-07
GC_11_290 b_11 NI_11 NS_290 0 -4.4144299263175144e-07
GC_11_291 b_11 NI_11 NS_291 0 -3.1825741658378627e-07
GC_11_292 b_11 NI_11 NS_292 0 3.1675254707177366e-07
GC_11_293 b_11 NI_11 NS_293 0 -5.0108235072919932e-07
GC_11_294 b_11 NI_11 NS_294 0 3.6711553667920874e-08
GC_11_295 b_11 NI_11 NS_295 0 -1.0041271910740457e-08
GC_11_296 b_11 NI_11 NS_296 0 6.2080184173308675e-08
GC_11_297 b_11 NI_11 NS_297 0 -3.2608850625598472e-12
GC_11_298 b_11 NI_11 NS_298 0 3.1978319502270015e-12
GC_11_299 b_11 NI_11 NS_299 0 -5.7750173960202934e-07
GC_11_300 b_11 NI_11 NS_300 0 4.5921289929588829e-08
GC_11_301 b_11 NI_11 NS_301 0 -2.9018156093857848e-07
GC_11_302 b_11 NI_11 NS_302 0 1.1752544804934037e-07
GC_11_303 b_11 NI_11 NS_303 0 -5.6680341832373164e-09
GC_11_304 b_11 NI_11 NS_304 0 -6.8755107841904587e-08
GC_11_305 b_11 NI_11 NS_305 0 -6.6097127022936146e-07
GC_11_306 b_11 NI_11 NS_306 0 1.3969830360393153e-07
GC_11_307 b_11 NI_11 NS_307 0 2.9822605481011705e-08
GC_11_308 b_11 NI_11 NS_308 0 1.2499650111728344e-07
GC_11_309 b_11 NI_11 NS_309 0 -6.1663280905059968e-11
GC_11_310 b_11 NI_11 NS_310 0 1.2835970580533626e-10
GC_11_311 b_11 NI_11 NS_311 0 -3.4930744681812283e-08
GC_11_312 b_11 NI_11 NS_312 0 1.9717738078563629e-07
GC_11_313 b_11 NI_11 NS_313 0 -3.6700067733485956e-07
GC_11_314 b_11 NI_11 NS_314 0 -4.4689709321370807e-08
GC_11_315 b_11 NI_11 NS_315 0 -1.8607422024236999e-07
GC_11_316 b_11 NI_11 NS_316 0 -2.7291584282352903e-09
GC_11_317 b_11 NI_11 NS_317 0 1.9304455733084556e-07
GC_11_318 b_11 NI_11 NS_318 0 8.1847720738231548e-08
GC_11_319 b_11 NI_11 NS_319 0 -2.6597640694369009e-07
GC_11_320 b_11 NI_11 NS_320 0 3.1322685401290108e-07
GC_11_321 b_11 NI_11 NS_321 0 1.2554885296802218e-07
GC_11_322 b_11 NI_11 NS_322 0 -1.4412638980752234e-07
GC_11_323 b_11 NI_11 NS_323 0 -5.8147603231669395e-08
GC_11_324 b_11 NI_11 NS_324 0 2.3784859634074377e-07
GC_11_325 b_11 NI_11 NS_325 0 -6.4297437901002878e-05
GC_11_326 b_11 NI_11 NS_326 0 3.5514238498082589e-12
GC_11_327 b_11 NI_11 NS_327 0 5.0206522290172771e-11
GC_11_328 b_11 NI_11 NS_328 0 -1.5827704276859361e-09
GC_11_329 b_11 NI_11 NS_329 0 -1.0722829845077973e-06
GC_11_330 b_11 NI_11 NS_330 0 -1.0608508874111980e-06
GC_11_331 b_11 NI_11 NS_331 0 4.1036061523746122e-07
GC_11_332 b_11 NI_11 NS_332 0 3.5893547448321589e-07
GC_11_333 b_11 NI_11 NS_333 0 -2.2645837197285659e-06
GC_11_334 b_11 NI_11 NS_334 0 2.1075511831342365e-06
GC_11_335 b_11 NI_11 NS_335 0 -2.5340144402830408e-06
GC_11_336 b_11 NI_11 NS_336 0 -1.2433713995259555e-06
GC_11_337 b_11 NI_11 NS_337 0 1.3995724520706924e-06
GC_11_338 b_11 NI_11 NS_338 0 1.0022095515951407e-06
GC_11_339 b_11 NI_11 NS_339 0 -1.1248422783415153e-06
GC_11_340 b_11 NI_11 NS_340 0 1.3421230198462376e-06
GC_11_341 b_11 NI_11 NS_341 0 7.2528837464812529e-07
GC_11_342 b_11 NI_11 NS_342 0 3.0434879858904896e-06
GC_11_343 b_11 NI_11 NS_343 0 -2.8542782669852104e-06
GC_11_344 b_11 NI_11 NS_344 0 4.6950421276918474e-07
GC_11_345 b_11 NI_11 NS_345 0 3.6961230921458044e-06
GC_11_346 b_11 NI_11 NS_346 0 -2.0128601172650411e-06
GC_11_347 b_11 NI_11 NS_347 0 -1.9025439131850111e-07
GC_11_348 b_11 NI_11 NS_348 0 2.5688281124282109e-06
GC_11_349 b_11 NI_11 NS_349 0 -4.0608163856820256e-06
GC_11_350 b_11 NI_11 NS_350 0 4.8420473864247660e-06
GC_11_351 b_11 NI_11 NS_351 0 6.4549017836934972e-07
GC_11_352 b_11 NI_11 NS_352 0 -1.5900720072032835e-06
GC_11_353 b_11 NI_11 NS_353 0 4.6200375869788088e-06
GC_11_354 b_11 NI_11 NS_354 0 9.9425459740750397e-06
GC_11_355 b_11 NI_11 NS_355 0 -1.1566840538016195e-07
GC_11_356 b_11 NI_11 NS_356 0 5.2796972049090199e-07
GC_11_357 b_11 NI_11 NS_357 0 -6.9198325102783251e-09
GC_11_358 b_11 NI_11 NS_358 0 -7.8936930054482656e-07
GC_11_359 b_11 NI_11 NS_359 0 5.3542029134805008e-06
GC_11_360 b_11 NI_11 NS_360 0 4.9601481586848411e-07
GC_11_361 b_11 NI_11 NS_361 0 8.4752671013929017e-07
GC_11_362 b_11 NI_11 NS_362 0 1.9215332074473240e-06
GC_11_363 b_11 NI_11 NS_363 0 3.1631193063712745e-08
GC_11_364 b_11 NI_11 NS_364 0 1.1340878556728844e-06
GC_11_365 b_11 NI_11 NS_365 0 5.8569823706211655e-07
GC_11_366 b_11 NI_11 NS_366 0 -1.1142341622619806e-06
GC_11_367 b_11 NI_11 NS_367 0 5.8308842629805595e-06
GC_11_368 b_11 NI_11 NS_368 0 4.0738797072866836e-06
GC_11_369 b_11 NI_11 NS_369 0 6.0565171129154814e-07
GC_11_370 b_11 NI_11 NS_370 0 8.6240411265903439e-07
GC_11_371 b_11 NI_11 NS_371 0 1.9671287350791000e-07
GC_11_372 b_11 NI_11 NS_372 0 2.4104682123336977e-07
GC_11_373 b_11 NI_11 NS_373 0 8.4506773754518199e-07
GC_11_374 b_11 NI_11 NS_374 0 -6.7479188876989936e-07
GC_11_375 b_11 NI_11 NS_375 0 6.6692136892953642e-06
GC_11_376 b_11 NI_11 NS_376 0 7.5282682322909765e-07
GC_11_377 b_11 NI_11 NS_377 0 7.7512335686447369e-07
GC_11_378 b_11 NI_11 NS_378 0 7.5176122584223821e-07
GC_11_379 b_11 NI_11 NS_379 0 6.6485231737631378e-07
GC_11_380 b_11 NI_11 NS_380 0 -6.6043462020637097e-08
GC_11_381 b_11 NI_11 NS_381 0 8.7117401296082778e-07
GC_11_382 b_11 NI_11 NS_382 0 -6.4327591127592566e-07
GC_11_383 b_11 NI_11 NS_383 0 5.7782970224983313e-06
GC_11_384 b_11 NI_11 NS_384 0 -1.5930787639181261e-06
GC_11_385 b_11 NI_11 NS_385 0 8.2495349562710594e-07
GC_11_386 b_11 NI_11 NS_386 0 5.6931957780991138e-07
GC_11_387 b_11 NI_11 NS_387 0 6.2573082926731346e-07
GC_11_388 b_11 NI_11 NS_388 0 -5.5367558781510452e-07
GC_11_389 b_11 NI_11 NS_389 0 9.3726424309104736e-07
GC_11_390 b_11 NI_11 NS_390 0 -4.4873357062558238e-07
GC_11_391 b_11 NI_11 NS_391 0 3.9054758422271746e-06
GC_11_392 b_11 NI_11 NS_392 0 -2.9926293450081277e-06
GC_11_393 b_11 NI_11 NS_393 0 8.9723586115500261e-07
GC_11_394 b_11 NI_11 NS_394 0 3.2914679275627296e-07
GC_11_395 b_11 NI_11 NS_395 0 2.1534418817498623e-07
GC_11_396 b_11 NI_11 NS_396 0 -7.9633368901714842e-07
GC_11_397 b_11 NI_11 NS_397 0 1.1591902965953778e-06
GC_11_398 b_11 NI_11 NS_398 0 -3.2770346759434548e-07
GC_11_399 b_11 NI_11 NS_399 0 1.6782755522506130e-06
GC_11_400 b_11 NI_11 NS_400 0 -3.0911767505389314e-06
GC_11_401 b_11 NI_11 NS_401 0 7.9264445503514927e-07
GC_11_402 b_11 NI_11 NS_402 0 -1.0570164290071468e-07
GC_11_403 b_11 NI_11 NS_403 0 -1.9831483591368102e-07
GC_11_404 b_11 NI_11 NS_404 0 -4.0881300698224303e-07
GC_11_405 b_11 NI_11 NS_405 0 8.5891446676145302e-12
GC_11_406 b_11 NI_11 NS_406 0 -1.5739889036957298e-11
GC_11_407 b_11 NI_11 NS_407 0 8.3767177938929471e-07
GC_11_408 b_11 NI_11 NS_408 0 -5.9585018647331949e-07
GC_11_409 b_11 NI_11 NS_409 0 4.9537203700649267e-07
GC_11_410 b_11 NI_11 NS_410 0 -3.5566005680104102e-08
GC_11_411 b_11 NI_11 NS_411 0 1.6374839311928927e-08
GC_11_412 b_11 NI_11 NS_412 0 -8.9213583652432756e-08
GC_11_413 b_11 NI_11 NS_413 0 5.2071533656906817e-07
GC_11_414 b_11 NI_11 NS_414 0 -1.9287830533793234e-08
GC_11_415 b_11 NI_11 NS_415 0 7.0590791211509430e-07
GC_11_416 b_11 NI_11 NS_416 0 -1.5618072848432789e-06
GC_11_417 b_11 NI_11 NS_417 0 4.0957995829789864e-10
GC_11_418 b_11 NI_11 NS_418 0 -5.8094713515743367e-10
GC_11_419 b_11 NI_11 NS_419 0 1.0094261239058910e-06
GC_11_420 b_11 NI_11 NS_420 0 -2.7418451570183223e-07
GC_11_421 b_11 NI_11 NS_421 0 3.5391575331011913e-07
GC_11_422 b_11 NI_11 NS_422 0 -1.7487895512836163e-07
GC_11_423 b_11 NI_11 NS_423 0 2.5449986409532842e-07
GC_11_424 b_11 NI_11 NS_424 0 2.6674221769231540e-08
GC_11_425 b_11 NI_11 NS_425 0 1.0861097661948931e-06
GC_11_426 b_11 NI_11 NS_426 0 -1.1751152210527382e-06
GC_11_427 b_11 NI_11 NS_427 0 6.5444234658491502e-07
GC_11_428 b_11 NI_11 NS_428 0 -3.3449257800913166e-07
GC_11_429 b_11 NI_11 NS_429 0 -2.1290010454039099e-07
GC_11_430 b_11 NI_11 NS_430 0 -9.8626427894762261e-08
GC_11_431 b_11 NI_11 NS_431 0 7.5675693958716067e-07
GC_11_432 b_11 NI_11 NS_432 0 3.2207292927148206e-07
GC_11_433 b_11 NI_11 NS_433 0 4.9622882787156384e-05
GC_11_434 b_11 NI_11 NS_434 0 3.6303600156571463e-12
GC_11_435 b_11 NI_11 NS_435 0 -4.1065549478614434e-12
GC_11_436 b_11 NI_11 NS_436 0 9.4552808742662489e-10
GC_11_437 b_11 NI_11 NS_437 0 -4.5592728708232096e-08
GC_11_438 b_11 NI_11 NS_438 0 2.5302100132000164e-07
GC_11_439 b_11 NI_11 NS_439 0 2.5930073472299552e-07
GC_11_440 b_11 NI_11 NS_440 0 4.0791655086969086e-07
GC_11_441 b_11 NI_11 NS_441 0 -1.3649528174905169e-07
GC_11_442 b_11 NI_11 NS_442 0 2.4393631439433393e-07
GC_11_443 b_11 NI_11 NS_443 0 7.8203509573192628e-07
GC_11_444 b_11 NI_11 NS_444 0 1.4417033179376424e-06
GC_11_445 b_11 NI_11 NS_445 0 1.0397082503838212e-06
GC_11_446 b_11 NI_11 NS_446 0 -5.2292447472922300e-07
GC_11_447 b_11 NI_11 NS_447 0 3.3637636171527303e-07
GC_11_448 b_11 NI_11 NS_448 0 8.8673917408017382e-07
GC_11_449 b_11 NI_11 NS_449 0 7.3264019038651572e-07
GC_11_450 b_11 NI_11 NS_450 0 -3.6972328883878880e-07
GC_11_451 b_11 NI_11 NS_451 0 4.3588547637149562e-06
GC_11_452 b_11 NI_11 NS_452 0 1.3805934521086804e-06
GC_11_453 b_11 NI_11 NS_453 0 -1.6438415195424687e-06
GC_11_454 b_11 NI_11 NS_454 0 -3.5789178768620875e-06
GC_11_455 b_11 NI_11 NS_455 0 2.4006556089394745e-07
GC_11_456 b_11 NI_11 NS_456 0 1.5509786147030545e-06
GC_11_457 b_11 NI_11 NS_457 0 2.9713800850411210e-06
GC_11_458 b_11 NI_11 NS_458 0 -4.7497990141087182e-06
GC_11_459 b_11 NI_11 NS_459 0 -7.7198179434637496e-07
GC_11_460 b_11 NI_11 NS_460 0 5.6526099645252183e-07
GC_11_461 b_11 NI_11 NS_461 0 5.5714198990255923e-06
GC_11_462 b_11 NI_11 NS_462 0 -5.8239750764943397e-06
GC_11_463 b_11 NI_11 NS_463 0 -3.3126921678249988e-06
GC_11_464 b_11 NI_11 NS_464 0 1.7946937549017728e-06
GC_11_465 b_11 NI_11 NS_465 0 8.6225842903552410e-07
GC_11_466 b_11 NI_11 NS_466 0 1.2280693091367326e-06
GC_11_467 b_11 NI_11 NS_467 0 1.5935582561200145e-06
GC_11_468 b_11 NI_11 NS_468 0 -4.1016190472119700e-06
GC_11_469 b_11 NI_11 NS_469 0 5.6918443162164791e-07
GC_11_470 b_11 NI_11 NS_470 0 1.9887015566480706e-07
GC_11_471 b_11 NI_11 NS_471 0 1.7374858153322994e-07
GC_11_472 b_11 NI_11 NS_472 0 -4.0365324601289513e-06
GC_11_473 b_11 NI_11 NS_473 0 -1.8756568644450529e-07
GC_11_474 b_11 NI_11 NS_474 0 1.6738463097983910e-07
GC_11_475 b_11 NI_11 NS_475 0 4.6371530286858279e-06
GC_11_476 b_11 NI_11 NS_476 0 -6.3342159582815935e-06
GC_11_477 b_11 NI_11 NS_477 0 -1.8279081944223418e-06
GC_11_478 b_11 NI_11 NS_478 0 -1.2891002214183870e-06
GC_11_479 b_11 NI_11 NS_479 0 1.3669284535156421e-06
GC_11_480 b_11 NI_11 NS_480 0 -1.1987253449247271e-06
GC_11_481 b_11 NI_11 NS_481 0 3.7640837927780634e-07
GC_11_482 b_11 NI_11 NS_482 0 -2.0979971433936187e-06
GC_11_483 b_11 NI_11 NS_483 0 -1.4883368417466387e-06
GC_11_484 b_11 NI_11 NS_484 0 -1.1766921777713626e-05
GC_11_485 b_11 NI_11 NS_485 0 -2.2685259448794451e-06
GC_11_486 b_11 NI_11 NS_486 0 -1.7028015921855590e-06
GC_11_487 b_11 NI_11 NS_487 0 -2.3846882858387197e-06
GC_11_488 b_11 NI_11 NS_488 0 -3.9900407805930374e-06
GC_11_489 b_11 NI_11 NS_489 0 -1.4877942094508706e-06
GC_11_490 b_11 NI_11 NS_490 0 -2.4193236661076112e-06
GC_11_491 b_11 NI_11 NS_491 0 -1.0718666766225755e-05
GC_11_492 b_11 NI_11 NS_492 0 -7.0858393718503260e-06
GC_11_493 b_11 NI_11 NS_493 0 -3.1913010058125985e-06
GC_11_494 b_11 NI_11 NS_494 0 -8.5705624233658506e-07
GC_11_495 b_11 NI_11 NS_495 0 -5.7484892881967566e-06
GC_11_496 b_11 NI_11 NS_496 0 -3.7009140035099367e-07
GC_11_497 b_11 NI_11 NS_497 0 -3.1247013239230615e-06
GC_11_498 b_11 NI_11 NS_498 0 -1.7467006971698380e-06
GC_11_499 b_11 NI_11 NS_499 0 -1.0620562918132085e-05
GC_11_500 b_11 NI_11 NS_500 0 3.3757038598658369e-06
GC_11_501 b_11 NI_11 NS_501 0 -3.6323500946349551e-06
GC_11_502 b_11 NI_11 NS_502 0 8.2990792999931142e-07
GC_11_503 b_11 NI_11 NS_503 0 -2.8726611817041039e-06
GC_11_504 b_11 NI_11 NS_504 0 3.9436375464279832e-06
GC_11_505 b_11 NI_11 NS_505 0 -4.3602279341257404e-06
GC_11_506 b_11 NI_11 NS_506 0 1.7215331639676934e-07
GC_11_507 b_11 NI_11 NS_507 0 -1.8596062245977610e-06
GC_11_508 b_11 NI_11 NS_508 0 7.2753444753164135e-06
GC_11_509 b_11 NI_11 NS_509 0 -1.5754108516182333e-06
GC_11_510 b_11 NI_11 NS_510 0 2.8117901311868006e-06
GC_11_511 b_11 NI_11 NS_511 0 9.3640991446373679e-07
GC_11_512 b_11 NI_11 NS_512 0 1.8342899553550661e-06
GC_11_513 b_11 NI_11 NS_513 0 -3.0126797300088598e-11
GC_11_514 b_11 NI_11 NS_514 0 -3.3795217410794132e-12
GC_11_515 b_11 NI_11 NS_515 0 -1.7324943137039587e-06
GC_11_516 b_11 NI_11 NS_516 0 2.1530117322134453e-06
GC_11_517 b_11 NI_11 NS_517 0 -3.2447797143416342e-07
GC_11_518 b_11 NI_11 NS_518 0 1.0585499699510950e-06
GC_11_519 b_11 NI_11 NS_519 0 1.4373513606786089e-07
GC_11_520 b_11 NI_11 NS_520 0 6.3907909761107501e-07
GC_11_521 b_11 NI_11 NS_521 0 -1.0432327218751568e-06
GC_11_522 b_11 NI_11 NS_522 0 1.2848490343861292e-06
GC_11_523 b_11 NI_11 NS_523 0 9.8805471319046219e-07
GC_11_524 b_11 NI_11 NS_524 0 1.8543066774958223e-06
GC_11_525 b_11 NI_11 NS_525 0 -1.5200210836308757e-09
GC_11_526 b_11 NI_11 NS_526 0 -7.6813237030151884e-10
GC_11_527 b_11 NI_11 NS_527 0 -4.6961215718338837e-07
GC_11_528 b_11 NI_11 NS_528 0 -2.3333868070758545e-08
GC_11_529 b_11 NI_11 NS_529 0 -3.1184749451633577e-07
GC_11_530 b_11 NI_11 NS_530 0 1.9127792178382423e-07
GC_11_531 b_11 NI_11 NS_531 0 -5.4919332832783691e-07
GC_11_532 b_11 NI_11 NS_532 0 1.5141534272166239e-07
GC_11_533 b_11 NI_11 NS_533 0 6.6185656069941749e-07
GC_11_534 b_11 NI_11 NS_534 0 8.3046362753867337e-07
GC_11_535 b_11 NI_11 NS_535 0 2.3283672177157386e-07
GC_11_536 b_11 NI_11 NS_536 0 7.0047496886630437e-07
GC_11_537 b_11 NI_11 NS_537 0 3.0952734196915788e-09
GC_11_538 b_11 NI_11 NS_538 0 -1.3231324142112723e-07
GC_11_539 b_11 NI_11 NS_539 0 -3.4727120514902818e-07
GC_11_540 b_11 NI_11 NS_540 0 2.9413081287928884e-07
GC_11_541 b_11 NI_11 NS_541 0 -9.0232958822447436e-05
GC_11_542 b_11 NI_11 NS_542 0 7.1467481412981950e-12
GC_11_543 b_11 NI_11 NS_543 0 -5.7273339924599885e-11
GC_11_544 b_11 NI_11 NS_544 0 3.3270946399318706e-10
GC_11_545 b_11 NI_11 NS_545 0 -1.5775940636582214e-06
GC_11_546 b_11 NI_11 NS_546 0 -1.5525976764956462e-06
GC_11_547 b_11 NI_11 NS_547 0 9.4591908790814787e-07
GC_11_548 b_11 NI_11 NS_548 0 7.1992430672776082e-07
GC_11_549 b_11 NI_11 NS_549 0 -2.7042603332488698e-06
GC_11_550 b_11 NI_11 NS_550 0 3.0432322761670964e-06
GC_11_551 b_11 NI_11 NS_551 0 -3.0477772176834282e-06
GC_11_552 b_11 NI_11 NS_552 0 -2.5663724414182445e-06
GC_11_553 b_11 NI_11 NS_553 0 1.5140825172942720e-06
GC_11_554 b_11 NI_11 NS_554 0 6.0867018694809266e-08
GC_11_555 b_11 NI_11 NS_555 0 -1.6616231581294326e-06
GC_11_556 b_11 NI_11 NS_556 0 1.7956744694072211e-06
GC_11_557 b_11 NI_11 NS_557 0 9.0473479384165556e-07
GC_11_558 b_11 NI_11 NS_558 0 4.1356157844988003e-06
GC_11_559 b_11 NI_11 NS_559 0 -4.2700514091212174e-06
GC_11_560 b_11 NI_11 NS_560 0 -2.0665758850166839e-06
GC_11_561 b_11 NI_11 NS_561 0 2.3210795955383609e-06
GC_11_562 b_11 NI_11 NS_562 0 -1.9750386438231130e-06
GC_11_563 b_11 NI_11 NS_563 0 -1.1664538130508150e-06
GC_11_564 b_11 NI_11 NS_564 0 3.2386767629894071e-06
GC_11_565 b_11 NI_11 NS_565 0 -8.4927506745991545e-06
GC_11_566 b_11 NI_11 NS_566 0 1.1257660829040442e-05
GC_11_567 b_11 NI_11 NS_567 0 1.2382795893328353e-06
GC_11_568 b_11 NI_11 NS_568 0 -1.6380387531913720e-06
GC_11_569 b_11 NI_11 NS_569 0 9.9626765032102678e-06
GC_11_570 b_11 NI_11 NS_570 0 1.7510982488004530e-05
GC_11_571 b_11 NI_11 NS_571 0 -6.2141816487791092e-07
GC_11_572 b_11 NI_11 NS_572 0 -5.7372126312971701e-07
GC_11_573 b_11 NI_11 NS_573 0 4.5338224715068441e-07
GC_11_574 b_11 NI_11 NS_574 0 -1.3531116996337299e-06
GC_11_575 b_11 NI_11 NS_575 0 7.0533250264044360e-06
GC_11_576 b_11 NI_11 NS_576 0 -2.6360793359115804e-07
GC_11_577 b_11 NI_11 NS_577 0 7.0541905670803150e-07
GC_11_578 b_11 NI_11 NS_578 0 2.9816718429036578e-06
GC_11_579 b_11 NI_11 NS_579 0 4.2391653745603082e-07
GC_11_580 b_11 NI_11 NS_580 0 2.9338710007094132e-06
GC_11_581 b_11 NI_11 NS_581 0 1.1537400576078313e-06
GC_11_582 b_11 NI_11 NS_582 0 -1.4005628041632435e-06
GC_11_583 b_11 NI_11 NS_583 0 9.4429358272955919e-06
GC_11_584 b_11 NI_11 NS_584 0 5.2402557332044533e-06
GC_11_585 b_11 NI_11 NS_585 0 5.8904435436093710e-07
GC_11_586 b_11 NI_11 NS_586 0 1.1278221302300017e-06
GC_11_587 b_11 NI_11 NS_587 0 5.5043726067740062e-08
GC_11_588 b_11 NI_11 NS_588 0 4.4723271984669972e-07
GC_11_589 b_11 NI_11 NS_589 0 1.2859226569548277e-06
GC_11_590 b_11 NI_11 NS_590 0 -8.4940678066574661e-07
GC_11_591 b_11 NI_11 NS_591 0 9.2174173445754635e-06
GC_11_592 b_11 NI_11 NS_592 0 6.4701247254571182e-07
GC_11_593 b_11 NI_11 NS_593 0 8.4642732474634886e-07
GC_11_594 b_11 NI_11 NS_594 0 1.4278802862336275e-06
GC_11_595 b_11 NI_11 NS_595 0 1.0142112816901291e-06
GC_11_596 b_11 NI_11 NS_596 0 5.9014854708266872e-07
GC_11_597 b_11 NI_11 NS_597 0 1.3671686378479497e-06
GC_11_598 b_11 NI_11 NS_598 0 -9.4667443677842930e-07
GC_11_599 b_11 NI_11 NS_599 0 8.0331064705082157e-06
GC_11_600 b_11 NI_11 NS_600 0 -2.1787352061490799e-06
GC_11_601 b_11 NI_11 NS_601 0 1.1742120462661293e-06
GC_11_602 b_11 NI_11 NS_602 0 1.5187607003737306e-06
GC_11_603 b_11 NI_11 NS_603 0 1.5706057400733682e-06
GC_11_604 b_11 NI_11 NS_604 0 -2.4568473491168452e-07
GC_11_605 b_11 NI_11 NS_605 0 1.3311101536014221e-06
GC_11_606 b_11 NI_11 NS_606 0 -9.9726164104524347e-07
GC_11_607 b_11 NI_11 NS_607 0 5.8014359417007884e-06
GC_11_608 b_11 NI_11 NS_608 0 -3.9293847873235988e-06
GC_11_609 b_11 NI_11 NS_609 0 1.8001485245925592e-06
GC_11_610 b_11 NI_11 NS_610 0 1.4046059612002007e-06
GC_11_611 b_11 NI_11 NS_611 0 1.0780206075756105e-06
GC_11_612 b_11 NI_11 NS_612 0 -1.3987218167396702e-06
GC_11_613 b_11 NI_11 NS_613 0 1.4203360183141213e-06
GC_11_614 b_11 NI_11 NS_614 0 -1.1295839060437586e-06
GC_11_615 b_11 NI_11 NS_615 0 2.9391206551260749e-06
GC_11_616 b_11 NI_11 NS_616 0 -4.1900422367294309e-06
GC_11_617 b_11 NI_11 NS_617 0 2.2053955854857455e-06
GC_11_618 b_11 NI_11 NS_618 0 2.9634962318712889e-07
GC_11_619 b_11 NI_11 NS_619 0 -3.3187066091815124e-07
GC_11_620 b_11 NI_11 NS_620 0 -1.1800080686615166e-06
GC_11_621 b_11 NI_11 NS_621 0 2.4885353982849419e-11
GC_11_622 b_11 NI_11 NS_622 0 -4.0917226468044085e-11
GC_11_623 b_11 NI_11 NS_623 0 7.9132784974973645e-07
GC_11_624 b_11 NI_11 NS_624 0 -1.5907635018577726e-06
GC_11_625 b_11 NI_11 NS_625 0 1.2547874403691662e-06
GC_11_626 b_11 NI_11 NS_626 0 2.2340425074141187e-07
GC_11_627 b_11 NI_11 NS_627 0 1.5908880298045186e-07
GC_11_628 b_11 NI_11 NS_628 0 -5.4772279036194644e-07
GC_11_629 b_11 NI_11 NS_629 0 5.4957143221997882e-07
GC_11_630 b_11 NI_11 NS_630 0 -8.9267308055882746e-07
GC_11_631 b_11 NI_11 NS_631 0 1.2802167678357862e-06
GC_11_632 b_11 NI_11 NS_632 0 -2.0630239483544660e-06
GC_11_633 b_11 NI_11 NS_633 0 4.7394939265746462e-10
GC_11_634 b_11 NI_11 NS_634 0 -1.2084252967943683e-09
GC_11_635 b_11 NI_11 NS_635 0 5.4791599554560016e-07
GC_11_636 b_11 NI_11 NS_636 0 -8.5973182684616817e-07
GC_11_637 b_11 NI_11 NS_637 0 7.1441927063736965e-07
GC_11_638 b_11 NI_11 NS_638 0 -9.5097433458538918e-07
GC_11_639 b_11 NI_11 NS_639 0 8.9079180881933475e-08
GC_11_640 b_11 NI_11 NS_640 0 5.0128481631672069e-08
GC_11_641 b_11 NI_11 NS_641 0 1.3250930802332785e-06
GC_11_642 b_11 NI_11 NS_642 0 -1.2292262761955437e-06
GC_11_643 b_11 NI_11 NS_643 0 1.6446052284193264e-06
GC_11_644 b_11 NI_11 NS_644 0 -2.9221591721822180e-07
GC_11_645 b_11 NI_11 NS_645 0 -2.2768043871951604e-07
GC_11_646 b_11 NI_11 NS_646 0 -7.3422419449116909e-07
GC_11_647 b_11 NI_11 NS_647 0 7.3335519895269940e-07
GC_11_648 b_11 NI_11 NS_648 0 2.8942338584147594e-07
GC_11_649 b_11 NI_11 NS_649 0 -5.1646798695687997e-05
GC_11_650 b_11 NI_11 NS_650 0 -7.9566427030670014e-12
GC_11_651 b_11 NI_11 NS_651 0 -2.0642376936136041e-10
GC_11_652 b_11 NI_11 NS_652 0 9.8399918745150515e-09
GC_11_653 b_11 NI_11 NS_653 0 5.5721847544480933e-07
GC_11_654 b_11 NI_11 NS_654 0 5.0159557898005750e-08
GC_11_655 b_11 NI_11 NS_655 0 2.9182992383992575e-06
GC_11_656 b_11 NI_11 NS_656 0 -1.4785626874605415e-06
GC_11_657 b_11 NI_11 NS_657 0 -3.1221352142645256e-06
GC_11_658 b_11 NI_11 NS_658 0 -2.6253130596995867e-06
GC_11_659 b_11 NI_11 NS_659 0 4.5600550102739252e-06
GC_11_660 b_11 NI_11 NS_660 0 -4.1953995852421246e-07
GC_11_661 b_11 NI_11 NS_661 0 -7.3317359573750682e-06
GC_11_662 b_11 NI_11 NS_662 0 -7.4847503239395851e-06
GC_11_663 b_11 NI_11 NS_663 0 -2.4481673741194443e-07
GC_11_664 b_11 NI_11 NS_664 0 -1.3835223270728539e-06
GC_11_665 b_11 NI_11 NS_665 0 -5.8631657947663872e-06
GC_11_666 b_11 NI_11 NS_666 0 2.4072496521457889e-06
GC_11_667 b_11 NI_11 NS_667 0 5.0674510783639878e-06
GC_11_668 b_11 NI_11 NS_668 0 -5.0233991665861474e-06
GC_11_669 b_11 NI_11 NS_669 0 -1.6437325812031853e-05
GC_11_670 b_11 NI_11 NS_670 0 4.9721645795789639e-06
GC_11_671 b_11 NI_11 NS_671 0 -1.1936073390886231e-06
GC_11_672 b_11 NI_11 NS_672 0 7.3470965657455894e-06
GC_11_673 b_11 NI_11 NS_673 0 -6.5660734996352732e-06
GC_11_674 b_11 NI_11 NS_674 0 -3.8974726674457829e-06
GC_11_675 b_11 NI_11 NS_675 0 -3.2508502689990759e-06
GC_11_676 b_11 NI_11 NS_676 0 8.1592787896994959e-06
GC_11_677 b_11 NI_11 NS_677 0 -1.3863283148517460e-06
GC_11_678 b_11 NI_11 NS_678 0 -3.8634305817366027e-06
GC_11_679 b_11 NI_11 NS_679 0 -3.9088389336375179e-06
GC_11_680 b_11 NI_11 NS_680 0 1.1192659970600639e-05
GC_11_681 b_11 NI_11 NS_681 0 -1.0533526163833406e-07
GC_11_682 b_11 NI_11 NS_682 0 7.4969856678526015e-06
GC_11_683 b_11 NI_11 NS_683 0 -3.5950148684621014e-06
GC_11_684 b_11 NI_11 NS_684 0 1.5343060687319634e-06
GC_11_685 b_11 NI_11 NS_685 0 -4.2006664695517802e-07
GC_11_686 b_11 NI_11 NS_686 0 8.2501961039146560e-06
GC_11_687 b_11 NI_11 NS_687 0 -5.3672269294246034e-07
GC_11_688 b_11 NI_11 NS_688 0 2.2139602226457790e-06
GC_11_689 b_11 NI_11 NS_689 0 -2.2958978944668313e-06
GC_11_690 b_11 NI_11 NS_690 0 8.3126795905288297e-06
GC_11_691 b_11 NI_11 NS_691 0 6.2644741480284979e-07
GC_11_692 b_11 NI_11 NS_692 0 9.9677232366416583e-06
GC_11_693 b_11 NI_11 NS_693 0 -6.6638618848404149e-07
GC_11_694 b_11 NI_11 NS_694 0 8.7834118357190500e-06
GC_11_695 b_11 NI_11 NS_695 0 -1.2310798051385836e-06
GC_11_696 b_11 NI_11 NS_696 0 4.0450382323175196e-06
GC_11_697 b_11 NI_11 NS_697 0 1.2531597097518103e-06
GC_11_698 b_11 NI_11 NS_698 0 1.2151059459829122e-05
GC_11_699 b_11 NI_11 NS_699 0 1.8598607082397892e-05
GC_11_700 b_11 NI_11 NS_700 0 1.6955555104137267e-05
GC_11_701 b_11 NI_11 NS_701 0 4.9927745479467939e-06
GC_11_702 b_11 NI_11 NS_702 0 7.7348604833023969e-06
GC_11_703 b_11 NI_11 NS_703 0 1.0287804763346166e-05
GC_11_704 b_11 NI_11 NS_704 0 3.8686390570116757e-06
GC_11_705 b_11 NI_11 NS_705 0 6.7815814395759931e-06
GC_11_706 b_11 NI_11 NS_706 0 1.0888476522568376e-05
GC_11_707 b_11 NI_11 NS_707 0 3.3297996583982408e-05
GC_11_708 b_11 NI_11 NS_708 0 -6.1160186097196134e-06
GC_11_709 b_11 NI_11 NS_709 0 8.1345732690543672e-06
GC_11_710 b_11 NI_11 NS_710 0 3.3940892912654208e-06
GC_11_711 b_11 NI_11 NS_711 0 1.1919583779267808e-05
GC_11_712 b_11 NI_11 NS_712 0 -1.0263713414075611e-05
GC_11_713 b_11 NI_11 NS_713 0 1.0740952229285949e-05
GC_11_714 b_11 NI_11 NS_714 0 6.4520281781210865e-06
GC_11_715 b_11 NI_11 NS_715 0 1.6864073006609370e-05
GC_11_716 b_11 NI_11 NS_716 0 -3.0725038689064046e-05
GC_11_717 b_11 NI_11 NS_717 0 8.0822545272638368e-06
GC_11_718 b_11 NI_11 NS_718 0 -2.9351845815070273e-06
GC_11_719 b_11 NI_11 NS_719 0 -3.2232091688073894e-06
GC_11_720 b_11 NI_11 NS_720 0 -1.6225074424539866e-05
GC_11_721 b_11 NI_11 NS_721 0 1.1764426851216578e-05
GC_11_722 b_11 NI_11 NS_722 0 -1.6046710627541997e-06
GC_11_723 b_11 NI_11 NS_723 0 -1.2697690406668576e-05
GC_11_724 b_11 NI_11 NS_724 0 -2.5038899439384442e-05
GC_11_725 b_11 NI_11 NS_725 0 -1.6043417862372891e-07
GC_11_726 b_11 NI_11 NS_726 0 -6.5987140136087396e-06
GC_11_727 b_11 NI_11 NS_727 0 -9.5600448251895806e-06
GC_11_728 b_11 NI_11 NS_728 0 -2.6183610899929098e-06
GC_11_729 b_11 NI_11 NS_729 0 1.0192255713336260e-10
GC_11_730 b_11 NI_11 NS_730 0 4.7260049302290456e-11
GC_11_731 b_11 NI_11 NS_731 0 1.4895148579373761e-06
GC_11_732 b_11 NI_11 NS_732 0 -4.6804882132483855e-06
GC_11_733 b_11 NI_11 NS_733 0 -1.3643762447735236e-06
GC_11_734 b_11 NI_11 NS_734 0 -1.3419853307157513e-06
GC_11_735 b_11 NI_11 NS_735 0 -4.8481160024181738e-06
GC_11_736 b_11 NI_11 NS_736 0 -9.9610103489413351e-07
GC_11_737 b_11 NI_11 NS_737 0 -1.1402780254133910e-06
GC_11_738 b_11 NI_11 NS_738 0 -2.7145518342428653e-06
GC_11_739 b_11 NI_11 NS_739 0 -9.9975792057213769e-06
GC_11_740 b_11 NI_11 NS_740 0 -4.0377362901655573e-06
GC_11_741 b_11 NI_11 NS_741 0 6.6624158169560194e-09
GC_11_742 b_11 NI_11 NS_742 0 5.4072847165811206e-09
GC_11_743 b_11 NI_11 NS_743 0 1.7619936142441860e-06
GC_11_744 b_11 NI_11 NS_744 0 4.8751324783396479e-07
GC_11_745 b_11 NI_11 NS_745 0 -1.6125717880839375e-06
GC_11_746 b_11 NI_11 NS_746 0 3.2218636426494935e-06
GC_11_747 b_11 NI_11 NS_747 0 -8.2907765394165729e-07
GC_11_748 b_11 NI_11 NS_748 0 6.9895331745570665e-07
GC_11_749 b_11 NI_11 NS_749 0 -7.6542251761156431e-06
GC_11_750 b_11 NI_11 NS_750 0 5.4120104464270793e-07
GC_11_751 b_11 NI_11 NS_751 0 -2.2205060223949395e-06
GC_11_752 b_11 NI_11 NS_752 0 1.9993207727952716e-06
GC_11_753 b_11 NI_11 NS_753 0 -2.0646060652252095e-06
GC_11_754 b_11 NI_11 NS_754 0 1.9702201187888038e-06
GC_11_755 b_11 NI_11 NS_755 0 1.2826140775434031e-06
GC_11_756 b_11 NI_11 NS_756 0 2.8349437389055445e-06
GC_11_757 b_11 NI_11 NS_757 0 -1.5116973209330250e-04
GC_11_758 b_11 NI_11 NS_758 0 3.7546598841752513e-11
GC_11_759 b_11 NI_11 NS_759 0 1.7615113257615672e-11
GC_11_760 b_11 NI_11 NS_760 0 8.7387846867973112e-10
GC_11_761 b_11 NI_11 NS_761 0 -2.3302531529100431e-06
GC_11_762 b_11 NI_11 NS_762 0 -1.6501620552439969e-06
GC_11_763 b_11 NI_11 NS_763 0 1.4540862361935820e-06
GC_11_764 b_11 NI_11 NS_764 0 3.8965308231188205e-06
GC_11_765 b_11 NI_11 NS_765 0 2.9654337140319574e-06
GC_11_766 b_11 NI_11 NS_766 0 5.4214123965398420e-06
GC_11_767 b_11 NI_11 NS_767 0 5.3772097822125401e-06
GC_11_768 b_11 NI_11 NS_768 0 -8.4804847490036109e-06
GC_11_769 b_11 NI_11 NS_769 0 -2.2508519049887351e-06
GC_11_770 b_11 NI_11 NS_770 0 -1.2662156659969794e-05
GC_11_771 b_11 NI_11 NS_771 0 -3.7274309588675667e-06
GC_11_772 b_11 NI_11 NS_772 0 2.7451147196257341e-06
GC_11_773 b_11 NI_11 NS_773 0 4.4942013687922807e-06
GC_11_774 b_11 NI_11 NS_774 0 1.5804074916351522e-06
GC_11_775 b_11 NI_11 NS_775 0 8.5384675981603366e-06
GC_11_776 b_11 NI_11 NS_776 0 -3.8252132085773118e-05
GC_11_777 b_11 NI_11 NS_777 0 -4.2843645921542235e-05
GC_11_778 b_11 NI_11 NS_778 0 -1.4538433936050804e-06
GC_11_779 b_11 NI_11 NS_779 0 -1.4647394371826490e-05
GC_11_780 b_11 NI_11 NS_780 0 -8.2775807264751092e-06
GC_11_781 b_11 NI_11 NS_781 0 -7.0243598634605752e-05
GC_11_782 b_11 NI_11 NS_782 0 7.5186044850558876e-05
GC_11_783 b_11 NI_11 NS_783 0 4.8693950976937240e-06
GC_11_784 b_11 NI_11 NS_784 0 1.3024168469148611e-05
GC_11_785 b_11 NI_11 NS_785 0 6.5219893047802443e-05
GC_11_786 b_11 NI_11 NS_786 0 1.2202210031326253e-04
GC_11_787 b_11 NI_11 NS_787 0 -2.7571748785179399e-07
GC_11_788 b_11 NI_11 NS_788 0 -3.7368889188360988e-05
GC_11_789 b_11 NI_11 NS_789 0 1.6806412904811804e-05
GC_11_790 b_11 NI_11 NS_790 0 4.1840162918711615e-06
GC_11_791 b_11 NI_11 NS_791 0 2.5159041336808370e-05
GC_11_792 b_11 NI_11 NS_792 0 -3.0985794573826693e-05
GC_11_793 b_11 NI_11 NS_793 0 -8.5163944408933128e-06
GC_11_794 b_11 NI_11 NS_794 0 -2.5732996889879336e-06
GC_11_795 b_11 NI_11 NS_795 0 -8.0803365949367260e-06
GC_11_796 b_11 NI_11 NS_796 0 2.4256748024574292e-05
GC_11_797 b_11 NI_11 NS_797 0 6.0403016307459326e-06
GC_11_798 b_11 NI_11 NS_798 0 8.3879441266226031e-06
GC_11_799 b_11 NI_11 NS_799 0 5.7351161438142023e-05
GC_11_800 b_11 NI_11 NS_800 0 2.3736651584561427e-05
GC_11_801 b_11 NI_11 NS_801 0 3.5347152603436151e-06
GC_11_802 b_11 NI_11 NS_802 0 -1.2244130836345103e-05
GC_11_803 b_11 NI_11 NS_803 0 -7.4154769599914765e-08
GC_11_804 b_11 NI_11 NS_804 0 -1.3740050856492290e-06
GC_11_805 b_11 NI_11 NS_805 0 7.1802735015736336e-06
GC_11_806 b_11 NI_11 NS_806 0 2.7779113231230720e-06
GC_11_807 b_11 NI_11 NS_807 0 4.2417158066958649e-05
GC_11_808 b_11 NI_11 NS_808 0 -1.9012475153000079e-05
GC_11_809 b_11 NI_11 NS_809 0 -2.5057075377338703e-06
GC_11_810 b_11 NI_11 NS_810 0 -7.6313017963550138e-06
GC_11_811 b_11 NI_11 NS_811 0 -2.8031620607922711e-06
GC_11_812 b_11 NI_11 NS_812 0 1.0883299557784438e-06
GC_11_813 b_11 NI_11 NS_813 0 9.8314179799252731e-06
GC_11_814 b_11 NI_11 NS_814 0 2.5417455252718137e-06
GC_11_815 b_11 NI_11 NS_815 0 2.2416089609475771e-05
GC_11_816 b_11 NI_11 NS_816 0 -3.3139475079304017e-05
GC_11_817 b_11 NI_11 NS_817 0 -5.7255553766850987e-06
GC_11_818 b_11 NI_11 NS_818 0 -4.2016025877016862e-06
GC_11_819 b_11 NI_11 NS_819 0 -8.8988219320295549e-07
GC_11_820 b_11 NI_11 NS_820 0 4.2524245129273106e-06
GC_11_821 b_11 NI_11 NS_821 0 1.2480231041174422e-05
GC_11_822 b_11 NI_11 NS_822 0 -2.7947895761401327e-07
GC_11_823 b_11 NI_11 NS_823 0 4.7407244122695477e-07
GC_11_824 b_11 NI_11 NS_824 0 -3.2834919002924451e-05
GC_11_825 b_11 NI_11 NS_825 0 -6.9267938707711222e-06
GC_11_826 b_11 NI_11 NS_826 0 4.0680033172104580e-07
GC_11_827 b_11 NI_11 NS_827 0 3.8410663650219147e-06
GC_11_828 b_11 NI_11 NS_828 0 3.5676051184222075e-06
GC_11_829 b_11 NI_11 NS_829 0 1.4108535310095255e-05
GC_11_830 b_11 NI_11 NS_830 0 -6.6872349083419219e-06
GC_11_831 b_11 NI_11 NS_831 0 -1.5604808656967535e-05
GC_11_832 b_11 NI_11 NS_832 0 -1.9003791943323888e-05
GC_11_833 b_11 NI_11 NS_833 0 -2.9951981074045067e-06
GC_11_834 b_11 NI_11 NS_834 0 5.1042286440047098e-06
GC_11_835 b_11 NI_11 NS_835 0 4.2096656210346286e-06
GC_11_836 b_11 NI_11 NS_836 0 -1.8810298573577995e-06
GC_11_837 b_11 NI_11 NS_837 0 -2.7916683932147865e-11
GC_11_838 b_11 NI_11 NS_838 0 5.8150864957441957e-12
GC_11_839 b_11 NI_11 NS_839 0 4.8699137466206950e-06
GC_11_840 b_11 NI_11 NS_840 0 -1.1668169836777485e-05
GC_11_841 b_11 NI_11 NS_841 0 -5.0904558426761730e-07
GC_11_842 b_11 NI_11 NS_842 0 2.7992314365992660e-06
GC_11_843 b_11 NI_11 NS_843 0 2.3509278632040767e-06
GC_11_844 b_11 NI_11 NS_844 0 -1.5716763864796212e-06
GC_11_845 b_11 NI_11 NS_845 0 2.1314585458344191e-06
GC_11_846 b_11 NI_11 NS_846 0 -9.8974505345331700e-06
GC_11_847 b_11 NI_11 NS_847 0 -1.0613671306170625e-05
GC_11_848 b_11 NI_11 NS_848 0 -3.5263816491703867e-06
GC_11_849 b_11 NI_11 NS_849 0 -2.3906760303211811e-10
GC_11_850 b_11 NI_11 NS_850 0 4.4559191400262564e-10
GC_11_851 b_11 NI_11 NS_851 0 -9.1766888296505710e-06
GC_11_852 b_11 NI_11 NS_852 0 -5.6138462667125024e-06
GC_11_853 b_11 NI_11 NS_853 0 1.9952310344206583e-06
GC_11_854 b_11 NI_11 NS_854 0 -6.7132344916335987e-06
GC_11_855 b_11 NI_11 NS_855 0 -3.3605892754247593e-06
GC_11_856 b_11 NI_11 NS_856 0 -1.7941591596821865e-07
GC_11_857 b_11 NI_11 NS_857 0 -8.5928703242071578e-06
GC_11_858 b_11 NI_11 NS_858 0 5.9552819158592037e-07
GC_11_859 b_11 NI_11 NS_859 0 2.6078615947019204e-06
GC_11_860 b_11 NI_11 NS_860 0 2.8392948884427544e-06
GC_11_861 b_11 NI_11 NS_861 0 9.9242080966193000e-07
GC_11_862 b_11 NI_11 NS_862 0 -3.6889661934158396e-06
GC_11_863 b_11 NI_11 NS_863 0 -5.4153669536808135e-06
GC_11_864 b_11 NI_11 NS_864 0 -4.2328094794469858e-06
GC_11_865 b_11 NI_11 NS_865 0 1.1804777683497181e-03
GC_11_866 b_11 NI_11 NS_866 0 -3.5559914947896637e-09
GC_11_867 b_11 NI_11 NS_867 0 -4.8002576918850535e-08
GC_11_868 b_11 NI_11 NS_868 0 -3.4752161331355564e-06
GC_11_869 b_11 NI_11 NS_869 0 -3.6812591732166331e-04
GC_11_870 b_11 NI_11 NS_870 0 1.3598228422270089e-04
GC_11_871 b_11 NI_11 NS_871 0 1.1297229504252978e-03
GC_11_872 b_11 NI_11 NS_872 0 1.9432474187168003e-03
GC_11_873 b_11 NI_11 NS_873 0 -6.5058703572620736e-05
GC_11_874 b_11 NI_11 NS_874 0 -3.4937467840565088e-03
GC_11_875 b_11 NI_11 NS_875 0 -1.5644000874451538e-03
GC_11_876 b_11 NI_11 NS_876 0 5.0906047862238199e-03
GC_11_877 b_11 NI_11 NS_877 0 4.2534009791018700e-03
GC_11_878 b_11 NI_11 NS_878 0 -4.9938043723831375e-03
GC_11_879 b_11 NI_11 NS_879 0 -1.0085534104762443e-03
GC_11_880 b_11 NI_11 NS_880 0 5.6397848515130035e-04
GC_11_881 b_11 NI_11 NS_881 0 -2.0807522902705146e-03
GC_11_882 b_11 NI_11 NS_882 0 -1.8633136559347693e-03
GC_11_883 b_11 NI_11 NS_883 0 3.6454404149434865e-03
GC_11_884 b_11 NI_11 NS_884 0 1.1647363854914255e-02
GC_11_885 b_11 NI_11 NS_885 0 -8.9814490637160941e-04
GC_11_886 b_11 NI_11 NS_886 0 -1.4854322467497044e-02
GC_11_887 b_11 NI_11 NS_887 0 -8.1235366917756912e-03
GC_11_888 b_11 NI_11 NS_888 0 1.9196054013952081e-03
GC_11_889 b_11 NI_11 NS_889 0 1.1263052262444843e-02
GC_11_890 b_11 NI_11 NS_890 0 -1.8122303811994292e-03
GC_11_891 b_11 NI_11 NS_891 0 -7.5672721671333461e-03
GC_11_892 b_11 NI_11 NS_892 0 -1.6811809006930984e-03
GC_11_893 b_11 NI_11 NS_893 0 1.5281711704015034e-02
GC_11_894 b_11 NI_11 NS_894 0 5.3008478715178909e-03
GC_11_895 b_11 NI_11 NS_895 0 -1.3082857193876184e-02
GC_11_896 b_11 NI_11 NS_896 0 -5.4612980857567540e-03
GC_11_897 b_11 NI_11 NS_897 0 -6.6370720068815170e-03
GC_11_898 b_11 NI_11 NS_898 0 3.4566941278901548e-03
GC_11_899 b_11 NI_11 NS_899 0 6.3616038437346398e-03
GC_11_900 b_11 NI_11 NS_900 0 -1.8793238139983908e-03
GC_11_901 b_11 NI_11 NS_901 0 -5.4737178432873960e-03
GC_11_902 b_11 NI_11 NS_902 0 2.1830275702704382e-03
GC_11_903 b_11 NI_11 NS_903 0 5.3937685500655376e-03
GC_11_904 b_11 NI_11 NS_904 0 -2.6324368439137264e-03
GC_11_905 b_11 NI_11 NS_905 0 -6.3064548530876573e-03
GC_11_906 b_11 NI_11 NS_906 0 -4.8381422322169357e-04
GC_11_907 b_11 NI_11 NS_907 0 7.6452813373800157e-03
GC_11_908 b_11 NI_11 NS_908 0 3.6298748801939355e-03
GC_11_909 b_11 NI_11 NS_909 0 -5.8336237575829153e-03
GC_11_910 b_11 NI_11 NS_910 0 -3.4645950540192071e-03
GC_11_911 b_11 NI_11 NS_911 0 2.9620064699018050e-04
GC_11_912 b_11 NI_11 NS_912 0 5.5810490949424437e-04
GC_11_913 b_11 NI_11 NS_913 0 -4.9270622018717019e-03
GC_11_914 b_11 NI_11 NS_914 0 8.9219844387939567e-04
GC_11_915 b_11 NI_11 NS_915 0 6.2063433395610559e-03
GC_11_916 b_11 NI_11 NS_916 0 6.8827280037008713e-04
GC_11_917 b_11 NI_11 NS_917 0 -5.3209627948281402e-03
GC_11_918 b_11 NI_11 NS_918 0 -4.8419034240276371e-04
GC_11_919 b_11 NI_11 NS_919 0 1.5503311578842901e-03
GC_11_920 b_11 NI_11 NS_920 0 -4.3208426471648005e-05
GC_11_921 b_11 NI_11 NS_921 0 -6.0223341909896623e-03
GC_11_922 b_11 NI_11 NS_922 0 1.9232416158411940e-03
GC_11_923 b_11 NI_11 NS_923 0 6.2616668284911419e-03
GC_11_924 b_11 NI_11 NS_924 0 2.1736512536827641e-04
GC_11_925 b_11 NI_11 NS_925 0 -5.0591977956354339e-03
GC_11_926 b_11 NI_11 NS_926 0 1.7016169638888457e-03
GC_11_927 b_11 NI_11 NS_927 0 2.4884743734153573e-03
GC_11_928 b_11 NI_11 NS_928 0 -9.5765186686157710e-04
GC_11_929 b_11 NI_11 NS_929 0 -6.5329624741576218e-03
GC_11_930 b_11 NI_11 NS_930 0 3.8846374153702077e-03
GC_11_931 b_11 NI_11 NS_931 0 7.4932671045410335e-03
GC_11_932 b_11 NI_11 NS_932 0 -1.0960284059472133e-03
GC_11_933 b_11 NI_11 NS_933 0 -3.9851195992949388e-03
GC_11_934 b_11 NI_11 NS_934 0 4.0409800184821251e-03
GC_11_935 b_11 NI_11 NS_935 0 2.8633259784485486e-03
GC_11_936 b_11 NI_11 NS_936 0 -3.0534881857054099e-03
GC_11_937 b_11 NI_11 NS_937 0 -6.0227294634721592e-03
GC_11_938 b_11 NI_11 NS_938 0 7.2373898824169046e-03
GC_11_939 b_11 NI_11 NS_939 0 7.9897123603499456e-03
GC_11_940 b_11 NI_11 NS_940 0 -4.8114592221880741e-03
GC_11_941 b_11 NI_11 NS_941 0 -5.3741854794193847e-04
GC_11_942 b_11 NI_11 NS_942 0 5.0204729911852179e-03
GC_11_943 b_11 NI_11 NS_943 0 2.4825585937043030e-04
GC_11_944 b_11 NI_11 NS_944 0 -4.7581979868240769e-03
GC_11_945 b_11 NI_11 NS_945 0 1.8109009045296763e-09
GC_11_946 b_11 NI_11 NS_946 0 3.2745350759719528e-09
GC_11_947 b_11 NI_11 NS_947 0 -1.4271956704142315e-03
GC_11_948 b_11 NI_11 NS_948 0 7.8707399222078898e-03
GC_11_949 b_11 NI_11 NS_949 0 -1.7997912138199010e-04
GC_11_950 b_11 NI_11 NS_950 0 3.0272438861498304e-03
GC_11_951 b_11 NI_11 NS_951 0 -1.3038560981469457e-04
GC_11_952 b_11 NI_11 NS_952 0 -3.3753040658697285e-03
GC_11_953 b_11 NI_11 NS_953 0 -8.7631227784924228e-04
GC_11_954 b_11 NI_11 NS_954 0 7.5304822482262241e-03
GC_11_955 b_11 NI_11 NS_955 0 3.7888078988001215e-03
GC_11_956 b_11 NI_11 NS_956 0 -6.1574217064608357e-03
GC_11_957 b_11 NI_11 NS_957 0 8.6236192411793657e-08
GC_11_958 b_11 NI_11 NS_958 0 -3.5294023117687628e-07
GC_11_959 b_11 NI_11 NS_959 0 6.7186800340163734e-03
GC_11_960 b_11 NI_11 NS_960 0 -5.3194114838276130e-03
GC_11_961 b_11 NI_11 NS_961 0 -2.6111717720343863e-03
GC_11_962 b_11 NI_11 NS_962 0 6.0542407261782701e-03
GC_11_963 b_11 NI_11 NS_963 0 -4.2922715109812602e-03
GC_11_964 b_11 NI_11 NS_964 0 1.4429442712241248e-05
GC_11_965 b_11 NI_11 NS_965 0 2.7173883569819230e-03
GC_11_966 b_11 NI_11 NS_966 0 -6.2040232047718353e-03
GC_11_967 b_11 NI_11 NS_967 0 2.0957197437900263e-03
GC_11_968 b_11 NI_11 NS_968 0 3.2562724655940652e-03
GC_11_969 b_11 NI_11 NS_969 0 -1.9700345763534401e-03
GC_11_970 b_11 NI_11 NS_970 0 -4.4205367865173236e-03
GC_11_971 b_11 NI_11 NS_971 0 2.8640861259799882e-03
GC_11_972 b_11 NI_11 NS_972 0 8.0083630266011251e-03
GC_11_973 b_11 NI_11 NS_973 0 -3.3036441655561540e-03
GC_11_974 b_11 NI_11 NS_974 0 1.8493853258671468e-09
GC_11_975 b_11 NI_11 NS_975 0 5.6032181502941214e-08
GC_11_976 b_11 NI_11 NS_976 0 1.8929694819886544e-06
GC_11_977 b_11 NI_11 NS_977 0 -9.1167728748561648e-05
GC_11_978 b_11 NI_11 NS_978 0 -5.7737931421662325e-05
GC_11_979 b_11 NI_11 NS_979 0 -1.2657732620225774e-03
GC_11_980 b_11 NI_11 NS_980 0 -2.9559391350491969e-04
GC_11_981 b_11 NI_11 NS_981 0 -1.6792134994910886e-03
GC_11_982 b_11 NI_11 NS_982 0 2.6464975804306005e-03
GC_11_983 b_11 NI_11 NS_983 0 5.1121163939702287e-04
GC_11_984 b_11 NI_11 NS_984 0 5.4276087175277295e-03
GC_11_985 b_11 NI_11 NS_985 0 7.1034879037031162e-03
GC_11_986 b_11 NI_11 NS_986 0 6.3629217883651721e-04
GC_11_987 b_11 NI_11 NS_987 0 6.4432949324230845e-04
GC_11_988 b_11 NI_11 NS_988 0 -6.6091957444520055e-04
GC_11_989 b_11 NI_11 NS_989 0 1.0576978459035833e-03
GC_11_990 b_11 NI_11 NS_990 0 1.5711412072036848e-03
GC_11_991 b_11 NI_11 NS_991 0 1.2687513992416433e-02
GC_11_992 b_11 NI_11 NS_992 0 1.3123213831239969e-02
GC_11_993 b_11 NI_11 NS_993 0 8.7187980180075206e-03
GC_11_994 b_11 NI_11 NS_994 0 -2.0392080760680484e-02
GC_11_995 b_11 NI_11 NS_995 0 8.3891007651850230e-03
GC_11_996 b_11 NI_11 NS_996 0 -2.9045258255855850e-03
GC_11_997 b_11 NI_11 NS_997 0 -1.2701289634500052e-02
GC_11_998 b_11 NI_11 NS_998 0 -3.8806698553382118e-02
GC_11_999 b_11 NI_11 NS_999 0 -7.2523391625196523e-03
GC_11_1000 b_11 NI_11 NS_1000 0 -2.1332749468762086e-03
GC_11_1001 b_11 NI_11 NS_1001 0 -5.2307199540881248e-02
GC_11_1002 b_11 NI_11 NS_1002 0 -1.7936156080951536e-03
GC_11_1003 b_11 NI_11 NS_1003 0 1.4914415710458489e-02
GC_11_1004 b_11 NI_11 NS_1004 0 8.6735766457814913e-03
GC_11_1005 b_11 NI_11 NS_1005 0 -5.9233530164824258e-03
GC_11_1006 b_11 NI_11 NS_1006 0 5.0044974736494444e-03
GC_11_1007 b_11 NI_11 NS_1007 0 8.3724199626970842e-03
GC_11_1008 b_11 NI_11 NS_1008 0 1.1688363049604611e-02
GC_11_1009 b_11 NI_11 NS_1009 0 4.5592638391056296e-03
GC_11_1010 b_11 NI_11 NS_1010 0 -2.9327411485256345e-03
GC_11_1011 b_11 NI_11 NS_1011 0 -7.8986738270046177e-03
GC_11_1012 b_11 NI_11 NS_1012 0 -8.1490651620074340e-03
GC_11_1013 b_11 NI_11 NS_1013 0 -5.6808140409970757e-03
GC_11_1014 b_11 NI_11 NS_1014 0 -6.1281001093603841e-04
GC_11_1015 b_11 NI_11 NS_1015 0 -1.8070850602408203e-02
GC_11_1016 b_11 NI_11 NS_1016 0 1.3578965346696208e-02
GC_11_1017 b_11 NI_11 NS_1017 0 4.7069865920809691e-03
GC_11_1018 b_11 NI_11 NS_1018 0 4.3794388563153158e-03
GC_11_1019 b_11 NI_11 NS_1019 0 6.5015827404072920e-04
GC_11_1020 b_11 NI_11 NS_1020 0 -1.0995438746514383e-04
GC_11_1021 b_11 NI_11 NS_1021 0 -3.7964000774214227e-03
GC_11_1022 b_11 NI_11 NS_1022 0 8.8498889360328519e-04
GC_11_1023 b_11 NI_11 NS_1023 0 -1.1178276372408385e-03
GC_11_1024 b_11 NI_11 NS_1024 0 1.6699689475247883e-02
GC_11_1025 b_11 NI_11 NS_1025 0 4.4472808477174306e-03
GC_11_1026 b_11 NI_11 NS_1026 0 7.0796447046562691e-04
GC_11_1027 b_11 NI_11 NS_1027 0 -5.1995804898919253e-04
GC_11_1028 b_11 NI_11 NS_1028 0 -2.2477509726368293e-03
GC_11_1029 b_11 NI_11 NS_1029 0 -4.9864557370828053e-03
GC_11_1030 b_11 NI_11 NS_1030 0 2.1108879669583429e-03
GC_11_1031 b_11 NI_11 NS_1031 0 7.3425285263141148e-03
GC_11_1032 b_11 NI_11 NS_1032 0 1.4345855708161765e-02
GC_11_1033 b_11 NI_11 NS_1033 0 4.1872276212500236e-03
GC_11_1034 b_11 NI_11 NS_1034 0 -1.6838583488149341e-03
GC_11_1035 b_11 NI_11 NS_1035 0 -3.3981244554010222e-03
GC_11_1036 b_11 NI_11 NS_1036 0 -2.1006228320542800e-03
GC_11_1037 b_11 NI_11 NS_1037 0 -5.4204253733874707e-03
GC_11_1038 b_11 NI_11 NS_1038 0 4.3817251711521727e-03
GC_11_1039 b_11 NI_11 NS_1039 0 1.3196874538179117e-02
GC_11_1040 b_11 NI_11 NS_1040 0 8.4333069183083319e-03
GC_11_1041 b_11 NI_11 NS_1041 0 2.8324343472100780e-03
GC_11_1042 b_11 NI_11 NS_1042 0 -4.1306062423332422e-03
GC_11_1043 b_11 NI_11 NS_1043 0 -5.3207858968504339e-03
GC_11_1044 b_11 NI_11 NS_1044 0 1.1381581027411509e-03
GC_11_1045 b_11 NI_11 NS_1045 0 -4.4310202425507025e-03
GC_11_1046 b_11 NI_11 NS_1046 0 8.3104314972415119e-03
GC_11_1047 b_11 NI_11 NS_1047 0 1.4612787213380439e-02
GC_11_1048 b_11 NI_11 NS_1048 0 -4.6824806816927431e-04
GC_11_1049 b_11 NI_11 NS_1049 0 -1.1845312440002421e-03
GC_11_1050 b_11 NI_11 NS_1050 0 -4.5473900572799413e-03
GC_11_1051 b_11 NI_11 NS_1051 0 -2.2825675113970932e-03
GC_11_1052 b_11 NI_11 NS_1052 0 4.3832539446405578e-03
GC_11_1053 b_11 NI_11 NS_1053 0 1.3571851004003309e-10
GC_11_1054 b_11 NI_11 NS_1054 0 -1.5466402002518953e-09
GC_11_1055 b_11 NI_11 NS_1055 0 1.4460267456937179e-03
GC_11_1056 b_11 NI_11 NS_1056 0 8.2165466663419381e-03
GC_11_1057 b_11 NI_11 NS_1057 0 -8.7895013012356360e-04
GC_11_1058 b_11 NI_11 NS_1058 0 -2.2072129540076082e-03
GC_11_1059 b_11 NI_11 NS_1059 0 -1.4679136789716657e-03
GC_11_1060 b_11 NI_11 NS_1060 0 2.7519856050621503e-03
GC_11_1061 b_11 NI_11 NS_1061 0 1.7320146213671026e-03
GC_11_1062 b_11 NI_11 NS_1062 0 7.6059320215133685e-03
GC_11_1063 b_11 NI_11 NS_1063 0 7.5874087826809603e-03
GC_11_1064 b_11 NI_11 NS_1064 0 -3.8276835702642916e-03
GC_11_1065 b_11 NI_11 NS_1065 0 -5.2101144615015857e-08
GC_11_1066 b_11 NI_11 NS_1066 0 -2.0817469170996233e-08
GC_11_1067 b_11 NI_11 NS_1067 0 1.1391243358446664e-02
GC_11_1068 b_11 NI_11 NS_1068 0 4.4700328420253276e-03
GC_11_1069 b_11 NI_11 NS_1069 0 -8.6185039051283544e-04
GC_11_1070 b_11 NI_11 NS_1070 0 6.4916224496049122e-03
GC_11_1071 b_11 NI_11 NS_1071 0 3.6263738653835504e-03
GC_11_1072 b_11 NI_11 NS_1072 0 4.0710465653183783e-04
GC_11_1073 b_11 NI_11 NS_1073 0 6.0525104791157311e-03
GC_11_1074 b_11 NI_11 NS_1074 0 -4.6635404975351779e-03
GC_11_1075 b_11 NI_11 NS_1075 0 -3.3929752426380532e-03
GC_11_1076 b_11 NI_11 NS_1076 0 -1.3533960203922261e-03
GC_11_1077 b_11 NI_11 NS_1077 0 1.1237969365618204e-04
GC_11_1078 b_11 NI_11 NS_1078 0 4.4958001859075371e-03
GC_11_1079 b_11 NI_11 NS_1079 0 7.2795569650201467e-03
GC_11_1080 b_11 NI_11 NS_1080 0 5.5305048439564432e-03
GC_11_1081 b_11 NI_11 NS_1081 0 -1.5530873157252996e-02
GC_11_1082 b_11 NI_11 NS_1082 0 6.4872979778679029e-09
GC_11_1083 b_11 NI_11 NS_1083 0 -1.0780989021983369e-06
GC_11_1084 b_11 NI_11 NS_1084 0 -2.3175273689931562e-05
GC_11_1085 b_11 NI_11 NS_1085 0 3.3380760691957014e-04
GC_11_1086 b_11 NI_11 NS_1086 0 -2.0548504348941833e-04
GC_11_1087 b_11 NI_11 NS_1087 0 -1.5862582016457861e-03
GC_11_1088 b_11 NI_11 NS_1088 0 -2.3361773046056472e-03
GC_11_1089 b_11 NI_11 NS_1089 0 -6.3216293149547171e-05
GC_11_1090 b_11 NI_11 NS_1090 0 4.3863824873940803e-03
GC_11_1091 b_11 NI_11 NS_1091 0 1.5399051133396923e-03
GC_11_1092 b_11 NI_11 NS_1092 0 -5.9456444705446613e-03
GC_11_1093 b_11 NI_11 NS_1093 0 -4.9710137011664303e-03
GC_11_1094 b_11 NI_11 NS_1094 0 6.5658936317762066e-03
GC_11_1095 b_11 NI_11 NS_1095 0 1.1033053449824549e-03
GC_11_1096 b_11 NI_11 NS_1096 0 -4.8869787764720108e-04
GC_11_1097 b_11 NI_11 NS_1097 0 2.8351196952451402e-03
GC_11_1098 b_11 NI_11 NS_1098 0 2.3742292490101288e-03
GC_11_1099 b_11 NI_11 NS_1099 0 -4.4219533089198074e-03
GC_11_1100 b_11 NI_11 NS_1100 0 -1.3476669330843538e-02
GC_11_1101 b_11 NI_11 NS_1101 0 1.7485556334057655e-03
GC_11_1102 b_11 NI_11 NS_1102 0 1.7702187650705983e-02
GC_11_1103 b_11 NI_11 NS_1103 0 9.8282590706879093e-03
GC_11_1104 b_11 NI_11 NS_1104 0 -2.3328384606742343e-03
GC_11_1105 b_11 NI_11 NS_1105 0 -1.3062251194868408e-02
GC_11_1106 b_11 NI_11 NS_1106 0 2.3406863257321997e-03
GC_11_1107 b_11 NI_11 NS_1107 0 9.2233755125555490e-03
GC_11_1108 b_11 NI_11 NS_1108 0 1.9112829960495400e-03
GC_11_1109 b_11 NI_11 NS_1109 0 -1.7997095729852034e-02
GC_11_1110 b_11 NI_11 NS_1110 0 -6.3438996795460324e-03
GC_11_1111 b_11 NI_11 NS_1111 0 1.5754262411181566e-02
GC_11_1112 b_11 NI_11 NS_1112 0 6.4095332590134611e-03
GC_11_1113 b_11 NI_11 NS_1113 0 8.1027179662440749e-03
GC_11_1114 b_11 NI_11 NS_1114 0 -4.2190607220787494e-03
GC_11_1115 b_11 NI_11 NS_1115 0 -7.4948905236186551e-03
GC_11_1116 b_11 NI_11 NS_1116 0 2.0941358803368412e-03
GC_11_1117 b_11 NI_11 NS_1117 0 6.7044806804505497e-03
GC_11_1118 b_11 NI_11 NS_1118 0 -2.7628598140632195e-03
GC_11_1119 b_11 NI_11 NS_1119 0 -6.5432384031292919e-03
GC_11_1120 b_11 NI_11 NS_1120 0 2.9299444241777501e-03
GC_11_1121 b_11 NI_11 NS_1121 0 7.6773811930028486e-03
GC_11_1122 b_11 NI_11 NS_1122 0 4.6375248856022570e-04
GC_11_1123 b_11 NI_11 NS_1123 0 -9.3401557078821532e-03
GC_11_1124 b_11 NI_11 NS_1124 0 -5.1079558757735387e-03
GC_11_1125 b_11 NI_11 NS_1125 0 6.8551899318492412e-03
GC_11_1126 b_11 NI_11 NS_1126 0 4.0869851681090037e-03
GC_11_1127 b_11 NI_11 NS_1127 0 -3.8349361445250114e-04
GC_11_1128 b_11 NI_11 NS_1128 0 -9.2299640121912643e-04
GC_11_1129 b_11 NI_11 NS_1129 0 5.6963380872604406e-03
GC_11_1130 b_11 NI_11 NS_1130 0 -1.3852984741729679e-03
GC_11_1131 b_11 NI_11 NS_1131 0 -9.1011003941192537e-03
GC_11_1132 b_11 NI_11 NS_1132 0 -1.2296022293431489e-03
GC_11_1133 b_11 NI_11 NS_1133 0 6.0201783816093016e-03
GC_11_1134 b_11 NI_11 NS_1134 0 7.1817207664889870e-04
GC_11_1135 b_11 NI_11 NS_1135 0 -2.6199034951045201e-03
GC_11_1136 b_11 NI_11 NS_1136 0 2.4600089255869586e-04
GC_11_1137 b_11 NI_11 NS_1137 0 6.7218306943104128e-03
GC_11_1138 b_11 NI_11 NS_1138 0 -2.2667468567521853e-03
GC_11_1139 b_11 NI_11 NS_1139 0 -9.2254224935980778e-03
GC_11_1140 b_11 NI_11 NS_1140 0 1.5046042797532922e-03
GC_11_1141 b_11 NI_11 NS_1141 0 5.7525380524021943e-03
GC_11_1142 b_11 NI_11 NS_1142 0 -1.5177994584734060e-03
GC_11_1143 b_11 NI_11 NS_1143 0 -3.2852559397145982e-03
GC_11_1144 b_11 NI_11 NS_1144 0 2.3899129607067352e-03
GC_11_1145 b_11 NI_11 NS_1145 0 7.2874261274710516e-03
GC_11_1146 b_11 NI_11 NS_1146 0 -4.1034637088346385e-03
GC_11_1147 b_11 NI_11 NS_1147 0 -8.5232818672608453e-03
GC_11_1148 b_11 NI_11 NS_1148 0 4.1574411160590413e-03
GC_11_1149 b_11 NI_11 NS_1149 0 4.8370640457207946e-03
GC_11_1150 b_11 NI_11 NS_1150 0 -3.8866661366854485e-03
GC_11_1151 b_11 NI_11 NS_1151 0 -2.3786683759336987e-03
GC_11_1152 b_11 NI_11 NS_1152 0 4.7281098936790599e-03
GC_11_1153 b_11 NI_11 NS_1153 0 7.0803227511905212e-03
GC_11_1154 b_11 NI_11 NS_1154 0 -7.3558597634443817e-03
GC_11_1155 b_11 NI_11 NS_1155 0 -7.0931606049231214e-03
GC_11_1156 b_11 NI_11 NS_1156 0 6.8359968044200683e-03
GC_11_1157 b_11 NI_11 NS_1157 0 1.6811452735812189e-03
GC_11_1158 b_11 NI_11 NS_1158 0 -5.3216374786754237e-03
GC_11_1159 b_11 NI_11 NS_1159 0 5.9853547441564932e-04
GC_11_1160 b_11 NI_11 NS_1160 0 5.4496391680694378e-03
GC_11_1161 b_11 NI_11 NS_1161 0 -4.1282284698505329e-09
GC_11_1162 b_11 NI_11 NS_1162 0 -1.3976315452962792e-08
GC_11_1163 b_11 NI_11 NS_1163 0 2.7262644697517518e-03
GC_11_1164 b_11 NI_11 NS_1164 0 -8.5984898986479295e-03
GC_11_1165 b_11 NI_11 NS_1165 0 8.7601838046849807e-04
GC_11_1166 b_11 NI_11 NS_1166 0 -3.4431550556227406e-03
GC_11_1167 b_11 NI_11 NS_1167 0 6.3792150906618727e-04
GC_11_1168 b_11 NI_11 NS_1168 0 4.0228568730467217e-03
GC_11_1169 b_11 NI_11 NS_1169 0 2.1875523767002363e-03
GC_11_1170 b_11 NI_11 NS_1170 0 -8.1664822243236544e-03
GC_11_1171 b_11 NI_11 NS_1171 0 -3.4772862845495302e-03
GC_11_1172 b_11 NI_11 NS_1172 0 6.9937176392018139e-03
GC_11_1173 b_11 NI_11 NS_1173 0 -8.5503704833711469e-08
GC_11_1174 b_11 NI_11 NS_1174 0 -3.1420277946797074e-07
GC_11_1175 b_11 NI_11 NS_1175 0 -7.9941562743269211e-03
GC_11_1176 b_11 NI_11 NS_1176 0 5.3784298215882745e-03
GC_11_1177 b_11 NI_11 NS_1177 0 4.1818213360578834e-03
GC_11_1178 b_11 NI_11 NS_1178 0 -6.8548439269165125e-03
GC_11_1179 b_11 NI_11 NS_1179 0 5.3337133249184909e-03
GC_11_1180 b_11 NI_11 NS_1180 0 7.4258456466223615e-04
GC_11_1181 b_11 NI_11 NS_1181 0 -2.3535041177445409e-03
GC_11_1182 b_11 NI_11 NS_1182 0 6.8399073945523744e-03
GC_11_1183 b_11 NI_11 NS_1183 0 -1.4841909516084726e-03
GC_11_1184 b_11 NI_11 NS_1184 0 -4.2255112741156082e-03
GC_11_1185 b_11 NI_11 NS_1185 0 2.3638870486139283e-03
GC_11_1186 b_11 NI_11 NS_1186 0 5.0284973850197104e-03
GC_11_1187 b_11 NI_11 NS_1187 0 -1.9828423316084615e-03
GC_11_1188 b_11 NI_11 NS_1188 0 -8.9598437125936823e-03
GC_11_1189 b_11 NI_11 NS_1189 0 -1.1185494524125716e-02
GC_11_1190 b_11 NI_11 NS_1190 0 8.4686186037579167e-09
GC_11_1191 b_11 NI_11 NS_1191 0 9.8720449475512484e-07
GC_11_1192 b_11 NI_11 NS_1192 0 3.6199551380031575e-05
GC_11_1193 b_11 NI_11 NS_1193 0 4.3663021223081496e-03
GC_11_1194 b_11 NI_11 NS_1194 0 -3.4896621308703429e-03
GC_11_1195 b_11 NI_11 NS_1195 0 -3.7149210583788529e-03
GC_11_1196 b_11 NI_11 NS_1196 0 6.2509193677475509e-03
GC_11_1197 b_11 NI_11 NS_1197 0 -8.7863563665941391e-03
GC_11_1198 b_11 NI_11 NS_1198 0 -5.9490013690354756e-03
GC_11_1199 b_11 NI_11 NS_1199 0 9.1761685454787908e-03
GC_11_1200 b_11 NI_11 NS_1200 0 -5.9808734151784778e-03
GC_11_1201 b_11 NI_11 NS_1201 0 7.1653413277863055e-03
GC_11_1202 b_11 NI_11 NS_1202 0 1.1911619373005486e-02
GC_11_1203 b_11 NI_11 NS_1203 0 -4.2323504151562316e-03
GC_11_1204 b_11 NI_11 NS_1204 0 -1.1251731252969932e-03
GC_11_1205 b_11 NI_11 NS_1205 0 -8.8793818740793614e-03
GC_11_1206 b_11 NI_11 NS_1206 0 -4.5103772678423419e-04
GC_11_1207 b_11 NI_11 NS_1207 0 1.4527710449907172e-02
GC_11_1208 b_11 NI_11 NS_1208 0 -1.0355589213584404e-02
GC_11_1209 b_11 NI_11 NS_1209 0 1.6511396692294768e-02
GC_11_1210 b_11 NI_11 NS_1210 0 4.0489420352340568e-03
GC_11_1211 b_11 NI_11 NS_1211 0 -1.1485124410396350e-02
GC_11_1212 b_11 NI_11 NS_1212 0 -1.9361272142187354e-04
GC_11_1213 b_11 NI_11 NS_1213 0 -1.6607747391134815e-02
GC_11_1214 b_11 NI_11 NS_1214 0 -4.4552720485059004e-02
GC_11_1215 b_11 NI_11 NS_1215 0 1.0667471198974914e-02
GC_11_1216 b_11 NI_11 NS_1216 0 1.0870814554198316e-03
GC_11_1217 b_11 NI_11 NS_1217 0 -4.8262938288978027e-02
GC_11_1218 b_11 NI_11 NS_1218 0 1.1004755311070350e-02
GC_11_1219 b_11 NI_11 NS_1219 0 -1.0464750274727421e-02
GC_11_1220 b_11 NI_11 NS_1220 0 5.4279680459603131e-04
GC_11_1221 b_11 NI_11 NS_1221 0 9.7653617581287856e-03
GC_11_1222 b_11 NI_11 NS_1222 0 -6.1129050456819572e-04
GC_11_1223 b_11 NI_11 NS_1223 0 4.5934349138384836e-03
GC_11_1224 b_11 NI_11 NS_1224 0 2.4194432162358351e-02
GC_11_1225 b_11 NI_11 NS_1225 0 -1.0736734333668318e-02
GC_11_1226 b_11 NI_11 NS_1226 0 1.9986348693273401e-03
GC_11_1227 b_11 NI_11 NS_1227 0 -8.4712998928282660e-03
GC_11_1228 b_11 NI_11 NS_1228 0 -1.3526363934167035e-02
GC_11_1229 b_11 NI_11 NS_1229 0 1.0155213247613265e-02
GC_11_1230 b_11 NI_11 NS_1230 0 9.6273171588178374e-04
GC_11_1231 b_11 NI_11 NS_1231 0 -1.9169420481953792e-02
GC_11_1232 b_11 NI_11 NS_1232 0 2.8673858330776330e-02
GC_11_1233 b_11 NI_11 NS_1233 0 -9.6256432137190474e-03
GC_11_1234 b_11 NI_11 NS_1234 0 -9.4348403335027487e-04
GC_11_1235 b_11 NI_11 NS_1235 0 1.8844340690093910e-03
GC_11_1236 b_11 NI_11 NS_1236 0 -1.3764811854074593e-03
GC_11_1237 b_11 NI_11 NS_1237 0 9.4635441062029240e-03
GC_11_1238 b_11 NI_11 NS_1238 0 -2.5486159515625452e-04
GC_11_1239 b_11 NI_11 NS_1239 0 -1.6535666022074881e-04
GC_11_1240 b_11 NI_11 NS_1240 0 3.0293307879733885e-02
GC_11_1241 b_11 NI_11 NS_1241 0 -8.5338141894666462e-03
GC_11_1242 b_11 NI_11 NS_1242 0 1.7750721830360841e-04
GC_11_1243 b_11 NI_11 NS_1243 0 2.1345391530945820e-04
GC_11_1244 b_11 NI_11 NS_1244 0 -5.4660285435324850e-03
GC_11_1245 b_11 NI_11 NS_1245 0 1.0030295022920585e-02
GC_11_1246 b_11 NI_11 NS_1246 0 -3.4496677931850393e-04
GC_11_1247 b_11 NI_11 NS_1247 0 8.9347314409424384e-03
GC_11_1248 b_11 NI_11 NS_1248 0 2.6406165044669118e-02
GC_11_1249 b_11 NI_11 NS_1249 0 -8.3546158718499301e-03
GC_11_1250 b_11 NI_11 NS_1250 0 1.4014780997477060e-03
GC_11_1251 b_11 NI_11 NS_1251 0 -2.5783439624136499e-03
GC_11_1252 b_11 NI_11 NS_1252 0 -7.3352797107030165e-03
GC_11_1253 b_11 NI_11 NS_1253 0 1.0543947422337586e-02
GC_11_1254 b_11 NI_11 NS_1254 0 -8.2792792755577666e-04
GC_11_1255 b_11 NI_11 NS_1255 0 1.4465689156419615e-02
GC_11_1256 b_11 NI_11 NS_1256 0 1.9992679090169524e-02
GC_11_1257 b_11 NI_11 NS_1257 0 -8.2668446234042160e-03
GC_11_1258 b_11 NI_11 NS_1258 0 2.9582400394920151e-03
GC_11_1259 b_11 NI_11 NS_1259 0 -5.5757319204505469e-03
GC_11_1260 b_11 NI_11 NS_1260 0 -6.9085922649490487e-03
GC_11_1261 b_11 NI_11 NS_1261 0 1.1230552140982300e-02
GC_11_1262 b_11 NI_11 NS_1262 0 -1.3725286175495623e-03
GC_11_1263 b_11 NI_11 NS_1263 0 1.5750291612864831e-02
GC_11_1264 b_11 NI_11 NS_1264 0 1.2967909579440683e-02
GC_11_1265 b_11 NI_11 NS_1265 0 -7.1659126163396156e-03
GC_11_1266 b_11 NI_11 NS_1266 0 5.1306008712621587e-03
GC_11_1267 b_11 NI_11 NS_1267 0 -6.8667054411296682e-03
GC_11_1268 b_11 NI_11 NS_1268 0 -4.8393396709037568e-03
GC_11_1269 b_11 NI_11 NS_1269 0 5.3089333333566265e-09
GC_11_1270 b_11 NI_11 NS_1270 0 4.4273840572322334e-08
GC_11_1271 b_11 NI_11 NS_1271 0 1.2002193431557647e-02
GC_11_1272 b_11 NI_11 NS_1272 0 -2.5686775917577857e-03
GC_11_1273 b_11 NI_11 NS_1273 0 -5.2367615751036196e-03
GC_11_1274 b_11 NI_11 NS_1274 0 4.7118182241628458e-03
GC_11_1275 b_11 NI_11 NS_1275 0 -6.1526710133823926e-03
GC_11_1276 b_11 NI_11 NS_1276 0 -4.3194207809051748e-03
GC_11_1277 b_11 NI_11 NS_1277 0 1.1768582397129714e-02
GC_11_1278 b_11 NI_11 NS_1278 0 -3.7146148516987903e-03
GC_11_1279 b_11 NI_11 NS_1279 0 1.3012629149799785e-02
GC_11_1280 b_11 NI_11 NS_1280 0 9.4653996569115679e-03
GC_11_1281 b_11 NI_11 NS_1281 0 3.9556754391074373e-06
GC_11_1282 b_11 NI_11 NS_1282 0 -9.4250559951816273e-07
GC_11_1283 b_11 NI_11 NS_1283 0 1.6124344536998774e-02
GC_11_1284 b_11 NI_11 NS_1284 0 1.6774826179895359e-02
GC_11_1285 b_11 NI_11 NS_1285 0 1.2055185343034550e-02
GC_11_1286 b_11 NI_11 NS_1286 0 -2.4727519594803819e-03
GC_11_1287 b_11 NI_11 NS_1287 0 -8.3469674952299389e-03
GC_11_1288 b_11 NI_11 NS_1288 0 8.5427821804031219e-05
GC_11_1289 b_11 NI_11 NS_1289 0 1.1349989965456296e-02
GC_11_1290 b_11 NI_11 NS_1290 0 7.3343074359889160e-03
GC_11_1291 b_11 NI_11 NS_1291 0 -4.6479068826677005e-03
GC_11_1292 b_11 NI_11 NS_1292 0 7.3636007418352552e-03
GC_11_1293 b_11 NI_11 NS_1293 0 -8.0750669090293783e-03
GC_11_1294 b_11 NI_11 NS_1294 0 -3.7254240451645485e-03
GC_11_1295 b_11 NI_11 NS_1295 0 1.5991411392139065e-02
GC_11_1296 b_11 NI_11 NS_1296 0 -7.7330084568801929e-03
GD_11_1 b_11 NI_11 NA_1 0 -2.2825069216537529e-06
GD_11_2 b_11 NI_11 NA_2 0 3.3590091094541810e-06
GD_11_3 b_11 NI_11 NA_3 0 -1.1565261946105435e-06
GD_11_4 b_11 NI_11 NA_4 0 8.8115152206316316e-06
GD_11_5 b_11 NI_11 NA_5 0 -2.9989183592912845e-06
GD_11_6 b_11 NI_11 NA_6 0 1.1439025780031576e-05
GD_11_7 b_11 NI_11 NA_7 0 3.1120406317218751e-06
GD_11_8 b_11 NI_11 NA_8 0 1.9066305826389776e-05
GD_11_9 b_11 NI_11 NA_9 0 1.0616252270114097e-02
GD_11_10 b_11 NI_11 NA_10 0 -1.1524162798605623e-03
GD_11_11 b_11 NI_11 NA_11 0 -1.0697627223894524e-02
GD_11_12 b_11 NI_11 NA_12 0 -4.9158970113934615e-03
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -2.9908308283269252e-05
GC_12_2 b_12 NI_12 NS_2 0 1.1048173540809494e-11
GC_12_3 b_12 NI_12 NS_3 0 -3.3938218059982685e-11
GC_12_4 b_12 NI_12 NS_4 0 2.1486379362083075e-10
GC_12_5 b_12 NI_12 NS_5 0 -4.0816364993404327e-07
GC_12_6 b_12 NI_12 NS_6 0 -2.7824141374906197e-07
GC_12_7 b_12 NI_12 NS_7 0 -1.0588668299743217e-07
GC_12_8 b_12 NI_12 NS_8 0 5.6550159263727485e-07
GC_12_9 b_12 NI_12 NS_9 0 2.3813316128924577e-07
GC_12_10 b_12 NI_12 NS_10 0 1.4039366221435538e-06
GC_12_11 b_12 NI_12 NS_11 0 1.1109692628170049e-06
GC_12_12 b_12 NI_12 NS_12 0 -3.7454403359547389e-07
GC_12_13 b_12 NI_12 NS_13 0 6.7784208369940567e-07
GC_12_14 b_12 NI_12 NS_14 0 -2.0281306696597115e-06
GC_12_15 b_12 NI_12 NS_15 0 -6.4680828222347754e-07
GC_12_16 b_12 NI_12 NS_16 0 2.8098249443086132e-07
GC_12_17 b_12 NI_12 NS_17 0 9.9940404903472908e-07
GC_12_18 b_12 NI_12 NS_18 0 6.6416435045734802e-07
GC_12_19 b_12 NI_12 NS_19 0 3.8974634508379906e-06
GC_12_20 b_12 NI_12 NS_20 0 -3.7311332574595683e-06
GC_12_21 b_12 NI_12 NS_21 0 -5.5969139605498052e-06
GC_12_22 b_12 NI_12 NS_22 0 -3.8629281967753817e-06
GC_12_23 b_12 NI_12 NS_23 0 -9.2017089514861276e-07
GC_12_24 b_12 NI_12 NS_24 0 -2.0450961424972531e-06
GC_12_25 b_12 NI_12 NS_25 0 -1.3600395241286685e-05
GC_12_26 b_12 NI_12 NS_26 0 5.3801221444912302e-06
GC_12_27 b_12 NI_12 NS_27 0 -5.3844130551922592e-07
GC_12_28 b_12 NI_12 NS_28 0 1.8937669959129984e-06
GC_12_29 b_12 NI_12 NS_29 0 7.8173254212640417e-07
GC_12_30 b_12 NI_12 NS_30 0 1.9309071374193838e-05
GC_12_31 b_12 NI_12 NS_31 0 2.7666945324019948e-06
GC_12_32 b_12 NI_12 NS_32 0 -4.5945379370158739e-06
GC_12_33 b_12 NI_12 NS_33 0 1.4653352659085446e-06
GC_12_34 b_12 NI_12 NS_34 0 1.7112794182573986e-06
GC_12_35 b_12 NI_12 NS_35 0 5.3166454903538502e-06
GC_12_36 b_12 NI_12 NS_36 0 -2.2410339501592307e-06
GC_12_37 b_12 NI_12 NS_37 0 -4.1276253296980854e-07
GC_12_38 b_12 NI_12 NS_38 0 -8.1224414459574651e-07
GC_12_39 b_12 NI_12 NS_39 0 -2.0565674354446983e-06
GC_12_40 b_12 NI_12 NS_40 0 2.3251974245262744e-06
GC_12_41 b_12 NI_12 NS_41 0 -3.0284610411362951e-08
GC_12_42 b_12 NI_12 NS_42 0 1.2397139387340766e-06
GC_12_43 b_12 NI_12 NS_43 0 5.2803295195043794e-06
GC_12_44 b_12 NI_12 NS_44 0 5.9467789494476427e-06
GC_12_45 b_12 NI_12 NS_45 0 1.4516661708037675e-06
GC_12_46 b_12 NI_12 NS_46 0 -1.0225314191849334e-06
GC_12_47 b_12 NI_12 NS_47 0 1.1386267894193876e-07
GC_12_48 b_12 NI_12 NS_48 0 -4.7253327233220491e-08
GC_12_49 b_12 NI_12 NS_49 0 5.0776027836679062e-07
GC_12_50 b_12 NI_12 NS_50 0 7.4654371741186156e-07
GC_12_51 b_12 NI_12 NS_51 0 6.0590689630892844e-06
GC_12_52 b_12 NI_12 NS_52 0 4.9646009212560059e-07
GC_12_53 b_12 NI_12 NS_53 0 5.5787748303254845e-07
GC_12_54 b_12 NI_12 NS_54 0 -8.6741898289039053e-07
GC_12_55 b_12 NI_12 NS_55 0 -1.2579210010159833e-07
GC_12_56 b_12 NI_12 NS_56 0 -3.6412120096354796e-08
GC_12_57 b_12 NI_12 NS_57 0 6.7967541992552200e-07
GC_12_58 b_12 NI_12 NS_58 0 8.5001181624839378e-07
GC_12_59 b_12 NI_12 NS_59 0 4.7885001273011068e-06
GC_12_60 b_12 NI_12 NS_60 0 -1.9381642210765248e-06
GC_12_61 b_12 NI_12 NS_61 0 1.3610293356760068e-07
GC_12_62 b_12 NI_12 NS_62 0 -7.2191733622202461e-07
GC_12_63 b_12 NI_12 NS_63 0 -1.2100901839712511e-07
GC_12_64 b_12 NI_12 NS_64 0 1.4828001789434197e-07
GC_12_65 b_12 NI_12 NS_65 0 9.4361580215653380e-07
GC_12_66 b_12 NI_12 NS_66 0 7.7731499327880812e-07
GC_12_67 b_12 NI_12 NS_67 0 2.7625393319042512e-06
GC_12_68 b_12 NI_12 NS_68 0 -3.0182467186098201e-06
GC_12_69 b_12 NI_12 NS_69 0 -1.0350699916584301e-07
GC_12_70 b_12 NI_12 NS_70 0 -4.8431896002293281e-07
GC_12_71 b_12 NI_12 NS_71 0 8.8977041661690617e-08
GC_12_72 b_12 NI_12 NS_72 0 2.0122410939866315e-07
GC_12_73 b_12 NI_12 NS_73 0 1.3138870181488878e-06
GC_12_74 b_12 NI_12 NS_74 0 5.1136158109649999e-07
GC_12_75 b_12 NI_12 NS_75 0 6.6546486260816715e-07
GC_12_76 b_12 NI_12 NS_76 0 -2.7705902449473729e-06
GC_12_77 b_12 NI_12 NS_77 0 -1.6499126488710237e-07
GC_12_78 b_12 NI_12 NS_78 0 -1.3966003970949140e-07
GC_12_79 b_12 NI_12 NS_79 0 2.2753950993271449e-07
GC_12_80 b_12 NI_12 NS_80 0 2.2630097424705945e-08
GC_12_81 b_12 NI_12 NS_81 0 1.6153036721853026e-12
GC_12_82 b_12 NI_12 NS_82 0 -6.1873191819603745e-12
GC_12_83 b_12 NI_12 NS_83 0 9.8103391432875826e-07
GC_12_84 b_12 NI_12 NS_84 0 -2.6426563813257424e-07
GC_12_85 b_12 NI_12 NS_85 0 -2.6851599613503260e-08
GC_12_86 b_12 NI_12 NS_86 0 4.9058529446703466e-08
GC_12_87 b_12 NI_12 NS_87 0 2.6314603700900798e-07
GC_12_88 b_12 NI_12 NS_88 0 1.1131715246372510e-08
GC_12_89 b_12 NI_12 NS_89 0 8.3328248479611782e-07
GC_12_90 b_12 NI_12 NS_90 0 -1.5920398283180220e-07
GC_12_91 b_12 NI_12 NS_91 0 -6.3068305813627861e-08
GC_12_92 b_12 NI_12 NS_92 0 -1.0947688784176443e-06
GC_12_93 b_12 NI_12 NS_93 0 7.6565874706255864e-11
GC_12_94 b_12 NI_12 NS_94 0 -1.9341066387631476e-10
GC_12_95 b_12 NI_12 NS_95 0 6.8042410224498655e-07
GC_12_96 b_12 NI_12 NS_96 0 -4.3030921083856372e-07
GC_12_97 b_12 NI_12 NS_97 0 4.2741780312399114e-07
GC_12_98 b_12 NI_12 NS_98 0 1.6120754430470254e-07
GC_12_99 b_12 NI_12 NS_99 0 1.4000314499101302e-07
GC_12_100 b_12 NI_12 NS_100 0 -8.2544234649855287e-08
GC_12_101 b_12 NI_12 NS_101 0 -1.4336330734690823e-07
GC_12_102 b_12 NI_12 NS_102 0 -6.7656483380121071e-07
GC_12_103 b_12 NI_12 NS_103 0 2.4259164645976997e-08
GC_12_104 b_12 NI_12 NS_104 0 2.3623504650132027e-07
GC_12_105 b_12 NI_12 NS_105 0 3.3298168142640307e-07
GC_12_106 b_12 NI_12 NS_106 0 -5.5339528610347338e-08
GC_12_107 b_12 NI_12 NS_107 0 4.0223423018619003e-07
GC_12_108 b_12 NI_12 NS_108 0 2.2651226649919812e-07
GC_12_109 b_12 NI_12 NS_109 0 1.0245384404630774e-05
GC_12_110 b_12 NI_12 NS_110 0 -4.7958086898930480e-12
GC_12_111 b_12 NI_12 NS_111 0 1.0352309461950196e-11
GC_12_112 b_12 NI_12 NS_112 0 3.7845449610601450e-10
GC_12_113 b_12 NI_12 NS_113 0 1.3513075199069558e-07
GC_12_114 b_12 NI_12 NS_114 0 1.0761869496418302e-07
GC_12_115 b_12 NI_12 NS_115 0 7.2008558191804797e-07
GC_12_116 b_12 NI_12 NS_116 0 -1.8726846770164046e-07
GC_12_117 b_12 NI_12 NS_117 0 -5.9812723150028692e-07
GC_12_118 b_12 NI_12 NS_118 0 -3.6307216105321621e-07
GC_12_119 b_12 NI_12 NS_119 0 1.3990038002423072e-06
GC_12_120 b_12 NI_12 NS_120 0 3.2530789789579805e-07
GC_12_121 b_12 NI_12 NS_121 0 -9.9970740420730507e-07
GC_12_122 b_12 NI_12 NS_122 0 -1.7789826492041437e-06
GC_12_123 b_12 NI_12 NS_123 0 2.5546169533659966e-07
GC_12_124 b_12 NI_12 NS_124 0 -5.4933178491233411e-09
GC_12_125 b_12 NI_12 NS_125 0 -8.7355623778937812e-07
GC_12_126 b_12 NI_12 NS_126 0 9.7895590821232403e-08
GC_12_127 b_12 NI_12 NS_127 0 2.5713369073814609e-06
GC_12_128 b_12 NI_12 NS_128 0 -1.1144097462074228e-06
GC_12_129 b_12 NI_12 NS_129 0 -3.9893100381186205e-06
GC_12_130 b_12 NI_12 NS_130 0 -2.3993359556128026e-07
GC_12_131 b_12 NI_12 NS_131 0 1.2124331027131517e-08
GC_12_132 b_12 NI_12 NS_132 0 1.6053661670610441e-06
GC_12_133 b_12 NI_12 NS_133 0 -8.3049194707182695e-07
GC_12_134 b_12 NI_12 NS_134 0 -2.6088802721510371e-06
GC_12_135 b_12 NI_12 NS_135 0 -7.8261936086596928e-07
GC_12_136 b_12 NI_12 NS_136 0 1.4932796965177986e-06
GC_12_137 b_12 NI_12 NS_137 0 5.8169705763869936e-07
GC_12_138 b_12 NI_12 NS_138 0 -3.0275525567298420e-06
GC_12_139 b_12 NI_12 NS_139 0 -1.4470917318015723e-06
GC_12_140 b_12 NI_12 NS_140 0 2.5662110033098771e-06
GC_12_141 b_12 NI_12 NS_141 0 2.3925480355137184e-07
GC_12_142 b_12 NI_12 NS_142 0 1.2705008299398183e-06
GC_12_143 b_12 NI_12 NS_143 0 -6.9734424876236944e-07
GC_12_144 b_12 NI_12 NS_144 0 -1.1693055761169895e-06
GC_12_145 b_12 NI_12 NS_145 0 -5.8085669477923509e-08
GC_12_146 b_12 NI_12 NS_146 0 1.0861710535558090e-06
GC_12_147 b_12 NI_12 NS_147 0 -6.5279075157651332e-07
GC_12_148 b_12 NI_12 NS_148 0 -7.6713158350068545e-07
GC_12_149 b_12 NI_12 NS_149 0 -5.1252986170164913e-07
GC_12_150 b_12 NI_12 NS_150 0 1.1060675340061559e-06
GC_12_151 b_12 NI_12 NS_151 0 4.4998916324480208e-08
GC_12_152 b_12 NI_12 NS_152 0 -8.8827920477425681e-07
GC_12_153 b_12 NI_12 NS_153 0 -9.1171402200195615e-07
GC_12_154 b_12 NI_12 NS_154 0 1.0678813774245165e-06
GC_12_155 b_12 NI_12 NS_155 0 -1.1158381734244404e-07
GC_12_156 b_12 NI_12 NS_156 0 7.9073132599578623e-09
GC_12_157 b_12 NI_12 NS_157 0 -3.3925157274094441e-07
GC_12_158 b_12 NI_12 NS_158 0 1.0187616796942840e-06
GC_12_159 b_12 NI_12 NS_159 0 -9.8166416343981874e-08
GC_12_160 b_12 NI_12 NS_160 0 1.1223304809720684e-07
GC_12_161 b_12 NI_12 NS_161 0 -3.0039650626792652e-07
GC_12_162 b_12 NI_12 NS_162 0 1.0059098579077405e-06
GC_12_163 b_12 NI_12 NS_163 0 8.0883148799485856e-08
GC_12_164 b_12 NI_12 NS_164 0 1.6439738303657139e-07
GC_12_165 b_12 NI_12 NS_165 0 -7.9044586517807623e-08
GC_12_166 b_12 NI_12 NS_166 0 1.1304480354768347e-06
GC_12_167 b_12 NI_12 NS_167 0 7.8461435070644521e-07
GC_12_168 b_12 NI_12 NS_168 0 -9.7572305952092197e-09
GC_12_169 b_12 NI_12 NS_169 0 8.4840744903802627e-08
GC_12_170 b_12 NI_12 NS_170 0 8.2101370224998685e-07
GC_12_171 b_12 NI_12 NS_171 0 3.1724417523711153e-07
GC_12_172 b_12 NI_12 NS_172 0 -1.9309453384819957e-07
GC_12_173 b_12 NI_12 NS_173 0 1.9072403262677129e-07
GC_12_174 b_12 NI_12 NS_174 0 1.0069310513740895e-06
GC_12_175 b_12 NI_12 NS_175 0 7.9530355784778524e-07
GC_12_176 b_12 NI_12 NS_176 0 -8.1778190577547437e-07
GC_12_177 b_12 NI_12 NS_177 0 3.2998220700329242e-07
GC_12_178 b_12 NI_12 NS_178 0 5.3262075283100538e-07
GC_12_179 b_12 NI_12 NS_179 0 -5.5954544162640607e-09
GC_12_180 b_12 NI_12 NS_180 0 -5.5296179046156724e-07
GC_12_181 b_12 NI_12 NS_181 0 4.5645173017769223e-07
GC_12_182 b_12 NI_12 NS_182 0 7.5300499817303438e-07
GC_12_183 b_12 NI_12 NS_183 0 -9.7866833983831847e-09
GC_12_184 b_12 NI_12 NS_184 0 -1.1013782684622823e-06
GC_12_185 b_12 NI_12 NS_185 0 3.1840043588340357e-07
GC_12_186 b_12 NI_12 NS_186 0 1.0305571075247319e-07
GC_12_187 b_12 NI_12 NS_187 0 -3.9308083154777316e-07
GC_12_188 b_12 NI_12 NS_188 0 -2.5353161545497120e-07
GC_12_189 b_12 NI_12 NS_189 0 1.4514761109395593e-12
GC_12_190 b_12 NI_12 NS_190 0 3.4002813665460301e-12
GC_12_191 b_12 NI_12 NS_191 0 3.9031448575710031e-07
GC_12_192 b_12 NI_12 NS_192 0 2.2952278612250100e-07
GC_12_193 b_12 NI_12 NS_193 0 1.1980138916968885e-07
GC_12_194 b_12 NI_12 NS_194 0 3.5452828361116567e-08
GC_12_195 b_12 NI_12 NS_195 0 -2.7884433894126043e-07
GC_12_196 b_12 NI_12 NS_196 0 -1.0897418227891816e-07
GC_12_197 b_12 NI_12 NS_197 0 3.2155753507775708e-07
GC_12_198 b_12 NI_12 NS_198 0 6.8216846624471697e-08
GC_12_199 b_12 NI_12 NS_199 0 -3.5584826363071270e-07
GC_12_200 b_12 NI_12 NS_200 0 -4.5135908231720298e-07
GC_12_201 b_12 NI_12 NS_201 0 -1.0584501395268609e-11
GC_12_202 b_12 NI_12 NS_202 0 3.2224644855529587e-10
GC_12_203 b_12 NI_12 NS_203 0 1.8885747801591307e-07
GC_12_204 b_12 NI_12 NS_204 0 -1.9033767453443507e-07
GC_12_205 b_12 NI_12 NS_205 0 -7.7180684285495896e-08
GC_12_206 b_12 NI_12 NS_206 0 3.9129239796736781e-07
GC_12_207 b_12 NI_12 NS_207 0 -1.7579626606763519e-07
GC_12_208 b_12 NI_12 NS_208 0 6.2408386104207005e-08
GC_12_209 b_12 NI_12 NS_209 0 -5.3348776636385670e-07
GC_12_210 b_12 NI_12 NS_210 0 -2.6042276745339723e-07
GC_12_211 b_12 NI_12 NS_211 0 5.9192787821755791e-08
GC_12_212 b_12 NI_12 NS_212 0 2.3074531720752467e-08
GC_12_213 b_12 NI_12 NS_213 0 -3.6617441544311378e-07
GC_12_214 b_12 NI_12 NS_214 0 6.6095576344680333e-08
GC_12_215 b_12 NI_12 NS_215 0 1.0697296130329235e-07
GC_12_216 b_12 NI_12 NS_216 0 3.2656863132434655e-07
GC_12_217 b_12 NI_12 NS_217 0 -6.4297366535075347e-05
GC_12_218 b_12 NI_12 NS_218 0 3.5514016371861566e-12
GC_12_219 b_12 NI_12 NS_219 0 5.0206553205357999e-11
GC_12_220 b_12 NI_12 NS_220 0 -1.5827692919046583e-09
GC_12_221 b_12 NI_12 NS_221 0 -1.0722886831006487e-06
GC_12_222 b_12 NI_12 NS_222 0 -1.0608543919763111e-06
GC_12_223 b_12 NI_12 NS_223 0 4.1036495344070129e-07
GC_12_224 b_12 NI_12 NS_224 0 3.5893531559271280e-07
GC_12_225 b_12 NI_12 NS_225 0 -2.2645987651145391e-06
GC_12_226 b_12 NI_12 NS_226 0 2.1075670721265009e-06
GC_12_227 b_12 NI_12 NS_227 0 -2.5340359916088536e-06
GC_12_228 b_12 NI_12 NS_228 0 -1.2433597079180271e-06
GC_12_229 b_12 NI_12 NS_229 0 1.3996057841419902e-06
GC_12_230 b_12 NI_12 NS_230 0 1.0022268169338159e-06
GC_12_231 b_12 NI_12 NS_231 0 -1.1248383720959314e-06
GC_12_232 b_12 NI_12 NS_232 0 1.3421367723413611e-06
GC_12_233 b_12 NI_12 NS_233 0 7.2530490180211072e-07
GC_12_234 b_12 NI_12 NS_234 0 3.0434984189872679e-06
GC_12_235 b_12 NI_12 NS_235 0 -2.8542570037330506e-06
GC_12_236 b_12 NI_12 NS_236 0 4.6955320129147800e-07
GC_12_237 b_12 NI_12 NS_237 0 3.6961788499331238e-06
GC_12_238 b_12 NI_12 NS_238 0 -2.0129350650978546e-06
GC_12_239 b_12 NI_12 NS_239 0 -1.9022140444644733e-07
GC_12_240 b_12 NI_12 NS_240 0 2.5688420718478661e-06
GC_12_241 b_12 NI_12 NS_241 0 -4.0608194886404184e-06
GC_12_242 b_12 NI_12 NS_242 0 4.8419302175124820e-06
GC_12_243 b_12 NI_12 NS_243 0 6.4547334345840213e-07
GC_12_244 b_12 NI_12 NS_244 0 -1.5900979692806419e-06
GC_12_245 b_12 NI_12 NS_245 0 4.6199372018076664e-06
GC_12_246 b_12 NI_12 NS_246 0 9.9424702866576212e-06
GC_12_247 b_12 NI_12 NS_247 0 -1.1565097154190526e-07
GC_12_248 b_12 NI_12 NS_248 0 5.2802458194921125e-07
GC_12_249 b_12 NI_12 NS_249 0 -6.9412657139212465e-09
GC_12_250 b_12 NI_12 NS_250 0 -7.8937892784184055e-07
GC_12_251 b_12 NI_12 NS_251 0 5.3542050048511507e-06
GC_12_252 b_12 NI_12 NS_252 0 4.9603750183075327e-07
GC_12_253 b_12 NI_12 NS_253 0 8.4753909293221891e-07
GC_12_254 b_12 NI_12 NS_254 0 1.9215375669305231e-06
GC_12_255 b_12 NI_12 NS_255 0 3.1609111135799572e-08
GC_12_256 b_12 NI_12 NS_256 0 1.1340689936498478e-06
GC_12_257 b_12 NI_12 NS_257 0 5.8568420727782189e-07
GC_12_258 b_12 NI_12 NS_258 0 -1.1142479091866034e-06
GC_12_259 b_12 NI_12 NS_259 0 5.8308363336396036e-06
GC_12_260 b_12 NI_12 NS_260 0 4.0738902138662810e-06
GC_12_261 b_12 NI_12 NS_261 0 6.0565364367944627e-07
GC_12_262 b_12 NI_12 NS_262 0 8.6242662587099552e-07
GC_12_263 b_12 NI_12 NS_263 0 1.9670984273352569e-07
GC_12_264 b_12 NI_12 NS_264 0 2.4104962017342846e-07
GC_12_265 b_12 NI_12 NS_265 0 8.4506095715150201e-07
GC_12_266 b_12 NI_12 NS_266 0 -6.7479285700615000e-07
GC_12_267 b_12 NI_12 NS_267 0 6.6692109803496671e-06
GC_12_268 b_12 NI_12 NS_268 0 7.5284978258272963e-07
GC_12_269 b_12 NI_12 NS_269 0 7.7512776237498446e-07
GC_12_270 b_12 NI_12 NS_270 0 7.5176623339266124e-07
GC_12_271 b_12 NI_12 NS_271 0 6.6484584739138983e-07
GC_12_272 b_12 NI_12 NS_272 0 -6.6045956142058920e-08
GC_12_273 b_12 NI_12 NS_273 0 8.7116245143633724e-07
GC_12_274 b_12 NI_12 NS_274 0 -6.4327720864918263e-07
GC_12_275 b_12 NI_12 NS_275 0 5.7782974674076393e-06
GC_12_276 b_12 NI_12 NS_276 0 -1.5930532474102947e-06
GC_12_277 b_12 NI_12 NS_277 0 8.2495561780508669e-07
GC_12_278 b_12 NI_12 NS_278 0 5.6932309669587052e-07
GC_12_279 b_12 NI_12 NS_279 0 6.2572602331385054e-07
GC_12_280 b_12 NI_12 NS_280 0 -5.5366802404506622e-07
GC_12_281 b_12 NI_12 NS_281 0 9.3725662648135485e-07
GC_12_282 b_12 NI_12 NS_282 0 -4.4872611125991253e-07
GC_12_283 b_12 NI_12 NS_283 0 3.9054998493424079e-06
GC_12_284 b_12 NI_12 NS_284 0 -2.9926146333458643e-06
GC_12_285 b_12 NI_12 NS_285 0 8.9724230469366842e-07
GC_12_286 b_12 NI_12 NS_286 0 3.2914693338498637e-07
GC_12_287 b_12 NI_12 NS_287 0 2.1534477383111749e-07
GC_12_288 b_12 NI_12 NS_288 0 -7.9633570207421885e-07
GC_12_289 b_12 NI_12 NS_289 0 1.1591912790832257e-06
GC_12_290 b_12 NI_12 NS_290 0 -3.2770069884350658e-07
GC_12_291 b_12 NI_12 NS_291 0 1.6782804201072562e-06
GC_12_292 b_12 NI_12 NS_292 0 -3.0911832874895768e-06
GC_12_293 b_12 NI_12 NS_293 0 7.9264169288315115e-07
GC_12_294 b_12 NI_12 NS_294 0 -1.0570353196085972e-07
GC_12_295 b_12 NI_12 NS_295 0 -1.9831590631654904e-07
GC_12_296 b_12 NI_12 NS_296 0 -4.0880849653195280e-07
GC_12_297 b_12 NI_12 NS_297 0 8.5890294943204728e-12
GC_12_298 b_12 NI_12 NS_298 0 -1.5740028401212552e-11
GC_12_299 b_12 NI_12 NS_299 0 8.3767168870467989e-07
GC_12_300 b_12 NI_12 NS_300 0 -5.9584682000669334e-07
GC_12_301 b_12 NI_12 NS_301 0 4.9537139012050847e-07
GC_12_302 b_12 NI_12 NS_302 0 -3.5565658234497431e-08
GC_12_303 b_12 NI_12 NS_303 0 1.6374995883127375e-08
GC_12_304 b_12 NI_12 NS_304 0 -8.9211613098687905e-08
GC_12_305 b_12 NI_12 NS_305 0 5.2071495002713678e-07
GC_12_306 b_12 NI_12 NS_306 0 -1.9284795423156731e-08
GC_12_307 b_12 NI_12 NS_307 0 7.0591054134169045e-07
GC_12_308 b_12 NI_12 NS_308 0 -1.5618082149018196e-06
GC_12_309 b_12 NI_12 NS_309 0 4.0958074137665253e-10
GC_12_310 b_12 NI_12 NS_310 0 -5.8094827353468171e-10
GC_12_311 b_12 NI_12 NS_311 0 1.0094277139276271e-06
GC_12_312 b_12 NI_12 NS_312 0 -2.7418518950582744e-07
GC_12_313 b_12 NI_12 NS_313 0 3.5391653606174067e-07
GC_12_314 b_12 NI_12 NS_314 0 -1.7487827155448464e-07
GC_12_315 b_12 NI_12 NS_315 0 2.5450016463877615e-07
GC_12_316 b_12 NI_12 NS_316 0 2.6674106577062691e-08
GC_12_317 b_12 NI_12 NS_317 0 1.0861129095685798e-06
GC_12_318 b_12 NI_12 NS_318 0 -1.1751149806845368e-06
GC_12_319 b_12 NI_12 NS_319 0 6.5444352488527654e-07
GC_12_320 b_12 NI_12 NS_320 0 -3.3449202110413264e-07
GC_12_321 b_12 NI_12 NS_321 0 -2.1289909954357518e-07
GC_12_322 b_12 NI_12 NS_322 0 -9.8626578360886055e-08
GC_12_323 b_12 NI_12 NS_323 0 7.5675761632252991e-07
GC_12_324 b_12 NI_12 NS_324 0 3.2207336586815541e-07
GC_12_325 b_12 NI_12 NS_325 0 8.6499750905509579e-06
GC_12_326 b_12 NI_12 NS_326 0 3.7611015403305126e-12
GC_12_327 b_12 NI_12 NS_327 0 -7.8508174662210827e-11
GC_12_328 b_12 NI_12 NS_328 0 2.5460397943689245e-09
GC_12_329 b_12 NI_12 NS_329 0 1.6514149959350005e-08
GC_12_330 b_12 NI_12 NS_330 0 -8.5494772205289571e-08
GC_12_331 b_12 NI_12 NS_331 0 -2.4857702652703282e-07
GC_12_332 b_12 NI_12 NS_332 0 2.6957995437593662e-07
GC_12_333 b_12 NI_12 NS_333 0 7.4441977713083533e-07
GC_12_334 b_12 NI_12 NS_334 0 -2.8507168972557434e-07
GC_12_335 b_12 NI_12 NS_335 0 -9.6886912610851696e-07
GC_12_336 b_12 NI_12 NS_336 0 -2.4196027924961805e-07
GC_12_337 b_12 NI_12 NS_337 0 1.0238386459143066e-06
GC_12_338 b_12 NI_12 NS_338 0 4.0092189553025757e-07
GC_12_339 b_12 NI_12 NS_339 0 -1.2005330360298715e-07
GC_12_340 b_12 NI_12 NS_340 0 -2.7540980813207535e-07
GC_12_341 b_12 NI_12 NS_341 0 1.0875946395573116e-07
GC_12_342 b_12 NI_12 NS_342 0 -5.1234282439472653e-07
GC_12_343 b_12 NI_12 NS_343 0 -2.0908859846863946e-06
GC_12_344 b_12 NI_12 NS_344 0 8.5580353729393054e-07
GC_12_345 b_12 NI_12 NS_345 0 2.4337653047647084e-06
GC_12_346 b_12 NI_12 NS_346 0 -6.0045401999150212e-07
GC_12_347 b_12 NI_12 NS_347 0 -6.6288728094609394e-07
GC_12_348 b_12 NI_12 NS_348 0 -1.4012568159388151e-06
GC_12_349 b_12 NI_12 NS_349 0 4.2235818713773959e-07
GC_12_350 b_12 NI_12 NS_350 0 1.8489189354920975e-06
GC_12_351 b_12 NI_12 NS_351 0 -2.9760479158494049e-08
GC_12_352 b_12 NI_12 NS_352 0 -1.3254972996615316e-06
GC_12_353 b_12 NI_12 NS_353 0 -6.4020217605116543e-07
GC_12_354 b_12 NI_12 NS_354 0 2.5950866871554369e-06
GC_12_355 b_12 NI_12 NS_355 0 4.5705238204427027e-07
GC_12_356 b_12 NI_12 NS_356 0 -2.2460566671006712e-06
GC_12_357 b_12 NI_12 NS_357 0 -8.0117684997280139e-07
GC_12_358 b_12 NI_12 NS_358 0 -9.3397538119556173e-07
GC_12_359 b_12 NI_12 NS_359 0 3.5739863394843955e-07
GC_12_360 b_12 NI_12 NS_360 0 9.1444699792138973e-07
GC_12_361 b_12 NI_12 NS_361 0 -5.5834208382291643e-07
GC_12_362 b_12 NI_12 NS_362 0 -7.2678592329864353e-07
GC_12_363 b_12 NI_12 NS_363 0 4.7648091226368444e-07
GC_12_364 b_12 NI_12 NS_364 0 7.4219337946451920e-07
GC_12_365 b_12 NI_12 NS_365 0 -1.7459565717520203e-07
GC_12_366 b_12 NI_12 NS_366 0 -8.7943210721328237e-07
GC_12_367 b_12 NI_12 NS_367 0 -3.4060706452077393e-07
GC_12_368 b_12 NI_12 NS_368 0 1.1609614368744585e-06
GC_12_369 b_12 NI_12 NS_369 0 2.5385915620619078e-07
GC_12_370 b_12 NI_12 NS_370 0 -8.4525457181816145e-07
GC_12_371 b_12 NI_12 NS_371 0 -6.5148053859937880e-08
GC_12_372 b_12 NI_12 NS_372 0 6.7372805652634027e-08
GC_12_373 b_12 NI_12 NS_373 0 -2.6093306733187101e-07
GC_12_374 b_12 NI_12 NS_374 0 -5.5061992718676064e-07
GC_12_375 b_12 NI_12 NS_375 0 1.8491359713220755e-07
GC_12_376 b_12 NI_12 NS_376 0 7.1949273911403835e-07
GC_12_377 b_12 NI_12 NS_377 0 -8.1165268854704649e-08
GC_12_378 b_12 NI_12 NS_378 0 -6.3616032831507521e-07
GC_12_379 b_12 NI_12 NS_379 0 1.0184239130584530e-07
GC_12_380 b_12 NI_12 NS_380 0 1.0497368746474568e-07
GC_12_381 b_12 NI_12 NS_381 0 -2.9217440263116187e-07
GC_12_382 b_12 NI_12 NS_382 0 -5.9433384797639111e-07
GC_12_383 b_12 NI_12 NS_383 0 1.6155156801861038e-07
GC_12_384 b_12 NI_12 NS_384 0 2.3346974633449267e-07
GC_12_385 b_12 NI_12 NS_385 0 -2.5774762587776436e-07
GC_12_386 b_12 NI_12 NS_386 0 -5.0844991012139482e-07
GC_12_387 b_12 NI_12 NS_387 0 4.9021996127565696e-08
GC_12_388 b_12 NI_12 NS_388 0 -4.9060950542413988e-08
GC_12_389 b_12 NI_12 NS_389 0 -3.6949400855706608e-07
GC_12_390 b_12 NI_12 NS_390 0 -5.5863817663682682e-07
GC_12_391 b_12 NI_12 NS_391 0 -2.3397526105808560e-07
GC_12_392 b_12 NI_12 NS_392 0 2.3114055522975372e-08
GC_12_393 b_12 NI_12 NS_393 0 -4.3492513332298083e-07
GC_12_394 b_12 NI_12 NS_394 0 -3.4101519234941691e-07
GC_12_395 b_12 NI_12 NS_395 0 -1.2370426229401057e-07
GC_12_396 b_12 NI_12 NS_396 0 1.7271131002047439e-08
GC_12_397 b_12 NI_12 NS_397 0 -5.6511190379415298e-07
GC_12_398 b_12 NI_12 NS_398 0 -4.3986477588015885e-07
GC_12_399 b_12 NI_12 NS_399 0 -3.1751829224933108e-07
GC_12_400 b_12 NI_12 NS_400 0 3.1817923197715301e-07
GC_12_401 b_12 NI_12 NS_401 0 -5.0074802986886245e-07
GC_12_402 b_12 NI_12 NS_402 0 3.7787371863318468e-08
GC_12_403 b_12 NI_12 NS_403 0 -9.9072370912194928e-09
GC_12_404 b_12 NI_12 NS_404 0 6.2428898920120466e-08
GC_12_405 b_12 NI_12 NS_405 0 -3.2503488151675524e-12
GC_12_406 b_12 NI_12 NS_406 0 3.2070824632223794e-12
GC_12_407 b_12 NI_12 NS_407 0 -5.7741464201701068e-07
GC_12_408 b_12 NI_12 NS_408 0 4.6881161072996694e-08
GC_12_409 b_12 NI_12 NS_409 0 -2.9017228092928781e-07
GC_12_410 b_12 NI_12 NS_410 0 1.1797448037049634e-07
GC_12_411 b_12 NI_12 NS_411 0 -5.7762078696505456e-09
GC_12_412 b_12 NI_12 NS_412 0 -6.8374782387117170e-08
GC_12_413 b_12 NI_12 NS_413 0 -6.6136356052261592e-07
GC_12_414 b_12 NI_12 NS_414 0 1.4039126896998428e-07
GC_12_415 b_12 NI_12 NS_415 0 2.9868784636110631e-08
GC_12_416 b_12 NI_12 NS_416 0 1.2538987198281494e-07
GC_12_417 b_12 NI_12 NS_417 0 -6.1347644169955822e-11
GC_12_418 b_12 NI_12 NS_418 0 1.2844592333419801e-10
GC_12_419 b_12 NI_12 NS_419 0 -3.4935746369590638e-08
GC_12_420 b_12 NI_12 NS_420 0 1.9709076046944075e-07
GC_12_421 b_12 NI_12 NS_421 0 -3.6685712436377348e-07
GC_12_422 b_12 NI_12 NS_422 0 -4.4445782515451381e-08
GC_12_423 b_12 NI_12 NS_423 0 -1.8614735962247023e-07
GC_12_424 b_12 NI_12 NS_424 0 -2.6651664039882905e-09
GC_12_425 b_12 NI_12 NS_425 0 1.9333591073637031e-07
GC_12_426 b_12 NI_12 NS_426 0 8.2524904397473680e-08
GC_12_427 b_12 NI_12 NS_427 0 -2.6572623231658500e-07
GC_12_428 b_12 NI_12 NS_428 0 3.1365984580018560e-07
GC_12_429 b_12 NI_12 NS_429 0 1.2571476804200631e-07
GC_12_430 b_12 NI_12 NS_430 0 -1.4398645116040895e-07
GC_12_431 b_12 NI_12 NS_431 0 -5.8257050425407554e-08
GC_12_432 b_12 NI_12 NS_432 0 2.3778824649861537e-07
GC_12_433 b_12 NI_12 NS_433 0 -9.0136355736544841e-05
GC_12_434 b_12 NI_12 NS_434 0 7.1502356229895023e-12
GC_12_435 b_12 NI_12 NS_435 0 -5.7297234131266524e-11
GC_12_436 b_12 NI_12 NS_436 0 3.3361240928755744e-10
GC_12_437 b_12 NI_12 NS_437 0 -1.5721768807573338e-06
GC_12_438 b_12 NI_12 NS_438 0 -1.5573916940731968e-06
GC_12_439 b_12 NI_12 NS_439 0 9.4297710286862335e-07
GC_12_440 b_12 NI_12 NS_440 0 7.2566155248078868e-07
GC_12_441 b_12 NI_12 NS_441 0 -2.7196321494779178e-06
GC_12_442 b_12 NI_12 NS_442 0 3.0307843604530503e-06
GC_12_443 b_12 NI_12 NS_443 0 -3.0496665386476411e-06
GC_12_444 b_12 NI_12 NS_444 0 -2.5769719569007695e-06
GC_12_445 b_12 NI_12 NS_445 0 1.5158942076104749e-06
GC_12_446 b_12 NI_12 NS_446 0 9.0896937247030561e-08
GC_12_447 b_12 NI_12 NS_447 0 -1.6657839818611221e-06
GC_12_448 b_12 NI_12 NS_448 0 1.7972661752921842e-06
GC_12_449 b_12 NI_12 NS_449 0 8.9123614654584304e-07
GC_12_450 b_12 NI_12 NS_450 0 4.1366233377629410e-06
GC_12_451 b_12 NI_12 NS_451 0 -4.2927705697191073e-06
GC_12_452 b_12 NI_12 NS_452 0 -2.0599950432792330e-06
GC_12_453 b_12 NI_12 NS_453 0 2.3787740707544206e-06
GC_12_454 b_12 NI_12 NS_454 0 -1.9358813155316805e-06
GC_12_455 b_12 NI_12 NS_455 0 -1.1788211007968489e-06
GC_12_456 b_12 NI_12 NS_456 0 3.2601449243831429e-06
GC_12_457 b_12 NI_12 NS_457 0 -8.4124028917054680e-06
GC_12_458 b_12 NI_12 NS_458 0 1.1213011411878179e-05
GC_12_459 b_12 NI_12 NS_459 0 1.2598105071922948e-06
GC_12_460 b_12 NI_12 NS_460 0 -1.6518676612093318e-06
GC_12_461 b_12 NI_12 NS_461 0 9.9604762727274718e-06
GC_12_462 b_12 NI_12 NS_462 0 1.7407376235673863e-05
GC_12_463 b_12 NI_12 NS_463 0 -6.6234990267550164e-07
GC_12_464 b_12 NI_12 NS_464 0 -5.4667126649048920e-07
GC_12_465 b_12 NI_12 NS_465 0 4.5572841082293303e-07
GC_12_466 b_12 NI_12 NS_466 0 -1.3700987618163008e-06
GC_12_467 b_12 NI_12 NS_467 0 7.0273663136345741e-06
GC_12_468 b_12 NI_12 NS_468 0 -2.3133444758448395e-07
GC_12_469 b_12 NI_12 NS_469 0 6.9999840924485819e-07
GC_12_470 b_12 NI_12 NS_470 0 2.9955124650599887e-06
GC_12_471 b_12 NI_12 NS_471 0 4.4109065986837420e-07
GC_12_472 b_12 NI_12 NS_472 0 2.9100582164222086e-06
GC_12_473 b_12 NI_12 NS_473 0 1.1671208981156471e-06
GC_12_474 b_12 NI_12 NS_474 0 -1.4115779126603250e-06
GC_12_475 b_12 NI_12 NS_475 0 9.4124698195029775e-06
GC_12_476 b_12 NI_12 NS_476 0 5.2153685051463780e-06
GC_12_477 b_12 NI_12 NS_477 0 5.7060036045163863e-07
GC_12_478 b_12 NI_12 NS_478 0 1.1337167597986733e-06
GC_12_479 b_12 NI_12 NS_479 0 5.6635909818430067e-08
GC_12_480 b_12 NI_12 NS_480 0 4.4780037014037347e-07
GC_12_481 b_12 NI_12 NS_481 0 1.2930178632400987e-06
GC_12_482 b_12 NI_12 NS_482 0 -8.5758347142630048e-07
GC_12_483 b_12 NI_12 NS_483 0 9.1863120105597734e-06
GC_12_484 b_12 NI_12 NS_484 0 6.5374887604811183e-07
GC_12_485 b_12 NI_12 NS_485 0 8.3835043995654953e-07
GC_12_486 b_12 NI_12 NS_486 0 1.4354656355013374e-06
GC_12_487 b_12 NI_12 NS_487 0 1.0193423026438046e-06
GC_12_488 b_12 NI_12 NS_488 0 5.8697996261425739e-07
GC_12_489 b_12 NI_12 NS_489 0 1.3710364091969658e-06
GC_12_490 b_12 NI_12 NS_490 0 -9.5622626157697716e-07
GC_12_491 b_12 NI_12 NS_491 0 8.0098216601307482e-06
GC_12_492 b_12 NI_12 NS_492 0 -2.1610559649359395e-06
GC_12_493 b_12 NI_12 NS_493 0 1.1721229921319296e-06
GC_12_494 b_12 NI_12 NS_494 0 1.5263091429408419e-06
GC_12_495 b_12 NI_12 NS_495 0 1.5749286378675025e-06
GC_12_496 b_12 NI_12 NS_496 0 -2.5368031413550410e-07
GC_12_497 b_12 NI_12 NS_497 0 1.3308034396931568e-06
GC_12_498 b_12 NI_12 NS_498 0 -1.0066192668787482e-06
GC_12_499 b_12 NI_12 NS_499 0 5.7892069274128987e-06
GC_12_500 b_12 NI_12 NS_500 0 -3.9086674630805704e-06
GC_12_501 b_12 NI_12 NS_501 0 1.8024564314863506e-06
GC_12_502 b_12 NI_12 NS_502 0 1.4095148117162175e-06
GC_12_503 b_12 NI_12 NS_503 0 1.0763945661744112e-06
GC_12_504 b_12 NI_12 NS_504 0 -1.4081499302208657e-06
GC_12_505 b_12 NI_12 NS_505 0 1.4146229366586583e-06
GC_12_506 b_12 NI_12 NS_506 0 -1.1369737720992846e-06
GC_12_507 b_12 NI_12 NS_507 0 2.9379405739425147e-06
GC_12_508 b_12 NI_12 NS_508 0 -4.1714562574521824e-06
GC_12_509 b_12 NI_12 NS_509 0 2.2085104875887723e-06
GC_12_510 b_12 NI_12 NS_510 0 2.9634361932213872e-07
GC_12_511 b_12 NI_12 NS_511 0 -3.3704327250260787e-07
GC_12_512 b_12 NI_12 NS_512 0 -1.1837413087423987e-06
GC_12_513 b_12 NI_12 NS_513 0 2.4875092887568648e-11
GC_12_514 b_12 NI_12 NS_514 0 -4.0913075593266720e-11
GC_12_515 b_12 NI_12 NS_515 0 7.8539226718749777e-07
GC_12_516 b_12 NI_12 NS_516 0 -1.5911469245474544e-06
GC_12_517 b_12 NI_12 NS_517 0 1.2557733139300301e-06
GC_12_518 b_12 NI_12 NS_518 0 2.2315349882104549e-07
GC_12_519 b_12 NI_12 NS_519 0 1.5659284056346824e-07
GC_12_520 b_12 NI_12 NS_520 0 -5.4948919021587329e-07
GC_12_521 b_12 NI_12 NS_521 0 5.4537294377017032e-07
GC_12_522 b_12 NI_12 NS_522 0 -8.9276766083096860e-07
GC_12_523 b_12 NI_12 NS_523 0 1.2830290295692675e-06
GC_12_524 b_12 NI_12 NS_524 0 -2.0549390827785975e-06
GC_12_525 b_12 NI_12 NS_525 0 4.7366014943532799e-10
GC_12_526 b_12 NI_12 NS_526 0 -1.2085632637236165e-09
GC_12_527 b_12 NI_12 NS_527 0 5.4539101365352945e-07
GC_12_528 b_12 NI_12 NS_528 0 -8.5655978748325295e-07
GC_12_529 b_12 NI_12 NS_529 0 7.1232724332121764e-07
GC_12_530 b_12 NI_12 NS_530 0 -9.5180860556408743e-07
GC_12_531 b_12 NI_12 NS_531 0 8.8751885403641791e-08
GC_12_532 b_12 NI_12 NS_532 0 5.0689002009894402e-08
GC_12_533 b_12 NI_12 NS_533 0 1.3271494380879537e-06
GC_12_534 b_12 NI_12 NS_534 0 -1.2248162895034914e-06
GC_12_535 b_12 NI_12 NS_535 0 1.6449393067482318e-06
GC_12_536 b_12 NI_12 NS_536 0 -2.9372198244700481e-07
GC_12_537 b_12 NI_12 NS_537 0 -2.3013047891115490e-07
GC_12_538 b_12 NI_12 NS_538 0 -7.3458698602084330e-07
GC_12_539 b_12 NI_12 NS_539 0 7.3260761873245616e-07
GC_12_540 b_12 NI_12 NS_540 0 2.8937259074941047e-07
GC_12_541 b_12 NI_12 NS_541 0 4.9610772991190690e-05
GC_12_542 b_12 NI_12 NS_542 0 3.6353664830597115e-12
GC_12_543 b_12 NI_12 NS_543 0 -4.1276395009054999e-12
GC_12_544 b_12 NI_12 NS_544 0 9.4606349821306945e-10
GC_12_545 b_12 NI_12 NS_545 0 -4.5694251452268520e-08
GC_12_546 b_12 NI_12 NS_546 0 2.5276731831868542e-07
GC_12_547 b_12 NI_12 NS_547 0 2.5906303270812556e-07
GC_12_548 b_12 NI_12 NS_548 0 4.0752877862473567e-07
GC_12_549 b_12 NI_12 NS_549 0 -1.3716172225583666e-07
GC_12_550 b_12 NI_12 NS_550 0 2.4384822143209491e-07
GC_12_551 b_12 NI_12 NS_551 0 7.8139033215938081e-07
GC_12_552 b_12 NI_12 NS_552 0 1.4415703339304654e-06
GC_12_553 b_12 NI_12 NS_553 0 1.0388734873020947e-06
GC_12_554 b_12 NI_12 NS_554 0 -5.2228256109397197e-07
GC_12_555 b_12 NI_12 NS_555 0 3.3588438046498606e-07
GC_12_556 b_12 NI_12 NS_556 0 8.8677771362843330e-07
GC_12_557 b_12 NI_12 NS_557 0 7.3258462884309236e-07
GC_12_558 b_12 NI_12 NS_558 0 -3.6895409723072375e-07
GC_12_559 b_12 NI_12 NS_559 0 4.3580342250138926e-06
GC_12_560 b_12 NI_12 NS_560 0 1.3814609905658436e-06
GC_12_561 b_12 NI_12 NS_561 0 -1.6431405652083291e-06
GC_12_562 b_12 NI_12 NS_562 0 -3.5781604831255004e-06
GC_12_563 b_12 NI_12 NS_563 0 2.3983175392115220e-07
GC_12_564 b_12 NI_12 NS_564 0 1.5513164709137411e-06
GC_12_565 b_12 NI_12 NS_565 0 2.9719512366106013e-06
GC_12_566 b_12 NI_12 NS_566 0 -4.7485561650445741e-06
GC_12_567 b_12 NI_12 NS_567 0 -7.7194418944309052e-07
GC_12_568 b_12 NI_12 NS_568 0 5.6548805772540601e-07
GC_12_569 b_12 NI_12 NS_569 0 5.5722032676964905e-06
GC_12_570 b_12 NI_12 NS_570 0 -5.8225121148156854e-06
GC_12_571 b_12 NI_12 NS_571 0 -3.3127674889955247e-06
GC_12_572 b_12 NI_12 NS_572 0 1.7944205544763977e-06
GC_12_573 b_12 NI_12 NS_573 0 8.6215747175261807e-07
GC_12_574 b_12 NI_12 NS_574 0 1.2284626993241903e-06
GC_12_575 b_12 NI_12 NS_575 0 1.5941355691815362e-06
GC_12_576 b_12 NI_12 NS_576 0 -4.1010708915559992e-06
GC_12_577 b_12 NI_12 NS_577 0 5.6926973522471065e-07
GC_12_578 b_12 NI_12 NS_578 0 1.9922709033500055e-07
GC_12_579 b_12 NI_12 NS_579 0 1.7434060426755545e-07
GC_12_580 b_12 NI_12 NS_580 0 -4.0363619344133091e-06
GC_12_581 b_12 NI_12 NS_581 0 -1.8756602397580504e-07
GC_12_582 b_12 NI_12 NS_582 0 1.6761042793530370e-07
GC_12_583 b_12 NI_12 NS_583 0 4.6377163291813014e-06
GC_12_584 b_12 NI_12 NS_584 0 -6.3334440459010014e-06
GC_12_585 b_12 NI_12 NS_585 0 -1.8278218709001165e-06
GC_12_586 b_12 NI_12 NS_586 0 -1.2890015002343846e-06
GC_12_587 b_12 NI_12 NS_587 0 1.3669191647901871e-06
GC_12_588 b_12 NI_12 NS_588 0 -1.1985547376084006e-06
GC_12_589 b_12 NI_12 NS_589 0 3.7643233251459044e-07
GC_12_590 b_12 NI_12 NS_590 0 -2.0976089175794464e-06
GC_12_591 b_12 NI_12 NS_591 0 -1.4875503157297784e-06
GC_12_592 b_12 NI_12 NS_592 0 -1.1765895605450919e-05
GC_12_593 b_12 NI_12 NS_593 0 -2.2683520541338000e-06
GC_12_594 b_12 NI_12 NS_594 0 -1.7024969218494275e-06
GC_12_595 b_12 NI_12 NS_595 0 -2.3842948597022922e-06
GC_12_596 b_12 NI_12 NS_596 0 -3.9896434485232935e-06
GC_12_597 b_12 NI_12 NS_597 0 -1.4876632363326576e-06
GC_12_598 b_12 NI_12 NS_598 0 -2.4187940708451609e-06
GC_12_599 b_12 NI_12 NS_599 0 -1.0716988022568635e-05
GC_12_600 b_12 NI_12 NS_600 0 -7.0850917053973754e-06
GC_12_601 b_12 NI_12 NS_601 0 -3.1909449457256600e-06
GC_12_602 b_12 NI_12 NS_602 0 -8.5674731283523207e-07
GC_12_603 b_12 NI_12 NS_603 0 -5.7476367963176025e-06
GC_12_604 b_12 NI_12 NS_604 0 -3.7004835247121932e-07
GC_12_605 b_12 NI_12 NS_605 0 -3.1243751808771300e-06
GC_12_606 b_12 NI_12 NS_606 0 -1.7461462864901344e-06
GC_12_607 b_12 NI_12 NS_607 0 -1.0618663952211215e-05
GC_12_608 b_12 NI_12 NS_608 0 3.3753559904398847e-06
GC_12_609 b_12 NI_12 NS_609 0 -3.6318005638369216e-06
GC_12_610 b_12 NI_12 NS_610 0 8.3009925602391878e-07
GC_12_611 b_12 NI_12 NS_611 0 -2.8719522352346491e-06
GC_12_612 b_12 NI_12 NS_612 0 3.9430648917234993e-06
GC_12_613 b_12 NI_12 NS_613 0 -4.3595837446973394e-06
GC_12_614 b_12 NI_12 NS_614 0 1.7264962895686570e-07
GC_12_615 b_12 NI_12 NS_615 0 -1.8585274569611680e-06
GC_12_616 b_12 NI_12 NS_616 0 7.2740539079145399e-06
GC_12_617 b_12 NI_12 NS_617 0 -1.5748465151681733e-06
GC_12_618 b_12 NI_12 NS_618 0 2.8115308990780342e-06
GC_12_619 b_12 NI_12 NS_619 0 9.3643768766641827e-07
GC_12_620 b_12 NI_12 NS_620 0 1.8337165857135626e-06
GC_12_621 b_12 NI_12 NS_621 0 -3.0124129187351162e-11
GC_12_622 b_12 NI_12 NS_622 0 -3.3889598368874748e-12
GC_12_623 b_12 NI_12 NS_623 0 -1.7319008600092636e-06
GC_12_624 b_12 NI_12 NS_624 0 2.1529089109536021e-06
GC_12_625 b_12 NI_12 NS_625 0 -3.2428003584426824e-07
GC_12_626 b_12 NI_12 NS_626 0 1.0583764812552100e-06
GC_12_627 b_12 NI_12 NS_627 0 1.4379982905042633e-07
GC_12_628 b_12 NI_12 NS_628 0 6.3880027744164973e-07
GC_12_629 b_12 NI_12 NS_629 0 -1.0428224717786430e-06
GC_12_630 b_12 NI_12 NS_630 0 1.2847613934193417e-06
GC_12_631 b_12 NI_12 NS_631 0 9.8816648844366813e-07
GC_12_632 b_12 NI_12 NS_632 0 1.8536024043615666e-06
GC_12_633 b_12 NI_12 NS_633 0 -1.5199212713091218e-09
GC_12_634 b_12 NI_12 NS_634 0 -7.6810695259631191e-10
GC_12_635 b_12 NI_12 NS_635 0 -4.6943524165553923e-07
GC_12_636 b_12 NI_12 NS_636 0 -2.3372168020445082e-08
GC_12_637 b_12 NI_12 NS_637 0 -3.1181052616124605e-07
GC_12_638 b_12 NI_12 NS_638 0 1.9126098523680625e-07
GC_12_639 b_12 NI_12 NS_639 0 -5.4910122087894835e-07
GC_12_640 b_12 NI_12 NS_640 0 1.5141087371644341e-07
GC_12_641 b_12 NI_12 NS_641 0 6.6188086543755849e-07
GC_12_642 b_12 NI_12 NS_642 0 8.2996781794545916e-07
GC_12_643 b_12 NI_12 NS_643 0 2.3288642134845893e-07
GC_12_644 b_12 NI_12 NS_644 0 7.0026481698283684e-07
GC_12_645 b_12 NI_12 NS_645 0 3.0418971802923238e-09
GC_12_646 b_12 NI_12 NS_646 0 -1.3243557842626220e-07
GC_12_647 b_12 NI_12 NS_647 0 -3.4705017391428955e-07
GC_12_648 b_12 NI_12 NS_648 0 2.9428872054585491e-07
GC_12_649 b_12 NI_12 NS_649 0 -1.5116580189751674e-04
GC_12_650 b_12 NI_12 NS_650 0 3.7546735532282108e-11
GC_12_651 b_12 NI_12 NS_651 0 1.7613934449061165e-11
GC_12_652 b_12 NI_12 NS_652 0 8.7391218009241016e-10
GC_12_653 b_12 NI_12 NS_653 0 -2.3302369757350062e-06
GC_12_654 b_12 NI_12 NS_654 0 -1.6501405067283550e-06
GC_12_655 b_12 NI_12 NS_655 0 1.4541335546261231e-06
GC_12_656 b_12 NI_12 NS_656 0 3.8965289544652495e-06
GC_12_657 b_12 NI_12 NS_657 0 2.9654767094117939e-06
GC_12_658 b_12 NI_12 NS_658 0 5.4214075951436729e-06
GC_12_659 b_12 NI_12 NS_659 0 5.3772560460992394e-06
GC_12_660 b_12 NI_12 NS_660 0 -8.4804540337924662e-06
GC_12_661 b_12 NI_12 NS_661 0 -2.2507456438285752e-06
GC_12_662 b_12 NI_12 NS_662 0 -1.2662236877763191e-05
GC_12_663 b_12 NI_12 NS_663 0 -3.7273752380533760e-06
GC_12_664 b_12 NI_12 NS_664 0 2.7450749092966887e-06
GC_12_665 b_12 NI_12 NS_665 0 4.4941459511111598e-06
GC_12_666 b_12 NI_12 NS_666 0 1.5803582194084578e-06
GC_12_667 b_12 NI_12 NS_667 0 8.5385434173206756e-06
GC_12_668 b_12 NI_12 NS_668 0 -3.8252066903542072e-05
GC_12_669 b_12 NI_12 NS_669 0 -4.2843508656223671e-05
GC_12_670 b_12 NI_12 NS_670 0 -1.4539742558933962e-06
GC_12_671 b_12 NI_12 NS_671 0 -1.4647321309074854e-05
GC_12_672 b_12 NI_12 NS_672 0 -8.2775498084624319e-06
GC_12_673 b_12 NI_12 NS_673 0 -7.0243420319279935e-05
GC_12_674 b_12 NI_12 NS_674 0 7.5185371357342547e-05
GC_12_675 b_12 NI_12 NS_675 0 4.8693902755918023e-06
GC_12_676 b_12 NI_12 NS_676 0 1.3024070501041624e-05
GC_12_677 b_12 NI_12 NS_677 0 6.5219383378212328e-05
GC_12_678 b_12 NI_12 NS_678 0 1.2202119243796634e-04
GC_12_679 b_12 NI_12 NS_679 0 -2.7583168732446691e-07
GC_12_680 b_12 NI_12 NS_680 0 -3.7368600931246176e-05
GC_12_681 b_12 NI_12 NS_681 0 1.6806379519788332e-05
GC_12_682 b_12 NI_12 NS_682 0 4.1838901649088106e-06
GC_12_683 b_12 NI_12 NS_683 0 2.5158697301376527e-05
GC_12_684 b_12 NI_12 NS_684 0 -3.0985672747469890e-05
GC_12_685 b_12 NI_12 NS_685 0 -8.5164695654003393e-06
GC_12_686 b_12 NI_12 NS_686 0 -2.5732801586015935e-06
GC_12_687 b_12 NI_12 NS_687 0 -8.0804278423976139e-06
GC_12_688 b_12 NI_12 NS_688 0 2.4256613197650361e-05
GC_12_689 b_12 NI_12 NS_689 0 6.0403100256736824e-06
GC_12_690 b_12 NI_12 NS_690 0 8.3878817749586490e-06
GC_12_691 b_12 NI_12 NS_691 0 5.7350643143454561e-05
GC_12_692 b_12 NI_12 NS_692 0 2.3736435898013009e-05
GC_12_693 b_12 NI_12 NS_693 0 3.5345631110172491e-06
GC_12_694 b_12 NI_12 NS_694 0 -1.2244041242765576e-05
GC_12_695 b_12 NI_12 NS_695 0 -7.4191807182478235e-08
GC_12_696 b_12 NI_12 NS_696 0 -1.3740256261155989e-06
GC_12_697 b_12 NI_12 NS_697 0 7.1802178399963440e-06
GC_12_698 b_12 NI_12 NS_698 0 2.7778757657677640e-06
GC_12_699 b_12 NI_12 NS_699 0 4.2416635209670570e-05
GC_12_700 b_12 NI_12 NS_700 0 -1.9012300122536442e-05
GC_12_701 b_12 NI_12 NS_701 0 -2.5057996356436424e-06
GC_12_702 b_12 NI_12 NS_702 0 -7.6312037372716200e-06
GC_12_703 b_12 NI_12 NS_703 0 -2.8031972039756903e-06
GC_12_704 b_12 NI_12 NS_704 0 1.0883876218637819e-06
GC_12_705 b_12 NI_12 NS_705 0 9.8313738412121503e-06
GC_12_706 b_12 NI_12 NS_706 0 2.5417304268863423e-06
GC_12_707 b_12 NI_12 NS_707 0 2.2415810106830317e-05
GC_12_708 b_12 NI_12 NS_708 0 -3.3139157740394737e-05
GC_12_709 b_12 NI_12 NS_709 0 -5.7255916214771250e-06
GC_12_710 b_12 NI_12 NS_710 0 -4.2015228867245712e-06
GC_12_711 b_12 NI_12 NS_711 0 -8.8987242265679047e-07
GC_12_712 b_12 NI_12 NS_712 0 4.2524741466772142e-06
GC_12_713 b_12 NI_12 NS_713 0 1.2480179638790574e-05
GC_12_714 b_12 NI_12 NS_714 0 -2.7949245562132882e-07
GC_12_715 b_12 NI_12 NS_715 0 4.7397689812219836e-07
GC_12_716 b_12 NI_12 NS_716 0 -3.2834666136422625e-05
GC_12_717 b_12 NI_12 NS_717 0 -6.9268143332932815e-06
GC_12_718 b_12 NI_12 NS_718 0 4.0684551534341532e-07
GC_12_719 b_12 NI_12 NS_719 0 3.8410641837752322e-06
GC_12_720 b_12 NI_12 NS_720 0 3.5676466391664066e-06
GC_12_721 b_12 NI_12 NS_721 0 1.4108458184621948e-05
GC_12_722 b_12 NI_12 NS_722 0 -6.6872354976167565e-06
GC_12_723 b_12 NI_12 NS_723 0 -1.5604808116486009e-05
GC_12_724 b_12 NI_12 NS_724 0 -1.9003616437865963e-05
GC_12_725 b_12 NI_12 NS_725 0 -2.9952205923727312e-06
GC_12_726 b_12 NI_12 NS_726 0 5.1042652612900051e-06
GC_12_727 b_12 NI_12 NS_727 0 4.2096732132719440e-06
GC_12_728 b_12 NI_12 NS_728 0 -1.8809864073347862e-06
GC_12_729 b_12 NI_12 NS_729 0 -2.7916018986279809e-11
GC_12_730 b_12 NI_12 NS_730 0 5.8155687346025427e-12
GC_12_731 b_12 NI_12 NS_731 0 4.8698610566326226e-06
GC_12_732 b_12 NI_12 NS_732 0 -1.1668132045165838e-05
GC_12_733 b_12 NI_12 NS_733 0 -5.0905717544445863e-07
GC_12_734 b_12 NI_12 NS_734 0 2.7992511672198080e-06
GC_12_735 b_12 NI_12 NS_735 0 2.3509245041519244e-06
GC_12_736 b_12 NI_12 NS_736 0 -1.5716519643993012e-06
GC_12_737 b_12 NI_12 NS_737 0 2.1314070655337414e-06
GC_12_738 b_12 NI_12 NS_738 0 -9.8974351507277158e-06
GC_12_739 b_12 NI_12 NS_739 0 -1.0613650039962233e-05
GC_12_740 b_12 NI_12 NS_740 0 -3.5263101205565950e-06
GC_12_741 b_12 NI_12 NS_741 0 -2.3906910207607486e-10
GC_12_742 b_12 NI_12 NS_742 0 4.4566872839277696e-10
GC_12_743 b_12 NI_12 NS_743 0 -9.1766900293513288e-06
GC_12_744 b_12 NI_12 NS_744 0 -5.6138367012930018e-06
GC_12_745 b_12 NI_12 NS_745 0 1.9952216093931757e-06
GC_12_746 b_12 NI_12 NS_746 0 -6.7132231771115170e-06
GC_12_747 b_12 NI_12 NS_747 0 -3.3605962762495165e-06
GC_12_748 b_12 NI_12 NS_748 0 -1.7941032037582419e-07
GC_12_749 b_12 NI_12 NS_749 0 -8.5928674021928665e-06
GC_12_750 b_12 NI_12 NS_750 0 5.9560157862968648e-07
GC_12_751 b_12 NI_12 NS_751 0 2.6078668501917944e-06
GC_12_752 b_12 NI_12 NS_752 0 2.8393330925832523e-06
GC_12_753 b_12 NI_12 NS_753 0 9.9244074338945146e-07
GC_12_754 b_12 NI_12 NS_754 0 -3.6889586077486844e-06
GC_12_755 b_12 NI_12 NS_755 0 -5.4153741128458496e-06
GC_12_756 b_12 NI_12 NS_756 0 -4.2328074415981151e-06
GC_12_757 b_12 NI_12 NS_757 0 -5.0477224990236760e-05
GC_12_758 b_12 NI_12 NS_758 0 -7.9794594858739323e-12
GC_12_759 b_12 NI_12 NS_759 0 -2.0628668851941627e-10
GC_12_760 b_12 NI_12 NS_760 0 9.8384587460819928e-09
GC_12_761 b_12 NI_12 NS_761 0 5.6375622735304104e-07
GC_12_762 b_12 NI_12 NS_762 0 4.4381100992507565e-08
GC_12_763 b_12 NI_12 NS_763 0 2.9366447764480328e-06
GC_12_764 b_12 NI_12 NS_764 0 -1.4886583502872263e-06
GC_12_765 b_12 NI_12 NS_765 0 -3.1321940489515177e-06
GC_12_766 b_12 NI_12 NS_766 0 -2.6552915101559059e-06
GC_12_767 b_12 NI_12 NS_767 0 4.5743595069604245e-06
GC_12_768 b_12 NI_12 NS_768 0 -4.2831837973759683e-07
GC_12_769 b_12 NI_12 NS_769 0 -7.3616118599736651e-06
GC_12_770 b_12 NI_12 NS_770 0 -7.5350579561300564e-06
GC_12_771 b_12 NI_12 NS_771 0 -2.4585698712454257e-07
GC_12_772 b_12 NI_12 NS_772 0 -1.3969578598961448e-06
GC_12_773 b_12 NI_12 NS_773 0 -5.8994749604602284e-06
GC_12_774 b_12 NI_12 NS_774 0 2.4069590451826504e-06
GC_12_775 b_12 NI_12 NS_775 0 5.0799360134779480e-06
GC_12_776 b_12 NI_12 NS_776 0 -5.0478328953330472e-06
GC_12_777 b_12 NI_12 NS_777 0 -1.6513908622818308e-05
GC_12_778 b_12 NI_12 NS_778 0 4.9731463204022417e-06
GC_12_779 b_12 NI_12 NS_779 0 -1.2104003762205426e-06
GC_12_780 b_12 NI_12 NS_780 0 7.3647400805812193e-06
GC_12_781 b_12 NI_12 NS_781 0 -6.6058685630754648e-06
GC_12_782 b_12 NI_12 NS_782 0 -3.9243502886197149e-06
GC_12_783 b_12 NI_12 NS_783 0 -3.2757672969867570e-06
GC_12_784 b_12 NI_12 NS_784 0 8.1805471743186158e-06
GC_12_785 b_12 NI_12 NS_785 0 -1.4123073047820192e-06
GC_12_786 b_12 NI_12 NS_786 0 -3.8938058832094629e-06
GC_12_787 b_12 NI_12 NS_787 0 -3.9336561887552849e-06
GC_12_788 b_12 NI_12 NS_788 0 1.1229367966197919e-05
GC_12_789 b_12 NI_12 NS_789 0 -1.1559733865314551e-07
GC_12_790 b_12 NI_12 NS_790 0 7.5148536127967341e-06
GC_12_791 b_12 NI_12 NS_791 0 -3.6231367195279675e-06
GC_12_792 b_12 NI_12 NS_792 0 1.5253183463075268e-06
GC_12_793 b_12 NI_12 NS_793 0 -4.3432151533410566e-07
GC_12_794 b_12 NI_12 NS_794 0 8.2698465669391085e-06
GC_12_795 b_12 NI_12 NS_795 0 -5.5569865868358855e-07
GC_12_796 b_12 NI_12 NS_796 0 2.2142468505688049e-06
GC_12_797 b_12 NI_12 NS_797 0 -2.3137636682240835e-06
GC_12_798 b_12 NI_12 NS_798 0 8.3308447631997505e-06
GC_12_799 b_12 NI_12 NS_799 0 6.0315811362608842e-07
GC_12_800 b_12 NI_12 NS_800 0 9.9619463653743308e-06
GC_12_801 b_12 NI_12 NS_801 0 -6.8797660924734196e-07
GC_12_802 b_12 NI_12 NS_802 0 8.8045969428012530e-06
GC_12_803 b_12 NI_12 NS_803 0 -1.2376792536153712e-06
GC_12_804 b_12 NI_12 NS_804 0 4.0443129405993464e-06
GC_12_805 b_12 NI_12 NS_805 0 1.2364273552953737e-06
GC_12_806 b_12 NI_12 NS_806 0 1.2169058281194751e-05
GC_12_807 b_12 NI_12 NS_807 0 1.8569136145298832e-05
GC_12_808 b_12 NI_12 NS_808 0 1.6970584950113438e-05
GC_12_809 b_12 NI_12 NS_809 0 4.9794872575574749e-06
GC_12_810 b_12 NI_12 NS_810 0 7.7555434494748196e-06
GC_12_811 b_12 NI_12 NS_811 0 1.0278855790236918e-05
GC_12_812 b_12 NI_12 NS_812 0 3.8769443413061608e-06
GC_12_813 b_12 NI_12 NS_813 0 6.7691299983564720e-06
GC_12_814 b_12 NI_12 NS_814 0 1.0908028789828267e-05
GC_12_815 b_12 NI_12 NS_815 0 3.3282822109837675e-05
GC_12_816 b_12 NI_12 NS_816 0 -6.0912175760129855e-06
GC_12_817 b_12 NI_12 NS_817 0 8.1276574980054853e-06
GC_12_818 b_12 NI_12 NS_818 0 3.4130676234755251e-06
GC_12_819 b_12 NI_12 NS_819 0 1.1915390257844165e-05
GC_12_820 b_12 NI_12 NS_820 0 -1.0252449413497727e-05
GC_12_821 b_12 NI_12 NS_821 0 1.0732664287981988e-05
GC_12_822 b_12 NI_12 NS_822 0 6.4703324989183926e-06
GC_12_823 b_12 NI_12 NS_823 0 1.6861235196635212e-05
GC_12_824 b_12 NI_12 NS_824 0 -3.0702835826055196e-05
GC_12_825 b_12 NI_12 NS_825 0 8.0800694418136213e-06
GC_12_826 b_12 NI_12 NS_826 0 -2.9184894814935855e-06
GC_12_827 b_12 NI_12 NS_827 0 -3.2230744049275240e-06
GC_12_828 b_12 NI_12 NS_828 0 -1.6215595292990598e-05
GC_12_829 b_12 NI_12 NS_829 0 1.1759403151291675e-05
GC_12_830 b_12 NI_12 NS_830 0 -1.5875023991893612e-06
GC_12_831 b_12 NI_12 NS_831 0 -1.2692758191451184e-05
GC_12_832 b_12 NI_12 NS_832 0 -2.5024419605443795e-05
GC_12_833 b_12 NI_12 NS_833 0 -1.5671333804302810e-07
GC_12_834 b_12 NI_12 NS_834 0 -6.5860905090269802e-06
GC_12_835 b_12 NI_12 NS_835 0 -9.5588616545545416e-06
GC_12_836 b_12 NI_12 NS_836 0 -2.6136597644367207e-06
GC_12_837 b_12 NI_12 NS_837 0 1.0214437706304764e-10
GC_12_838 b_12 NI_12 NS_838 0 4.7347227039197555e-11
GC_12_839 b_12 NI_12 NS_839 0 1.4916302373562935e-06
GC_12_840 b_12 NI_12 NS_840 0 -4.6685481192171217e-06
GC_12_841 b_12 NI_12 NS_841 0 -1.3624857815388159e-06
GC_12_842 b_12 NI_12 NS_842 0 -1.3366693981292788e-06
GC_12_843 b_12 NI_12 NS_843 0 -4.8492450391466567e-06
GC_12_844 b_12 NI_12 NS_844 0 -9.9200195884019749e-07
GC_12_845 b_12 NI_12 NS_845 0 -1.1407273786350301e-06
GC_12_846 b_12 NI_12 NS_846 0 -2.7064160119493670e-06
GC_12_847 b_12 NI_12 NS_847 0 -9.9964601616103598e-06
GC_12_848 b_12 NI_12 NS_848 0 -4.0330068116233057e-06
GC_12_849 b_12 NI_12 NS_849 0 6.6625987038664061e-09
GC_12_850 b_12 NI_12 NS_850 0 5.4065805906042634e-09
GC_12_851 b_12 NI_12 NS_851 0 1.7627792955653998e-06
GC_12_852 b_12 NI_12 NS_852 0 4.8652332682072880e-07
GC_12_853 b_12 NI_12 NS_853 0 -1.6104309631664033e-06
GC_12_854 b_12 NI_12 NS_854 0 3.2255923626683964e-06
GC_12_855 b_12 NI_12 NS_855 0 -8.2940683922477161e-07
GC_12_856 b_12 NI_12 NS_856 0 7.0026345154566696e-07
GC_12_857 b_12 NI_12 NS_857 0 -7.6527107937888097e-06
GC_12_858 b_12 NI_12 NS_858 0 5.4683765790791451e-07
GC_12_859 b_12 NI_12 NS_859 0 -2.2162359597433271e-06
GC_12_860 b_12 NI_12 NS_860 0 2.0035047733763996e-06
GC_12_861 b_12 NI_12 NS_861 0 -2.0640124554414139e-06
GC_12_862 b_12 NI_12 NS_862 0 1.9717473922586412e-06
GC_12_863 b_12 NI_12 NS_863 0 1.2832743856719176e-06
GC_12_864 b_12 NI_12 NS_864 0 2.8361930426589573e-06
GC_12_865 b_12 NI_12 NS_865 0 -3.3036468990326707e-03
GC_12_866 b_12 NI_12 NS_866 0 1.8493852318561979e-09
GC_12_867 b_12 NI_12 NS_867 0 5.6032182859234192e-08
GC_12_868 b_12 NI_12 NS_868 0 1.8929694299607495e-06
GC_12_869 b_12 NI_12 NS_869 0 -9.1167742619689853e-05
GC_12_870 b_12 NI_12 NS_870 0 -5.7737889504323747e-05
GC_12_871 b_12 NI_12 NS_871 0 -1.2657732945403817e-03
GC_12_872 b_12 NI_12 NS_872 0 -2.9559375648287089e-04
GC_12_873 b_12 NI_12 NS_873 0 -1.6792132369024414e-03
GC_12_874 b_12 NI_12 NS_874 0 2.6464978351653022e-03
GC_12_875 b_12 NI_12 NS_875 0 5.1121225987294080e-04
GC_12_876 b_12 NI_12 NS_876 0 5.4276091317546783e-03
GC_12_877 b_12 NI_12 NS_877 0 7.1034890038042938e-03
GC_12_878 b_12 NI_12 NS_878 0 6.3629119994814971e-04
GC_12_879 b_12 NI_12 NS_879 0 6.4433018680413502e-04
GC_12_880 b_12 NI_12 NS_880 0 -6.6092006917636511e-04
GC_12_881 b_12 NI_12 NS_881 0 1.0576972016031383e-03
GC_12_882 b_12 NI_12 NS_882 0 1.5711403184788966e-03
GC_12_883 b_12 NI_12 NS_883 0 1.2687514766286465e-02
GC_12_884 b_12 NI_12 NS_884 0 1.3123212030775322e-02
GC_12_885 b_12 NI_12 NS_885 0 8.7187958199708669e-03
GC_12_886 b_12 NI_12 NS_886 0 -2.0392081355487007e-02
GC_12_887 b_12 NI_12 NS_887 0 8.3891006226464206e-03
GC_12_888 b_12 NI_12 NS_888 0 -2.9045267711130173e-03
GC_12_889 b_12 NI_12 NS_889 0 -1.2701294089145948e-02
GC_12_890 b_12 NI_12 NS_890 0 -3.8806698439854195e-02
GC_12_891 b_12 NI_12 NS_891 0 -7.2523396002941148e-03
GC_12_892 b_12 NI_12 NS_892 0 -2.1332744475554112e-03
GC_12_893 b_12 NI_12 NS_893 0 -5.2307204259538852e-02
GC_12_894 b_12 NI_12 NS_894 0 -1.7936127206527892e-03
GC_12_895 b_12 NI_12 NS_895 0 1.4914417223305046e-02
GC_12_896 b_12 NI_12 NS_896 0 8.6735768624812831e-03
GC_12_897 b_12 NI_12 NS_897 0 -5.9233541172649647e-03
GC_12_898 b_12 NI_12 NS_898 0 5.0044976579553665e-03
GC_12_899 b_12 NI_12 NS_899 0 8.3724192690853710e-03
GC_12_900 b_12 NI_12 NS_900 0 1.1688366950464338e-02
GC_12_901 b_12 NI_12 NS_901 0 4.5592638711198889e-03
GC_12_902 b_12 NI_12 NS_902 0 -2.9327397603978885e-03
GC_12_903 b_12 NI_12 NS_903 0 -7.8986718195548436e-03
GC_12_904 b_12 NI_12 NS_904 0 -8.1490630826487106e-03
GC_12_905 b_12 NI_12 NS_905 0 -5.6808135805708846e-03
GC_12_906 b_12 NI_12 NS_906 0 -6.1280929445905812e-04
GC_12_907 b_12 NI_12 NS_907 0 -1.8070847598322795e-02
GC_12_908 b_12 NI_12 NS_908 0 1.3578968420272484e-02
GC_12_909 b_12 NI_12 NS_909 0 4.7069876755458503e-03
GC_12_910 b_12 NI_12 NS_910 0 4.3794382397135019e-03
GC_12_911 b_12 NI_12 NS_911 0 6.5015896044742533e-04
GC_12_912 b_12 NI_12 NS_912 0 -1.0995413337265865e-04
GC_12_913 b_12 NI_12 NS_913 0 -3.7963992716311219e-03
GC_12_914 b_12 NI_12 NS_914 0 8.8498855781905990e-04
GC_12_915 b_12 NI_12 NS_915 0 -1.1178265682942274e-03
GC_12_916 b_12 NI_12 NS_916 0 1.6699689301459816e-02
GC_12_917 b_12 NI_12 NS_917 0 4.4472810509516214e-03
GC_12_918 b_12 NI_12 NS_918 0 7.0796490958417106e-04
GC_12_919 b_12 NI_12 NS_919 0 -5.1995707412455983e-04
GC_12_920 b_12 NI_12 NS_920 0 -2.2477503351890533e-03
GC_12_921 b_12 NI_12 NS_921 0 -4.9864550089647689e-03
GC_12_922 b_12 NI_12 NS_922 0 2.1108885097515504e-03
GC_12_923 b_12 NI_12 NS_923 0 7.3425321006322479e-03
GC_12_924 b_12 NI_12 NS_924 0 1.4345855443076415e-02
GC_12_925 b_12 NI_12 NS_925 0 4.1872288107967209e-03
GC_12_926 b_12 NI_12 NS_926 0 -1.6838584160417899e-03
GC_12_927 b_12 NI_12 NS_927 0 -3.3981227897296822e-03
GC_12_928 b_12 NI_12 NS_928 0 -2.1006244636292029e-03
GC_12_929 b_12 NI_12 NS_929 0 -5.4204239089510747e-03
GC_12_930 b_12 NI_12 NS_930 0 4.3817247906773760e-03
GC_12_931 b_12 NI_12 NS_931 0 1.3196875147406119e-02
GC_12_932 b_12 NI_12 NS_932 0 8.4333026005832326e-03
GC_12_933 b_12 NI_12 NS_933 0 2.8324347532634299e-03
GC_12_934 b_12 NI_12 NS_934 0 -4.1306074030110912e-03
GC_12_935 b_12 NI_12 NS_935 0 -5.3207869913107549e-03
GC_12_936 b_12 NI_12 NS_936 0 1.1381564703151451e-03
GC_12_937 b_12 NI_12 NS_937 0 -4.4310195680555232e-03
GC_12_938 b_12 NI_12 NS_938 0 8.3104298943740846e-03
GC_12_939 b_12 NI_12 NS_939 0 1.4612784024007959e-02
GC_12_940 b_12 NI_12 NS_940 0 -4.6824940608539638e-04
GC_12_941 b_12 NI_12 NS_941 0 -1.1845324052724595e-03
GC_12_942 b_12 NI_12 NS_942 0 -4.5473906493801149e-03
GC_12_943 b_12 NI_12 NS_943 0 -2.2825683634537870e-03
GC_12_944 b_12 NI_12 NS_944 0 4.3832546954991865e-03
GC_12_945 b_12 NI_12 NS_945 0 1.3572124102703460e-10
GC_12_946 b_12 NI_12 NS_946 0 -1.5466290572752125e-09
GC_12_947 b_12 NI_12 NS_947 0 1.4460258736973335e-03
GC_12_948 b_12 NI_12 NS_948 0 8.2165464986437287e-03
GC_12_949 b_12 NI_12 NS_949 0 -8.7895028726767686e-04
GC_12_950 b_12 NI_12 NS_950 0 -2.2072127790473605e-03
GC_12_951 b_12 NI_12 NS_951 0 -1.4679137060319611e-03
GC_12_952 b_12 NI_12 NS_952 0 2.7519857599257336e-03
GC_12_953 b_12 NI_12 NS_953 0 1.7320144499257471e-03
GC_12_954 b_12 NI_12 NS_954 0 7.6059319536920245e-03
GC_12_955 b_12 NI_12 NS_955 0 7.5874083949251389e-03
GC_12_956 b_12 NI_12 NS_956 0 -3.8276827678557735e-03
GC_12_957 b_12 NI_12 NS_957 0 -5.2101119164686736e-08
GC_12_958 b_12 NI_12 NS_958 0 -2.0817340503786414e-08
GC_12_959 b_12 NI_12 NS_959 0 1.1391243302509154e-02
GC_12_960 b_12 NI_12 NS_960 0 4.4700329663060479e-03
GC_12_961 b_12 NI_12 NS_961 0 -8.6185047910623510e-04
GC_12_962 b_12 NI_12 NS_962 0 6.4916224701406103e-03
GC_12_963 b_12 NI_12 NS_963 0 3.6263738520309163e-03
GC_12_964 b_12 NI_12 NS_964 0 4.0710467498280965e-04
GC_12_965 b_12 NI_12 NS_965 0 6.0525103063653893e-03
GC_12_966 b_12 NI_12 NS_966 0 -4.6635403202262343e-03
GC_12_967 b_12 NI_12 NS_967 0 -3.3929753841016306e-03
GC_12_968 b_12 NI_12 NS_968 0 -1.3533959425933650e-03
GC_12_969 b_12 NI_12 NS_969 0 1.1237967062708607e-04
GC_12_970 b_12 NI_12 NS_970 0 4.4958003009575656e-03
GC_12_971 b_12 NI_12 NS_971 0 7.2795569197375903e-03
GC_12_972 b_12 NI_12 NS_972 0 5.5305048218879807e-03
GC_12_973 b_12 NI_12 NS_973 0 1.1808601739319220e-03
GC_12_974 b_12 NI_12 NS_974 0 -3.5561504517945821e-09
GC_12_975 b_12 NI_12 NS_975 0 -4.8002201619163657e-08
GC_12_976 b_12 NI_12 NS_976 0 -3.4752337930990040e-06
GC_12_977 b_12 NI_12 NS_977 0 -3.6811894665243013e-04
GC_12_978 b_12 NI_12 NS_978 0 1.3598159843515961e-04
GC_12_979 b_12 NI_12 NS_979 0 1.1297148004086840e-03
GC_12_980 b_12 NI_12 NS_980 0 1.9432455940075590e-03
GC_12_981 b_12 NI_12 NS_981 0 -6.5025362219072046e-05
GC_12_982 b_12 NI_12 NS_982 0 -3.4937339203137611e-03
GC_12_983 b_12 NI_12 NS_983 0 -1.5644030835217774e-03
GC_12_984 b_12 NI_12 NS_984 0 5.0905614508096010e-03
GC_12_985 b_12 NI_12 NS_985 0 4.2534104358232464e-03
GC_12_986 b_12 NI_12 NS_986 0 -4.9937797865621447e-03
GC_12_987 b_12 NI_12 NS_987 0 -1.0085420667726996e-03
GC_12_988 b_12 NI_12 NS_988 0 5.6396308343244705e-04
GC_12_989 b_12 NI_12 NS_989 0 -2.0807418986297311e-03
GC_12_990 b_12 NI_12 NS_990 0 -1.8633296175921356e-03
GC_12_991 b_12 NI_12 NS_991 0 3.6453743243146774e-03
GC_12_992 b_12 NI_12 NS_992 0 1.1647299721461085e-02
GC_12_993 b_12 NI_12 NS_993 0 -8.9809376412843488e-04
GC_12_994 b_12 NI_12 NS_994 0 -1.4854264015549646e-02
GC_12_995 b_12 NI_12 NS_995 0 -8.1235082744216432e-03
GC_12_996 b_12 NI_12 NS_996 0 1.9195541370244569e-03
GC_12_997 b_12 NI_12 NS_997 0 1.1262993899966090e-02
GC_12_998 b_12 NI_12 NS_998 0 -1.8122030646772218e-03
GC_12_999 b_12 NI_12 NS_999 0 -7.5672396693017606e-03
GC_12_1000 b_12 NI_12 NS_1000 0 -1.6812110656907549e-03
GC_12_1001 b_12 NI_12 NS_1001 0 1.5281607338987278e-02
GC_12_1002 b_12 NI_12 NS_1002 0 5.3008467150273903e-03
GC_12_1003 b_12 NI_12 NS_1003 0 -1.3082790601246154e-02
GC_12_1004 b_12 NI_12 NS_1004 0 -5.4613195741109637e-03
GC_12_1005 b_12 NI_12 NS_1005 0 -6.6370644341744271e-03
GC_12_1006 b_12 NI_12 NS_1006 0 3.4566491501496514e-03
GC_12_1007 b_12 NI_12 NS_1007 0 6.3615686418213172e-03
GC_12_1008 b_12 NI_12 NS_1008 0 -1.8793111909254903e-03
GC_12_1009 b_12 NI_12 NS_1009 0 -5.4737174823898177e-03
GC_12_1010 b_12 NI_12 NS_1010 0 2.1829945210678388e-03
GC_12_1011 b_12 NI_12 NS_1011 0 5.3937402484608467e-03
GC_12_1012 b_12 NI_12 NS_1012 0 -2.6324139397165690e-03
GC_12_1013 b_12 NI_12 NS_1013 0 -6.3064434681043878e-03
GC_12_1014 b_12 NI_12 NS_1014 0 -4.8383766170777655e-04
GC_12_1015 b_12 NI_12 NS_1015 0 7.6452212090595811e-03
GC_12_1016 b_12 NI_12 NS_1016 0 3.6298699377665497e-03
GC_12_1017 b_12 NI_12 NS_1017 0 -5.8336100716466169e-03
GC_12_1018 b_12 NI_12 NS_1018 0 -3.4646020589867298e-03
GC_12_1019 b_12 NI_12 NS_1019 0 2.9619270154025620e-04
GC_12_1020 b_12 NI_12 NS_1020 0 5.5809921323429345e-04
GC_12_1021 b_12 NI_12 NS_1021 0 -4.9270674088370799e-03
GC_12_1022 b_12 NI_12 NS_1022 0 8.9217933472842174e-04
GC_12_1023 b_12 NI_12 NS_1023 0 6.2062906001030139e-03
GC_12_1024 b_12 NI_12 NS_1024 0 6.8829116828050992e-04
GC_12_1025 b_12 NI_12 NS_1025 0 -5.3209606423649377e-03
GC_12_1026 b_12 NI_12 NS_1026 0 -4.8420041089505106e-04
GC_12_1027 b_12 NI_12 NS_1027 0 1.5503170145524344e-03
GC_12_1028 b_12 NI_12 NS_1028 0 -4.3200389211267897e-05
GC_12_1029 b_12 NI_12 NS_1029 0 -6.0223399978072524e-03
GC_12_1030 b_12 NI_12 NS_1030 0 1.9232230871373194e-03
GC_12_1031 b_12 NI_12 NS_1031 0 6.2616320411049732e-03
GC_12_1032 b_12 NI_12 NS_1032 0 2.1740092674779455e-04
GC_12_1033 b_12 NI_12 NS_1033 0 -5.0592004869657922e-03
GC_12_1034 b_12 NI_12 NS_1034 0 1.7016082211230125e-03
GC_12_1035 b_12 NI_12 NS_1035 0 2.4884719812638349e-03
GC_12_1036 b_12 NI_12 NS_1036 0 -9.5763486206148422e-04
GC_12_1037 b_12 NI_12 NS_1037 0 -6.5329668169026266e-03
GC_12_1038 b_12 NI_12 NS_1038 0 3.8846211805321270e-03
GC_12_1039 b_12 NI_12 NS_1039 0 7.4932612544993046e-03
GC_12_1040 b_12 NI_12 NS_1040 0 -1.0960049926956419e-03
GC_12_1041 b_12 NI_12 NS_1041 0 -3.9851227910626215e-03
GC_12_1042 b_12 NI_12 NS_1042 0 4.0409663137632142e-03
GC_12_1043 b_12 NI_12 NS_1043 0 2.8633248923086063e-03
GC_12_1044 b_12 NI_12 NS_1044 0 -3.0534840298027258e-03
GC_12_1045 b_12 NI_12 NS_1045 0 -6.0227358976723934e-03
GC_12_1046 b_12 NI_12 NS_1046 0 7.2373634148458037e-03
GC_12_1047 b_12 NI_12 NS_1047 0 7.9896911475288469e-03
GC_12_1048 b_12 NI_12 NS_1048 0 -4.8114454952553906e-03
GC_12_1049 b_12 NI_12 NS_1049 0 -5.3743564158304381e-04
GC_12_1050 b_12 NI_12 NS_1050 0 5.0204611318347952e-03
GC_12_1051 b_12 NI_12 NS_1051 0 2.4825046595663427e-04
GC_12_1052 b_12 NI_12 NS_1052 0 -4.7581887208287092e-03
GC_12_1053 b_12 NI_12 NS_1053 0 1.8107928901071105e-09
GC_12_1054 b_12 NI_12 NS_1054 0 3.2741501040531965e-09
GC_12_1055 b_12 NI_12 NS_1055 0 -1.4272198943199761e-03
GC_12_1056 b_12 NI_12 NS_1056 0 7.8707210220527232e-03
GC_12_1057 b_12 NI_12 NS_1057 0 -1.7999304571087379e-04
GC_12_1058 b_12 NI_12 NS_1058 0 3.0272429820566481e-03
GC_12_1059 b_12 NI_12 NS_1059 0 -1.3039321363529172e-04
GC_12_1060 b_12 NI_12 NS_1060 0 -3.3752920552105946e-03
GC_12_1061 b_12 NI_12 NS_1061 0 -8.7633793226000469e-04
GC_12_1062 b_12 NI_12 NS_1062 0 7.5304798544569389e-03
GC_12_1063 b_12 NI_12 NS_1063 0 3.7887923511290950e-03
GC_12_1064 b_12 NI_12 NS_1064 0 -6.1573981675864739e-03
GC_12_1065 b_12 NI_12 NS_1065 0 8.6224200991924421e-08
GC_12_1066 b_12 NI_12 NS_1066 0 -3.5295605187751478e-07
GC_12_1067 b_12 NI_12 NS_1067 0 6.7186821084001622e-03
GC_12_1068 b_12 NI_12 NS_1068 0 -5.3194058456996441e-03
GC_12_1069 b_12 NI_12 NS_1069 0 -2.6111750021721738e-03
GC_12_1070 b_12 NI_12 NS_1070 0 6.0542434733270355e-03
GC_12_1071 b_12 NI_12 NS_1071 0 -4.2922721003970940e-03
GC_12_1072 b_12 NI_12 NS_1072 0 1.4428546680421502e-05
GC_12_1073 b_12 NI_12 NS_1073 0 2.7173858195240711e-03
GC_12_1074 b_12 NI_12 NS_1074 0 -6.2039927976014929e-03
GC_12_1075 b_12 NI_12 NS_1075 0 2.0957202069938567e-03
GC_12_1076 b_12 NI_12 NS_1076 0 3.2562858946081318e-03
GC_12_1077 b_12 NI_12 NS_1077 0 -1.9700288888947369e-03
GC_12_1078 b_12 NI_12 NS_1078 0 -4.4205336936085741e-03
GC_12_1079 b_12 NI_12 NS_1079 0 2.8640819012434445e-03
GC_12_1080 b_12 NI_12 NS_1080 0 8.0083594488233774e-03
GC_12_1081 b_12 NI_12 NS_1081 0 -1.1185279376495169e-02
GC_12_1082 b_12 NI_12 NS_1082 0 8.4685599379781664e-09
GC_12_1083 b_12 NI_12 NS_1083 0 9.8720479039848735e-07
GC_12_1084 b_12 NI_12 NS_1084 0 3.6199545496263432e-05
GC_12_1085 b_12 NI_12 NS_1085 0 4.3662912875136670e-03
GC_12_1086 b_12 NI_12 NS_1086 0 -3.4896484630100102e-03
GC_12_1087 b_12 NI_12 NS_1087 0 -3.7149060354284510e-03
GC_12_1088 b_12 NI_12 NS_1088 0 6.2509109946303019e-03
GC_12_1089 b_12 NI_12 NS_1089 0 -8.7863142414627803e-03
GC_12_1090 b_12 NI_12 NS_1090 0 -5.9489752875886487e-03
GC_12_1091 b_12 NI_12 NS_1091 0 9.1761797798189416e-03
GC_12_1092 b_12 NI_12 NS_1092 0 -5.9808517457276252e-03
GC_12_1093 b_12 NI_12 NS_1093 0 7.1653526999403971e-03
GC_12_1094 b_12 NI_12 NS_1094 0 1.1911537129995464e-02
GC_12_1095 b_12 NI_12 NS_1095 0 -4.2323324249870925e-03
GC_12_1096 b_12 NI_12 NS_1096 0 -1.1251858155896866e-03
GC_12_1097 b_12 NI_12 NS_1097 0 -8.8793679314604166e-03
GC_12_1098 b_12 NI_12 NS_1098 0 -4.5104630038791677e-04
GC_12_1099 b_12 NI_12 NS_1099 0 1.4527755321812922e-02
GC_12_1100 b_12 NI_12 NS_1100 0 -1.0355613445957331e-02
GC_12_1101 b_12 NI_12 NS_1101 0 1.6511277364412210e-02
GC_12_1102 b_12 NI_12 NS_1102 0 4.0488541992527664e-03
GC_12_1103 b_12 NI_12 NS_1103 0 -1.1485096904880397e-02
GC_12_1104 b_12 NI_12 NS_1104 0 -1.9365551308907661e-04
GC_12_1105 b_12 NI_12 NS_1105 0 -1.6607928795363734e-02
GC_12_1106 b_12 NI_12 NS_1106 0 -4.4552658492506662e-02
GC_12_1107 b_12 NI_12 NS_1107 0 1.0667428746024298e-02
GC_12_1108 b_12 NI_12 NS_1108 0 1.0871065886580041e-03
GC_12_1109 b_12 NI_12 NS_1109 0 -4.8262941139429354e-02
GC_12_1110 b_12 NI_12 NS_1110 0 1.1004960874499078e-02
GC_12_1111 b_12 NI_12 NS_1111 0 -1.0464675764068629e-02
GC_12_1112 b_12 NI_12 NS_1112 0 5.4274358073734118e-04
GC_12_1113 b_12 NI_12 NS_1113 0 9.7653670045278022e-03
GC_12_1114 b_12 NI_12 NS_1114 0 -6.1125908729398179e-04
GC_12_1115 b_12 NI_12 NS_1115 0 4.5935001210853678e-03
GC_12_1116 b_12 NI_12 NS_1116 0 2.4194352017548298e-02
GC_12_1117 b_12 NI_12 NS_1117 0 -1.0736723882076676e-02
GC_12_1118 b_12 NI_12 NS_1118 0 1.9985970886217562e-03
GC_12_1119 b_12 NI_12 NS_1119 0 -8.4713551750907144e-03
GC_12_1120 b_12 NI_12 NS_1120 0 -1.3526350664748565e-02
GC_12_1121 b_12 NI_12 NS_1121 0 1.0155187241942214e-02
GC_12_1122 b_12 NI_12 NS_1122 0 9.6274154049786850e-04
GC_12_1123 b_12 NI_12 NS_1123 0 -1.9169415519194162e-02
GC_12_1124 b_12 NI_12 NS_1124 0 2.8673875820675206e-02
GC_12_1125 b_12 NI_12 NS_1125 0 -9.6256271575944768e-03
GC_12_1126 b_12 NI_12 NS_1126 0 -9.4348130219993459e-04
GC_12_1127 b_12 NI_12 NS_1127 0 1.8844253103819108e-03
GC_12_1128 b_12 NI_12 NS_1128 0 -1.3764834336368447e-03
GC_12_1129 b_12 NI_12 NS_1129 0 9.4635237704808906e-03
GC_12_1130 b_12 NI_12 NS_1130 0 -2.5484784349157470e-04
GC_12_1131 b_12 NI_12 NS_1131 0 -1.6533832552837591e-04
GC_12_1132 b_12 NI_12 NS_1132 0 3.0293333407721498e-02
GC_12_1133 b_12 NI_12 NS_1133 0 -8.5338011500219208e-03
GC_12_1134 b_12 NI_12 NS_1134 0 1.7751168612594313e-04
GC_12_1135 b_12 NI_12 NS_1135 0 2.1345969456636597e-04
GC_12_1136 b_12 NI_12 NS_1136 0 -5.4660073177406282e-03
GC_12_1137 b_12 NI_12 NS_1137 0 1.0030303273366429e-02
GC_12_1138 b_12 NI_12 NS_1138 0 -3.4494237350455714e-04
GC_12_1139 b_12 NI_12 NS_1139 0 8.9348145095483889e-03
GC_12_1140 b_12 NI_12 NS_1140 0 2.6406119584732265e-02
GC_12_1141 b_12 NI_12 NS_1141 0 -8.3546000991697872e-03
GC_12_1142 b_12 NI_12 NS_1142 0 1.4014563641278649e-03
GC_12_1143 b_12 NI_12 NS_1143 0 -2.5783439599642252e-03
GC_12_1144 b_12 NI_12 NS_1144 0 -7.3353039518004011e-03
GC_12_1145 b_12 NI_12 NS_1145 0 1.0543965173685813e-02
GC_12_1146 b_12 NI_12 NS_1146 0 -8.2793970013570947e-04
GC_12_1147 b_12 NI_12 NS_1147 0 1.4465642920805419e-02
GC_12_1148 b_12 NI_12 NS_1148 0 1.9992583304367269e-02
GC_12_1149 b_12 NI_12 NS_1149 0 -8.2668735491135646e-03
GC_12_1150 b_12 NI_12 NS_1150 0 2.9582086887172151e-03
GC_12_1151 b_12 NI_12 NS_1151 0 -5.5757779430508358e-03
GC_12_1152 b_12 NI_12 NS_1152 0 -6.9085578495300375e-03
GC_12_1153 b_12 NI_12 NS_1153 0 1.1230527511867252e-02
GC_12_1154 b_12 NI_12 NS_1154 0 -1.3725268963395662e-03
GC_12_1155 b_12 NI_12 NS_1155 0 1.5750276386525788e-02
GC_12_1156 b_12 NI_12 NS_1156 0 1.2967935418100509e-02
GC_12_1157 b_12 NI_12 NS_1157 0 -7.1659215694945006e-03
GC_12_1158 b_12 NI_12 NS_1158 0 5.1306122149715003e-03
GC_12_1159 b_12 NI_12 NS_1159 0 -6.8666947950799303e-03
GC_12_1160 b_12 NI_12 NS_1160 0 -4.8393286791391325e-03
GC_12_1161 b_12 NI_12 NS_1161 0 5.3071452032256577e-09
GC_12_1162 b_12 NI_12 NS_1162 0 4.4270338912678590e-08
GC_12_1163 b_12 NI_12 NS_1163 0 1.2002195621242695e-02
GC_12_1164 b_12 NI_12 NS_1164 0 -2.5686794927881423e-03
GC_12_1165 b_12 NI_12 NS_1165 0 -5.2367704422840956e-03
GC_12_1166 b_12 NI_12 NS_1166 0 4.7118192201663842e-03
GC_12_1167 b_12 NI_12 NS_1167 0 -6.1526742979980875e-03
GC_12_1168 b_12 NI_12 NS_1168 0 -4.3194119094503028e-03
GC_12_1169 b_12 NI_12 NS_1169 0 1.1768575557949313e-02
GC_12_1170 b_12 NI_12 NS_1170 0 -3.7146120562839462e-03
GC_12_1171 b_12 NI_12 NS_1171 0 1.3012617293798103e-02
GC_12_1172 b_12 NI_12 NS_1172 0 9.4653948492795688e-03
GC_12_1173 b_12 NI_12 NS_1173 0 3.9556737042503774e-06
GC_12_1174 b_12 NI_12 NS_1174 0 -9.4249395502127373e-07
GC_12_1175 b_12 NI_12 NS_1175 0 1.6124343467209465e-02
GC_12_1176 b_12 NI_12 NS_1176 0 1.6774829947488624e-02
GC_12_1177 b_12 NI_12 NS_1177 0 1.2055182474557113e-02
GC_12_1178 b_12 NI_12 NS_1178 0 -2.4727508758171472e-03
GC_12_1179 b_12 NI_12 NS_1179 0 -8.3469679066029319e-03
GC_12_1180 b_12 NI_12 NS_1180 0 8.5428313336857812e-05
GC_12_1181 b_12 NI_12 NS_1181 0 1.1349989885884905e-02
GC_12_1182 b_12 NI_12 NS_1182 0 7.3343135227424746e-03
GC_12_1183 b_12 NI_12 NS_1183 0 -4.6479092972973278e-03
GC_12_1184 b_12 NI_12 NS_1184 0 7.3636033677158359e-03
GC_12_1185 b_12 NI_12 NS_1185 0 -8.0750671336778223e-03
GC_12_1186 b_12 NI_12 NS_1186 0 -3.7254214076016812e-03
GC_12_1187 b_12 NI_12 NS_1187 0 1.5991409503421278e-02
GC_12_1188 b_12 NI_12 NS_1188 0 -7.7330097246568908e-03
GC_12_1189 b_12 NI_12 NS_1189 0 -1.5530873157256113e-02
GC_12_1190 b_12 NI_12 NS_1190 0 6.4872979778632533e-09
GC_12_1191 b_12 NI_12 NS_1191 0 -1.0780989021982944e-06
GC_12_1192 b_12 NI_12 NS_1192 0 -2.3175273689931599e-05
GC_12_1193 b_12 NI_12 NS_1193 0 3.3380760691955003e-04
GC_12_1194 b_12 NI_12 NS_1194 0 -2.0548504348944253e-04
GC_12_1195 b_12 NI_12 NS_1195 0 -1.5862582016457952e-03
GC_12_1196 b_12 NI_12 NS_1196 0 -2.3361773046056797e-03
GC_12_1197 b_12 NI_12 NS_1197 0 -6.3216293149614229e-05
GC_12_1198 b_12 NI_12 NS_1198 0 4.3863824873940594e-03
GC_12_1199 b_12 NI_12 NS_1199 0 1.5399051133395962e-03
GC_12_1200 b_12 NI_12 NS_1200 0 -5.9456444705446978e-03
GC_12_1201 b_12 NI_12 NS_1201 0 -4.9710137011665561e-03
GC_12_1202 b_12 NI_12 NS_1202 0 6.5658936317763202e-03
GC_12_1203 b_12 NI_12 NS_1203 0 1.1033053449823658e-03
GC_12_1204 b_12 NI_12 NS_1204 0 -4.8869787764716714e-04
GC_12_1205 b_12 NI_12 NS_1205 0 2.8351196952451992e-03
GC_12_1206 b_12 NI_12 NS_1206 0 2.3742292490102563e-03
GC_12_1207 b_12 NI_12 NS_1207 0 -4.4219533089198430e-03
GC_12_1208 b_12 NI_12 NS_1208 0 -1.3476669330843342e-02
GC_12_1209 b_12 NI_12 NS_1209 0 1.7485556334059275e-03
GC_12_1210 b_12 NI_12 NS_1210 0 1.7702187650705945e-02
GC_12_1211 b_12 NI_12 NS_1211 0 9.8282590706878763e-03
GC_12_1212 b_12 NI_12 NS_1212 0 -2.3328384606742291e-03
GC_12_1213 b_12 NI_12 NS_1213 0 -1.3062251194868316e-02
GC_12_1214 b_12 NI_12 NS_1214 0 2.3406863257323415e-03
GC_12_1215 b_12 NI_12 NS_1215 0 9.2233755125555681e-03
GC_12_1216 b_12 NI_12 NS_1216 0 1.9112829960495541e-03
GC_12_1217 b_12 NI_12 NS_1217 0 -1.7997095729851826e-02
GC_12_1218 b_12 NI_12 NS_1218 0 -6.3438996795458615e-03
GC_12_1219 b_12 NI_12 NS_1219 0 1.5754262411181545e-02
GC_12_1220 b_12 NI_12 NS_1220 0 6.4095332590133830e-03
GC_12_1221 b_12 NI_12 NS_1221 0 8.1027179662440992e-03
GC_12_1222 b_12 NI_12 NS_1222 0 -4.2190607220787164e-03
GC_12_1223 b_12 NI_12 NS_1223 0 -7.4948905236185085e-03
GC_12_1224 b_12 NI_12 NS_1224 0 2.0941358803367991e-03
GC_12_1225 b_12 NI_12 NS_1225 0 6.7044806804505879e-03
GC_12_1226 b_12 NI_12 NS_1226 0 -2.7628598140632416e-03
GC_12_1227 b_12 NI_12 NS_1227 0 -6.5432384031292529e-03
GC_12_1228 b_12 NI_12 NS_1228 0 2.9299444241776256e-03
GC_12_1229 b_12 NI_12 NS_1229 0 7.6773811930028564e-03
GC_12_1230 b_12 NI_12 NS_1230 0 4.6375248856018488e-04
GC_12_1231 b_12 NI_12 NS_1231 0 -9.3401557078821688e-03
GC_12_1232 b_12 NI_12 NS_1232 0 -5.1079558757738163e-03
GC_12_1233 b_12 NI_12 NS_1233 0 6.8551899318491484e-03
GC_12_1234 b_12 NI_12 NS_1234 0 4.0869851681089604e-03
GC_12_1235 b_12 NI_12 NS_1235 0 -3.8349361445254288e-04
GC_12_1236 b_12 NI_12 NS_1236 0 -9.2299640121921479e-04
GC_12_1237 b_12 NI_12 NS_1237 0 5.6963380872603313e-03
GC_12_1238 b_12 NI_12 NS_1238 0 -1.3852984741730473e-03
GC_12_1239 b_12 NI_12 NS_1239 0 -9.1011003941197949e-03
GC_12_1240 b_12 NI_12 NS_1240 0 -1.2296022293431818e-03
GC_12_1241 b_12 NI_12 NS_1241 0 6.0201783816091706e-03
GC_12_1242 b_12 NI_12 NS_1242 0 7.1817207664895530e-04
GC_12_1243 b_12 NI_12 NS_1243 0 -2.6199034951047465e-03
GC_12_1244 b_12 NI_12 NS_1244 0 2.4600089255879100e-04
GC_12_1245 b_12 NI_12 NS_1245 0 6.7218306943101968e-03
GC_12_1246 b_12 NI_12 NS_1246 0 -2.2667468567521419e-03
GC_12_1247 b_12 NI_12 NS_1247 0 -9.2254224935984924e-03
GC_12_1248 b_12 NI_12 NS_1248 0 1.5046042797539642e-03
GC_12_1249 b_12 NI_12 NS_1249 0 5.7525380524020868e-03
GC_12_1250 b_12 NI_12 NS_1250 0 -1.5177994584732273e-03
GC_12_1251 b_12 NI_12 NS_1251 0 -3.2852559397146433e-03
GC_12_1252 b_12 NI_12 NS_1252 0 2.3899129607071442e-03
GC_12_1253 b_12 NI_12 NS_1253 0 7.2874261274708156e-03
GC_12_1254 b_12 NI_12 NS_1254 0 -4.1034637088344286e-03
GC_12_1255 b_12 NI_12 NS_1255 0 -8.5232818672604828e-03
GC_12_1256 b_12 NI_12 NS_1256 0 4.1574411160600483e-03
GC_12_1257 b_12 NI_12 NS_1257 0 4.8370640457208024e-03
GC_12_1258 b_12 NI_12 NS_1258 0 -3.8866661366850882e-03
GC_12_1259 b_12 NI_12 NS_1259 0 -2.3786683759331839e-03
GC_12_1260 b_12 NI_12 NS_1260 0 4.7281098936793825e-03
GC_12_1261 b_12 NI_12 NS_1261 0 7.0803227511904709e-03
GC_12_1262 b_12 NI_12 NS_1262 0 -7.3558597634438084e-03
GC_12_1263 b_12 NI_12 NS_1263 0 -7.0931606049218924e-03
GC_12_1264 b_12 NI_12 NS_1264 0 6.8359968044201871e-03
GC_12_1265 b_12 NI_12 NS_1265 0 1.6811452735816942e-03
GC_12_1266 b_12 NI_12 NS_1266 0 -5.3216374786752658e-03
GC_12_1267 b_12 NI_12 NS_1267 0 5.9853547441598542e-04
GC_12_1268 b_12 NI_12 NS_1268 0 5.4496391680691003e-03
GC_12_1269 b_12 NI_12 NS_1269 0 -4.1282284699775118e-09
GC_12_1270 b_12 NI_12 NS_1270 0 -1.3976315452979372e-08
GC_12_1271 b_12 NI_12 NS_1271 0 2.7262644697522149e-03
GC_12_1272 b_12 NI_12 NS_1272 0 -8.5984898986478132e-03
GC_12_1273 b_12 NI_12 NS_1273 0 8.7601838046867284e-04
GC_12_1274 b_12 NI_12 NS_1274 0 -3.4431550556228369e-03
GC_12_1275 b_12 NI_12 NS_1275 0 6.3792150906627975e-04
GC_12_1276 b_12 NI_12 NS_1276 0 4.0228568730465413e-03
GC_12_1277 b_12 NI_12 NS_1277 0 2.1875523767005286e-03
GC_12_1278 b_12 NI_12 NS_1278 0 -8.1664822243236838e-03
GC_12_1279 b_12 NI_12 NS_1279 0 -3.4772862845492357e-03
GC_12_1280 b_12 NI_12 NS_1280 0 6.9937176392013498e-03
GC_12_1281 b_12 NI_12 NS_1281 0 -8.5503704833925107e-08
GC_12_1282 b_12 NI_12 NS_1282 0 -3.1420277946804829e-07
GC_12_1283 b_12 NI_12 NS_1283 0 -7.9941562743269280e-03
GC_12_1284 b_12 NI_12 NS_1284 0 5.3784298215881756e-03
GC_12_1285 b_12 NI_12 NS_1285 0 4.1818213360579363e-03
GC_12_1286 b_12 NI_12 NS_1286 0 -6.8548439269165663e-03
GC_12_1287 b_12 NI_12 NS_1287 0 5.3337133249184970e-03
GC_12_1288 b_12 NI_12 NS_1288 0 7.4258456466222737e-04
GC_12_1289 b_12 NI_12 NS_1289 0 -2.3535041177444858e-03
GC_12_1290 b_12 NI_12 NS_1290 0 6.8399073945520404e-03
GC_12_1291 b_12 NI_12 NS_1291 0 -1.4841909516084190e-03
GC_12_1292 b_12 NI_12 NS_1292 0 -4.2255112741157704e-03
GC_12_1293 b_12 NI_12 NS_1293 0 2.3638870486138758e-03
GC_12_1294 b_12 NI_12 NS_1294 0 5.0284973850196150e-03
GC_12_1295 b_12 NI_12 NS_1295 0 -1.9828423316084190e-03
GC_12_1296 b_12 NI_12 NS_1296 0 -8.9598437125936545e-03
GD_12_1 b_12 NI_12 NA_1 0 3.3591008775674810e-06
GD_12_2 b_12 NI_12 NA_2 0 -2.2825700879504667e-06
GD_12_3 b_12 NI_12 NA_3 0 8.8115117030140447e-06
GD_12_4 b_12 NI_12 NA_4 0 -1.1882829028417722e-06
GD_12_5 b_12 NI_12 NA_5 0 1.1430792612964073e-05
GD_12_6 b_12 NI_12 NA_6 0 -3.0002492543132885e-06
GD_12_7 b_12 NI_12 NA_7 0 1.9065700481093511e-05
GD_12_8 b_12 NI_12 NA_8 0 2.6760852083171124e-06
GD_12_9 b_12 NI_12 NA_9 0 -1.1524163930707564e-03
GD_12_10 b_12 NI_12 NA_10 0 1.0616351945255224e-02
GD_12_11 b_12 NI_12 NA_11 0 -4.9159271056684424e-03
GD_12_12 b_12 NI_12 NA_12 0 -1.0697627223894317e-02
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 3.8329546824379270e+00
GS_1_1 0 NS_1 NA_1 0 4.7428518688027549e-01
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 1.0843846705160875e+04
GS_2_1 0 NS_2 NA_1 0 4.7428518688027549e-01
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 3.3457029134706481e+03
GS_3_1 0 NS_3 NA_1 0 4.7428518688027549e-01
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 5.4313394337993634e+02
GS_4_1 0 NS_4 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 2.0342898045173075e+02
RS_6 NS_6 0 2.0342898045173075e+02
GL_5 0 NS_5 NS_6 0 2.5883098202682536e-01
GL_6 0 NS_6 NS_5 0 -2.5883098202682536e-01
GS_5_1 0 NS_5 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 1.2739936959261519e+02
RS_8 NS_8 0 1.2739936959261519e+02
GL_7 0 NS_7 NS_8 0 2.5122204303896745e-01
GL_8 0 NS_8 NS_7 0 -2.5122204303896745e-01
GS_7_1 0 NS_7 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 1.1105129555360161e+02
RS_10 NS_10 0 1.1105129555360161e+02
GL_9 0 NS_9 NS_10 0 2.4643422119526687e-01
GL_10 0 NS_10 NS_9 0 -2.4643422119526687e-01
GS_9_1 0 NS_9 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 1.0856580972218713e+02
RS_12 NS_12 0 1.0856580972218713e+02
GL_11 0 NS_11 NS_12 0 2.4007148694878275e-01
GL_12 0 NS_12 NS_11 0 -2.4007148694878275e-01
GS_11_1 0 NS_11 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 1.0135860176893434e+02
RS_14 NS_14 0 1.0135860176893435e+02
GL_13 0 NS_13 NS_14 0 2.3570758371916220e-01
GL_14 0 NS_14 NS_13 0 -2.3570758371916220e-01
GS_13_1 0 NS_13 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 1.2858526276753685e+02
RS_16 NS_16 0 1.2858526276753685e+02
GL_15 0 NS_15 NS_16 0 2.2966634995600790e-01
GL_16 0 NS_16 NS_15 0 -2.2966634995600790e-01
GS_15_1 0 NS_15 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 1.1773437593549667e+02
RS_18 NS_18 0 1.1773437593549667e+02
GL_17 0 NS_17 NS_18 0 2.2732609444056490e-01
GL_18 0 NS_18 NS_17 0 -2.2732609444056490e-01
GS_17_1 0 NS_17 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 9.8170265044265946e+01
RS_20 NS_20 0 9.8170265044265932e+01
GL_19 0 NS_19 NS_20 0 2.2031598117475365e-01
GL_20 0 NS_20 NS_19 0 -2.2031598117475365e-01
GS_19_1 0 NS_19 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 9.5355901421613709e+01
RS_22 NS_22 0 9.5355901421613694e+01
GL_21 0 NS_21 NS_22 0 2.1739680820836188e-01
GL_22 0 NS_22 NS_21 0 -2.1739680820836188e-01
GS_21_1 0 NS_21 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 1.0859722031634941e+02
RS_24 NS_24 0 1.0859722031634941e+02
GL_23 0 NS_23 NS_24 0 2.0887403840929383e-01
GL_24 0 NS_24 NS_23 0 -2.0887403840929383e-01
GS_23_1 0 NS_23 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 7.7959989808728068e+01
RS_26 NS_26 0 7.7959989808728054e+01
GL_25 0 NS_25 NS_26 0 2.0447808896343445e-01
GL_26 0 NS_26 NS_25 0 -2.0447808896343445e-01
GS_25_1 0 NS_25 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 1.1088851678406323e+02
RS_28 NS_28 0 1.1088851678406321e+02
GL_27 0 NS_27 NS_28 0 1.9843399276071924e-01
GL_28 0 NS_28 NS_27 0 -1.9843399276071924e-01
GS_27_1 0 NS_27 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 8.1179760966262847e+01
RS_30 NS_30 0 8.1179760966262847e+01
GL_29 0 NS_29 NS_30 0 1.8978022990658949e-01
GL_30 0 NS_30 NS_29 0 -1.8978022990658949e-01
GS_29_1 0 NS_29 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 1.0523970815054612e+02
RS_32 NS_32 0 1.0523970815054612e+02
GL_31 0 NS_31 NS_32 0 1.8836779078363333e-01
GL_32 0 NS_32 NS_31 0 -1.8836779078363333e-01
GS_31_1 0 NS_31 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 1.1208834663822537e+02
RS_34 NS_34 0 1.1208834663822537e+02
GL_33 0 NS_33 NS_34 0 1.7925451755127267e-01
GL_34 0 NS_34 NS_33 0 -1.7925451755127267e-01
GS_33_1 0 NS_33 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 9.2475617668062213e+01
RS_36 NS_36 0 9.2475617668062199e+01
GL_35 0 NS_35 NS_36 0 1.7507216970358189e-01
GL_36 0 NS_36 NS_35 0 -1.7507216970358189e-01
GS_35_1 0 NS_35 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 1.1555782965375326e+02
RS_38 NS_38 0 1.1555782965375326e+02
GL_37 0 NS_37 NS_38 0 1.6918904340923188e-01
GL_38 0 NS_38 NS_37 0 -1.6918904340923188e-01
GS_37_1 0 NS_37 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 9.6856782813111039e+01
RS_40 NS_40 0 9.6856782813111039e+01
GL_39 0 NS_39 NS_40 0 1.6488898173469207e-01
GL_40 0 NS_40 NS_39 0 -1.6488898173469207e-01
GS_39_1 0 NS_39 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 1.1717534841017003e+02
RS_42 NS_42 0 1.1717534841017003e+02
GL_41 0 NS_41 NS_42 0 1.5866517390841936e-01
GL_42 0 NS_42 NS_41 0 -1.5866517390841936e-01
GS_41_1 0 NS_41 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 8.8607873746940697e+01
RS_44 NS_44 0 8.8607873746940697e+01
GL_43 0 NS_43 NS_44 0 1.5214737618207635e-01
GL_44 0 NS_44 NS_43 0 -1.5214737618207635e-01
GS_43_1 0 NS_43 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 1.1741456484283673e+02
RS_46 NS_46 0 1.1741456484283673e+02
GL_45 0 NS_45 NS_46 0 1.4829748860889613e-01
GL_46 0 NS_46 NS_45 0 -1.4829748860889613e-01
GS_45_1 0 NS_45 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 1.3292289814180702e+02
RS_48 NS_48 0 1.3292289814180702e+02
GL_47 0 NS_47 NS_48 0 1.4243056778188259e-01
GL_48 0 NS_48 NS_47 0 -1.4243056778188259e-01
GS_47_1 0 NS_47 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 1.2325134819531741e+02
RS_50 NS_50 0 1.2325134819531739e+02
GL_49 0 NS_49 NS_50 0 1.3890785074828846e-01
GL_50 0 NS_50 NS_49 0 -1.3890785074828846e-01
GS_49_1 0 NS_49 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 9.1909059882883227e+01
RS_52 NS_52 0 9.1909059882883227e+01
GL_51 0 NS_51 NS_52 0 1.3373879533989103e-01
GL_52 0 NS_52 NS_51 0 -1.3373879533989103e-01
GS_51_1 0 NS_51 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 1.2276824880349510e+02
RS_54 NS_54 0 1.2276824880349510e+02
GL_53 0 NS_53 NS_54 0 1.2885409674522977e-01
GL_54 0 NS_54 NS_53 0 -1.2885409674522977e-01
GS_53_1 0 NS_53 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 1.1612442076026501e+02
RS_56 NS_56 0 1.1612442076026501e+02
GL_55 0 NS_55 NS_56 0 1.2417838026896348e-01
GL_56 0 NS_56 NS_55 0 -1.2417838026896348e-01
GS_55_1 0 NS_55 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 1.2130204223875414e+02
RS_58 NS_58 0 1.2130204223875414e+02
GL_57 0 NS_57 NS_58 0 1.1919240021970828e-01
GL_58 0 NS_58 NS_57 0 -1.1919240021970828e-01
GS_57_1 0 NS_57 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 9.3083309227260045e+01
RS_60 NS_60 0 9.3083309227260045e+01
GL_59 0 NS_59 NS_60 0 1.1485268189050464e-01
GL_60 0 NS_60 NS_59 0 -1.1485268189050464e-01
GS_59_1 0 NS_59 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 1.2387094149263906e+02
RS_62 NS_62 0 1.2387094149263908e+02
GL_61 0 NS_61 NS_62 0 1.0935451806229070e-01
GL_62 0 NS_62 NS_61 0 -1.0935451806229070e-01
GS_61_1 0 NS_61 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 1.1186020221520803e+02
RS_64 NS_64 0 1.1186020221520802e+02
GL_63 0 NS_63 NS_64 0 1.0538242730807947e-01
GL_64 0 NS_64 NS_63 0 -1.0538242730807947e-01
GS_63_1 0 NS_63 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 1.2031265815570148e+02
RS_66 NS_66 0 1.2031265815570150e+02
GL_65 0 NS_65 NS_66 0 9.9497602364102364e-02
GL_66 0 NS_66 NS_65 0 -9.9497602364102364e-02
GS_65_1 0 NS_65 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 9.6254518048655143e+01
RS_68 NS_68 0 9.6254518048655143e+01
GL_67 0 NS_67 NS_68 0 9.5930770757699110e-02
GL_68 0 NS_68 NS_67 0 -9.5930770757699110e-02
GS_67_1 0 NS_67 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 1.2318640771018909e+02
RS_70 NS_70 0 1.2318640771018909e+02
GL_69 0 NS_69 NS_70 0 8.9880619653662355e-02
GL_70 0 NS_70 NS_69 0 -8.9880619653662355e-02
GS_69_1 0 NS_69 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 1.1312630346155738e+02
RS_72 NS_72 0 1.1312630346155738e+02
GL_71 0 NS_71 NS_72 0 8.6534434501560398e-02
GL_72 0 NS_72 NS_71 0 -8.6534434501560398e-02
GS_71_1 0 NS_71 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 1.1831504703984019e+02
RS_74 NS_74 0 1.1831504703984019e+02
GL_73 0 NS_73 NS_74 0 7.9864296724202116e-02
GL_74 0 NS_74 NS_73 0 -7.9864296724202116e-02
GS_73_1 0 NS_73 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 1.0281987486447559e+02
RS_76 NS_76 0 1.0281987486447559e+02
GL_75 0 NS_75 NS_76 0 7.6950339194481784e-02
GL_76 0 NS_76 NS_75 0 -7.6950339194481784e-02
GS_75_1 0 NS_75 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 1.2230186914382300e+02
RS_78 NS_78 0 1.2230186914382300e+02
GL_77 0 NS_77 NS_78 0 7.0709298709435750e-02
GL_78 0 NS_78 NS_77 0 -7.0709298709435750e-02
GS_77_1 0 NS_77 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 1.2215699953322022e+02
RS_80 NS_80 0 1.2215699953322020e+02
GL_79 0 NS_79 NS_80 0 6.7518227185671367e-02
GL_80 0 NS_80 NS_79 0 -6.7518227185671367e-02
GS_79_1 0 NS_79 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 3.4305564408226764e+03
RS_82 NS_82 0 3.4305564408226769e+03
GL_81 0 NS_81 NS_82 0 5.4396471187208063e-02
GL_82 0 NS_82 NS_81 0 -5.4396471187208063e-02
GS_81_1 0 NS_81 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 1.1894859826238778e+02
RS_84 NS_84 0 1.1894859826238779e+02
GL_83 0 NS_83 NS_84 0 6.0591569497719031e-02
GL_84 0 NS_84 NS_83 0 -6.0591569497719031e-02
GS_83_1 0 NS_83 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 1.3537641711503298e+02
RS_86 NS_86 0 1.3537641711503298e+02
GL_85 0 NS_85 NS_86 0 5.1190778164089609e-02
GL_86 0 NS_86 NS_85 0 -5.1190778164089609e-02
GS_85_1 0 NS_85 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 1.3105452427659637e+02
RS_88 NS_88 0 1.3105452427659637e+02
GL_87 0 NS_87 NS_88 0 4.7418984574880592e-02
GL_88 0 NS_88 NS_87 0 -4.7418984574880592e-02
GS_87_1 0 NS_87 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 1.2170234397098790e+02
RS_90 NS_90 0 1.2170234397098790e+02
GL_89 0 NS_89 NS_90 0 4.0778813929127578e-02
GL_90 0 NS_90 NS_89 0 -4.0778813929127578e-02
GS_89_1 0 NS_89 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 1.1550510326517782e+02
RS_92 NS_92 0 1.1550510326517782e+02
GL_91 0 NS_91 NS_92 0 5.7236026076957713e-02
GL_92 0 NS_92 NS_91 0 -5.7236026076957713e-02
GS_91_1 0 NS_91 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 6.2039157456337159e+02
RS_94 NS_94 0 6.2039157456337159e+02
GL_93 0 NS_93 NS_94 0 1.9354364738401211e-02
GL_94 0 NS_94 NS_93 0 -1.9354364738401211e-02
GS_93_1 0 NS_93 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 1.1050313240441588e+02
RS_96 NS_96 0 1.1050313240441587e+02
GL_95 0 NS_95 NS_96 0 1.6472588786558075e-02
GL_96 0 NS_96 NS_95 0 -1.6472588786558075e-02
GS_95_1 0 NS_95 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 1.2869119986945731e+02
RS_98 NS_98 0 1.2869119986945731e+02
GL_97 0 NS_97 NS_98 0 2.0888592987579706e-02
GL_98 0 NS_98 NS_97 0 -2.0888592987579706e-02
GS_97_1 0 NS_97 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 1.4314560950270646e+02
RS_100 NS_100 0 1.4314560950270646e+02
GL_99 0 NS_99 NS_100 0 9.7871236580563716e-03
GL_100 0 NS_100 NS_99 0 -9.7871236580563716e-03
GS_99_1 0 NS_99 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 1.1863004336811436e+02
RS_102 NS_102 0 1.1863004336811436e+02
GL_101 0 NS_101 NS_102 0 3.7627463994326378e-02
GL_102 0 NS_102 NS_101 0 -3.7627463994326378e-02
GS_101_1 0 NS_101 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 1.2686172273444870e+02
RS_104 NS_104 0 1.2686172273444869e+02
GL_103 0 NS_103 NS_104 0 3.1975218188091938e-02
GL_104 0 NS_104 NS_103 0 -3.1975218188091938e-02
GS_103_1 0 NS_103 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 1.3141621772977734e+02
RS_106 NS_106 0 1.3141621772977737e+02
GL_105 0 NS_105 NS_106 0 2.8228381102665165e-02
GL_106 0 NS_106 NS_105 0 -2.8228381102665165e-02
GS_105_1 0 NS_105 NA_1 0 4.7428518688027549e-01
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 1.2452833644614726e+02
RS_108 NS_108 0 1.2452833644614726e+02
GL_107 0 NS_107 NS_108 0 2.1457325426059259e-03
GL_108 0 NS_108 NS_107 0 -2.1457325426059259e-03
GS_107_1 0 NS_107 NA_1 0 4.7428518688027549e-01
*
* Real pole n. 109
CS_109 NS_109 0 9.9999999999999998e-13
RS_109 NS_109 0 3.8329546824379270e+00
GS_109_2 0 NS_109 NA_2 0 4.7428518688027549e-01
*
* Real pole n. 110
CS_110 NS_110 0 9.9999999999999998e-13
RS_110 NS_110 0 1.0843846705160875e+04
GS_110_2 0 NS_110 NA_2 0 4.7428518688027549e-01
*
* Real pole n. 111
CS_111 NS_111 0 9.9999999999999998e-13
RS_111 NS_111 0 3.3457029134706481e+03
GS_111_2 0 NS_111 NA_2 0 4.7428518688027549e-01
*
* Real pole n. 112
CS_112 NS_112 0 9.9999999999999998e-13
RS_112 NS_112 0 5.4313394337993634e+02
GS_112_2 0 NS_112 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 2.0342898045173075e+02
RS_114 NS_114 0 2.0342898045173075e+02
GL_113 0 NS_113 NS_114 0 2.5883098202682536e-01
GL_114 0 NS_114 NS_113 0 -2.5883098202682536e-01
GS_113_2 0 NS_113 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 1.2739936959261519e+02
RS_116 NS_116 0 1.2739936959261519e+02
GL_115 0 NS_115 NS_116 0 2.5122204303896745e-01
GL_116 0 NS_116 NS_115 0 -2.5122204303896745e-01
GS_115_2 0 NS_115 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 1.1105129555360161e+02
RS_118 NS_118 0 1.1105129555360161e+02
GL_117 0 NS_117 NS_118 0 2.4643422119526687e-01
GL_118 0 NS_118 NS_117 0 -2.4643422119526687e-01
GS_117_2 0 NS_117 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 1.0856580972218713e+02
RS_120 NS_120 0 1.0856580972218713e+02
GL_119 0 NS_119 NS_120 0 2.4007148694878275e-01
GL_120 0 NS_120 NS_119 0 -2.4007148694878275e-01
GS_119_2 0 NS_119 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 1.0135860176893434e+02
RS_122 NS_122 0 1.0135860176893435e+02
GL_121 0 NS_121 NS_122 0 2.3570758371916220e-01
GL_122 0 NS_122 NS_121 0 -2.3570758371916220e-01
GS_121_2 0 NS_121 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 1.2858526276753685e+02
RS_124 NS_124 0 1.2858526276753685e+02
GL_123 0 NS_123 NS_124 0 2.2966634995600790e-01
GL_124 0 NS_124 NS_123 0 -2.2966634995600790e-01
GS_123_2 0 NS_123 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 1.1773437593549667e+02
RS_126 NS_126 0 1.1773437593549667e+02
GL_125 0 NS_125 NS_126 0 2.2732609444056490e-01
GL_126 0 NS_126 NS_125 0 -2.2732609444056490e-01
GS_125_2 0 NS_125 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 9.8170265044265946e+01
RS_128 NS_128 0 9.8170265044265932e+01
GL_127 0 NS_127 NS_128 0 2.2031598117475365e-01
GL_128 0 NS_128 NS_127 0 -2.2031598117475365e-01
GS_127_2 0 NS_127 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 9.5355901421613709e+01
RS_130 NS_130 0 9.5355901421613694e+01
GL_129 0 NS_129 NS_130 0 2.1739680820836188e-01
GL_130 0 NS_130 NS_129 0 -2.1739680820836188e-01
GS_129_2 0 NS_129 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 1.0859722031634941e+02
RS_132 NS_132 0 1.0859722031634941e+02
GL_131 0 NS_131 NS_132 0 2.0887403840929383e-01
GL_132 0 NS_132 NS_131 0 -2.0887403840929383e-01
GS_131_2 0 NS_131 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 133/134
CS_133 NS_133 0 9.9999999999999998e-13
CS_134 NS_134 0 9.9999999999999998e-13
RS_133 NS_133 0 7.7959989808728068e+01
RS_134 NS_134 0 7.7959989808728054e+01
GL_133 0 NS_133 NS_134 0 2.0447808896343445e-01
GL_134 0 NS_134 NS_133 0 -2.0447808896343445e-01
GS_133_2 0 NS_133 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 1.1088851678406323e+02
RS_136 NS_136 0 1.1088851678406321e+02
GL_135 0 NS_135 NS_136 0 1.9843399276071924e-01
GL_136 0 NS_136 NS_135 0 -1.9843399276071924e-01
GS_135_2 0 NS_135 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 8.1179760966262847e+01
RS_138 NS_138 0 8.1179760966262847e+01
GL_137 0 NS_137 NS_138 0 1.8978022990658949e-01
GL_138 0 NS_138 NS_137 0 -1.8978022990658949e-01
GS_137_2 0 NS_137 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 1.0523970815054612e+02
RS_140 NS_140 0 1.0523970815054612e+02
GL_139 0 NS_139 NS_140 0 1.8836779078363333e-01
GL_140 0 NS_140 NS_139 0 -1.8836779078363333e-01
GS_139_2 0 NS_139 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 1.1208834663822537e+02
RS_142 NS_142 0 1.1208834663822537e+02
GL_141 0 NS_141 NS_142 0 1.7925451755127267e-01
GL_142 0 NS_142 NS_141 0 -1.7925451755127267e-01
GS_141_2 0 NS_141 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 9.2475617668062213e+01
RS_144 NS_144 0 9.2475617668062199e+01
GL_143 0 NS_143 NS_144 0 1.7507216970358189e-01
GL_144 0 NS_144 NS_143 0 -1.7507216970358189e-01
GS_143_2 0 NS_143 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 1.1555782965375326e+02
RS_146 NS_146 0 1.1555782965375326e+02
GL_145 0 NS_145 NS_146 0 1.6918904340923188e-01
GL_146 0 NS_146 NS_145 0 -1.6918904340923188e-01
GS_145_2 0 NS_145 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 9.6856782813111039e+01
RS_148 NS_148 0 9.6856782813111039e+01
GL_147 0 NS_147 NS_148 0 1.6488898173469207e-01
GL_148 0 NS_148 NS_147 0 -1.6488898173469207e-01
GS_147_2 0 NS_147 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 1.1717534841017003e+02
RS_150 NS_150 0 1.1717534841017003e+02
GL_149 0 NS_149 NS_150 0 1.5866517390841936e-01
GL_150 0 NS_150 NS_149 0 -1.5866517390841936e-01
GS_149_2 0 NS_149 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 8.8607873746940697e+01
RS_152 NS_152 0 8.8607873746940697e+01
GL_151 0 NS_151 NS_152 0 1.5214737618207635e-01
GL_152 0 NS_152 NS_151 0 -1.5214737618207635e-01
GS_151_2 0 NS_151 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 1.1741456484283673e+02
RS_154 NS_154 0 1.1741456484283673e+02
GL_153 0 NS_153 NS_154 0 1.4829748860889613e-01
GL_154 0 NS_154 NS_153 0 -1.4829748860889613e-01
GS_153_2 0 NS_153 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 1.3292289814180702e+02
RS_156 NS_156 0 1.3292289814180702e+02
GL_155 0 NS_155 NS_156 0 1.4243056778188259e-01
GL_156 0 NS_156 NS_155 0 -1.4243056778188259e-01
GS_155_2 0 NS_155 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 1.2325134819531741e+02
RS_158 NS_158 0 1.2325134819531739e+02
GL_157 0 NS_157 NS_158 0 1.3890785074828846e-01
GL_158 0 NS_158 NS_157 0 -1.3890785074828846e-01
GS_157_2 0 NS_157 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 9.1909059882883227e+01
RS_160 NS_160 0 9.1909059882883227e+01
GL_159 0 NS_159 NS_160 0 1.3373879533989103e-01
GL_160 0 NS_160 NS_159 0 -1.3373879533989103e-01
GS_159_2 0 NS_159 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 1.2276824880349510e+02
RS_162 NS_162 0 1.2276824880349510e+02
GL_161 0 NS_161 NS_162 0 1.2885409674522977e-01
GL_162 0 NS_162 NS_161 0 -1.2885409674522977e-01
GS_161_2 0 NS_161 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 163/164
CS_163 NS_163 0 9.9999999999999998e-13
CS_164 NS_164 0 9.9999999999999998e-13
RS_163 NS_163 0 1.1612442076026501e+02
RS_164 NS_164 0 1.1612442076026501e+02
GL_163 0 NS_163 NS_164 0 1.2417838026896348e-01
GL_164 0 NS_164 NS_163 0 -1.2417838026896348e-01
GS_163_2 0 NS_163 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 1.2130204223875414e+02
RS_166 NS_166 0 1.2130204223875414e+02
GL_165 0 NS_165 NS_166 0 1.1919240021970828e-01
GL_166 0 NS_166 NS_165 0 -1.1919240021970828e-01
GS_165_2 0 NS_165 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 9.3083309227260045e+01
RS_168 NS_168 0 9.3083309227260045e+01
GL_167 0 NS_167 NS_168 0 1.1485268189050464e-01
GL_168 0 NS_168 NS_167 0 -1.1485268189050464e-01
GS_167_2 0 NS_167 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 1.2387094149263906e+02
RS_170 NS_170 0 1.2387094149263908e+02
GL_169 0 NS_169 NS_170 0 1.0935451806229070e-01
GL_170 0 NS_170 NS_169 0 -1.0935451806229070e-01
GS_169_2 0 NS_169 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 1.1186020221520803e+02
RS_172 NS_172 0 1.1186020221520802e+02
GL_171 0 NS_171 NS_172 0 1.0538242730807947e-01
GL_172 0 NS_172 NS_171 0 -1.0538242730807947e-01
GS_171_2 0 NS_171 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 1.2031265815570148e+02
RS_174 NS_174 0 1.2031265815570150e+02
GL_173 0 NS_173 NS_174 0 9.9497602364102364e-02
GL_174 0 NS_174 NS_173 0 -9.9497602364102364e-02
GS_173_2 0 NS_173 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 9.6254518048655143e+01
RS_176 NS_176 0 9.6254518048655143e+01
GL_175 0 NS_175 NS_176 0 9.5930770757699110e-02
GL_176 0 NS_176 NS_175 0 -9.5930770757699110e-02
GS_175_2 0 NS_175 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 1.2318640771018909e+02
RS_178 NS_178 0 1.2318640771018909e+02
GL_177 0 NS_177 NS_178 0 8.9880619653662355e-02
GL_178 0 NS_178 NS_177 0 -8.9880619653662355e-02
GS_177_2 0 NS_177 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 1.1312630346155738e+02
RS_180 NS_180 0 1.1312630346155738e+02
GL_179 0 NS_179 NS_180 0 8.6534434501560398e-02
GL_180 0 NS_180 NS_179 0 -8.6534434501560398e-02
GS_179_2 0 NS_179 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 181/182
CS_181 NS_181 0 9.9999999999999998e-13
CS_182 NS_182 0 9.9999999999999998e-13
RS_181 NS_181 0 1.1831504703984019e+02
RS_182 NS_182 0 1.1831504703984019e+02
GL_181 0 NS_181 NS_182 0 7.9864296724202116e-02
GL_182 0 NS_182 NS_181 0 -7.9864296724202116e-02
GS_181_2 0 NS_181 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 183/184
CS_183 NS_183 0 9.9999999999999998e-13
CS_184 NS_184 0 9.9999999999999998e-13
RS_183 NS_183 0 1.0281987486447559e+02
RS_184 NS_184 0 1.0281987486447559e+02
GL_183 0 NS_183 NS_184 0 7.6950339194481784e-02
GL_184 0 NS_184 NS_183 0 -7.6950339194481784e-02
GS_183_2 0 NS_183 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 1.2230186914382300e+02
RS_186 NS_186 0 1.2230186914382300e+02
GL_185 0 NS_185 NS_186 0 7.0709298709435750e-02
GL_186 0 NS_186 NS_185 0 -7.0709298709435750e-02
GS_185_2 0 NS_185 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 1.2215699953322022e+02
RS_188 NS_188 0 1.2215699953322020e+02
GL_187 0 NS_187 NS_188 0 6.7518227185671367e-02
GL_188 0 NS_188 NS_187 0 -6.7518227185671367e-02
GS_187_2 0 NS_187 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 3.4305564408226764e+03
RS_190 NS_190 0 3.4305564408226769e+03
GL_189 0 NS_189 NS_190 0 5.4396471187208063e-02
GL_190 0 NS_190 NS_189 0 -5.4396471187208063e-02
GS_189_2 0 NS_189 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 1.1894859826238778e+02
RS_192 NS_192 0 1.1894859826238779e+02
GL_191 0 NS_191 NS_192 0 6.0591569497719031e-02
GL_192 0 NS_192 NS_191 0 -6.0591569497719031e-02
GS_191_2 0 NS_191 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 1.3537641711503298e+02
RS_194 NS_194 0 1.3537641711503298e+02
GL_193 0 NS_193 NS_194 0 5.1190778164089609e-02
GL_194 0 NS_194 NS_193 0 -5.1190778164089609e-02
GS_193_2 0 NS_193 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 1.3105452427659637e+02
RS_196 NS_196 0 1.3105452427659637e+02
GL_195 0 NS_195 NS_196 0 4.7418984574880592e-02
GL_196 0 NS_196 NS_195 0 -4.7418984574880592e-02
GS_195_2 0 NS_195 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 1.2170234397098790e+02
RS_198 NS_198 0 1.2170234397098790e+02
GL_197 0 NS_197 NS_198 0 4.0778813929127578e-02
GL_198 0 NS_198 NS_197 0 -4.0778813929127578e-02
GS_197_2 0 NS_197 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 1.1550510326517782e+02
RS_200 NS_200 0 1.1550510326517782e+02
GL_199 0 NS_199 NS_200 0 5.7236026076957713e-02
GL_200 0 NS_200 NS_199 0 -5.7236026076957713e-02
GS_199_2 0 NS_199 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 201/202
CS_201 NS_201 0 9.9999999999999998e-13
CS_202 NS_202 0 9.9999999999999998e-13
RS_201 NS_201 0 6.2039157456337159e+02
RS_202 NS_202 0 6.2039157456337159e+02
GL_201 0 NS_201 NS_202 0 1.9354364738401211e-02
GL_202 0 NS_202 NS_201 0 -1.9354364738401211e-02
GS_201_2 0 NS_201 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 203/204
CS_203 NS_203 0 9.9999999999999998e-13
CS_204 NS_204 0 9.9999999999999998e-13
RS_203 NS_203 0 1.1050313240441588e+02
RS_204 NS_204 0 1.1050313240441587e+02
GL_203 0 NS_203 NS_204 0 1.6472588786558075e-02
GL_204 0 NS_204 NS_203 0 -1.6472588786558075e-02
GS_203_2 0 NS_203 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 1.2869119986945731e+02
RS_206 NS_206 0 1.2869119986945731e+02
GL_205 0 NS_205 NS_206 0 2.0888592987579706e-02
GL_206 0 NS_206 NS_205 0 -2.0888592987579706e-02
GS_205_2 0 NS_205 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 1.4314560950270646e+02
RS_208 NS_208 0 1.4314560950270646e+02
GL_207 0 NS_207 NS_208 0 9.7871236580563716e-03
GL_208 0 NS_208 NS_207 0 -9.7871236580563716e-03
GS_207_2 0 NS_207 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 1.1863004336811436e+02
RS_210 NS_210 0 1.1863004336811436e+02
GL_209 0 NS_209 NS_210 0 3.7627463994326378e-02
GL_210 0 NS_210 NS_209 0 -3.7627463994326378e-02
GS_209_2 0 NS_209 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 1.2686172273444870e+02
RS_212 NS_212 0 1.2686172273444869e+02
GL_211 0 NS_211 NS_212 0 3.1975218188091938e-02
GL_212 0 NS_212 NS_211 0 -3.1975218188091938e-02
GS_211_2 0 NS_211 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 1.3141621772977734e+02
RS_214 NS_214 0 1.3141621772977737e+02
GL_213 0 NS_213 NS_214 0 2.8228381102665165e-02
GL_214 0 NS_214 NS_213 0 -2.8228381102665165e-02
GS_213_2 0 NS_213 NA_2 0 4.7428518688027549e-01
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 1.2452833644614726e+02
RS_216 NS_216 0 1.2452833644614726e+02
GL_215 0 NS_215 NS_216 0 2.1457325426059259e-03
GL_216 0 NS_216 NS_215 0 -2.1457325426059259e-03
GS_215_2 0 NS_215 NA_2 0 4.7428518688027549e-01
*
* Real pole n. 217
CS_217 NS_217 0 9.9999999999999998e-13
RS_217 NS_217 0 3.8329546824379270e+00
GS_217_3 0 NS_217 NA_3 0 4.7428518688027549e-01
*
* Real pole n. 218
CS_218 NS_218 0 9.9999999999999998e-13
RS_218 NS_218 0 1.0843846705160875e+04
GS_218_3 0 NS_218 NA_3 0 4.7428518688027549e-01
*
* Real pole n. 219
CS_219 NS_219 0 9.9999999999999998e-13
RS_219 NS_219 0 3.3457029134706481e+03
GS_219_3 0 NS_219 NA_3 0 4.7428518688027549e-01
*
* Real pole n. 220
CS_220 NS_220 0 9.9999999999999998e-13
RS_220 NS_220 0 5.4313394337993634e+02
GS_220_3 0 NS_220 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 221/222
CS_221 NS_221 0 9.9999999999999998e-13
CS_222 NS_222 0 9.9999999999999998e-13
RS_221 NS_221 0 2.0342898045173075e+02
RS_222 NS_222 0 2.0342898045173075e+02
GL_221 0 NS_221 NS_222 0 2.5883098202682536e-01
GL_222 0 NS_222 NS_221 0 -2.5883098202682536e-01
GS_221_3 0 NS_221 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 223/224
CS_223 NS_223 0 9.9999999999999998e-13
CS_224 NS_224 0 9.9999999999999998e-13
RS_223 NS_223 0 1.2739936959261519e+02
RS_224 NS_224 0 1.2739936959261519e+02
GL_223 0 NS_223 NS_224 0 2.5122204303896745e-01
GL_224 0 NS_224 NS_223 0 -2.5122204303896745e-01
GS_223_3 0 NS_223 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 225/226
CS_225 NS_225 0 9.9999999999999998e-13
CS_226 NS_226 0 9.9999999999999998e-13
RS_225 NS_225 0 1.1105129555360161e+02
RS_226 NS_226 0 1.1105129555360161e+02
GL_225 0 NS_225 NS_226 0 2.4643422119526687e-01
GL_226 0 NS_226 NS_225 0 -2.4643422119526687e-01
GS_225_3 0 NS_225 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 1.0856580972218713e+02
RS_228 NS_228 0 1.0856580972218713e+02
GL_227 0 NS_227 NS_228 0 2.4007148694878275e-01
GL_228 0 NS_228 NS_227 0 -2.4007148694878275e-01
GS_227_3 0 NS_227 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 229/230
CS_229 NS_229 0 9.9999999999999998e-13
CS_230 NS_230 0 9.9999999999999998e-13
RS_229 NS_229 0 1.0135860176893434e+02
RS_230 NS_230 0 1.0135860176893435e+02
GL_229 0 NS_229 NS_230 0 2.3570758371916220e-01
GL_230 0 NS_230 NS_229 0 -2.3570758371916220e-01
GS_229_3 0 NS_229 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 1.2858526276753685e+02
RS_232 NS_232 0 1.2858526276753685e+02
GL_231 0 NS_231 NS_232 0 2.2966634995600790e-01
GL_232 0 NS_232 NS_231 0 -2.2966634995600790e-01
GS_231_3 0 NS_231 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 1.1773437593549667e+02
RS_234 NS_234 0 1.1773437593549667e+02
GL_233 0 NS_233 NS_234 0 2.2732609444056490e-01
GL_234 0 NS_234 NS_233 0 -2.2732609444056490e-01
GS_233_3 0 NS_233 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 9.8170265044265946e+01
RS_236 NS_236 0 9.8170265044265932e+01
GL_235 0 NS_235 NS_236 0 2.2031598117475365e-01
GL_236 0 NS_236 NS_235 0 -2.2031598117475365e-01
GS_235_3 0 NS_235 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 9.5355901421613709e+01
RS_238 NS_238 0 9.5355901421613694e+01
GL_237 0 NS_237 NS_238 0 2.1739680820836188e-01
GL_238 0 NS_238 NS_237 0 -2.1739680820836188e-01
GS_237_3 0 NS_237 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 1.0859722031634941e+02
RS_240 NS_240 0 1.0859722031634941e+02
GL_239 0 NS_239 NS_240 0 2.0887403840929383e-01
GL_240 0 NS_240 NS_239 0 -2.0887403840929383e-01
GS_239_3 0 NS_239 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 241/242
CS_241 NS_241 0 9.9999999999999998e-13
CS_242 NS_242 0 9.9999999999999998e-13
RS_241 NS_241 0 7.7959989808728068e+01
RS_242 NS_242 0 7.7959989808728054e+01
GL_241 0 NS_241 NS_242 0 2.0447808896343445e-01
GL_242 0 NS_242 NS_241 0 -2.0447808896343445e-01
GS_241_3 0 NS_241 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 243/244
CS_243 NS_243 0 9.9999999999999998e-13
CS_244 NS_244 0 9.9999999999999998e-13
RS_243 NS_243 0 1.1088851678406323e+02
RS_244 NS_244 0 1.1088851678406321e+02
GL_243 0 NS_243 NS_244 0 1.9843399276071924e-01
GL_244 0 NS_244 NS_243 0 -1.9843399276071924e-01
GS_243_3 0 NS_243 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 245/246
CS_245 NS_245 0 9.9999999999999998e-13
CS_246 NS_246 0 9.9999999999999998e-13
RS_245 NS_245 0 8.1179760966262847e+01
RS_246 NS_246 0 8.1179760966262847e+01
GL_245 0 NS_245 NS_246 0 1.8978022990658949e-01
GL_246 0 NS_246 NS_245 0 -1.8978022990658949e-01
GS_245_3 0 NS_245 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 247/248
CS_247 NS_247 0 9.9999999999999998e-13
CS_248 NS_248 0 9.9999999999999998e-13
RS_247 NS_247 0 1.0523970815054612e+02
RS_248 NS_248 0 1.0523970815054612e+02
GL_247 0 NS_247 NS_248 0 1.8836779078363333e-01
GL_248 0 NS_248 NS_247 0 -1.8836779078363333e-01
GS_247_3 0 NS_247 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 249/250
CS_249 NS_249 0 9.9999999999999998e-13
CS_250 NS_250 0 9.9999999999999998e-13
RS_249 NS_249 0 1.1208834663822537e+02
RS_250 NS_250 0 1.1208834663822537e+02
GL_249 0 NS_249 NS_250 0 1.7925451755127267e-01
GL_250 0 NS_250 NS_249 0 -1.7925451755127267e-01
GS_249_3 0 NS_249 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 251/252
CS_251 NS_251 0 9.9999999999999998e-13
CS_252 NS_252 0 9.9999999999999998e-13
RS_251 NS_251 0 9.2475617668062213e+01
RS_252 NS_252 0 9.2475617668062199e+01
GL_251 0 NS_251 NS_252 0 1.7507216970358189e-01
GL_252 0 NS_252 NS_251 0 -1.7507216970358189e-01
GS_251_3 0 NS_251 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 253/254
CS_253 NS_253 0 9.9999999999999998e-13
CS_254 NS_254 0 9.9999999999999998e-13
RS_253 NS_253 0 1.1555782965375326e+02
RS_254 NS_254 0 1.1555782965375326e+02
GL_253 0 NS_253 NS_254 0 1.6918904340923188e-01
GL_254 0 NS_254 NS_253 0 -1.6918904340923188e-01
GS_253_3 0 NS_253 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 255/256
CS_255 NS_255 0 9.9999999999999998e-13
CS_256 NS_256 0 9.9999999999999998e-13
RS_255 NS_255 0 9.6856782813111039e+01
RS_256 NS_256 0 9.6856782813111039e+01
GL_255 0 NS_255 NS_256 0 1.6488898173469207e-01
GL_256 0 NS_256 NS_255 0 -1.6488898173469207e-01
GS_255_3 0 NS_255 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 257/258
CS_257 NS_257 0 9.9999999999999998e-13
CS_258 NS_258 0 9.9999999999999998e-13
RS_257 NS_257 0 1.1717534841017003e+02
RS_258 NS_258 0 1.1717534841017003e+02
GL_257 0 NS_257 NS_258 0 1.5866517390841936e-01
GL_258 0 NS_258 NS_257 0 -1.5866517390841936e-01
GS_257_3 0 NS_257 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 259/260
CS_259 NS_259 0 9.9999999999999998e-13
CS_260 NS_260 0 9.9999999999999998e-13
RS_259 NS_259 0 8.8607873746940697e+01
RS_260 NS_260 0 8.8607873746940697e+01
GL_259 0 NS_259 NS_260 0 1.5214737618207635e-01
GL_260 0 NS_260 NS_259 0 -1.5214737618207635e-01
GS_259_3 0 NS_259 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 261/262
CS_261 NS_261 0 9.9999999999999998e-13
CS_262 NS_262 0 9.9999999999999998e-13
RS_261 NS_261 0 1.1741456484283673e+02
RS_262 NS_262 0 1.1741456484283673e+02
GL_261 0 NS_261 NS_262 0 1.4829748860889613e-01
GL_262 0 NS_262 NS_261 0 -1.4829748860889613e-01
GS_261_3 0 NS_261 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 263/264
CS_263 NS_263 0 9.9999999999999998e-13
CS_264 NS_264 0 9.9999999999999998e-13
RS_263 NS_263 0 1.3292289814180702e+02
RS_264 NS_264 0 1.3292289814180702e+02
GL_263 0 NS_263 NS_264 0 1.4243056778188259e-01
GL_264 0 NS_264 NS_263 0 -1.4243056778188259e-01
GS_263_3 0 NS_263 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 265/266
CS_265 NS_265 0 9.9999999999999998e-13
CS_266 NS_266 0 9.9999999999999998e-13
RS_265 NS_265 0 1.2325134819531741e+02
RS_266 NS_266 0 1.2325134819531739e+02
GL_265 0 NS_265 NS_266 0 1.3890785074828846e-01
GL_266 0 NS_266 NS_265 0 -1.3890785074828846e-01
GS_265_3 0 NS_265 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 267/268
CS_267 NS_267 0 9.9999999999999998e-13
CS_268 NS_268 0 9.9999999999999998e-13
RS_267 NS_267 0 9.1909059882883227e+01
RS_268 NS_268 0 9.1909059882883227e+01
GL_267 0 NS_267 NS_268 0 1.3373879533989103e-01
GL_268 0 NS_268 NS_267 0 -1.3373879533989103e-01
GS_267_3 0 NS_267 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 269/270
CS_269 NS_269 0 9.9999999999999998e-13
CS_270 NS_270 0 9.9999999999999998e-13
RS_269 NS_269 0 1.2276824880349510e+02
RS_270 NS_270 0 1.2276824880349510e+02
GL_269 0 NS_269 NS_270 0 1.2885409674522977e-01
GL_270 0 NS_270 NS_269 0 -1.2885409674522977e-01
GS_269_3 0 NS_269 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 271/272
CS_271 NS_271 0 9.9999999999999998e-13
CS_272 NS_272 0 9.9999999999999998e-13
RS_271 NS_271 0 1.1612442076026501e+02
RS_272 NS_272 0 1.1612442076026501e+02
GL_271 0 NS_271 NS_272 0 1.2417838026896348e-01
GL_272 0 NS_272 NS_271 0 -1.2417838026896348e-01
GS_271_3 0 NS_271 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 273/274
CS_273 NS_273 0 9.9999999999999998e-13
CS_274 NS_274 0 9.9999999999999998e-13
RS_273 NS_273 0 1.2130204223875414e+02
RS_274 NS_274 0 1.2130204223875414e+02
GL_273 0 NS_273 NS_274 0 1.1919240021970828e-01
GL_274 0 NS_274 NS_273 0 -1.1919240021970828e-01
GS_273_3 0 NS_273 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 275/276
CS_275 NS_275 0 9.9999999999999998e-13
CS_276 NS_276 0 9.9999999999999998e-13
RS_275 NS_275 0 9.3083309227260045e+01
RS_276 NS_276 0 9.3083309227260045e+01
GL_275 0 NS_275 NS_276 0 1.1485268189050464e-01
GL_276 0 NS_276 NS_275 0 -1.1485268189050464e-01
GS_275_3 0 NS_275 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 277/278
CS_277 NS_277 0 9.9999999999999998e-13
CS_278 NS_278 0 9.9999999999999998e-13
RS_277 NS_277 0 1.2387094149263906e+02
RS_278 NS_278 0 1.2387094149263908e+02
GL_277 0 NS_277 NS_278 0 1.0935451806229070e-01
GL_278 0 NS_278 NS_277 0 -1.0935451806229070e-01
GS_277_3 0 NS_277 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 279/280
CS_279 NS_279 0 9.9999999999999998e-13
CS_280 NS_280 0 9.9999999999999998e-13
RS_279 NS_279 0 1.1186020221520803e+02
RS_280 NS_280 0 1.1186020221520802e+02
GL_279 0 NS_279 NS_280 0 1.0538242730807947e-01
GL_280 0 NS_280 NS_279 0 -1.0538242730807947e-01
GS_279_3 0 NS_279 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 281/282
CS_281 NS_281 0 9.9999999999999998e-13
CS_282 NS_282 0 9.9999999999999998e-13
RS_281 NS_281 0 1.2031265815570148e+02
RS_282 NS_282 0 1.2031265815570150e+02
GL_281 0 NS_281 NS_282 0 9.9497602364102364e-02
GL_282 0 NS_282 NS_281 0 -9.9497602364102364e-02
GS_281_3 0 NS_281 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 283/284
CS_283 NS_283 0 9.9999999999999998e-13
CS_284 NS_284 0 9.9999999999999998e-13
RS_283 NS_283 0 9.6254518048655143e+01
RS_284 NS_284 0 9.6254518048655143e+01
GL_283 0 NS_283 NS_284 0 9.5930770757699110e-02
GL_284 0 NS_284 NS_283 0 -9.5930770757699110e-02
GS_283_3 0 NS_283 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 285/286
CS_285 NS_285 0 9.9999999999999998e-13
CS_286 NS_286 0 9.9999999999999998e-13
RS_285 NS_285 0 1.2318640771018909e+02
RS_286 NS_286 0 1.2318640771018909e+02
GL_285 0 NS_285 NS_286 0 8.9880619653662355e-02
GL_286 0 NS_286 NS_285 0 -8.9880619653662355e-02
GS_285_3 0 NS_285 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 287/288
CS_287 NS_287 0 9.9999999999999998e-13
CS_288 NS_288 0 9.9999999999999998e-13
RS_287 NS_287 0 1.1312630346155738e+02
RS_288 NS_288 0 1.1312630346155738e+02
GL_287 0 NS_287 NS_288 0 8.6534434501560398e-02
GL_288 0 NS_288 NS_287 0 -8.6534434501560398e-02
GS_287_3 0 NS_287 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 289/290
CS_289 NS_289 0 9.9999999999999998e-13
CS_290 NS_290 0 9.9999999999999998e-13
RS_289 NS_289 0 1.1831504703984019e+02
RS_290 NS_290 0 1.1831504703984019e+02
GL_289 0 NS_289 NS_290 0 7.9864296724202116e-02
GL_290 0 NS_290 NS_289 0 -7.9864296724202116e-02
GS_289_3 0 NS_289 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 291/292
CS_291 NS_291 0 9.9999999999999998e-13
CS_292 NS_292 0 9.9999999999999998e-13
RS_291 NS_291 0 1.0281987486447559e+02
RS_292 NS_292 0 1.0281987486447559e+02
GL_291 0 NS_291 NS_292 0 7.6950339194481784e-02
GL_292 0 NS_292 NS_291 0 -7.6950339194481784e-02
GS_291_3 0 NS_291 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 293/294
CS_293 NS_293 0 9.9999999999999998e-13
CS_294 NS_294 0 9.9999999999999998e-13
RS_293 NS_293 0 1.2230186914382300e+02
RS_294 NS_294 0 1.2230186914382300e+02
GL_293 0 NS_293 NS_294 0 7.0709298709435750e-02
GL_294 0 NS_294 NS_293 0 -7.0709298709435750e-02
GS_293_3 0 NS_293 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 295/296
CS_295 NS_295 0 9.9999999999999998e-13
CS_296 NS_296 0 9.9999999999999998e-13
RS_295 NS_295 0 1.2215699953322022e+02
RS_296 NS_296 0 1.2215699953322020e+02
GL_295 0 NS_295 NS_296 0 6.7518227185671367e-02
GL_296 0 NS_296 NS_295 0 -6.7518227185671367e-02
GS_295_3 0 NS_295 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 297/298
CS_297 NS_297 0 9.9999999999999998e-13
CS_298 NS_298 0 9.9999999999999998e-13
RS_297 NS_297 0 3.4305564408226764e+03
RS_298 NS_298 0 3.4305564408226769e+03
GL_297 0 NS_297 NS_298 0 5.4396471187208063e-02
GL_298 0 NS_298 NS_297 0 -5.4396471187208063e-02
GS_297_3 0 NS_297 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 299/300
CS_299 NS_299 0 9.9999999999999998e-13
CS_300 NS_300 0 9.9999999999999998e-13
RS_299 NS_299 0 1.1894859826238778e+02
RS_300 NS_300 0 1.1894859826238779e+02
GL_299 0 NS_299 NS_300 0 6.0591569497719031e-02
GL_300 0 NS_300 NS_299 0 -6.0591569497719031e-02
GS_299_3 0 NS_299 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 301/302
CS_301 NS_301 0 9.9999999999999998e-13
CS_302 NS_302 0 9.9999999999999998e-13
RS_301 NS_301 0 1.3537641711503298e+02
RS_302 NS_302 0 1.3537641711503298e+02
GL_301 0 NS_301 NS_302 0 5.1190778164089609e-02
GL_302 0 NS_302 NS_301 0 -5.1190778164089609e-02
GS_301_3 0 NS_301 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 303/304
CS_303 NS_303 0 9.9999999999999998e-13
CS_304 NS_304 0 9.9999999999999998e-13
RS_303 NS_303 0 1.3105452427659637e+02
RS_304 NS_304 0 1.3105452427659637e+02
GL_303 0 NS_303 NS_304 0 4.7418984574880592e-02
GL_304 0 NS_304 NS_303 0 -4.7418984574880592e-02
GS_303_3 0 NS_303 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 305/306
CS_305 NS_305 0 9.9999999999999998e-13
CS_306 NS_306 0 9.9999999999999998e-13
RS_305 NS_305 0 1.2170234397098790e+02
RS_306 NS_306 0 1.2170234397098790e+02
GL_305 0 NS_305 NS_306 0 4.0778813929127578e-02
GL_306 0 NS_306 NS_305 0 -4.0778813929127578e-02
GS_305_3 0 NS_305 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 307/308
CS_307 NS_307 0 9.9999999999999998e-13
CS_308 NS_308 0 9.9999999999999998e-13
RS_307 NS_307 0 1.1550510326517782e+02
RS_308 NS_308 0 1.1550510326517782e+02
GL_307 0 NS_307 NS_308 0 5.7236026076957713e-02
GL_308 0 NS_308 NS_307 0 -5.7236026076957713e-02
GS_307_3 0 NS_307 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 309/310
CS_309 NS_309 0 9.9999999999999998e-13
CS_310 NS_310 0 9.9999999999999998e-13
RS_309 NS_309 0 6.2039157456337159e+02
RS_310 NS_310 0 6.2039157456337159e+02
GL_309 0 NS_309 NS_310 0 1.9354364738401211e-02
GL_310 0 NS_310 NS_309 0 -1.9354364738401211e-02
GS_309_3 0 NS_309 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 311/312
CS_311 NS_311 0 9.9999999999999998e-13
CS_312 NS_312 0 9.9999999999999998e-13
RS_311 NS_311 0 1.1050313240441588e+02
RS_312 NS_312 0 1.1050313240441587e+02
GL_311 0 NS_311 NS_312 0 1.6472588786558075e-02
GL_312 0 NS_312 NS_311 0 -1.6472588786558075e-02
GS_311_3 0 NS_311 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 313/314
CS_313 NS_313 0 9.9999999999999998e-13
CS_314 NS_314 0 9.9999999999999998e-13
RS_313 NS_313 0 1.2869119986945731e+02
RS_314 NS_314 0 1.2869119986945731e+02
GL_313 0 NS_313 NS_314 0 2.0888592987579706e-02
GL_314 0 NS_314 NS_313 0 -2.0888592987579706e-02
GS_313_3 0 NS_313 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 315/316
CS_315 NS_315 0 9.9999999999999998e-13
CS_316 NS_316 0 9.9999999999999998e-13
RS_315 NS_315 0 1.4314560950270646e+02
RS_316 NS_316 0 1.4314560950270646e+02
GL_315 0 NS_315 NS_316 0 9.7871236580563716e-03
GL_316 0 NS_316 NS_315 0 -9.7871236580563716e-03
GS_315_3 0 NS_315 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 317/318
CS_317 NS_317 0 9.9999999999999998e-13
CS_318 NS_318 0 9.9999999999999998e-13
RS_317 NS_317 0 1.1863004336811436e+02
RS_318 NS_318 0 1.1863004336811436e+02
GL_317 0 NS_317 NS_318 0 3.7627463994326378e-02
GL_318 0 NS_318 NS_317 0 -3.7627463994326378e-02
GS_317_3 0 NS_317 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 319/320
CS_319 NS_319 0 9.9999999999999998e-13
CS_320 NS_320 0 9.9999999999999998e-13
RS_319 NS_319 0 1.2686172273444870e+02
RS_320 NS_320 0 1.2686172273444869e+02
GL_319 0 NS_319 NS_320 0 3.1975218188091938e-02
GL_320 0 NS_320 NS_319 0 -3.1975218188091938e-02
GS_319_3 0 NS_319 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 321/322
CS_321 NS_321 0 9.9999999999999998e-13
CS_322 NS_322 0 9.9999999999999998e-13
RS_321 NS_321 0 1.3141621772977734e+02
RS_322 NS_322 0 1.3141621772977737e+02
GL_321 0 NS_321 NS_322 0 2.8228381102665165e-02
GL_322 0 NS_322 NS_321 0 -2.8228381102665165e-02
GS_321_3 0 NS_321 NA_3 0 4.7428518688027549e-01
*
* Complex pair n. 323/324
CS_323 NS_323 0 9.9999999999999998e-13
CS_324 NS_324 0 9.9999999999999998e-13
RS_323 NS_323 0 1.2452833644614726e+02
RS_324 NS_324 0 1.2452833644614726e+02
GL_323 0 NS_323 NS_324 0 2.1457325426059259e-03
GL_324 0 NS_324 NS_323 0 -2.1457325426059259e-03
GS_323_3 0 NS_323 NA_3 0 4.7428518688027549e-01
*
* Real pole n. 325
CS_325 NS_325 0 9.9999999999999998e-13
RS_325 NS_325 0 3.8329546824379270e+00
GS_325_4 0 NS_325 NA_4 0 4.7428518688027549e-01
*
* Real pole n. 326
CS_326 NS_326 0 9.9999999999999998e-13
RS_326 NS_326 0 1.0843846705160875e+04
GS_326_4 0 NS_326 NA_4 0 4.7428518688027549e-01
*
* Real pole n. 327
CS_327 NS_327 0 9.9999999999999998e-13
RS_327 NS_327 0 3.3457029134706481e+03
GS_327_4 0 NS_327 NA_4 0 4.7428518688027549e-01
*
* Real pole n. 328
CS_328 NS_328 0 9.9999999999999998e-13
RS_328 NS_328 0 5.4313394337993634e+02
GS_328_4 0 NS_328 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 329/330
CS_329 NS_329 0 9.9999999999999998e-13
CS_330 NS_330 0 9.9999999999999998e-13
RS_329 NS_329 0 2.0342898045173075e+02
RS_330 NS_330 0 2.0342898045173075e+02
GL_329 0 NS_329 NS_330 0 2.5883098202682536e-01
GL_330 0 NS_330 NS_329 0 -2.5883098202682536e-01
GS_329_4 0 NS_329 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 331/332
CS_331 NS_331 0 9.9999999999999998e-13
CS_332 NS_332 0 9.9999999999999998e-13
RS_331 NS_331 0 1.2739936959261519e+02
RS_332 NS_332 0 1.2739936959261519e+02
GL_331 0 NS_331 NS_332 0 2.5122204303896745e-01
GL_332 0 NS_332 NS_331 0 -2.5122204303896745e-01
GS_331_4 0 NS_331 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 333/334
CS_333 NS_333 0 9.9999999999999998e-13
CS_334 NS_334 0 9.9999999999999998e-13
RS_333 NS_333 0 1.1105129555360161e+02
RS_334 NS_334 0 1.1105129555360161e+02
GL_333 0 NS_333 NS_334 0 2.4643422119526687e-01
GL_334 0 NS_334 NS_333 0 -2.4643422119526687e-01
GS_333_4 0 NS_333 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 335/336
CS_335 NS_335 0 9.9999999999999998e-13
CS_336 NS_336 0 9.9999999999999998e-13
RS_335 NS_335 0 1.0856580972218713e+02
RS_336 NS_336 0 1.0856580972218713e+02
GL_335 0 NS_335 NS_336 0 2.4007148694878275e-01
GL_336 0 NS_336 NS_335 0 -2.4007148694878275e-01
GS_335_4 0 NS_335 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 337/338
CS_337 NS_337 0 9.9999999999999998e-13
CS_338 NS_338 0 9.9999999999999998e-13
RS_337 NS_337 0 1.0135860176893434e+02
RS_338 NS_338 0 1.0135860176893435e+02
GL_337 0 NS_337 NS_338 0 2.3570758371916220e-01
GL_338 0 NS_338 NS_337 0 -2.3570758371916220e-01
GS_337_4 0 NS_337 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 339/340
CS_339 NS_339 0 9.9999999999999998e-13
CS_340 NS_340 0 9.9999999999999998e-13
RS_339 NS_339 0 1.2858526276753685e+02
RS_340 NS_340 0 1.2858526276753685e+02
GL_339 0 NS_339 NS_340 0 2.2966634995600790e-01
GL_340 0 NS_340 NS_339 0 -2.2966634995600790e-01
GS_339_4 0 NS_339 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 341/342
CS_341 NS_341 0 9.9999999999999998e-13
CS_342 NS_342 0 9.9999999999999998e-13
RS_341 NS_341 0 1.1773437593549667e+02
RS_342 NS_342 0 1.1773437593549667e+02
GL_341 0 NS_341 NS_342 0 2.2732609444056490e-01
GL_342 0 NS_342 NS_341 0 -2.2732609444056490e-01
GS_341_4 0 NS_341 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 343/344
CS_343 NS_343 0 9.9999999999999998e-13
CS_344 NS_344 0 9.9999999999999998e-13
RS_343 NS_343 0 9.8170265044265946e+01
RS_344 NS_344 0 9.8170265044265932e+01
GL_343 0 NS_343 NS_344 0 2.2031598117475365e-01
GL_344 0 NS_344 NS_343 0 -2.2031598117475365e-01
GS_343_4 0 NS_343 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 345/346
CS_345 NS_345 0 9.9999999999999998e-13
CS_346 NS_346 0 9.9999999999999998e-13
RS_345 NS_345 0 9.5355901421613709e+01
RS_346 NS_346 0 9.5355901421613694e+01
GL_345 0 NS_345 NS_346 0 2.1739680820836188e-01
GL_346 0 NS_346 NS_345 0 -2.1739680820836188e-01
GS_345_4 0 NS_345 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 347/348
CS_347 NS_347 0 9.9999999999999998e-13
CS_348 NS_348 0 9.9999999999999998e-13
RS_347 NS_347 0 1.0859722031634941e+02
RS_348 NS_348 0 1.0859722031634941e+02
GL_347 0 NS_347 NS_348 0 2.0887403840929383e-01
GL_348 0 NS_348 NS_347 0 -2.0887403840929383e-01
GS_347_4 0 NS_347 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 349/350
CS_349 NS_349 0 9.9999999999999998e-13
CS_350 NS_350 0 9.9999999999999998e-13
RS_349 NS_349 0 7.7959989808728068e+01
RS_350 NS_350 0 7.7959989808728054e+01
GL_349 0 NS_349 NS_350 0 2.0447808896343445e-01
GL_350 0 NS_350 NS_349 0 -2.0447808896343445e-01
GS_349_4 0 NS_349 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 351/352
CS_351 NS_351 0 9.9999999999999998e-13
CS_352 NS_352 0 9.9999999999999998e-13
RS_351 NS_351 0 1.1088851678406323e+02
RS_352 NS_352 0 1.1088851678406321e+02
GL_351 0 NS_351 NS_352 0 1.9843399276071924e-01
GL_352 0 NS_352 NS_351 0 -1.9843399276071924e-01
GS_351_4 0 NS_351 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 353/354
CS_353 NS_353 0 9.9999999999999998e-13
CS_354 NS_354 0 9.9999999999999998e-13
RS_353 NS_353 0 8.1179760966262847e+01
RS_354 NS_354 0 8.1179760966262847e+01
GL_353 0 NS_353 NS_354 0 1.8978022990658949e-01
GL_354 0 NS_354 NS_353 0 -1.8978022990658949e-01
GS_353_4 0 NS_353 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 355/356
CS_355 NS_355 0 9.9999999999999998e-13
CS_356 NS_356 0 9.9999999999999998e-13
RS_355 NS_355 0 1.0523970815054612e+02
RS_356 NS_356 0 1.0523970815054612e+02
GL_355 0 NS_355 NS_356 0 1.8836779078363333e-01
GL_356 0 NS_356 NS_355 0 -1.8836779078363333e-01
GS_355_4 0 NS_355 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 357/358
CS_357 NS_357 0 9.9999999999999998e-13
CS_358 NS_358 0 9.9999999999999998e-13
RS_357 NS_357 0 1.1208834663822537e+02
RS_358 NS_358 0 1.1208834663822537e+02
GL_357 0 NS_357 NS_358 0 1.7925451755127267e-01
GL_358 0 NS_358 NS_357 0 -1.7925451755127267e-01
GS_357_4 0 NS_357 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 359/360
CS_359 NS_359 0 9.9999999999999998e-13
CS_360 NS_360 0 9.9999999999999998e-13
RS_359 NS_359 0 9.2475617668062213e+01
RS_360 NS_360 0 9.2475617668062199e+01
GL_359 0 NS_359 NS_360 0 1.7507216970358189e-01
GL_360 0 NS_360 NS_359 0 -1.7507216970358189e-01
GS_359_4 0 NS_359 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 361/362
CS_361 NS_361 0 9.9999999999999998e-13
CS_362 NS_362 0 9.9999999999999998e-13
RS_361 NS_361 0 1.1555782965375326e+02
RS_362 NS_362 0 1.1555782965375326e+02
GL_361 0 NS_361 NS_362 0 1.6918904340923188e-01
GL_362 0 NS_362 NS_361 0 -1.6918904340923188e-01
GS_361_4 0 NS_361 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 363/364
CS_363 NS_363 0 9.9999999999999998e-13
CS_364 NS_364 0 9.9999999999999998e-13
RS_363 NS_363 0 9.6856782813111039e+01
RS_364 NS_364 0 9.6856782813111039e+01
GL_363 0 NS_363 NS_364 0 1.6488898173469207e-01
GL_364 0 NS_364 NS_363 0 -1.6488898173469207e-01
GS_363_4 0 NS_363 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 365/366
CS_365 NS_365 0 9.9999999999999998e-13
CS_366 NS_366 0 9.9999999999999998e-13
RS_365 NS_365 0 1.1717534841017003e+02
RS_366 NS_366 0 1.1717534841017003e+02
GL_365 0 NS_365 NS_366 0 1.5866517390841936e-01
GL_366 0 NS_366 NS_365 0 -1.5866517390841936e-01
GS_365_4 0 NS_365 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 367/368
CS_367 NS_367 0 9.9999999999999998e-13
CS_368 NS_368 0 9.9999999999999998e-13
RS_367 NS_367 0 8.8607873746940697e+01
RS_368 NS_368 0 8.8607873746940697e+01
GL_367 0 NS_367 NS_368 0 1.5214737618207635e-01
GL_368 0 NS_368 NS_367 0 -1.5214737618207635e-01
GS_367_4 0 NS_367 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 369/370
CS_369 NS_369 0 9.9999999999999998e-13
CS_370 NS_370 0 9.9999999999999998e-13
RS_369 NS_369 0 1.1741456484283673e+02
RS_370 NS_370 0 1.1741456484283673e+02
GL_369 0 NS_369 NS_370 0 1.4829748860889613e-01
GL_370 0 NS_370 NS_369 0 -1.4829748860889613e-01
GS_369_4 0 NS_369 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 371/372
CS_371 NS_371 0 9.9999999999999998e-13
CS_372 NS_372 0 9.9999999999999998e-13
RS_371 NS_371 0 1.3292289814180702e+02
RS_372 NS_372 0 1.3292289814180702e+02
GL_371 0 NS_371 NS_372 0 1.4243056778188259e-01
GL_372 0 NS_372 NS_371 0 -1.4243056778188259e-01
GS_371_4 0 NS_371 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 373/374
CS_373 NS_373 0 9.9999999999999998e-13
CS_374 NS_374 0 9.9999999999999998e-13
RS_373 NS_373 0 1.2325134819531741e+02
RS_374 NS_374 0 1.2325134819531739e+02
GL_373 0 NS_373 NS_374 0 1.3890785074828846e-01
GL_374 0 NS_374 NS_373 0 -1.3890785074828846e-01
GS_373_4 0 NS_373 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 375/376
CS_375 NS_375 0 9.9999999999999998e-13
CS_376 NS_376 0 9.9999999999999998e-13
RS_375 NS_375 0 9.1909059882883227e+01
RS_376 NS_376 0 9.1909059882883227e+01
GL_375 0 NS_375 NS_376 0 1.3373879533989103e-01
GL_376 0 NS_376 NS_375 0 -1.3373879533989103e-01
GS_375_4 0 NS_375 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 377/378
CS_377 NS_377 0 9.9999999999999998e-13
CS_378 NS_378 0 9.9999999999999998e-13
RS_377 NS_377 0 1.2276824880349510e+02
RS_378 NS_378 0 1.2276824880349510e+02
GL_377 0 NS_377 NS_378 0 1.2885409674522977e-01
GL_378 0 NS_378 NS_377 0 -1.2885409674522977e-01
GS_377_4 0 NS_377 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 379/380
CS_379 NS_379 0 9.9999999999999998e-13
CS_380 NS_380 0 9.9999999999999998e-13
RS_379 NS_379 0 1.1612442076026501e+02
RS_380 NS_380 0 1.1612442076026501e+02
GL_379 0 NS_379 NS_380 0 1.2417838026896348e-01
GL_380 0 NS_380 NS_379 0 -1.2417838026896348e-01
GS_379_4 0 NS_379 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 381/382
CS_381 NS_381 0 9.9999999999999998e-13
CS_382 NS_382 0 9.9999999999999998e-13
RS_381 NS_381 0 1.2130204223875414e+02
RS_382 NS_382 0 1.2130204223875414e+02
GL_381 0 NS_381 NS_382 0 1.1919240021970828e-01
GL_382 0 NS_382 NS_381 0 -1.1919240021970828e-01
GS_381_4 0 NS_381 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 383/384
CS_383 NS_383 0 9.9999999999999998e-13
CS_384 NS_384 0 9.9999999999999998e-13
RS_383 NS_383 0 9.3083309227260045e+01
RS_384 NS_384 0 9.3083309227260045e+01
GL_383 0 NS_383 NS_384 0 1.1485268189050464e-01
GL_384 0 NS_384 NS_383 0 -1.1485268189050464e-01
GS_383_4 0 NS_383 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 385/386
CS_385 NS_385 0 9.9999999999999998e-13
CS_386 NS_386 0 9.9999999999999998e-13
RS_385 NS_385 0 1.2387094149263906e+02
RS_386 NS_386 0 1.2387094149263908e+02
GL_385 0 NS_385 NS_386 0 1.0935451806229070e-01
GL_386 0 NS_386 NS_385 0 -1.0935451806229070e-01
GS_385_4 0 NS_385 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 387/388
CS_387 NS_387 0 9.9999999999999998e-13
CS_388 NS_388 0 9.9999999999999998e-13
RS_387 NS_387 0 1.1186020221520803e+02
RS_388 NS_388 0 1.1186020221520802e+02
GL_387 0 NS_387 NS_388 0 1.0538242730807947e-01
GL_388 0 NS_388 NS_387 0 -1.0538242730807947e-01
GS_387_4 0 NS_387 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 389/390
CS_389 NS_389 0 9.9999999999999998e-13
CS_390 NS_390 0 9.9999999999999998e-13
RS_389 NS_389 0 1.2031265815570148e+02
RS_390 NS_390 0 1.2031265815570150e+02
GL_389 0 NS_389 NS_390 0 9.9497602364102364e-02
GL_390 0 NS_390 NS_389 0 -9.9497602364102364e-02
GS_389_4 0 NS_389 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 391/392
CS_391 NS_391 0 9.9999999999999998e-13
CS_392 NS_392 0 9.9999999999999998e-13
RS_391 NS_391 0 9.6254518048655143e+01
RS_392 NS_392 0 9.6254518048655143e+01
GL_391 0 NS_391 NS_392 0 9.5930770757699110e-02
GL_392 0 NS_392 NS_391 0 -9.5930770757699110e-02
GS_391_4 0 NS_391 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 393/394
CS_393 NS_393 0 9.9999999999999998e-13
CS_394 NS_394 0 9.9999999999999998e-13
RS_393 NS_393 0 1.2318640771018909e+02
RS_394 NS_394 0 1.2318640771018909e+02
GL_393 0 NS_393 NS_394 0 8.9880619653662355e-02
GL_394 0 NS_394 NS_393 0 -8.9880619653662355e-02
GS_393_4 0 NS_393 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 395/396
CS_395 NS_395 0 9.9999999999999998e-13
CS_396 NS_396 0 9.9999999999999998e-13
RS_395 NS_395 0 1.1312630346155738e+02
RS_396 NS_396 0 1.1312630346155738e+02
GL_395 0 NS_395 NS_396 0 8.6534434501560398e-02
GL_396 0 NS_396 NS_395 0 -8.6534434501560398e-02
GS_395_4 0 NS_395 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 397/398
CS_397 NS_397 0 9.9999999999999998e-13
CS_398 NS_398 0 9.9999999999999998e-13
RS_397 NS_397 0 1.1831504703984019e+02
RS_398 NS_398 0 1.1831504703984019e+02
GL_397 0 NS_397 NS_398 0 7.9864296724202116e-02
GL_398 0 NS_398 NS_397 0 -7.9864296724202116e-02
GS_397_4 0 NS_397 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 399/400
CS_399 NS_399 0 9.9999999999999998e-13
CS_400 NS_400 0 9.9999999999999998e-13
RS_399 NS_399 0 1.0281987486447559e+02
RS_400 NS_400 0 1.0281987486447559e+02
GL_399 0 NS_399 NS_400 0 7.6950339194481784e-02
GL_400 0 NS_400 NS_399 0 -7.6950339194481784e-02
GS_399_4 0 NS_399 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 401/402
CS_401 NS_401 0 9.9999999999999998e-13
CS_402 NS_402 0 9.9999999999999998e-13
RS_401 NS_401 0 1.2230186914382300e+02
RS_402 NS_402 0 1.2230186914382300e+02
GL_401 0 NS_401 NS_402 0 7.0709298709435750e-02
GL_402 0 NS_402 NS_401 0 -7.0709298709435750e-02
GS_401_4 0 NS_401 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 403/404
CS_403 NS_403 0 9.9999999999999998e-13
CS_404 NS_404 0 9.9999999999999998e-13
RS_403 NS_403 0 1.2215699953322022e+02
RS_404 NS_404 0 1.2215699953322020e+02
GL_403 0 NS_403 NS_404 0 6.7518227185671367e-02
GL_404 0 NS_404 NS_403 0 -6.7518227185671367e-02
GS_403_4 0 NS_403 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 405/406
CS_405 NS_405 0 9.9999999999999998e-13
CS_406 NS_406 0 9.9999999999999998e-13
RS_405 NS_405 0 3.4305564408226764e+03
RS_406 NS_406 0 3.4305564408226769e+03
GL_405 0 NS_405 NS_406 0 5.4396471187208063e-02
GL_406 0 NS_406 NS_405 0 -5.4396471187208063e-02
GS_405_4 0 NS_405 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 407/408
CS_407 NS_407 0 9.9999999999999998e-13
CS_408 NS_408 0 9.9999999999999998e-13
RS_407 NS_407 0 1.1894859826238778e+02
RS_408 NS_408 0 1.1894859826238779e+02
GL_407 0 NS_407 NS_408 0 6.0591569497719031e-02
GL_408 0 NS_408 NS_407 0 -6.0591569497719031e-02
GS_407_4 0 NS_407 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 409/410
CS_409 NS_409 0 9.9999999999999998e-13
CS_410 NS_410 0 9.9999999999999998e-13
RS_409 NS_409 0 1.3537641711503298e+02
RS_410 NS_410 0 1.3537641711503298e+02
GL_409 0 NS_409 NS_410 0 5.1190778164089609e-02
GL_410 0 NS_410 NS_409 0 -5.1190778164089609e-02
GS_409_4 0 NS_409 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 411/412
CS_411 NS_411 0 9.9999999999999998e-13
CS_412 NS_412 0 9.9999999999999998e-13
RS_411 NS_411 0 1.3105452427659637e+02
RS_412 NS_412 0 1.3105452427659637e+02
GL_411 0 NS_411 NS_412 0 4.7418984574880592e-02
GL_412 0 NS_412 NS_411 0 -4.7418984574880592e-02
GS_411_4 0 NS_411 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 413/414
CS_413 NS_413 0 9.9999999999999998e-13
CS_414 NS_414 0 9.9999999999999998e-13
RS_413 NS_413 0 1.2170234397098790e+02
RS_414 NS_414 0 1.2170234397098790e+02
GL_413 0 NS_413 NS_414 0 4.0778813929127578e-02
GL_414 0 NS_414 NS_413 0 -4.0778813929127578e-02
GS_413_4 0 NS_413 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 415/416
CS_415 NS_415 0 9.9999999999999998e-13
CS_416 NS_416 0 9.9999999999999998e-13
RS_415 NS_415 0 1.1550510326517782e+02
RS_416 NS_416 0 1.1550510326517782e+02
GL_415 0 NS_415 NS_416 0 5.7236026076957713e-02
GL_416 0 NS_416 NS_415 0 -5.7236026076957713e-02
GS_415_4 0 NS_415 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 417/418
CS_417 NS_417 0 9.9999999999999998e-13
CS_418 NS_418 0 9.9999999999999998e-13
RS_417 NS_417 0 6.2039157456337159e+02
RS_418 NS_418 0 6.2039157456337159e+02
GL_417 0 NS_417 NS_418 0 1.9354364738401211e-02
GL_418 0 NS_418 NS_417 0 -1.9354364738401211e-02
GS_417_4 0 NS_417 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 419/420
CS_419 NS_419 0 9.9999999999999998e-13
CS_420 NS_420 0 9.9999999999999998e-13
RS_419 NS_419 0 1.1050313240441588e+02
RS_420 NS_420 0 1.1050313240441587e+02
GL_419 0 NS_419 NS_420 0 1.6472588786558075e-02
GL_420 0 NS_420 NS_419 0 -1.6472588786558075e-02
GS_419_4 0 NS_419 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 421/422
CS_421 NS_421 0 9.9999999999999998e-13
CS_422 NS_422 0 9.9999999999999998e-13
RS_421 NS_421 0 1.2869119986945731e+02
RS_422 NS_422 0 1.2869119986945731e+02
GL_421 0 NS_421 NS_422 0 2.0888592987579706e-02
GL_422 0 NS_422 NS_421 0 -2.0888592987579706e-02
GS_421_4 0 NS_421 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 423/424
CS_423 NS_423 0 9.9999999999999998e-13
CS_424 NS_424 0 9.9999999999999998e-13
RS_423 NS_423 0 1.4314560950270646e+02
RS_424 NS_424 0 1.4314560950270646e+02
GL_423 0 NS_423 NS_424 0 9.7871236580563716e-03
GL_424 0 NS_424 NS_423 0 -9.7871236580563716e-03
GS_423_4 0 NS_423 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 425/426
CS_425 NS_425 0 9.9999999999999998e-13
CS_426 NS_426 0 9.9999999999999998e-13
RS_425 NS_425 0 1.1863004336811436e+02
RS_426 NS_426 0 1.1863004336811436e+02
GL_425 0 NS_425 NS_426 0 3.7627463994326378e-02
GL_426 0 NS_426 NS_425 0 -3.7627463994326378e-02
GS_425_4 0 NS_425 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 427/428
CS_427 NS_427 0 9.9999999999999998e-13
CS_428 NS_428 0 9.9999999999999998e-13
RS_427 NS_427 0 1.2686172273444870e+02
RS_428 NS_428 0 1.2686172273444869e+02
GL_427 0 NS_427 NS_428 0 3.1975218188091938e-02
GL_428 0 NS_428 NS_427 0 -3.1975218188091938e-02
GS_427_4 0 NS_427 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 429/430
CS_429 NS_429 0 9.9999999999999998e-13
CS_430 NS_430 0 9.9999999999999998e-13
RS_429 NS_429 0 1.3141621772977734e+02
RS_430 NS_430 0 1.3141621772977737e+02
GL_429 0 NS_429 NS_430 0 2.8228381102665165e-02
GL_430 0 NS_430 NS_429 0 -2.8228381102665165e-02
GS_429_4 0 NS_429 NA_4 0 4.7428518688027549e-01
*
* Complex pair n. 431/432
CS_431 NS_431 0 9.9999999999999998e-13
CS_432 NS_432 0 9.9999999999999998e-13
RS_431 NS_431 0 1.2452833644614726e+02
RS_432 NS_432 0 1.2452833644614726e+02
GL_431 0 NS_431 NS_432 0 2.1457325426059259e-03
GL_432 0 NS_432 NS_431 0 -2.1457325426059259e-03
GS_431_4 0 NS_431 NA_4 0 4.7428518688027549e-01
*
* Real pole n. 433
CS_433 NS_433 0 9.9999999999999998e-13
RS_433 NS_433 0 3.8329546824379270e+00
GS_433_5 0 NS_433 NA_5 0 4.7428518688027549e-01
*
* Real pole n. 434
CS_434 NS_434 0 9.9999999999999998e-13
RS_434 NS_434 0 1.0843846705160875e+04
GS_434_5 0 NS_434 NA_5 0 4.7428518688027549e-01
*
* Real pole n. 435
CS_435 NS_435 0 9.9999999999999998e-13
RS_435 NS_435 0 3.3457029134706481e+03
GS_435_5 0 NS_435 NA_5 0 4.7428518688027549e-01
*
* Real pole n. 436
CS_436 NS_436 0 9.9999999999999998e-13
RS_436 NS_436 0 5.4313394337993634e+02
GS_436_5 0 NS_436 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 437/438
CS_437 NS_437 0 9.9999999999999998e-13
CS_438 NS_438 0 9.9999999999999998e-13
RS_437 NS_437 0 2.0342898045173075e+02
RS_438 NS_438 0 2.0342898045173075e+02
GL_437 0 NS_437 NS_438 0 2.5883098202682536e-01
GL_438 0 NS_438 NS_437 0 -2.5883098202682536e-01
GS_437_5 0 NS_437 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 439/440
CS_439 NS_439 0 9.9999999999999998e-13
CS_440 NS_440 0 9.9999999999999998e-13
RS_439 NS_439 0 1.2739936959261519e+02
RS_440 NS_440 0 1.2739936959261519e+02
GL_439 0 NS_439 NS_440 0 2.5122204303896745e-01
GL_440 0 NS_440 NS_439 0 -2.5122204303896745e-01
GS_439_5 0 NS_439 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 441/442
CS_441 NS_441 0 9.9999999999999998e-13
CS_442 NS_442 0 9.9999999999999998e-13
RS_441 NS_441 0 1.1105129555360161e+02
RS_442 NS_442 0 1.1105129555360161e+02
GL_441 0 NS_441 NS_442 0 2.4643422119526687e-01
GL_442 0 NS_442 NS_441 0 -2.4643422119526687e-01
GS_441_5 0 NS_441 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 443/444
CS_443 NS_443 0 9.9999999999999998e-13
CS_444 NS_444 0 9.9999999999999998e-13
RS_443 NS_443 0 1.0856580972218713e+02
RS_444 NS_444 0 1.0856580972218713e+02
GL_443 0 NS_443 NS_444 0 2.4007148694878275e-01
GL_444 0 NS_444 NS_443 0 -2.4007148694878275e-01
GS_443_5 0 NS_443 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 445/446
CS_445 NS_445 0 9.9999999999999998e-13
CS_446 NS_446 0 9.9999999999999998e-13
RS_445 NS_445 0 1.0135860176893434e+02
RS_446 NS_446 0 1.0135860176893435e+02
GL_445 0 NS_445 NS_446 0 2.3570758371916220e-01
GL_446 0 NS_446 NS_445 0 -2.3570758371916220e-01
GS_445_5 0 NS_445 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 447/448
CS_447 NS_447 0 9.9999999999999998e-13
CS_448 NS_448 0 9.9999999999999998e-13
RS_447 NS_447 0 1.2858526276753685e+02
RS_448 NS_448 0 1.2858526276753685e+02
GL_447 0 NS_447 NS_448 0 2.2966634995600790e-01
GL_448 0 NS_448 NS_447 0 -2.2966634995600790e-01
GS_447_5 0 NS_447 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 449/450
CS_449 NS_449 0 9.9999999999999998e-13
CS_450 NS_450 0 9.9999999999999998e-13
RS_449 NS_449 0 1.1773437593549667e+02
RS_450 NS_450 0 1.1773437593549667e+02
GL_449 0 NS_449 NS_450 0 2.2732609444056490e-01
GL_450 0 NS_450 NS_449 0 -2.2732609444056490e-01
GS_449_5 0 NS_449 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 451/452
CS_451 NS_451 0 9.9999999999999998e-13
CS_452 NS_452 0 9.9999999999999998e-13
RS_451 NS_451 0 9.8170265044265946e+01
RS_452 NS_452 0 9.8170265044265932e+01
GL_451 0 NS_451 NS_452 0 2.2031598117475365e-01
GL_452 0 NS_452 NS_451 0 -2.2031598117475365e-01
GS_451_5 0 NS_451 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 453/454
CS_453 NS_453 0 9.9999999999999998e-13
CS_454 NS_454 0 9.9999999999999998e-13
RS_453 NS_453 0 9.5355901421613709e+01
RS_454 NS_454 0 9.5355901421613694e+01
GL_453 0 NS_453 NS_454 0 2.1739680820836188e-01
GL_454 0 NS_454 NS_453 0 -2.1739680820836188e-01
GS_453_5 0 NS_453 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 455/456
CS_455 NS_455 0 9.9999999999999998e-13
CS_456 NS_456 0 9.9999999999999998e-13
RS_455 NS_455 0 1.0859722031634941e+02
RS_456 NS_456 0 1.0859722031634941e+02
GL_455 0 NS_455 NS_456 0 2.0887403840929383e-01
GL_456 0 NS_456 NS_455 0 -2.0887403840929383e-01
GS_455_5 0 NS_455 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 457/458
CS_457 NS_457 0 9.9999999999999998e-13
CS_458 NS_458 0 9.9999999999999998e-13
RS_457 NS_457 0 7.7959989808728068e+01
RS_458 NS_458 0 7.7959989808728054e+01
GL_457 0 NS_457 NS_458 0 2.0447808896343445e-01
GL_458 0 NS_458 NS_457 0 -2.0447808896343445e-01
GS_457_5 0 NS_457 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 459/460
CS_459 NS_459 0 9.9999999999999998e-13
CS_460 NS_460 0 9.9999999999999998e-13
RS_459 NS_459 0 1.1088851678406323e+02
RS_460 NS_460 0 1.1088851678406321e+02
GL_459 0 NS_459 NS_460 0 1.9843399276071924e-01
GL_460 0 NS_460 NS_459 0 -1.9843399276071924e-01
GS_459_5 0 NS_459 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 461/462
CS_461 NS_461 0 9.9999999999999998e-13
CS_462 NS_462 0 9.9999999999999998e-13
RS_461 NS_461 0 8.1179760966262847e+01
RS_462 NS_462 0 8.1179760966262847e+01
GL_461 0 NS_461 NS_462 0 1.8978022990658949e-01
GL_462 0 NS_462 NS_461 0 -1.8978022990658949e-01
GS_461_5 0 NS_461 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 463/464
CS_463 NS_463 0 9.9999999999999998e-13
CS_464 NS_464 0 9.9999999999999998e-13
RS_463 NS_463 0 1.0523970815054612e+02
RS_464 NS_464 0 1.0523970815054612e+02
GL_463 0 NS_463 NS_464 0 1.8836779078363333e-01
GL_464 0 NS_464 NS_463 0 -1.8836779078363333e-01
GS_463_5 0 NS_463 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 465/466
CS_465 NS_465 0 9.9999999999999998e-13
CS_466 NS_466 0 9.9999999999999998e-13
RS_465 NS_465 0 1.1208834663822537e+02
RS_466 NS_466 0 1.1208834663822537e+02
GL_465 0 NS_465 NS_466 0 1.7925451755127267e-01
GL_466 0 NS_466 NS_465 0 -1.7925451755127267e-01
GS_465_5 0 NS_465 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 467/468
CS_467 NS_467 0 9.9999999999999998e-13
CS_468 NS_468 0 9.9999999999999998e-13
RS_467 NS_467 0 9.2475617668062213e+01
RS_468 NS_468 0 9.2475617668062199e+01
GL_467 0 NS_467 NS_468 0 1.7507216970358189e-01
GL_468 0 NS_468 NS_467 0 -1.7507216970358189e-01
GS_467_5 0 NS_467 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 469/470
CS_469 NS_469 0 9.9999999999999998e-13
CS_470 NS_470 0 9.9999999999999998e-13
RS_469 NS_469 0 1.1555782965375326e+02
RS_470 NS_470 0 1.1555782965375326e+02
GL_469 0 NS_469 NS_470 0 1.6918904340923188e-01
GL_470 0 NS_470 NS_469 0 -1.6918904340923188e-01
GS_469_5 0 NS_469 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 471/472
CS_471 NS_471 0 9.9999999999999998e-13
CS_472 NS_472 0 9.9999999999999998e-13
RS_471 NS_471 0 9.6856782813111039e+01
RS_472 NS_472 0 9.6856782813111039e+01
GL_471 0 NS_471 NS_472 0 1.6488898173469207e-01
GL_472 0 NS_472 NS_471 0 -1.6488898173469207e-01
GS_471_5 0 NS_471 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 473/474
CS_473 NS_473 0 9.9999999999999998e-13
CS_474 NS_474 0 9.9999999999999998e-13
RS_473 NS_473 0 1.1717534841017003e+02
RS_474 NS_474 0 1.1717534841017003e+02
GL_473 0 NS_473 NS_474 0 1.5866517390841936e-01
GL_474 0 NS_474 NS_473 0 -1.5866517390841936e-01
GS_473_5 0 NS_473 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 475/476
CS_475 NS_475 0 9.9999999999999998e-13
CS_476 NS_476 0 9.9999999999999998e-13
RS_475 NS_475 0 8.8607873746940697e+01
RS_476 NS_476 0 8.8607873746940697e+01
GL_475 0 NS_475 NS_476 0 1.5214737618207635e-01
GL_476 0 NS_476 NS_475 0 -1.5214737618207635e-01
GS_475_5 0 NS_475 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 477/478
CS_477 NS_477 0 9.9999999999999998e-13
CS_478 NS_478 0 9.9999999999999998e-13
RS_477 NS_477 0 1.1741456484283673e+02
RS_478 NS_478 0 1.1741456484283673e+02
GL_477 0 NS_477 NS_478 0 1.4829748860889613e-01
GL_478 0 NS_478 NS_477 0 -1.4829748860889613e-01
GS_477_5 0 NS_477 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 479/480
CS_479 NS_479 0 9.9999999999999998e-13
CS_480 NS_480 0 9.9999999999999998e-13
RS_479 NS_479 0 1.3292289814180702e+02
RS_480 NS_480 0 1.3292289814180702e+02
GL_479 0 NS_479 NS_480 0 1.4243056778188259e-01
GL_480 0 NS_480 NS_479 0 -1.4243056778188259e-01
GS_479_5 0 NS_479 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 481/482
CS_481 NS_481 0 9.9999999999999998e-13
CS_482 NS_482 0 9.9999999999999998e-13
RS_481 NS_481 0 1.2325134819531741e+02
RS_482 NS_482 0 1.2325134819531739e+02
GL_481 0 NS_481 NS_482 0 1.3890785074828846e-01
GL_482 0 NS_482 NS_481 0 -1.3890785074828846e-01
GS_481_5 0 NS_481 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 483/484
CS_483 NS_483 0 9.9999999999999998e-13
CS_484 NS_484 0 9.9999999999999998e-13
RS_483 NS_483 0 9.1909059882883227e+01
RS_484 NS_484 0 9.1909059882883227e+01
GL_483 0 NS_483 NS_484 0 1.3373879533989103e-01
GL_484 0 NS_484 NS_483 0 -1.3373879533989103e-01
GS_483_5 0 NS_483 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 485/486
CS_485 NS_485 0 9.9999999999999998e-13
CS_486 NS_486 0 9.9999999999999998e-13
RS_485 NS_485 0 1.2276824880349510e+02
RS_486 NS_486 0 1.2276824880349510e+02
GL_485 0 NS_485 NS_486 0 1.2885409674522977e-01
GL_486 0 NS_486 NS_485 0 -1.2885409674522977e-01
GS_485_5 0 NS_485 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 487/488
CS_487 NS_487 0 9.9999999999999998e-13
CS_488 NS_488 0 9.9999999999999998e-13
RS_487 NS_487 0 1.1612442076026501e+02
RS_488 NS_488 0 1.1612442076026501e+02
GL_487 0 NS_487 NS_488 0 1.2417838026896348e-01
GL_488 0 NS_488 NS_487 0 -1.2417838026896348e-01
GS_487_5 0 NS_487 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 489/490
CS_489 NS_489 0 9.9999999999999998e-13
CS_490 NS_490 0 9.9999999999999998e-13
RS_489 NS_489 0 1.2130204223875414e+02
RS_490 NS_490 0 1.2130204223875414e+02
GL_489 0 NS_489 NS_490 0 1.1919240021970828e-01
GL_490 0 NS_490 NS_489 0 -1.1919240021970828e-01
GS_489_5 0 NS_489 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 491/492
CS_491 NS_491 0 9.9999999999999998e-13
CS_492 NS_492 0 9.9999999999999998e-13
RS_491 NS_491 0 9.3083309227260045e+01
RS_492 NS_492 0 9.3083309227260045e+01
GL_491 0 NS_491 NS_492 0 1.1485268189050464e-01
GL_492 0 NS_492 NS_491 0 -1.1485268189050464e-01
GS_491_5 0 NS_491 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 493/494
CS_493 NS_493 0 9.9999999999999998e-13
CS_494 NS_494 0 9.9999999999999998e-13
RS_493 NS_493 0 1.2387094149263906e+02
RS_494 NS_494 0 1.2387094149263908e+02
GL_493 0 NS_493 NS_494 0 1.0935451806229070e-01
GL_494 0 NS_494 NS_493 0 -1.0935451806229070e-01
GS_493_5 0 NS_493 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 495/496
CS_495 NS_495 0 9.9999999999999998e-13
CS_496 NS_496 0 9.9999999999999998e-13
RS_495 NS_495 0 1.1186020221520803e+02
RS_496 NS_496 0 1.1186020221520802e+02
GL_495 0 NS_495 NS_496 0 1.0538242730807947e-01
GL_496 0 NS_496 NS_495 0 -1.0538242730807947e-01
GS_495_5 0 NS_495 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 497/498
CS_497 NS_497 0 9.9999999999999998e-13
CS_498 NS_498 0 9.9999999999999998e-13
RS_497 NS_497 0 1.2031265815570148e+02
RS_498 NS_498 0 1.2031265815570150e+02
GL_497 0 NS_497 NS_498 0 9.9497602364102364e-02
GL_498 0 NS_498 NS_497 0 -9.9497602364102364e-02
GS_497_5 0 NS_497 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 499/500
CS_499 NS_499 0 9.9999999999999998e-13
CS_500 NS_500 0 9.9999999999999998e-13
RS_499 NS_499 0 9.6254518048655143e+01
RS_500 NS_500 0 9.6254518048655143e+01
GL_499 0 NS_499 NS_500 0 9.5930770757699110e-02
GL_500 0 NS_500 NS_499 0 -9.5930770757699110e-02
GS_499_5 0 NS_499 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 501/502
CS_501 NS_501 0 9.9999999999999998e-13
CS_502 NS_502 0 9.9999999999999998e-13
RS_501 NS_501 0 1.2318640771018909e+02
RS_502 NS_502 0 1.2318640771018909e+02
GL_501 0 NS_501 NS_502 0 8.9880619653662355e-02
GL_502 0 NS_502 NS_501 0 -8.9880619653662355e-02
GS_501_5 0 NS_501 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 503/504
CS_503 NS_503 0 9.9999999999999998e-13
CS_504 NS_504 0 9.9999999999999998e-13
RS_503 NS_503 0 1.1312630346155738e+02
RS_504 NS_504 0 1.1312630346155738e+02
GL_503 0 NS_503 NS_504 0 8.6534434501560398e-02
GL_504 0 NS_504 NS_503 0 -8.6534434501560398e-02
GS_503_5 0 NS_503 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 505/506
CS_505 NS_505 0 9.9999999999999998e-13
CS_506 NS_506 0 9.9999999999999998e-13
RS_505 NS_505 0 1.1831504703984019e+02
RS_506 NS_506 0 1.1831504703984019e+02
GL_505 0 NS_505 NS_506 0 7.9864296724202116e-02
GL_506 0 NS_506 NS_505 0 -7.9864296724202116e-02
GS_505_5 0 NS_505 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 507/508
CS_507 NS_507 0 9.9999999999999998e-13
CS_508 NS_508 0 9.9999999999999998e-13
RS_507 NS_507 0 1.0281987486447559e+02
RS_508 NS_508 0 1.0281987486447559e+02
GL_507 0 NS_507 NS_508 0 7.6950339194481784e-02
GL_508 0 NS_508 NS_507 0 -7.6950339194481784e-02
GS_507_5 0 NS_507 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 509/510
CS_509 NS_509 0 9.9999999999999998e-13
CS_510 NS_510 0 9.9999999999999998e-13
RS_509 NS_509 0 1.2230186914382300e+02
RS_510 NS_510 0 1.2230186914382300e+02
GL_509 0 NS_509 NS_510 0 7.0709298709435750e-02
GL_510 0 NS_510 NS_509 0 -7.0709298709435750e-02
GS_509_5 0 NS_509 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 511/512
CS_511 NS_511 0 9.9999999999999998e-13
CS_512 NS_512 0 9.9999999999999998e-13
RS_511 NS_511 0 1.2215699953322022e+02
RS_512 NS_512 0 1.2215699953322020e+02
GL_511 0 NS_511 NS_512 0 6.7518227185671367e-02
GL_512 0 NS_512 NS_511 0 -6.7518227185671367e-02
GS_511_5 0 NS_511 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 513/514
CS_513 NS_513 0 9.9999999999999998e-13
CS_514 NS_514 0 9.9999999999999998e-13
RS_513 NS_513 0 3.4305564408226764e+03
RS_514 NS_514 0 3.4305564408226769e+03
GL_513 0 NS_513 NS_514 0 5.4396471187208063e-02
GL_514 0 NS_514 NS_513 0 -5.4396471187208063e-02
GS_513_5 0 NS_513 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 515/516
CS_515 NS_515 0 9.9999999999999998e-13
CS_516 NS_516 0 9.9999999999999998e-13
RS_515 NS_515 0 1.1894859826238778e+02
RS_516 NS_516 0 1.1894859826238779e+02
GL_515 0 NS_515 NS_516 0 6.0591569497719031e-02
GL_516 0 NS_516 NS_515 0 -6.0591569497719031e-02
GS_515_5 0 NS_515 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 517/518
CS_517 NS_517 0 9.9999999999999998e-13
CS_518 NS_518 0 9.9999999999999998e-13
RS_517 NS_517 0 1.3537641711503298e+02
RS_518 NS_518 0 1.3537641711503298e+02
GL_517 0 NS_517 NS_518 0 5.1190778164089609e-02
GL_518 0 NS_518 NS_517 0 -5.1190778164089609e-02
GS_517_5 0 NS_517 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 519/520
CS_519 NS_519 0 9.9999999999999998e-13
CS_520 NS_520 0 9.9999999999999998e-13
RS_519 NS_519 0 1.3105452427659637e+02
RS_520 NS_520 0 1.3105452427659637e+02
GL_519 0 NS_519 NS_520 0 4.7418984574880592e-02
GL_520 0 NS_520 NS_519 0 -4.7418984574880592e-02
GS_519_5 0 NS_519 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 521/522
CS_521 NS_521 0 9.9999999999999998e-13
CS_522 NS_522 0 9.9999999999999998e-13
RS_521 NS_521 0 1.2170234397098790e+02
RS_522 NS_522 0 1.2170234397098790e+02
GL_521 0 NS_521 NS_522 0 4.0778813929127578e-02
GL_522 0 NS_522 NS_521 0 -4.0778813929127578e-02
GS_521_5 0 NS_521 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 523/524
CS_523 NS_523 0 9.9999999999999998e-13
CS_524 NS_524 0 9.9999999999999998e-13
RS_523 NS_523 0 1.1550510326517782e+02
RS_524 NS_524 0 1.1550510326517782e+02
GL_523 0 NS_523 NS_524 0 5.7236026076957713e-02
GL_524 0 NS_524 NS_523 0 -5.7236026076957713e-02
GS_523_5 0 NS_523 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 525/526
CS_525 NS_525 0 9.9999999999999998e-13
CS_526 NS_526 0 9.9999999999999998e-13
RS_525 NS_525 0 6.2039157456337159e+02
RS_526 NS_526 0 6.2039157456337159e+02
GL_525 0 NS_525 NS_526 0 1.9354364738401211e-02
GL_526 0 NS_526 NS_525 0 -1.9354364738401211e-02
GS_525_5 0 NS_525 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 527/528
CS_527 NS_527 0 9.9999999999999998e-13
CS_528 NS_528 0 9.9999999999999998e-13
RS_527 NS_527 0 1.1050313240441588e+02
RS_528 NS_528 0 1.1050313240441587e+02
GL_527 0 NS_527 NS_528 0 1.6472588786558075e-02
GL_528 0 NS_528 NS_527 0 -1.6472588786558075e-02
GS_527_5 0 NS_527 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 529/530
CS_529 NS_529 0 9.9999999999999998e-13
CS_530 NS_530 0 9.9999999999999998e-13
RS_529 NS_529 0 1.2869119986945731e+02
RS_530 NS_530 0 1.2869119986945731e+02
GL_529 0 NS_529 NS_530 0 2.0888592987579706e-02
GL_530 0 NS_530 NS_529 0 -2.0888592987579706e-02
GS_529_5 0 NS_529 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 531/532
CS_531 NS_531 0 9.9999999999999998e-13
CS_532 NS_532 0 9.9999999999999998e-13
RS_531 NS_531 0 1.4314560950270646e+02
RS_532 NS_532 0 1.4314560950270646e+02
GL_531 0 NS_531 NS_532 0 9.7871236580563716e-03
GL_532 0 NS_532 NS_531 0 -9.7871236580563716e-03
GS_531_5 0 NS_531 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 533/534
CS_533 NS_533 0 9.9999999999999998e-13
CS_534 NS_534 0 9.9999999999999998e-13
RS_533 NS_533 0 1.1863004336811436e+02
RS_534 NS_534 0 1.1863004336811436e+02
GL_533 0 NS_533 NS_534 0 3.7627463994326378e-02
GL_534 0 NS_534 NS_533 0 -3.7627463994326378e-02
GS_533_5 0 NS_533 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 535/536
CS_535 NS_535 0 9.9999999999999998e-13
CS_536 NS_536 0 9.9999999999999998e-13
RS_535 NS_535 0 1.2686172273444870e+02
RS_536 NS_536 0 1.2686172273444869e+02
GL_535 0 NS_535 NS_536 0 3.1975218188091938e-02
GL_536 0 NS_536 NS_535 0 -3.1975218188091938e-02
GS_535_5 0 NS_535 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 537/538
CS_537 NS_537 0 9.9999999999999998e-13
CS_538 NS_538 0 9.9999999999999998e-13
RS_537 NS_537 0 1.3141621772977734e+02
RS_538 NS_538 0 1.3141621772977737e+02
GL_537 0 NS_537 NS_538 0 2.8228381102665165e-02
GL_538 0 NS_538 NS_537 0 -2.8228381102665165e-02
GS_537_5 0 NS_537 NA_5 0 4.7428518688027549e-01
*
* Complex pair n. 539/540
CS_539 NS_539 0 9.9999999999999998e-13
CS_540 NS_540 0 9.9999999999999998e-13
RS_539 NS_539 0 1.2452833644614726e+02
RS_540 NS_540 0 1.2452833644614726e+02
GL_539 0 NS_539 NS_540 0 2.1457325426059259e-03
GL_540 0 NS_540 NS_539 0 -2.1457325426059259e-03
GS_539_5 0 NS_539 NA_5 0 4.7428518688027549e-01
*
* Real pole n. 541
CS_541 NS_541 0 9.9999999999999998e-13
RS_541 NS_541 0 3.8329546824379270e+00
GS_541_6 0 NS_541 NA_6 0 4.7428518688027549e-01
*
* Real pole n. 542
CS_542 NS_542 0 9.9999999999999998e-13
RS_542 NS_542 0 1.0843846705160875e+04
GS_542_6 0 NS_542 NA_6 0 4.7428518688027549e-01
*
* Real pole n. 543
CS_543 NS_543 0 9.9999999999999998e-13
RS_543 NS_543 0 3.3457029134706481e+03
GS_543_6 0 NS_543 NA_6 0 4.7428518688027549e-01
*
* Real pole n. 544
CS_544 NS_544 0 9.9999999999999998e-13
RS_544 NS_544 0 5.4313394337993634e+02
GS_544_6 0 NS_544 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 545/546
CS_545 NS_545 0 9.9999999999999998e-13
CS_546 NS_546 0 9.9999999999999998e-13
RS_545 NS_545 0 2.0342898045173075e+02
RS_546 NS_546 0 2.0342898045173075e+02
GL_545 0 NS_545 NS_546 0 2.5883098202682536e-01
GL_546 0 NS_546 NS_545 0 -2.5883098202682536e-01
GS_545_6 0 NS_545 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 547/548
CS_547 NS_547 0 9.9999999999999998e-13
CS_548 NS_548 0 9.9999999999999998e-13
RS_547 NS_547 0 1.2739936959261519e+02
RS_548 NS_548 0 1.2739936959261519e+02
GL_547 0 NS_547 NS_548 0 2.5122204303896745e-01
GL_548 0 NS_548 NS_547 0 -2.5122204303896745e-01
GS_547_6 0 NS_547 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 549/550
CS_549 NS_549 0 9.9999999999999998e-13
CS_550 NS_550 0 9.9999999999999998e-13
RS_549 NS_549 0 1.1105129555360161e+02
RS_550 NS_550 0 1.1105129555360161e+02
GL_549 0 NS_549 NS_550 0 2.4643422119526687e-01
GL_550 0 NS_550 NS_549 0 -2.4643422119526687e-01
GS_549_6 0 NS_549 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 551/552
CS_551 NS_551 0 9.9999999999999998e-13
CS_552 NS_552 0 9.9999999999999998e-13
RS_551 NS_551 0 1.0856580972218713e+02
RS_552 NS_552 0 1.0856580972218713e+02
GL_551 0 NS_551 NS_552 0 2.4007148694878275e-01
GL_552 0 NS_552 NS_551 0 -2.4007148694878275e-01
GS_551_6 0 NS_551 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 553/554
CS_553 NS_553 0 9.9999999999999998e-13
CS_554 NS_554 0 9.9999999999999998e-13
RS_553 NS_553 0 1.0135860176893434e+02
RS_554 NS_554 0 1.0135860176893435e+02
GL_553 0 NS_553 NS_554 0 2.3570758371916220e-01
GL_554 0 NS_554 NS_553 0 -2.3570758371916220e-01
GS_553_6 0 NS_553 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 555/556
CS_555 NS_555 0 9.9999999999999998e-13
CS_556 NS_556 0 9.9999999999999998e-13
RS_555 NS_555 0 1.2858526276753685e+02
RS_556 NS_556 0 1.2858526276753685e+02
GL_555 0 NS_555 NS_556 0 2.2966634995600790e-01
GL_556 0 NS_556 NS_555 0 -2.2966634995600790e-01
GS_555_6 0 NS_555 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 557/558
CS_557 NS_557 0 9.9999999999999998e-13
CS_558 NS_558 0 9.9999999999999998e-13
RS_557 NS_557 0 1.1773437593549667e+02
RS_558 NS_558 0 1.1773437593549667e+02
GL_557 0 NS_557 NS_558 0 2.2732609444056490e-01
GL_558 0 NS_558 NS_557 0 -2.2732609444056490e-01
GS_557_6 0 NS_557 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 559/560
CS_559 NS_559 0 9.9999999999999998e-13
CS_560 NS_560 0 9.9999999999999998e-13
RS_559 NS_559 0 9.8170265044265946e+01
RS_560 NS_560 0 9.8170265044265932e+01
GL_559 0 NS_559 NS_560 0 2.2031598117475365e-01
GL_560 0 NS_560 NS_559 0 -2.2031598117475365e-01
GS_559_6 0 NS_559 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 561/562
CS_561 NS_561 0 9.9999999999999998e-13
CS_562 NS_562 0 9.9999999999999998e-13
RS_561 NS_561 0 9.5355901421613709e+01
RS_562 NS_562 0 9.5355901421613694e+01
GL_561 0 NS_561 NS_562 0 2.1739680820836188e-01
GL_562 0 NS_562 NS_561 0 -2.1739680820836188e-01
GS_561_6 0 NS_561 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 563/564
CS_563 NS_563 0 9.9999999999999998e-13
CS_564 NS_564 0 9.9999999999999998e-13
RS_563 NS_563 0 1.0859722031634941e+02
RS_564 NS_564 0 1.0859722031634941e+02
GL_563 0 NS_563 NS_564 0 2.0887403840929383e-01
GL_564 0 NS_564 NS_563 0 -2.0887403840929383e-01
GS_563_6 0 NS_563 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 565/566
CS_565 NS_565 0 9.9999999999999998e-13
CS_566 NS_566 0 9.9999999999999998e-13
RS_565 NS_565 0 7.7959989808728068e+01
RS_566 NS_566 0 7.7959989808728054e+01
GL_565 0 NS_565 NS_566 0 2.0447808896343445e-01
GL_566 0 NS_566 NS_565 0 -2.0447808896343445e-01
GS_565_6 0 NS_565 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 567/568
CS_567 NS_567 0 9.9999999999999998e-13
CS_568 NS_568 0 9.9999999999999998e-13
RS_567 NS_567 0 1.1088851678406323e+02
RS_568 NS_568 0 1.1088851678406321e+02
GL_567 0 NS_567 NS_568 0 1.9843399276071924e-01
GL_568 0 NS_568 NS_567 0 -1.9843399276071924e-01
GS_567_6 0 NS_567 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 569/570
CS_569 NS_569 0 9.9999999999999998e-13
CS_570 NS_570 0 9.9999999999999998e-13
RS_569 NS_569 0 8.1179760966262847e+01
RS_570 NS_570 0 8.1179760966262847e+01
GL_569 0 NS_569 NS_570 0 1.8978022990658949e-01
GL_570 0 NS_570 NS_569 0 -1.8978022990658949e-01
GS_569_6 0 NS_569 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 571/572
CS_571 NS_571 0 9.9999999999999998e-13
CS_572 NS_572 0 9.9999999999999998e-13
RS_571 NS_571 0 1.0523970815054612e+02
RS_572 NS_572 0 1.0523970815054612e+02
GL_571 0 NS_571 NS_572 0 1.8836779078363333e-01
GL_572 0 NS_572 NS_571 0 -1.8836779078363333e-01
GS_571_6 0 NS_571 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 573/574
CS_573 NS_573 0 9.9999999999999998e-13
CS_574 NS_574 0 9.9999999999999998e-13
RS_573 NS_573 0 1.1208834663822537e+02
RS_574 NS_574 0 1.1208834663822537e+02
GL_573 0 NS_573 NS_574 0 1.7925451755127267e-01
GL_574 0 NS_574 NS_573 0 -1.7925451755127267e-01
GS_573_6 0 NS_573 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 575/576
CS_575 NS_575 0 9.9999999999999998e-13
CS_576 NS_576 0 9.9999999999999998e-13
RS_575 NS_575 0 9.2475617668062213e+01
RS_576 NS_576 0 9.2475617668062199e+01
GL_575 0 NS_575 NS_576 0 1.7507216970358189e-01
GL_576 0 NS_576 NS_575 0 -1.7507216970358189e-01
GS_575_6 0 NS_575 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 577/578
CS_577 NS_577 0 9.9999999999999998e-13
CS_578 NS_578 0 9.9999999999999998e-13
RS_577 NS_577 0 1.1555782965375326e+02
RS_578 NS_578 0 1.1555782965375326e+02
GL_577 0 NS_577 NS_578 0 1.6918904340923188e-01
GL_578 0 NS_578 NS_577 0 -1.6918904340923188e-01
GS_577_6 0 NS_577 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 579/580
CS_579 NS_579 0 9.9999999999999998e-13
CS_580 NS_580 0 9.9999999999999998e-13
RS_579 NS_579 0 9.6856782813111039e+01
RS_580 NS_580 0 9.6856782813111039e+01
GL_579 0 NS_579 NS_580 0 1.6488898173469207e-01
GL_580 0 NS_580 NS_579 0 -1.6488898173469207e-01
GS_579_6 0 NS_579 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 581/582
CS_581 NS_581 0 9.9999999999999998e-13
CS_582 NS_582 0 9.9999999999999998e-13
RS_581 NS_581 0 1.1717534841017003e+02
RS_582 NS_582 0 1.1717534841017003e+02
GL_581 0 NS_581 NS_582 0 1.5866517390841936e-01
GL_582 0 NS_582 NS_581 0 -1.5866517390841936e-01
GS_581_6 0 NS_581 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 583/584
CS_583 NS_583 0 9.9999999999999998e-13
CS_584 NS_584 0 9.9999999999999998e-13
RS_583 NS_583 0 8.8607873746940697e+01
RS_584 NS_584 0 8.8607873746940697e+01
GL_583 0 NS_583 NS_584 0 1.5214737618207635e-01
GL_584 0 NS_584 NS_583 0 -1.5214737618207635e-01
GS_583_6 0 NS_583 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 585/586
CS_585 NS_585 0 9.9999999999999998e-13
CS_586 NS_586 0 9.9999999999999998e-13
RS_585 NS_585 0 1.1741456484283673e+02
RS_586 NS_586 0 1.1741456484283673e+02
GL_585 0 NS_585 NS_586 0 1.4829748860889613e-01
GL_586 0 NS_586 NS_585 0 -1.4829748860889613e-01
GS_585_6 0 NS_585 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 587/588
CS_587 NS_587 0 9.9999999999999998e-13
CS_588 NS_588 0 9.9999999999999998e-13
RS_587 NS_587 0 1.3292289814180702e+02
RS_588 NS_588 0 1.3292289814180702e+02
GL_587 0 NS_587 NS_588 0 1.4243056778188259e-01
GL_588 0 NS_588 NS_587 0 -1.4243056778188259e-01
GS_587_6 0 NS_587 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 589/590
CS_589 NS_589 0 9.9999999999999998e-13
CS_590 NS_590 0 9.9999999999999998e-13
RS_589 NS_589 0 1.2325134819531741e+02
RS_590 NS_590 0 1.2325134819531739e+02
GL_589 0 NS_589 NS_590 0 1.3890785074828846e-01
GL_590 0 NS_590 NS_589 0 -1.3890785074828846e-01
GS_589_6 0 NS_589 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 591/592
CS_591 NS_591 0 9.9999999999999998e-13
CS_592 NS_592 0 9.9999999999999998e-13
RS_591 NS_591 0 9.1909059882883227e+01
RS_592 NS_592 0 9.1909059882883227e+01
GL_591 0 NS_591 NS_592 0 1.3373879533989103e-01
GL_592 0 NS_592 NS_591 0 -1.3373879533989103e-01
GS_591_6 0 NS_591 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 593/594
CS_593 NS_593 0 9.9999999999999998e-13
CS_594 NS_594 0 9.9999999999999998e-13
RS_593 NS_593 0 1.2276824880349510e+02
RS_594 NS_594 0 1.2276824880349510e+02
GL_593 0 NS_593 NS_594 0 1.2885409674522977e-01
GL_594 0 NS_594 NS_593 0 -1.2885409674522977e-01
GS_593_6 0 NS_593 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 595/596
CS_595 NS_595 0 9.9999999999999998e-13
CS_596 NS_596 0 9.9999999999999998e-13
RS_595 NS_595 0 1.1612442076026501e+02
RS_596 NS_596 0 1.1612442076026501e+02
GL_595 0 NS_595 NS_596 0 1.2417838026896348e-01
GL_596 0 NS_596 NS_595 0 -1.2417838026896348e-01
GS_595_6 0 NS_595 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 597/598
CS_597 NS_597 0 9.9999999999999998e-13
CS_598 NS_598 0 9.9999999999999998e-13
RS_597 NS_597 0 1.2130204223875414e+02
RS_598 NS_598 0 1.2130204223875414e+02
GL_597 0 NS_597 NS_598 0 1.1919240021970828e-01
GL_598 0 NS_598 NS_597 0 -1.1919240021970828e-01
GS_597_6 0 NS_597 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 599/600
CS_599 NS_599 0 9.9999999999999998e-13
CS_600 NS_600 0 9.9999999999999998e-13
RS_599 NS_599 0 9.3083309227260045e+01
RS_600 NS_600 0 9.3083309227260045e+01
GL_599 0 NS_599 NS_600 0 1.1485268189050464e-01
GL_600 0 NS_600 NS_599 0 -1.1485268189050464e-01
GS_599_6 0 NS_599 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 601/602
CS_601 NS_601 0 9.9999999999999998e-13
CS_602 NS_602 0 9.9999999999999998e-13
RS_601 NS_601 0 1.2387094149263906e+02
RS_602 NS_602 0 1.2387094149263908e+02
GL_601 0 NS_601 NS_602 0 1.0935451806229070e-01
GL_602 0 NS_602 NS_601 0 -1.0935451806229070e-01
GS_601_6 0 NS_601 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 603/604
CS_603 NS_603 0 9.9999999999999998e-13
CS_604 NS_604 0 9.9999999999999998e-13
RS_603 NS_603 0 1.1186020221520803e+02
RS_604 NS_604 0 1.1186020221520802e+02
GL_603 0 NS_603 NS_604 0 1.0538242730807947e-01
GL_604 0 NS_604 NS_603 0 -1.0538242730807947e-01
GS_603_6 0 NS_603 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 605/606
CS_605 NS_605 0 9.9999999999999998e-13
CS_606 NS_606 0 9.9999999999999998e-13
RS_605 NS_605 0 1.2031265815570148e+02
RS_606 NS_606 0 1.2031265815570150e+02
GL_605 0 NS_605 NS_606 0 9.9497602364102364e-02
GL_606 0 NS_606 NS_605 0 -9.9497602364102364e-02
GS_605_6 0 NS_605 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 607/608
CS_607 NS_607 0 9.9999999999999998e-13
CS_608 NS_608 0 9.9999999999999998e-13
RS_607 NS_607 0 9.6254518048655143e+01
RS_608 NS_608 0 9.6254518048655143e+01
GL_607 0 NS_607 NS_608 0 9.5930770757699110e-02
GL_608 0 NS_608 NS_607 0 -9.5930770757699110e-02
GS_607_6 0 NS_607 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 609/610
CS_609 NS_609 0 9.9999999999999998e-13
CS_610 NS_610 0 9.9999999999999998e-13
RS_609 NS_609 0 1.2318640771018909e+02
RS_610 NS_610 0 1.2318640771018909e+02
GL_609 0 NS_609 NS_610 0 8.9880619653662355e-02
GL_610 0 NS_610 NS_609 0 -8.9880619653662355e-02
GS_609_6 0 NS_609 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 611/612
CS_611 NS_611 0 9.9999999999999998e-13
CS_612 NS_612 0 9.9999999999999998e-13
RS_611 NS_611 0 1.1312630346155738e+02
RS_612 NS_612 0 1.1312630346155738e+02
GL_611 0 NS_611 NS_612 0 8.6534434501560398e-02
GL_612 0 NS_612 NS_611 0 -8.6534434501560398e-02
GS_611_6 0 NS_611 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 613/614
CS_613 NS_613 0 9.9999999999999998e-13
CS_614 NS_614 0 9.9999999999999998e-13
RS_613 NS_613 0 1.1831504703984019e+02
RS_614 NS_614 0 1.1831504703984019e+02
GL_613 0 NS_613 NS_614 0 7.9864296724202116e-02
GL_614 0 NS_614 NS_613 0 -7.9864296724202116e-02
GS_613_6 0 NS_613 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 615/616
CS_615 NS_615 0 9.9999999999999998e-13
CS_616 NS_616 0 9.9999999999999998e-13
RS_615 NS_615 0 1.0281987486447559e+02
RS_616 NS_616 0 1.0281987486447559e+02
GL_615 0 NS_615 NS_616 0 7.6950339194481784e-02
GL_616 0 NS_616 NS_615 0 -7.6950339194481784e-02
GS_615_6 0 NS_615 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 617/618
CS_617 NS_617 0 9.9999999999999998e-13
CS_618 NS_618 0 9.9999999999999998e-13
RS_617 NS_617 0 1.2230186914382300e+02
RS_618 NS_618 0 1.2230186914382300e+02
GL_617 0 NS_617 NS_618 0 7.0709298709435750e-02
GL_618 0 NS_618 NS_617 0 -7.0709298709435750e-02
GS_617_6 0 NS_617 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 619/620
CS_619 NS_619 0 9.9999999999999998e-13
CS_620 NS_620 0 9.9999999999999998e-13
RS_619 NS_619 0 1.2215699953322022e+02
RS_620 NS_620 0 1.2215699953322020e+02
GL_619 0 NS_619 NS_620 0 6.7518227185671367e-02
GL_620 0 NS_620 NS_619 0 -6.7518227185671367e-02
GS_619_6 0 NS_619 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 621/622
CS_621 NS_621 0 9.9999999999999998e-13
CS_622 NS_622 0 9.9999999999999998e-13
RS_621 NS_621 0 3.4305564408226764e+03
RS_622 NS_622 0 3.4305564408226769e+03
GL_621 0 NS_621 NS_622 0 5.4396471187208063e-02
GL_622 0 NS_622 NS_621 0 -5.4396471187208063e-02
GS_621_6 0 NS_621 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 623/624
CS_623 NS_623 0 9.9999999999999998e-13
CS_624 NS_624 0 9.9999999999999998e-13
RS_623 NS_623 0 1.1894859826238778e+02
RS_624 NS_624 0 1.1894859826238779e+02
GL_623 0 NS_623 NS_624 0 6.0591569497719031e-02
GL_624 0 NS_624 NS_623 0 -6.0591569497719031e-02
GS_623_6 0 NS_623 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 625/626
CS_625 NS_625 0 9.9999999999999998e-13
CS_626 NS_626 0 9.9999999999999998e-13
RS_625 NS_625 0 1.3537641711503298e+02
RS_626 NS_626 0 1.3537641711503298e+02
GL_625 0 NS_625 NS_626 0 5.1190778164089609e-02
GL_626 0 NS_626 NS_625 0 -5.1190778164089609e-02
GS_625_6 0 NS_625 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 627/628
CS_627 NS_627 0 9.9999999999999998e-13
CS_628 NS_628 0 9.9999999999999998e-13
RS_627 NS_627 0 1.3105452427659637e+02
RS_628 NS_628 0 1.3105452427659637e+02
GL_627 0 NS_627 NS_628 0 4.7418984574880592e-02
GL_628 0 NS_628 NS_627 0 -4.7418984574880592e-02
GS_627_6 0 NS_627 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 629/630
CS_629 NS_629 0 9.9999999999999998e-13
CS_630 NS_630 0 9.9999999999999998e-13
RS_629 NS_629 0 1.2170234397098790e+02
RS_630 NS_630 0 1.2170234397098790e+02
GL_629 0 NS_629 NS_630 0 4.0778813929127578e-02
GL_630 0 NS_630 NS_629 0 -4.0778813929127578e-02
GS_629_6 0 NS_629 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 631/632
CS_631 NS_631 0 9.9999999999999998e-13
CS_632 NS_632 0 9.9999999999999998e-13
RS_631 NS_631 0 1.1550510326517782e+02
RS_632 NS_632 0 1.1550510326517782e+02
GL_631 0 NS_631 NS_632 0 5.7236026076957713e-02
GL_632 0 NS_632 NS_631 0 -5.7236026076957713e-02
GS_631_6 0 NS_631 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 633/634
CS_633 NS_633 0 9.9999999999999998e-13
CS_634 NS_634 0 9.9999999999999998e-13
RS_633 NS_633 0 6.2039157456337159e+02
RS_634 NS_634 0 6.2039157456337159e+02
GL_633 0 NS_633 NS_634 0 1.9354364738401211e-02
GL_634 0 NS_634 NS_633 0 -1.9354364738401211e-02
GS_633_6 0 NS_633 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 635/636
CS_635 NS_635 0 9.9999999999999998e-13
CS_636 NS_636 0 9.9999999999999998e-13
RS_635 NS_635 0 1.1050313240441588e+02
RS_636 NS_636 0 1.1050313240441587e+02
GL_635 0 NS_635 NS_636 0 1.6472588786558075e-02
GL_636 0 NS_636 NS_635 0 -1.6472588786558075e-02
GS_635_6 0 NS_635 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 637/638
CS_637 NS_637 0 9.9999999999999998e-13
CS_638 NS_638 0 9.9999999999999998e-13
RS_637 NS_637 0 1.2869119986945731e+02
RS_638 NS_638 0 1.2869119986945731e+02
GL_637 0 NS_637 NS_638 0 2.0888592987579706e-02
GL_638 0 NS_638 NS_637 0 -2.0888592987579706e-02
GS_637_6 0 NS_637 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 639/640
CS_639 NS_639 0 9.9999999999999998e-13
CS_640 NS_640 0 9.9999999999999998e-13
RS_639 NS_639 0 1.4314560950270646e+02
RS_640 NS_640 0 1.4314560950270646e+02
GL_639 0 NS_639 NS_640 0 9.7871236580563716e-03
GL_640 0 NS_640 NS_639 0 -9.7871236580563716e-03
GS_639_6 0 NS_639 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 641/642
CS_641 NS_641 0 9.9999999999999998e-13
CS_642 NS_642 0 9.9999999999999998e-13
RS_641 NS_641 0 1.1863004336811436e+02
RS_642 NS_642 0 1.1863004336811436e+02
GL_641 0 NS_641 NS_642 0 3.7627463994326378e-02
GL_642 0 NS_642 NS_641 0 -3.7627463994326378e-02
GS_641_6 0 NS_641 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 643/644
CS_643 NS_643 0 9.9999999999999998e-13
CS_644 NS_644 0 9.9999999999999998e-13
RS_643 NS_643 0 1.2686172273444870e+02
RS_644 NS_644 0 1.2686172273444869e+02
GL_643 0 NS_643 NS_644 0 3.1975218188091938e-02
GL_644 0 NS_644 NS_643 0 -3.1975218188091938e-02
GS_643_6 0 NS_643 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 645/646
CS_645 NS_645 0 9.9999999999999998e-13
CS_646 NS_646 0 9.9999999999999998e-13
RS_645 NS_645 0 1.3141621772977734e+02
RS_646 NS_646 0 1.3141621772977737e+02
GL_645 0 NS_645 NS_646 0 2.8228381102665165e-02
GL_646 0 NS_646 NS_645 0 -2.8228381102665165e-02
GS_645_6 0 NS_645 NA_6 0 4.7428518688027549e-01
*
* Complex pair n. 647/648
CS_647 NS_647 0 9.9999999999999998e-13
CS_648 NS_648 0 9.9999999999999998e-13
RS_647 NS_647 0 1.2452833644614726e+02
RS_648 NS_648 0 1.2452833644614726e+02
GL_647 0 NS_647 NS_648 0 2.1457325426059259e-03
GL_648 0 NS_648 NS_647 0 -2.1457325426059259e-03
GS_647_6 0 NS_647 NA_6 0 4.7428518688027549e-01
*
* Real pole n. 649
CS_649 NS_649 0 9.9999999999999998e-13
RS_649 NS_649 0 3.8329546824379270e+00
GS_649_7 0 NS_649 NA_7 0 4.7428518688027549e-01
*
* Real pole n. 650
CS_650 NS_650 0 9.9999999999999998e-13
RS_650 NS_650 0 1.0843846705160875e+04
GS_650_7 0 NS_650 NA_7 0 4.7428518688027549e-01
*
* Real pole n. 651
CS_651 NS_651 0 9.9999999999999998e-13
RS_651 NS_651 0 3.3457029134706481e+03
GS_651_7 0 NS_651 NA_7 0 4.7428518688027549e-01
*
* Real pole n. 652
CS_652 NS_652 0 9.9999999999999998e-13
RS_652 NS_652 0 5.4313394337993634e+02
GS_652_7 0 NS_652 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 653/654
CS_653 NS_653 0 9.9999999999999998e-13
CS_654 NS_654 0 9.9999999999999998e-13
RS_653 NS_653 0 2.0342898045173075e+02
RS_654 NS_654 0 2.0342898045173075e+02
GL_653 0 NS_653 NS_654 0 2.5883098202682536e-01
GL_654 0 NS_654 NS_653 0 -2.5883098202682536e-01
GS_653_7 0 NS_653 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 655/656
CS_655 NS_655 0 9.9999999999999998e-13
CS_656 NS_656 0 9.9999999999999998e-13
RS_655 NS_655 0 1.2739936959261519e+02
RS_656 NS_656 0 1.2739936959261519e+02
GL_655 0 NS_655 NS_656 0 2.5122204303896745e-01
GL_656 0 NS_656 NS_655 0 -2.5122204303896745e-01
GS_655_7 0 NS_655 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 657/658
CS_657 NS_657 0 9.9999999999999998e-13
CS_658 NS_658 0 9.9999999999999998e-13
RS_657 NS_657 0 1.1105129555360161e+02
RS_658 NS_658 0 1.1105129555360161e+02
GL_657 0 NS_657 NS_658 0 2.4643422119526687e-01
GL_658 0 NS_658 NS_657 0 -2.4643422119526687e-01
GS_657_7 0 NS_657 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 659/660
CS_659 NS_659 0 9.9999999999999998e-13
CS_660 NS_660 0 9.9999999999999998e-13
RS_659 NS_659 0 1.0856580972218713e+02
RS_660 NS_660 0 1.0856580972218713e+02
GL_659 0 NS_659 NS_660 0 2.4007148694878275e-01
GL_660 0 NS_660 NS_659 0 -2.4007148694878275e-01
GS_659_7 0 NS_659 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 661/662
CS_661 NS_661 0 9.9999999999999998e-13
CS_662 NS_662 0 9.9999999999999998e-13
RS_661 NS_661 0 1.0135860176893434e+02
RS_662 NS_662 0 1.0135860176893435e+02
GL_661 0 NS_661 NS_662 0 2.3570758371916220e-01
GL_662 0 NS_662 NS_661 0 -2.3570758371916220e-01
GS_661_7 0 NS_661 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 663/664
CS_663 NS_663 0 9.9999999999999998e-13
CS_664 NS_664 0 9.9999999999999998e-13
RS_663 NS_663 0 1.2858526276753685e+02
RS_664 NS_664 0 1.2858526276753685e+02
GL_663 0 NS_663 NS_664 0 2.2966634995600790e-01
GL_664 0 NS_664 NS_663 0 -2.2966634995600790e-01
GS_663_7 0 NS_663 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 665/666
CS_665 NS_665 0 9.9999999999999998e-13
CS_666 NS_666 0 9.9999999999999998e-13
RS_665 NS_665 0 1.1773437593549667e+02
RS_666 NS_666 0 1.1773437593549667e+02
GL_665 0 NS_665 NS_666 0 2.2732609444056490e-01
GL_666 0 NS_666 NS_665 0 -2.2732609444056490e-01
GS_665_7 0 NS_665 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 667/668
CS_667 NS_667 0 9.9999999999999998e-13
CS_668 NS_668 0 9.9999999999999998e-13
RS_667 NS_667 0 9.8170265044265946e+01
RS_668 NS_668 0 9.8170265044265932e+01
GL_667 0 NS_667 NS_668 0 2.2031598117475365e-01
GL_668 0 NS_668 NS_667 0 -2.2031598117475365e-01
GS_667_7 0 NS_667 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 669/670
CS_669 NS_669 0 9.9999999999999998e-13
CS_670 NS_670 0 9.9999999999999998e-13
RS_669 NS_669 0 9.5355901421613709e+01
RS_670 NS_670 0 9.5355901421613694e+01
GL_669 0 NS_669 NS_670 0 2.1739680820836188e-01
GL_670 0 NS_670 NS_669 0 -2.1739680820836188e-01
GS_669_7 0 NS_669 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 671/672
CS_671 NS_671 0 9.9999999999999998e-13
CS_672 NS_672 0 9.9999999999999998e-13
RS_671 NS_671 0 1.0859722031634941e+02
RS_672 NS_672 0 1.0859722031634941e+02
GL_671 0 NS_671 NS_672 0 2.0887403840929383e-01
GL_672 0 NS_672 NS_671 0 -2.0887403840929383e-01
GS_671_7 0 NS_671 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 673/674
CS_673 NS_673 0 9.9999999999999998e-13
CS_674 NS_674 0 9.9999999999999998e-13
RS_673 NS_673 0 7.7959989808728068e+01
RS_674 NS_674 0 7.7959989808728054e+01
GL_673 0 NS_673 NS_674 0 2.0447808896343445e-01
GL_674 0 NS_674 NS_673 0 -2.0447808896343445e-01
GS_673_7 0 NS_673 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 675/676
CS_675 NS_675 0 9.9999999999999998e-13
CS_676 NS_676 0 9.9999999999999998e-13
RS_675 NS_675 0 1.1088851678406323e+02
RS_676 NS_676 0 1.1088851678406321e+02
GL_675 0 NS_675 NS_676 0 1.9843399276071924e-01
GL_676 0 NS_676 NS_675 0 -1.9843399276071924e-01
GS_675_7 0 NS_675 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 677/678
CS_677 NS_677 0 9.9999999999999998e-13
CS_678 NS_678 0 9.9999999999999998e-13
RS_677 NS_677 0 8.1179760966262847e+01
RS_678 NS_678 0 8.1179760966262847e+01
GL_677 0 NS_677 NS_678 0 1.8978022990658949e-01
GL_678 0 NS_678 NS_677 0 -1.8978022990658949e-01
GS_677_7 0 NS_677 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 679/680
CS_679 NS_679 0 9.9999999999999998e-13
CS_680 NS_680 0 9.9999999999999998e-13
RS_679 NS_679 0 1.0523970815054612e+02
RS_680 NS_680 0 1.0523970815054612e+02
GL_679 0 NS_679 NS_680 0 1.8836779078363333e-01
GL_680 0 NS_680 NS_679 0 -1.8836779078363333e-01
GS_679_7 0 NS_679 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 681/682
CS_681 NS_681 0 9.9999999999999998e-13
CS_682 NS_682 0 9.9999999999999998e-13
RS_681 NS_681 0 1.1208834663822537e+02
RS_682 NS_682 0 1.1208834663822537e+02
GL_681 0 NS_681 NS_682 0 1.7925451755127267e-01
GL_682 0 NS_682 NS_681 0 -1.7925451755127267e-01
GS_681_7 0 NS_681 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 683/684
CS_683 NS_683 0 9.9999999999999998e-13
CS_684 NS_684 0 9.9999999999999998e-13
RS_683 NS_683 0 9.2475617668062213e+01
RS_684 NS_684 0 9.2475617668062199e+01
GL_683 0 NS_683 NS_684 0 1.7507216970358189e-01
GL_684 0 NS_684 NS_683 0 -1.7507216970358189e-01
GS_683_7 0 NS_683 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 685/686
CS_685 NS_685 0 9.9999999999999998e-13
CS_686 NS_686 0 9.9999999999999998e-13
RS_685 NS_685 0 1.1555782965375326e+02
RS_686 NS_686 0 1.1555782965375326e+02
GL_685 0 NS_685 NS_686 0 1.6918904340923188e-01
GL_686 0 NS_686 NS_685 0 -1.6918904340923188e-01
GS_685_7 0 NS_685 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 687/688
CS_687 NS_687 0 9.9999999999999998e-13
CS_688 NS_688 0 9.9999999999999998e-13
RS_687 NS_687 0 9.6856782813111039e+01
RS_688 NS_688 0 9.6856782813111039e+01
GL_687 0 NS_687 NS_688 0 1.6488898173469207e-01
GL_688 0 NS_688 NS_687 0 -1.6488898173469207e-01
GS_687_7 0 NS_687 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 689/690
CS_689 NS_689 0 9.9999999999999998e-13
CS_690 NS_690 0 9.9999999999999998e-13
RS_689 NS_689 0 1.1717534841017003e+02
RS_690 NS_690 0 1.1717534841017003e+02
GL_689 0 NS_689 NS_690 0 1.5866517390841936e-01
GL_690 0 NS_690 NS_689 0 -1.5866517390841936e-01
GS_689_7 0 NS_689 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 691/692
CS_691 NS_691 0 9.9999999999999998e-13
CS_692 NS_692 0 9.9999999999999998e-13
RS_691 NS_691 0 8.8607873746940697e+01
RS_692 NS_692 0 8.8607873746940697e+01
GL_691 0 NS_691 NS_692 0 1.5214737618207635e-01
GL_692 0 NS_692 NS_691 0 -1.5214737618207635e-01
GS_691_7 0 NS_691 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 693/694
CS_693 NS_693 0 9.9999999999999998e-13
CS_694 NS_694 0 9.9999999999999998e-13
RS_693 NS_693 0 1.1741456484283673e+02
RS_694 NS_694 0 1.1741456484283673e+02
GL_693 0 NS_693 NS_694 0 1.4829748860889613e-01
GL_694 0 NS_694 NS_693 0 -1.4829748860889613e-01
GS_693_7 0 NS_693 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 695/696
CS_695 NS_695 0 9.9999999999999998e-13
CS_696 NS_696 0 9.9999999999999998e-13
RS_695 NS_695 0 1.3292289814180702e+02
RS_696 NS_696 0 1.3292289814180702e+02
GL_695 0 NS_695 NS_696 0 1.4243056778188259e-01
GL_696 0 NS_696 NS_695 0 -1.4243056778188259e-01
GS_695_7 0 NS_695 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 697/698
CS_697 NS_697 0 9.9999999999999998e-13
CS_698 NS_698 0 9.9999999999999998e-13
RS_697 NS_697 0 1.2325134819531741e+02
RS_698 NS_698 0 1.2325134819531739e+02
GL_697 0 NS_697 NS_698 0 1.3890785074828846e-01
GL_698 0 NS_698 NS_697 0 -1.3890785074828846e-01
GS_697_7 0 NS_697 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 699/700
CS_699 NS_699 0 9.9999999999999998e-13
CS_700 NS_700 0 9.9999999999999998e-13
RS_699 NS_699 0 9.1909059882883227e+01
RS_700 NS_700 0 9.1909059882883227e+01
GL_699 0 NS_699 NS_700 0 1.3373879533989103e-01
GL_700 0 NS_700 NS_699 0 -1.3373879533989103e-01
GS_699_7 0 NS_699 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 701/702
CS_701 NS_701 0 9.9999999999999998e-13
CS_702 NS_702 0 9.9999999999999998e-13
RS_701 NS_701 0 1.2276824880349510e+02
RS_702 NS_702 0 1.2276824880349510e+02
GL_701 0 NS_701 NS_702 0 1.2885409674522977e-01
GL_702 0 NS_702 NS_701 0 -1.2885409674522977e-01
GS_701_7 0 NS_701 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 703/704
CS_703 NS_703 0 9.9999999999999998e-13
CS_704 NS_704 0 9.9999999999999998e-13
RS_703 NS_703 0 1.1612442076026501e+02
RS_704 NS_704 0 1.1612442076026501e+02
GL_703 0 NS_703 NS_704 0 1.2417838026896348e-01
GL_704 0 NS_704 NS_703 0 -1.2417838026896348e-01
GS_703_7 0 NS_703 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 705/706
CS_705 NS_705 0 9.9999999999999998e-13
CS_706 NS_706 0 9.9999999999999998e-13
RS_705 NS_705 0 1.2130204223875414e+02
RS_706 NS_706 0 1.2130204223875414e+02
GL_705 0 NS_705 NS_706 0 1.1919240021970828e-01
GL_706 0 NS_706 NS_705 0 -1.1919240021970828e-01
GS_705_7 0 NS_705 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 707/708
CS_707 NS_707 0 9.9999999999999998e-13
CS_708 NS_708 0 9.9999999999999998e-13
RS_707 NS_707 0 9.3083309227260045e+01
RS_708 NS_708 0 9.3083309227260045e+01
GL_707 0 NS_707 NS_708 0 1.1485268189050464e-01
GL_708 0 NS_708 NS_707 0 -1.1485268189050464e-01
GS_707_7 0 NS_707 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 709/710
CS_709 NS_709 0 9.9999999999999998e-13
CS_710 NS_710 0 9.9999999999999998e-13
RS_709 NS_709 0 1.2387094149263906e+02
RS_710 NS_710 0 1.2387094149263908e+02
GL_709 0 NS_709 NS_710 0 1.0935451806229070e-01
GL_710 0 NS_710 NS_709 0 -1.0935451806229070e-01
GS_709_7 0 NS_709 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 711/712
CS_711 NS_711 0 9.9999999999999998e-13
CS_712 NS_712 0 9.9999999999999998e-13
RS_711 NS_711 0 1.1186020221520803e+02
RS_712 NS_712 0 1.1186020221520802e+02
GL_711 0 NS_711 NS_712 0 1.0538242730807947e-01
GL_712 0 NS_712 NS_711 0 -1.0538242730807947e-01
GS_711_7 0 NS_711 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 713/714
CS_713 NS_713 0 9.9999999999999998e-13
CS_714 NS_714 0 9.9999999999999998e-13
RS_713 NS_713 0 1.2031265815570148e+02
RS_714 NS_714 0 1.2031265815570150e+02
GL_713 0 NS_713 NS_714 0 9.9497602364102364e-02
GL_714 0 NS_714 NS_713 0 -9.9497602364102364e-02
GS_713_7 0 NS_713 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 715/716
CS_715 NS_715 0 9.9999999999999998e-13
CS_716 NS_716 0 9.9999999999999998e-13
RS_715 NS_715 0 9.6254518048655143e+01
RS_716 NS_716 0 9.6254518048655143e+01
GL_715 0 NS_715 NS_716 0 9.5930770757699110e-02
GL_716 0 NS_716 NS_715 0 -9.5930770757699110e-02
GS_715_7 0 NS_715 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 717/718
CS_717 NS_717 0 9.9999999999999998e-13
CS_718 NS_718 0 9.9999999999999998e-13
RS_717 NS_717 0 1.2318640771018909e+02
RS_718 NS_718 0 1.2318640771018909e+02
GL_717 0 NS_717 NS_718 0 8.9880619653662355e-02
GL_718 0 NS_718 NS_717 0 -8.9880619653662355e-02
GS_717_7 0 NS_717 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 719/720
CS_719 NS_719 0 9.9999999999999998e-13
CS_720 NS_720 0 9.9999999999999998e-13
RS_719 NS_719 0 1.1312630346155738e+02
RS_720 NS_720 0 1.1312630346155738e+02
GL_719 0 NS_719 NS_720 0 8.6534434501560398e-02
GL_720 0 NS_720 NS_719 0 -8.6534434501560398e-02
GS_719_7 0 NS_719 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 721/722
CS_721 NS_721 0 9.9999999999999998e-13
CS_722 NS_722 0 9.9999999999999998e-13
RS_721 NS_721 0 1.1831504703984019e+02
RS_722 NS_722 0 1.1831504703984019e+02
GL_721 0 NS_721 NS_722 0 7.9864296724202116e-02
GL_722 0 NS_722 NS_721 0 -7.9864296724202116e-02
GS_721_7 0 NS_721 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 723/724
CS_723 NS_723 0 9.9999999999999998e-13
CS_724 NS_724 0 9.9999999999999998e-13
RS_723 NS_723 0 1.0281987486447559e+02
RS_724 NS_724 0 1.0281987486447559e+02
GL_723 0 NS_723 NS_724 0 7.6950339194481784e-02
GL_724 0 NS_724 NS_723 0 -7.6950339194481784e-02
GS_723_7 0 NS_723 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 725/726
CS_725 NS_725 0 9.9999999999999998e-13
CS_726 NS_726 0 9.9999999999999998e-13
RS_725 NS_725 0 1.2230186914382300e+02
RS_726 NS_726 0 1.2230186914382300e+02
GL_725 0 NS_725 NS_726 0 7.0709298709435750e-02
GL_726 0 NS_726 NS_725 0 -7.0709298709435750e-02
GS_725_7 0 NS_725 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 727/728
CS_727 NS_727 0 9.9999999999999998e-13
CS_728 NS_728 0 9.9999999999999998e-13
RS_727 NS_727 0 1.2215699953322022e+02
RS_728 NS_728 0 1.2215699953322020e+02
GL_727 0 NS_727 NS_728 0 6.7518227185671367e-02
GL_728 0 NS_728 NS_727 0 -6.7518227185671367e-02
GS_727_7 0 NS_727 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 729/730
CS_729 NS_729 0 9.9999999999999998e-13
CS_730 NS_730 0 9.9999999999999998e-13
RS_729 NS_729 0 3.4305564408226764e+03
RS_730 NS_730 0 3.4305564408226769e+03
GL_729 0 NS_729 NS_730 0 5.4396471187208063e-02
GL_730 0 NS_730 NS_729 0 -5.4396471187208063e-02
GS_729_7 0 NS_729 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 731/732
CS_731 NS_731 0 9.9999999999999998e-13
CS_732 NS_732 0 9.9999999999999998e-13
RS_731 NS_731 0 1.1894859826238778e+02
RS_732 NS_732 0 1.1894859826238779e+02
GL_731 0 NS_731 NS_732 0 6.0591569497719031e-02
GL_732 0 NS_732 NS_731 0 -6.0591569497719031e-02
GS_731_7 0 NS_731 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 733/734
CS_733 NS_733 0 9.9999999999999998e-13
CS_734 NS_734 0 9.9999999999999998e-13
RS_733 NS_733 0 1.3537641711503298e+02
RS_734 NS_734 0 1.3537641711503298e+02
GL_733 0 NS_733 NS_734 0 5.1190778164089609e-02
GL_734 0 NS_734 NS_733 0 -5.1190778164089609e-02
GS_733_7 0 NS_733 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 735/736
CS_735 NS_735 0 9.9999999999999998e-13
CS_736 NS_736 0 9.9999999999999998e-13
RS_735 NS_735 0 1.3105452427659637e+02
RS_736 NS_736 0 1.3105452427659637e+02
GL_735 0 NS_735 NS_736 0 4.7418984574880592e-02
GL_736 0 NS_736 NS_735 0 -4.7418984574880592e-02
GS_735_7 0 NS_735 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 737/738
CS_737 NS_737 0 9.9999999999999998e-13
CS_738 NS_738 0 9.9999999999999998e-13
RS_737 NS_737 0 1.2170234397098790e+02
RS_738 NS_738 0 1.2170234397098790e+02
GL_737 0 NS_737 NS_738 0 4.0778813929127578e-02
GL_738 0 NS_738 NS_737 0 -4.0778813929127578e-02
GS_737_7 0 NS_737 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 739/740
CS_739 NS_739 0 9.9999999999999998e-13
CS_740 NS_740 0 9.9999999999999998e-13
RS_739 NS_739 0 1.1550510326517782e+02
RS_740 NS_740 0 1.1550510326517782e+02
GL_739 0 NS_739 NS_740 0 5.7236026076957713e-02
GL_740 0 NS_740 NS_739 0 -5.7236026076957713e-02
GS_739_7 0 NS_739 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 741/742
CS_741 NS_741 0 9.9999999999999998e-13
CS_742 NS_742 0 9.9999999999999998e-13
RS_741 NS_741 0 6.2039157456337159e+02
RS_742 NS_742 0 6.2039157456337159e+02
GL_741 0 NS_741 NS_742 0 1.9354364738401211e-02
GL_742 0 NS_742 NS_741 0 -1.9354364738401211e-02
GS_741_7 0 NS_741 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 743/744
CS_743 NS_743 0 9.9999999999999998e-13
CS_744 NS_744 0 9.9999999999999998e-13
RS_743 NS_743 0 1.1050313240441588e+02
RS_744 NS_744 0 1.1050313240441587e+02
GL_743 0 NS_743 NS_744 0 1.6472588786558075e-02
GL_744 0 NS_744 NS_743 0 -1.6472588786558075e-02
GS_743_7 0 NS_743 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 745/746
CS_745 NS_745 0 9.9999999999999998e-13
CS_746 NS_746 0 9.9999999999999998e-13
RS_745 NS_745 0 1.2869119986945731e+02
RS_746 NS_746 0 1.2869119986945731e+02
GL_745 0 NS_745 NS_746 0 2.0888592987579706e-02
GL_746 0 NS_746 NS_745 0 -2.0888592987579706e-02
GS_745_7 0 NS_745 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 747/748
CS_747 NS_747 0 9.9999999999999998e-13
CS_748 NS_748 0 9.9999999999999998e-13
RS_747 NS_747 0 1.4314560950270646e+02
RS_748 NS_748 0 1.4314560950270646e+02
GL_747 0 NS_747 NS_748 0 9.7871236580563716e-03
GL_748 0 NS_748 NS_747 0 -9.7871236580563716e-03
GS_747_7 0 NS_747 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 749/750
CS_749 NS_749 0 9.9999999999999998e-13
CS_750 NS_750 0 9.9999999999999998e-13
RS_749 NS_749 0 1.1863004336811436e+02
RS_750 NS_750 0 1.1863004336811436e+02
GL_749 0 NS_749 NS_750 0 3.7627463994326378e-02
GL_750 0 NS_750 NS_749 0 -3.7627463994326378e-02
GS_749_7 0 NS_749 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 751/752
CS_751 NS_751 0 9.9999999999999998e-13
CS_752 NS_752 0 9.9999999999999998e-13
RS_751 NS_751 0 1.2686172273444870e+02
RS_752 NS_752 0 1.2686172273444869e+02
GL_751 0 NS_751 NS_752 0 3.1975218188091938e-02
GL_752 0 NS_752 NS_751 0 -3.1975218188091938e-02
GS_751_7 0 NS_751 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 753/754
CS_753 NS_753 0 9.9999999999999998e-13
CS_754 NS_754 0 9.9999999999999998e-13
RS_753 NS_753 0 1.3141621772977734e+02
RS_754 NS_754 0 1.3141621772977737e+02
GL_753 0 NS_753 NS_754 0 2.8228381102665165e-02
GL_754 0 NS_754 NS_753 0 -2.8228381102665165e-02
GS_753_7 0 NS_753 NA_7 0 4.7428518688027549e-01
*
* Complex pair n. 755/756
CS_755 NS_755 0 9.9999999999999998e-13
CS_756 NS_756 0 9.9999999999999998e-13
RS_755 NS_755 0 1.2452833644614726e+02
RS_756 NS_756 0 1.2452833644614726e+02
GL_755 0 NS_755 NS_756 0 2.1457325426059259e-03
GL_756 0 NS_756 NS_755 0 -2.1457325426059259e-03
GS_755_7 0 NS_755 NA_7 0 4.7428518688027549e-01
*
* Real pole n. 757
CS_757 NS_757 0 9.9999999999999998e-13
RS_757 NS_757 0 3.8329546824379270e+00
GS_757_8 0 NS_757 NA_8 0 4.7428518688027549e-01
*
* Real pole n. 758
CS_758 NS_758 0 9.9999999999999998e-13
RS_758 NS_758 0 1.0843846705160875e+04
GS_758_8 0 NS_758 NA_8 0 4.7428518688027549e-01
*
* Real pole n. 759
CS_759 NS_759 0 9.9999999999999998e-13
RS_759 NS_759 0 3.3457029134706481e+03
GS_759_8 0 NS_759 NA_8 0 4.7428518688027549e-01
*
* Real pole n. 760
CS_760 NS_760 0 9.9999999999999998e-13
RS_760 NS_760 0 5.4313394337993634e+02
GS_760_8 0 NS_760 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 761/762
CS_761 NS_761 0 9.9999999999999998e-13
CS_762 NS_762 0 9.9999999999999998e-13
RS_761 NS_761 0 2.0342898045173075e+02
RS_762 NS_762 0 2.0342898045173075e+02
GL_761 0 NS_761 NS_762 0 2.5883098202682536e-01
GL_762 0 NS_762 NS_761 0 -2.5883098202682536e-01
GS_761_8 0 NS_761 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 763/764
CS_763 NS_763 0 9.9999999999999998e-13
CS_764 NS_764 0 9.9999999999999998e-13
RS_763 NS_763 0 1.2739936959261519e+02
RS_764 NS_764 0 1.2739936959261519e+02
GL_763 0 NS_763 NS_764 0 2.5122204303896745e-01
GL_764 0 NS_764 NS_763 0 -2.5122204303896745e-01
GS_763_8 0 NS_763 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 765/766
CS_765 NS_765 0 9.9999999999999998e-13
CS_766 NS_766 0 9.9999999999999998e-13
RS_765 NS_765 0 1.1105129555360161e+02
RS_766 NS_766 0 1.1105129555360161e+02
GL_765 0 NS_765 NS_766 0 2.4643422119526687e-01
GL_766 0 NS_766 NS_765 0 -2.4643422119526687e-01
GS_765_8 0 NS_765 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 767/768
CS_767 NS_767 0 9.9999999999999998e-13
CS_768 NS_768 0 9.9999999999999998e-13
RS_767 NS_767 0 1.0856580972218713e+02
RS_768 NS_768 0 1.0856580972218713e+02
GL_767 0 NS_767 NS_768 0 2.4007148694878275e-01
GL_768 0 NS_768 NS_767 0 -2.4007148694878275e-01
GS_767_8 0 NS_767 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 769/770
CS_769 NS_769 0 9.9999999999999998e-13
CS_770 NS_770 0 9.9999999999999998e-13
RS_769 NS_769 0 1.0135860176893434e+02
RS_770 NS_770 0 1.0135860176893435e+02
GL_769 0 NS_769 NS_770 0 2.3570758371916220e-01
GL_770 0 NS_770 NS_769 0 -2.3570758371916220e-01
GS_769_8 0 NS_769 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 771/772
CS_771 NS_771 0 9.9999999999999998e-13
CS_772 NS_772 0 9.9999999999999998e-13
RS_771 NS_771 0 1.2858526276753685e+02
RS_772 NS_772 0 1.2858526276753685e+02
GL_771 0 NS_771 NS_772 0 2.2966634995600790e-01
GL_772 0 NS_772 NS_771 0 -2.2966634995600790e-01
GS_771_8 0 NS_771 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 773/774
CS_773 NS_773 0 9.9999999999999998e-13
CS_774 NS_774 0 9.9999999999999998e-13
RS_773 NS_773 0 1.1773437593549667e+02
RS_774 NS_774 0 1.1773437593549667e+02
GL_773 0 NS_773 NS_774 0 2.2732609444056490e-01
GL_774 0 NS_774 NS_773 0 -2.2732609444056490e-01
GS_773_8 0 NS_773 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 775/776
CS_775 NS_775 0 9.9999999999999998e-13
CS_776 NS_776 0 9.9999999999999998e-13
RS_775 NS_775 0 9.8170265044265946e+01
RS_776 NS_776 0 9.8170265044265932e+01
GL_775 0 NS_775 NS_776 0 2.2031598117475365e-01
GL_776 0 NS_776 NS_775 0 -2.2031598117475365e-01
GS_775_8 0 NS_775 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 777/778
CS_777 NS_777 0 9.9999999999999998e-13
CS_778 NS_778 0 9.9999999999999998e-13
RS_777 NS_777 0 9.5355901421613709e+01
RS_778 NS_778 0 9.5355901421613694e+01
GL_777 0 NS_777 NS_778 0 2.1739680820836188e-01
GL_778 0 NS_778 NS_777 0 -2.1739680820836188e-01
GS_777_8 0 NS_777 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 779/780
CS_779 NS_779 0 9.9999999999999998e-13
CS_780 NS_780 0 9.9999999999999998e-13
RS_779 NS_779 0 1.0859722031634941e+02
RS_780 NS_780 0 1.0859722031634941e+02
GL_779 0 NS_779 NS_780 0 2.0887403840929383e-01
GL_780 0 NS_780 NS_779 0 -2.0887403840929383e-01
GS_779_8 0 NS_779 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 781/782
CS_781 NS_781 0 9.9999999999999998e-13
CS_782 NS_782 0 9.9999999999999998e-13
RS_781 NS_781 0 7.7959989808728068e+01
RS_782 NS_782 0 7.7959989808728054e+01
GL_781 0 NS_781 NS_782 0 2.0447808896343445e-01
GL_782 0 NS_782 NS_781 0 -2.0447808896343445e-01
GS_781_8 0 NS_781 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 783/784
CS_783 NS_783 0 9.9999999999999998e-13
CS_784 NS_784 0 9.9999999999999998e-13
RS_783 NS_783 0 1.1088851678406323e+02
RS_784 NS_784 0 1.1088851678406321e+02
GL_783 0 NS_783 NS_784 0 1.9843399276071924e-01
GL_784 0 NS_784 NS_783 0 -1.9843399276071924e-01
GS_783_8 0 NS_783 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 785/786
CS_785 NS_785 0 9.9999999999999998e-13
CS_786 NS_786 0 9.9999999999999998e-13
RS_785 NS_785 0 8.1179760966262847e+01
RS_786 NS_786 0 8.1179760966262847e+01
GL_785 0 NS_785 NS_786 0 1.8978022990658949e-01
GL_786 0 NS_786 NS_785 0 -1.8978022990658949e-01
GS_785_8 0 NS_785 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 787/788
CS_787 NS_787 0 9.9999999999999998e-13
CS_788 NS_788 0 9.9999999999999998e-13
RS_787 NS_787 0 1.0523970815054612e+02
RS_788 NS_788 0 1.0523970815054612e+02
GL_787 0 NS_787 NS_788 0 1.8836779078363333e-01
GL_788 0 NS_788 NS_787 0 -1.8836779078363333e-01
GS_787_8 0 NS_787 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 789/790
CS_789 NS_789 0 9.9999999999999998e-13
CS_790 NS_790 0 9.9999999999999998e-13
RS_789 NS_789 0 1.1208834663822537e+02
RS_790 NS_790 0 1.1208834663822537e+02
GL_789 0 NS_789 NS_790 0 1.7925451755127267e-01
GL_790 0 NS_790 NS_789 0 -1.7925451755127267e-01
GS_789_8 0 NS_789 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 791/792
CS_791 NS_791 0 9.9999999999999998e-13
CS_792 NS_792 0 9.9999999999999998e-13
RS_791 NS_791 0 9.2475617668062213e+01
RS_792 NS_792 0 9.2475617668062199e+01
GL_791 0 NS_791 NS_792 0 1.7507216970358189e-01
GL_792 0 NS_792 NS_791 0 -1.7507216970358189e-01
GS_791_8 0 NS_791 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 793/794
CS_793 NS_793 0 9.9999999999999998e-13
CS_794 NS_794 0 9.9999999999999998e-13
RS_793 NS_793 0 1.1555782965375326e+02
RS_794 NS_794 0 1.1555782965375326e+02
GL_793 0 NS_793 NS_794 0 1.6918904340923188e-01
GL_794 0 NS_794 NS_793 0 -1.6918904340923188e-01
GS_793_8 0 NS_793 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 795/796
CS_795 NS_795 0 9.9999999999999998e-13
CS_796 NS_796 0 9.9999999999999998e-13
RS_795 NS_795 0 9.6856782813111039e+01
RS_796 NS_796 0 9.6856782813111039e+01
GL_795 0 NS_795 NS_796 0 1.6488898173469207e-01
GL_796 0 NS_796 NS_795 0 -1.6488898173469207e-01
GS_795_8 0 NS_795 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 797/798
CS_797 NS_797 0 9.9999999999999998e-13
CS_798 NS_798 0 9.9999999999999998e-13
RS_797 NS_797 0 1.1717534841017003e+02
RS_798 NS_798 0 1.1717534841017003e+02
GL_797 0 NS_797 NS_798 0 1.5866517390841936e-01
GL_798 0 NS_798 NS_797 0 -1.5866517390841936e-01
GS_797_8 0 NS_797 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 799/800
CS_799 NS_799 0 9.9999999999999998e-13
CS_800 NS_800 0 9.9999999999999998e-13
RS_799 NS_799 0 8.8607873746940697e+01
RS_800 NS_800 0 8.8607873746940697e+01
GL_799 0 NS_799 NS_800 0 1.5214737618207635e-01
GL_800 0 NS_800 NS_799 0 -1.5214737618207635e-01
GS_799_8 0 NS_799 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 801/802
CS_801 NS_801 0 9.9999999999999998e-13
CS_802 NS_802 0 9.9999999999999998e-13
RS_801 NS_801 0 1.1741456484283673e+02
RS_802 NS_802 0 1.1741456484283673e+02
GL_801 0 NS_801 NS_802 0 1.4829748860889613e-01
GL_802 0 NS_802 NS_801 0 -1.4829748860889613e-01
GS_801_8 0 NS_801 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 803/804
CS_803 NS_803 0 9.9999999999999998e-13
CS_804 NS_804 0 9.9999999999999998e-13
RS_803 NS_803 0 1.3292289814180702e+02
RS_804 NS_804 0 1.3292289814180702e+02
GL_803 0 NS_803 NS_804 0 1.4243056778188259e-01
GL_804 0 NS_804 NS_803 0 -1.4243056778188259e-01
GS_803_8 0 NS_803 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 805/806
CS_805 NS_805 0 9.9999999999999998e-13
CS_806 NS_806 0 9.9999999999999998e-13
RS_805 NS_805 0 1.2325134819531741e+02
RS_806 NS_806 0 1.2325134819531739e+02
GL_805 0 NS_805 NS_806 0 1.3890785074828846e-01
GL_806 0 NS_806 NS_805 0 -1.3890785074828846e-01
GS_805_8 0 NS_805 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 807/808
CS_807 NS_807 0 9.9999999999999998e-13
CS_808 NS_808 0 9.9999999999999998e-13
RS_807 NS_807 0 9.1909059882883227e+01
RS_808 NS_808 0 9.1909059882883227e+01
GL_807 0 NS_807 NS_808 0 1.3373879533989103e-01
GL_808 0 NS_808 NS_807 0 -1.3373879533989103e-01
GS_807_8 0 NS_807 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 809/810
CS_809 NS_809 0 9.9999999999999998e-13
CS_810 NS_810 0 9.9999999999999998e-13
RS_809 NS_809 0 1.2276824880349510e+02
RS_810 NS_810 0 1.2276824880349510e+02
GL_809 0 NS_809 NS_810 0 1.2885409674522977e-01
GL_810 0 NS_810 NS_809 0 -1.2885409674522977e-01
GS_809_8 0 NS_809 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 811/812
CS_811 NS_811 0 9.9999999999999998e-13
CS_812 NS_812 0 9.9999999999999998e-13
RS_811 NS_811 0 1.1612442076026501e+02
RS_812 NS_812 0 1.1612442076026501e+02
GL_811 0 NS_811 NS_812 0 1.2417838026896348e-01
GL_812 0 NS_812 NS_811 0 -1.2417838026896348e-01
GS_811_8 0 NS_811 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 813/814
CS_813 NS_813 0 9.9999999999999998e-13
CS_814 NS_814 0 9.9999999999999998e-13
RS_813 NS_813 0 1.2130204223875414e+02
RS_814 NS_814 0 1.2130204223875414e+02
GL_813 0 NS_813 NS_814 0 1.1919240021970828e-01
GL_814 0 NS_814 NS_813 0 -1.1919240021970828e-01
GS_813_8 0 NS_813 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 815/816
CS_815 NS_815 0 9.9999999999999998e-13
CS_816 NS_816 0 9.9999999999999998e-13
RS_815 NS_815 0 9.3083309227260045e+01
RS_816 NS_816 0 9.3083309227260045e+01
GL_815 0 NS_815 NS_816 0 1.1485268189050464e-01
GL_816 0 NS_816 NS_815 0 -1.1485268189050464e-01
GS_815_8 0 NS_815 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 817/818
CS_817 NS_817 0 9.9999999999999998e-13
CS_818 NS_818 0 9.9999999999999998e-13
RS_817 NS_817 0 1.2387094149263906e+02
RS_818 NS_818 0 1.2387094149263908e+02
GL_817 0 NS_817 NS_818 0 1.0935451806229070e-01
GL_818 0 NS_818 NS_817 0 -1.0935451806229070e-01
GS_817_8 0 NS_817 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 819/820
CS_819 NS_819 0 9.9999999999999998e-13
CS_820 NS_820 0 9.9999999999999998e-13
RS_819 NS_819 0 1.1186020221520803e+02
RS_820 NS_820 0 1.1186020221520802e+02
GL_819 0 NS_819 NS_820 0 1.0538242730807947e-01
GL_820 0 NS_820 NS_819 0 -1.0538242730807947e-01
GS_819_8 0 NS_819 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 821/822
CS_821 NS_821 0 9.9999999999999998e-13
CS_822 NS_822 0 9.9999999999999998e-13
RS_821 NS_821 0 1.2031265815570148e+02
RS_822 NS_822 0 1.2031265815570150e+02
GL_821 0 NS_821 NS_822 0 9.9497602364102364e-02
GL_822 0 NS_822 NS_821 0 -9.9497602364102364e-02
GS_821_8 0 NS_821 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 823/824
CS_823 NS_823 0 9.9999999999999998e-13
CS_824 NS_824 0 9.9999999999999998e-13
RS_823 NS_823 0 9.6254518048655143e+01
RS_824 NS_824 0 9.6254518048655143e+01
GL_823 0 NS_823 NS_824 0 9.5930770757699110e-02
GL_824 0 NS_824 NS_823 0 -9.5930770757699110e-02
GS_823_8 0 NS_823 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 825/826
CS_825 NS_825 0 9.9999999999999998e-13
CS_826 NS_826 0 9.9999999999999998e-13
RS_825 NS_825 0 1.2318640771018909e+02
RS_826 NS_826 0 1.2318640771018909e+02
GL_825 0 NS_825 NS_826 0 8.9880619653662355e-02
GL_826 0 NS_826 NS_825 0 -8.9880619653662355e-02
GS_825_8 0 NS_825 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 827/828
CS_827 NS_827 0 9.9999999999999998e-13
CS_828 NS_828 0 9.9999999999999998e-13
RS_827 NS_827 0 1.1312630346155738e+02
RS_828 NS_828 0 1.1312630346155738e+02
GL_827 0 NS_827 NS_828 0 8.6534434501560398e-02
GL_828 0 NS_828 NS_827 0 -8.6534434501560398e-02
GS_827_8 0 NS_827 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 829/830
CS_829 NS_829 0 9.9999999999999998e-13
CS_830 NS_830 0 9.9999999999999998e-13
RS_829 NS_829 0 1.1831504703984019e+02
RS_830 NS_830 0 1.1831504703984019e+02
GL_829 0 NS_829 NS_830 0 7.9864296724202116e-02
GL_830 0 NS_830 NS_829 0 -7.9864296724202116e-02
GS_829_8 0 NS_829 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 831/832
CS_831 NS_831 0 9.9999999999999998e-13
CS_832 NS_832 0 9.9999999999999998e-13
RS_831 NS_831 0 1.0281987486447559e+02
RS_832 NS_832 0 1.0281987486447559e+02
GL_831 0 NS_831 NS_832 0 7.6950339194481784e-02
GL_832 0 NS_832 NS_831 0 -7.6950339194481784e-02
GS_831_8 0 NS_831 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 833/834
CS_833 NS_833 0 9.9999999999999998e-13
CS_834 NS_834 0 9.9999999999999998e-13
RS_833 NS_833 0 1.2230186914382300e+02
RS_834 NS_834 0 1.2230186914382300e+02
GL_833 0 NS_833 NS_834 0 7.0709298709435750e-02
GL_834 0 NS_834 NS_833 0 -7.0709298709435750e-02
GS_833_8 0 NS_833 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 835/836
CS_835 NS_835 0 9.9999999999999998e-13
CS_836 NS_836 0 9.9999999999999998e-13
RS_835 NS_835 0 1.2215699953322022e+02
RS_836 NS_836 0 1.2215699953322020e+02
GL_835 0 NS_835 NS_836 0 6.7518227185671367e-02
GL_836 0 NS_836 NS_835 0 -6.7518227185671367e-02
GS_835_8 0 NS_835 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 837/838
CS_837 NS_837 0 9.9999999999999998e-13
CS_838 NS_838 0 9.9999999999999998e-13
RS_837 NS_837 0 3.4305564408226764e+03
RS_838 NS_838 0 3.4305564408226769e+03
GL_837 0 NS_837 NS_838 0 5.4396471187208063e-02
GL_838 0 NS_838 NS_837 0 -5.4396471187208063e-02
GS_837_8 0 NS_837 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 839/840
CS_839 NS_839 0 9.9999999999999998e-13
CS_840 NS_840 0 9.9999999999999998e-13
RS_839 NS_839 0 1.1894859826238778e+02
RS_840 NS_840 0 1.1894859826238779e+02
GL_839 0 NS_839 NS_840 0 6.0591569497719031e-02
GL_840 0 NS_840 NS_839 0 -6.0591569497719031e-02
GS_839_8 0 NS_839 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 841/842
CS_841 NS_841 0 9.9999999999999998e-13
CS_842 NS_842 0 9.9999999999999998e-13
RS_841 NS_841 0 1.3537641711503298e+02
RS_842 NS_842 0 1.3537641711503298e+02
GL_841 0 NS_841 NS_842 0 5.1190778164089609e-02
GL_842 0 NS_842 NS_841 0 -5.1190778164089609e-02
GS_841_8 0 NS_841 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 843/844
CS_843 NS_843 0 9.9999999999999998e-13
CS_844 NS_844 0 9.9999999999999998e-13
RS_843 NS_843 0 1.3105452427659637e+02
RS_844 NS_844 0 1.3105452427659637e+02
GL_843 0 NS_843 NS_844 0 4.7418984574880592e-02
GL_844 0 NS_844 NS_843 0 -4.7418984574880592e-02
GS_843_8 0 NS_843 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 845/846
CS_845 NS_845 0 9.9999999999999998e-13
CS_846 NS_846 0 9.9999999999999998e-13
RS_845 NS_845 0 1.2170234397098790e+02
RS_846 NS_846 0 1.2170234397098790e+02
GL_845 0 NS_845 NS_846 0 4.0778813929127578e-02
GL_846 0 NS_846 NS_845 0 -4.0778813929127578e-02
GS_845_8 0 NS_845 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 847/848
CS_847 NS_847 0 9.9999999999999998e-13
CS_848 NS_848 0 9.9999999999999998e-13
RS_847 NS_847 0 1.1550510326517782e+02
RS_848 NS_848 0 1.1550510326517782e+02
GL_847 0 NS_847 NS_848 0 5.7236026076957713e-02
GL_848 0 NS_848 NS_847 0 -5.7236026076957713e-02
GS_847_8 0 NS_847 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 849/850
CS_849 NS_849 0 9.9999999999999998e-13
CS_850 NS_850 0 9.9999999999999998e-13
RS_849 NS_849 0 6.2039157456337159e+02
RS_850 NS_850 0 6.2039157456337159e+02
GL_849 0 NS_849 NS_850 0 1.9354364738401211e-02
GL_850 0 NS_850 NS_849 0 -1.9354364738401211e-02
GS_849_8 0 NS_849 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 851/852
CS_851 NS_851 0 9.9999999999999998e-13
CS_852 NS_852 0 9.9999999999999998e-13
RS_851 NS_851 0 1.1050313240441588e+02
RS_852 NS_852 0 1.1050313240441587e+02
GL_851 0 NS_851 NS_852 0 1.6472588786558075e-02
GL_852 0 NS_852 NS_851 0 -1.6472588786558075e-02
GS_851_8 0 NS_851 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 853/854
CS_853 NS_853 0 9.9999999999999998e-13
CS_854 NS_854 0 9.9999999999999998e-13
RS_853 NS_853 0 1.2869119986945731e+02
RS_854 NS_854 0 1.2869119986945731e+02
GL_853 0 NS_853 NS_854 0 2.0888592987579706e-02
GL_854 0 NS_854 NS_853 0 -2.0888592987579706e-02
GS_853_8 0 NS_853 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 855/856
CS_855 NS_855 0 9.9999999999999998e-13
CS_856 NS_856 0 9.9999999999999998e-13
RS_855 NS_855 0 1.4314560950270646e+02
RS_856 NS_856 0 1.4314560950270646e+02
GL_855 0 NS_855 NS_856 0 9.7871236580563716e-03
GL_856 0 NS_856 NS_855 0 -9.7871236580563716e-03
GS_855_8 0 NS_855 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 857/858
CS_857 NS_857 0 9.9999999999999998e-13
CS_858 NS_858 0 9.9999999999999998e-13
RS_857 NS_857 0 1.1863004336811436e+02
RS_858 NS_858 0 1.1863004336811436e+02
GL_857 0 NS_857 NS_858 0 3.7627463994326378e-02
GL_858 0 NS_858 NS_857 0 -3.7627463994326378e-02
GS_857_8 0 NS_857 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 859/860
CS_859 NS_859 0 9.9999999999999998e-13
CS_860 NS_860 0 9.9999999999999998e-13
RS_859 NS_859 0 1.2686172273444870e+02
RS_860 NS_860 0 1.2686172273444869e+02
GL_859 0 NS_859 NS_860 0 3.1975218188091938e-02
GL_860 0 NS_860 NS_859 0 -3.1975218188091938e-02
GS_859_8 0 NS_859 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 861/862
CS_861 NS_861 0 9.9999999999999998e-13
CS_862 NS_862 0 9.9999999999999998e-13
RS_861 NS_861 0 1.3141621772977734e+02
RS_862 NS_862 0 1.3141621772977737e+02
GL_861 0 NS_861 NS_862 0 2.8228381102665165e-02
GL_862 0 NS_862 NS_861 0 -2.8228381102665165e-02
GS_861_8 0 NS_861 NA_8 0 4.7428518688027549e-01
*
* Complex pair n. 863/864
CS_863 NS_863 0 9.9999999999999998e-13
CS_864 NS_864 0 9.9999999999999998e-13
RS_863 NS_863 0 1.2452833644614726e+02
RS_864 NS_864 0 1.2452833644614726e+02
GL_863 0 NS_863 NS_864 0 2.1457325426059259e-03
GL_864 0 NS_864 NS_863 0 -2.1457325426059259e-03
GS_863_8 0 NS_863 NA_8 0 4.7428518688027549e-01
*
* Real pole n. 865
CS_865 NS_865 0 9.9999999999999998e-13
RS_865 NS_865 0 3.8329546824379270e+00
GS_865_9 0 NS_865 NA_9 0 4.7428518688027549e-01
*
* Real pole n. 866
CS_866 NS_866 0 9.9999999999999998e-13
RS_866 NS_866 0 1.0843846705160875e+04
GS_866_9 0 NS_866 NA_9 0 4.7428518688027549e-01
*
* Real pole n. 867
CS_867 NS_867 0 9.9999999999999998e-13
RS_867 NS_867 0 3.3457029134706481e+03
GS_867_9 0 NS_867 NA_9 0 4.7428518688027549e-01
*
* Real pole n. 868
CS_868 NS_868 0 9.9999999999999998e-13
RS_868 NS_868 0 5.4313394337993634e+02
GS_868_9 0 NS_868 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 869/870
CS_869 NS_869 0 9.9999999999999998e-13
CS_870 NS_870 0 9.9999999999999998e-13
RS_869 NS_869 0 2.0342898045173075e+02
RS_870 NS_870 0 2.0342898045173075e+02
GL_869 0 NS_869 NS_870 0 2.5883098202682536e-01
GL_870 0 NS_870 NS_869 0 -2.5883098202682536e-01
GS_869_9 0 NS_869 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 871/872
CS_871 NS_871 0 9.9999999999999998e-13
CS_872 NS_872 0 9.9999999999999998e-13
RS_871 NS_871 0 1.2739936959261519e+02
RS_872 NS_872 0 1.2739936959261519e+02
GL_871 0 NS_871 NS_872 0 2.5122204303896745e-01
GL_872 0 NS_872 NS_871 0 -2.5122204303896745e-01
GS_871_9 0 NS_871 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 873/874
CS_873 NS_873 0 9.9999999999999998e-13
CS_874 NS_874 0 9.9999999999999998e-13
RS_873 NS_873 0 1.1105129555360161e+02
RS_874 NS_874 0 1.1105129555360161e+02
GL_873 0 NS_873 NS_874 0 2.4643422119526687e-01
GL_874 0 NS_874 NS_873 0 -2.4643422119526687e-01
GS_873_9 0 NS_873 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 875/876
CS_875 NS_875 0 9.9999999999999998e-13
CS_876 NS_876 0 9.9999999999999998e-13
RS_875 NS_875 0 1.0856580972218713e+02
RS_876 NS_876 0 1.0856580972218713e+02
GL_875 0 NS_875 NS_876 0 2.4007148694878275e-01
GL_876 0 NS_876 NS_875 0 -2.4007148694878275e-01
GS_875_9 0 NS_875 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 877/878
CS_877 NS_877 0 9.9999999999999998e-13
CS_878 NS_878 0 9.9999999999999998e-13
RS_877 NS_877 0 1.0135860176893434e+02
RS_878 NS_878 0 1.0135860176893435e+02
GL_877 0 NS_877 NS_878 0 2.3570758371916220e-01
GL_878 0 NS_878 NS_877 0 -2.3570758371916220e-01
GS_877_9 0 NS_877 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 879/880
CS_879 NS_879 0 9.9999999999999998e-13
CS_880 NS_880 0 9.9999999999999998e-13
RS_879 NS_879 0 1.2858526276753685e+02
RS_880 NS_880 0 1.2858526276753685e+02
GL_879 0 NS_879 NS_880 0 2.2966634995600790e-01
GL_880 0 NS_880 NS_879 0 -2.2966634995600790e-01
GS_879_9 0 NS_879 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 881/882
CS_881 NS_881 0 9.9999999999999998e-13
CS_882 NS_882 0 9.9999999999999998e-13
RS_881 NS_881 0 1.1773437593549667e+02
RS_882 NS_882 0 1.1773437593549667e+02
GL_881 0 NS_881 NS_882 0 2.2732609444056490e-01
GL_882 0 NS_882 NS_881 0 -2.2732609444056490e-01
GS_881_9 0 NS_881 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 883/884
CS_883 NS_883 0 9.9999999999999998e-13
CS_884 NS_884 0 9.9999999999999998e-13
RS_883 NS_883 0 9.8170265044265946e+01
RS_884 NS_884 0 9.8170265044265932e+01
GL_883 0 NS_883 NS_884 0 2.2031598117475365e-01
GL_884 0 NS_884 NS_883 0 -2.2031598117475365e-01
GS_883_9 0 NS_883 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 885/886
CS_885 NS_885 0 9.9999999999999998e-13
CS_886 NS_886 0 9.9999999999999998e-13
RS_885 NS_885 0 9.5355901421613709e+01
RS_886 NS_886 0 9.5355901421613694e+01
GL_885 0 NS_885 NS_886 0 2.1739680820836188e-01
GL_886 0 NS_886 NS_885 0 -2.1739680820836188e-01
GS_885_9 0 NS_885 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 887/888
CS_887 NS_887 0 9.9999999999999998e-13
CS_888 NS_888 0 9.9999999999999998e-13
RS_887 NS_887 0 1.0859722031634941e+02
RS_888 NS_888 0 1.0859722031634941e+02
GL_887 0 NS_887 NS_888 0 2.0887403840929383e-01
GL_888 0 NS_888 NS_887 0 -2.0887403840929383e-01
GS_887_9 0 NS_887 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 889/890
CS_889 NS_889 0 9.9999999999999998e-13
CS_890 NS_890 0 9.9999999999999998e-13
RS_889 NS_889 0 7.7959989808728068e+01
RS_890 NS_890 0 7.7959989808728054e+01
GL_889 0 NS_889 NS_890 0 2.0447808896343445e-01
GL_890 0 NS_890 NS_889 0 -2.0447808896343445e-01
GS_889_9 0 NS_889 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 891/892
CS_891 NS_891 0 9.9999999999999998e-13
CS_892 NS_892 0 9.9999999999999998e-13
RS_891 NS_891 0 1.1088851678406323e+02
RS_892 NS_892 0 1.1088851678406321e+02
GL_891 0 NS_891 NS_892 0 1.9843399276071924e-01
GL_892 0 NS_892 NS_891 0 -1.9843399276071924e-01
GS_891_9 0 NS_891 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 893/894
CS_893 NS_893 0 9.9999999999999998e-13
CS_894 NS_894 0 9.9999999999999998e-13
RS_893 NS_893 0 8.1179760966262847e+01
RS_894 NS_894 0 8.1179760966262847e+01
GL_893 0 NS_893 NS_894 0 1.8978022990658949e-01
GL_894 0 NS_894 NS_893 0 -1.8978022990658949e-01
GS_893_9 0 NS_893 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 895/896
CS_895 NS_895 0 9.9999999999999998e-13
CS_896 NS_896 0 9.9999999999999998e-13
RS_895 NS_895 0 1.0523970815054612e+02
RS_896 NS_896 0 1.0523970815054612e+02
GL_895 0 NS_895 NS_896 0 1.8836779078363333e-01
GL_896 0 NS_896 NS_895 0 -1.8836779078363333e-01
GS_895_9 0 NS_895 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 897/898
CS_897 NS_897 0 9.9999999999999998e-13
CS_898 NS_898 0 9.9999999999999998e-13
RS_897 NS_897 0 1.1208834663822537e+02
RS_898 NS_898 0 1.1208834663822537e+02
GL_897 0 NS_897 NS_898 0 1.7925451755127267e-01
GL_898 0 NS_898 NS_897 0 -1.7925451755127267e-01
GS_897_9 0 NS_897 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 899/900
CS_899 NS_899 0 9.9999999999999998e-13
CS_900 NS_900 0 9.9999999999999998e-13
RS_899 NS_899 0 9.2475617668062213e+01
RS_900 NS_900 0 9.2475617668062199e+01
GL_899 0 NS_899 NS_900 0 1.7507216970358189e-01
GL_900 0 NS_900 NS_899 0 -1.7507216970358189e-01
GS_899_9 0 NS_899 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 901/902
CS_901 NS_901 0 9.9999999999999998e-13
CS_902 NS_902 0 9.9999999999999998e-13
RS_901 NS_901 0 1.1555782965375326e+02
RS_902 NS_902 0 1.1555782965375326e+02
GL_901 0 NS_901 NS_902 0 1.6918904340923188e-01
GL_902 0 NS_902 NS_901 0 -1.6918904340923188e-01
GS_901_9 0 NS_901 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 903/904
CS_903 NS_903 0 9.9999999999999998e-13
CS_904 NS_904 0 9.9999999999999998e-13
RS_903 NS_903 0 9.6856782813111039e+01
RS_904 NS_904 0 9.6856782813111039e+01
GL_903 0 NS_903 NS_904 0 1.6488898173469207e-01
GL_904 0 NS_904 NS_903 0 -1.6488898173469207e-01
GS_903_9 0 NS_903 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 905/906
CS_905 NS_905 0 9.9999999999999998e-13
CS_906 NS_906 0 9.9999999999999998e-13
RS_905 NS_905 0 1.1717534841017003e+02
RS_906 NS_906 0 1.1717534841017003e+02
GL_905 0 NS_905 NS_906 0 1.5866517390841936e-01
GL_906 0 NS_906 NS_905 0 -1.5866517390841936e-01
GS_905_9 0 NS_905 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 907/908
CS_907 NS_907 0 9.9999999999999998e-13
CS_908 NS_908 0 9.9999999999999998e-13
RS_907 NS_907 0 8.8607873746940697e+01
RS_908 NS_908 0 8.8607873746940697e+01
GL_907 0 NS_907 NS_908 0 1.5214737618207635e-01
GL_908 0 NS_908 NS_907 0 -1.5214737618207635e-01
GS_907_9 0 NS_907 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 909/910
CS_909 NS_909 0 9.9999999999999998e-13
CS_910 NS_910 0 9.9999999999999998e-13
RS_909 NS_909 0 1.1741456484283673e+02
RS_910 NS_910 0 1.1741456484283673e+02
GL_909 0 NS_909 NS_910 0 1.4829748860889613e-01
GL_910 0 NS_910 NS_909 0 -1.4829748860889613e-01
GS_909_9 0 NS_909 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 911/912
CS_911 NS_911 0 9.9999999999999998e-13
CS_912 NS_912 0 9.9999999999999998e-13
RS_911 NS_911 0 1.3292289814180702e+02
RS_912 NS_912 0 1.3292289814180702e+02
GL_911 0 NS_911 NS_912 0 1.4243056778188259e-01
GL_912 0 NS_912 NS_911 0 -1.4243056778188259e-01
GS_911_9 0 NS_911 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 913/914
CS_913 NS_913 0 9.9999999999999998e-13
CS_914 NS_914 0 9.9999999999999998e-13
RS_913 NS_913 0 1.2325134819531741e+02
RS_914 NS_914 0 1.2325134819531739e+02
GL_913 0 NS_913 NS_914 0 1.3890785074828846e-01
GL_914 0 NS_914 NS_913 0 -1.3890785074828846e-01
GS_913_9 0 NS_913 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 915/916
CS_915 NS_915 0 9.9999999999999998e-13
CS_916 NS_916 0 9.9999999999999998e-13
RS_915 NS_915 0 9.1909059882883227e+01
RS_916 NS_916 0 9.1909059882883227e+01
GL_915 0 NS_915 NS_916 0 1.3373879533989103e-01
GL_916 0 NS_916 NS_915 0 -1.3373879533989103e-01
GS_915_9 0 NS_915 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 917/918
CS_917 NS_917 0 9.9999999999999998e-13
CS_918 NS_918 0 9.9999999999999998e-13
RS_917 NS_917 0 1.2276824880349510e+02
RS_918 NS_918 0 1.2276824880349510e+02
GL_917 0 NS_917 NS_918 0 1.2885409674522977e-01
GL_918 0 NS_918 NS_917 0 -1.2885409674522977e-01
GS_917_9 0 NS_917 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 919/920
CS_919 NS_919 0 9.9999999999999998e-13
CS_920 NS_920 0 9.9999999999999998e-13
RS_919 NS_919 0 1.1612442076026501e+02
RS_920 NS_920 0 1.1612442076026501e+02
GL_919 0 NS_919 NS_920 0 1.2417838026896348e-01
GL_920 0 NS_920 NS_919 0 -1.2417838026896348e-01
GS_919_9 0 NS_919 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 921/922
CS_921 NS_921 0 9.9999999999999998e-13
CS_922 NS_922 0 9.9999999999999998e-13
RS_921 NS_921 0 1.2130204223875414e+02
RS_922 NS_922 0 1.2130204223875414e+02
GL_921 0 NS_921 NS_922 0 1.1919240021970828e-01
GL_922 0 NS_922 NS_921 0 -1.1919240021970828e-01
GS_921_9 0 NS_921 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 923/924
CS_923 NS_923 0 9.9999999999999998e-13
CS_924 NS_924 0 9.9999999999999998e-13
RS_923 NS_923 0 9.3083309227260045e+01
RS_924 NS_924 0 9.3083309227260045e+01
GL_923 0 NS_923 NS_924 0 1.1485268189050464e-01
GL_924 0 NS_924 NS_923 0 -1.1485268189050464e-01
GS_923_9 0 NS_923 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 925/926
CS_925 NS_925 0 9.9999999999999998e-13
CS_926 NS_926 0 9.9999999999999998e-13
RS_925 NS_925 0 1.2387094149263906e+02
RS_926 NS_926 0 1.2387094149263908e+02
GL_925 0 NS_925 NS_926 0 1.0935451806229070e-01
GL_926 0 NS_926 NS_925 0 -1.0935451806229070e-01
GS_925_9 0 NS_925 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 927/928
CS_927 NS_927 0 9.9999999999999998e-13
CS_928 NS_928 0 9.9999999999999998e-13
RS_927 NS_927 0 1.1186020221520803e+02
RS_928 NS_928 0 1.1186020221520802e+02
GL_927 0 NS_927 NS_928 0 1.0538242730807947e-01
GL_928 0 NS_928 NS_927 0 -1.0538242730807947e-01
GS_927_9 0 NS_927 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 929/930
CS_929 NS_929 0 9.9999999999999998e-13
CS_930 NS_930 0 9.9999999999999998e-13
RS_929 NS_929 0 1.2031265815570148e+02
RS_930 NS_930 0 1.2031265815570150e+02
GL_929 0 NS_929 NS_930 0 9.9497602364102364e-02
GL_930 0 NS_930 NS_929 0 -9.9497602364102364e-02
GS_929_9 0 NS_929 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 931/932
CS_931 NS_931 0 9.9999999999999998e-13
CS_932 NS_932 0 9.9999999999999998e-13
RS_931 NS_931 0 9.6254518048655143e+01
RS_932 NS_932 0 9.6254518048655143e+01
GL_931 0 NS_931 NS_932 0 9.5930770757699110e-02
GL_932 0 NS_932 NS_931 0 -9.5930770757699110e-02
GS_931_9 0 NS_931 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 933/934
CS_933 NS_933 0 9.9999999999999998e-13
CS_934 NS_934 0 9.9999999999999998e-13
RS_933 NS_933 0 1.2318640771018909e+02
RS_934 NS_934 0 1.2318640771018909e+02
GL_933 0 NS_933 NS_934 0 8.9880619653662355e-02
GL_934 0 NS_934 NS_933 0 -8.9880619653662355e-02
GS_933_9 0 NS_933 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 935/936
CS_935 NS_935 0 9.9999999999999998e-13
CS_936 NS_936 0 9.9999999999999998e-13
RS_935 NS_935 0 1.1312630346155738e+02
RS_936 NS_936 0 1.1312630346155738e+02
GL_935 0 NS_935 NS_936 0 8.6534434501560398e-02
GL_936 0 NS_936 NS_935 0 -8.6534434501560398e-02
GS_935_9 0 NS_935 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 937/938
CS_937 NS_937 0 9.9999999999999998e-13
CS_938 NS_938 0 9.9999999999999998e-13
RS_937 NS_937 0 1.1831504703984019e+02
RS_938 NS_938 0 1.1831504703984019e+02
GL_937 0 NS_937 NS_938 0 7.9864296724202116e-02
GL_938 0 NS_938 NS_937 0 -7.9864296724202116e-02
GS_937_9 0 NS_937 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 939/940
CS_939 NS_939 0 9.9999999999999998e-13
CS_940 NS_940 0 9.9999999999999998e-13
RS_939 NS_939 0 1.0281987486447559e+02
RS_940 NS_940 0 1.0281987486447559e+02
GL_939 0 NS_939 NS_940 0 7.6950339194481784e-02
GL_940 0 NS_940 NS_939 0 -7.6950339194481784e-02
GS_939_9 0 NS_939 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 941/942
CS_941 NS_941 0 9.9999999999999998e-13
CS_942 NS_942 0 9.9999999999999998e-13
RS_941 NS_941 0 1.2230186914382300e+02
RS_942 NS_942 0 1.2230186914382300e+02
GL_941 0 NS_941 NS_942 0 7.0709298709435750e-02
GL_942 0 NS_942 NS_941 0 -7.0709298709435750e-02
GS_941_9 0 NS_941 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 943/944
CS_943 NS_943 0 9.9999999999999998e-13
CS_944 NS_944 0 9.9999999999999998e-13
RS_943 NS_943 0 1.2215699953322022e+02
RS_944 NS_944 0 1.2215699953322020e+02
GL_943 0 NS_943 NS_944 0 6.7518227185671367e-02
GL_944 0 NS_944 NS_943 0 -6.7518227185671367e-02
GS_943_9 0 NS_943 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 945/946
CS_945 NS_945 0 9.9999999999999998e-13
CS_946 NS_946 0 9.9999999999999998e-13
RS_945 NS_945 0 3.4305564408226764e+03
RS_946 NS_946 0 3.4305564408226769e+03
GL_945 0 NS_945 NS_946 0 5.4396471187208063e-02
GL_946 0 NS_946 NS_945 0 -5.4396471187208063e-02
GS_945_9 0 NS_945 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 947/948
CS_947 NS_947 0 9.9999999999999998e-13
CS_948 NS_948 0 9.9999999999999998e-13
RS_947 NS_947 0 1.1894859826238778e+02
RS_948 NS_948 0 1.1894859826238779e+02
GL_947 0 NS_947 NS_948 0 6.0591569497719031e-02
GL_948 0 NS_948 NS_947 0 -6.0591569497719031e-02
GS_947_9 0 NS_947 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 949/950
CS_949 NS_949 0 9.9999999999999998e-13
CS_950 NS_950 0 9.9999999999999998e-13
RS_949 NS_949 0 1.3537641711503298e+02
RS_950 NS_950 0 1.3537641711503298e+02
GL_949 0 NS_949 NS_950 0 5.1190778164089609e-02
GL_950 0 NS_950 NS_949 0 -5.1190778164089609e-02
GS_949_9 0 NS_949 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 951/952
CS_951 NS_951 0 9.9999999999999998e-13
CS_952 NS_952 0 9.9999999999999998e-13
RS_951 NS_951 0 1.3105452427659637e+02
RS_952 NS_952 0 1.3105452427659637e+02
GL_951 0 NS_951 NS_952 0 4.7418984574880592e-02
GL_952 0 NS_952 NS_951 0 -4.7418984574880592e-02
GS_951_9 0 NS_951 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 953/954
CS_953 NS_953 0 9.9999999999999998e-13
CS_954 NS_954 0 9.9999999999999998e-13
RS_953 NS_953 0 1.2170234397098790e+02
RS_954 NS_954 0 1.2170234397098790e+02
GL_953 0 NS_953 NS_954 0 4.0778813929127578e-02
GL_954 0 NS_954 NS_953 0 -4.0778813929127578e-02
GS_953_9 0 NS_953 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 955/956
CS_955 NS_955 0 9.9999999999999998e-13
CS_956 NS_956 0 9.9999999999999998e-13
RS_955 NS_955 0 1.1550510326517782e+02
RS_956 NS_956 0 1.1550510326517782e+02
GL_955 0 NS_955 NS_956 0 5.7236026076957713e-02
GL_956 0 NS_956 NS_955 0 -5.7236026076957713e-02
GS_955_9 0 NS_955 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 957/958
CS_957 NS_957 0 9.9999999999999998e-13
CS_958 NS_958 0 9.9999999999999998e-13
RS_957 NS_957 0 6.2039157456337159e+02
RS_958 NS_958 0 6.2039157456337159e+02
GL_957 0 NS_957 NS_958 0 1.9354364738401211e-02
GL_958 0 NS_958 NS_957 0 -1.9354364738401211e-02
GS_957_9 0 NS_957 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 959/960
CS_959 NS_959 0 9.9999999999999998e-13
CS_960 NS_960 0 9.9999999999999998e-13
RS_959 NS_959 0 1.1050313240441588e+02
RS_960 NS_960 0 1.1050313240441587e+02
GL_959 0 NS_959 NS_960 0 1.6472588786558075e-02
GL_960 0 NS_960 NS_959 0 -1.6472588786558075e-02
GS_959_9 0 NS_959 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 961/962
CS_961 NS_961 0 9.9999999999999998e-13
CS_962 NS_962 0 9.9999999999999998e-13
RS_961 NS_961 0 1.2869119986945731e+02
RS_962 NS_962 0 1.2869119986945731e+02
GL_961 0 NS_961 NS_962 0 2.0888592987579706e-02
GL_962 0 NS_962 NS_961 0 -2.0888592987579706e-02
GS_961_9 0 NS_961 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 963/964
CS_963 NS_963 0 9.9999999999999998e-13
CS_964 NS_964 0 9.9999999999999998e-13
RS_963 NS_963 0 1.4314560950270646e+02
RS_964 NS_964 0 1.4314560950270646e+02
GL_963 0 NS_963 NS_964 0 9.7871236580563716e-03
GL_964 0 NS_964 NS_963 0 -9.7871236580563716e-03
GS_963_9 0 NS_963 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 965/966
CS_965 NS_965 0 9.9999999999999998e-13
CS_966 NS_966 0 9.9999999999999998e-13
RS_965 NS_965 0 1.1863004336811436e+02
RS_966 NS_966 0 1.1863004336811436e+02
GL_965 0 NS_965 NS_966 0 3.7627463994326378e-02
GL_966 0 NS_966 NS_965 0 -3.7627463994326378e-02
GS_965_9 0 NS_965 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 967/968
CS_967 NS_967 0 9.9999999999999998e-13
CS_968 NS_968 0 9.9999999999999998e-13
RS_967 NS_967 0 1.2686172273444870e+02
RS_968 NS_968 0 1.2686172273444869e+02
GL_967 0 NS_967 NS_968 0 3.1975218188091938e-02
GL_968 0 NS_968 NS_967 0 -3.1975218188091938e-02
GS_967_9 0 NS_967 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 969/970
CS_969 NS_969 0 9.9999999999999998e-13
CS_970 NS_970 0 9.9999999999999998e-13
RS_969 NS_969 0 1.3141621772977734e+02
RS_970 NS_970 0 1.3141621772977737e+02
GL_969 0 NS_969 NS_970 0 2.8228381102665165e-02
GL_970 0 NS_970 NS_969 0 -2.8228381102665165e-02
GS_969_9 0 NS_969 NA_9 0 4.7428518688027549e-01
*
* Complex pair n. 971/972
CS_971 NS_971 0 9.9999999999999998e-13
CS_972 NS_972 0 9.9999999999999998e-13
RS_971 NS_971 0 1.2452833644614726e+02
RS_972 NS_972 0 1.2452833644614726e+02
GL_971 0 NS_971 NS_972 0 2.1457325426059259e-03
GL_972 0 NS_972 NS_971 0 -2.1457325426059259e-03
GS_971_9 0 NS_971 NA_9 0 4.7428518688027549e-01
*
* Real pole n. 973
CS_973 NS_973 0 9.9999999999999998e-13
RS_973 NS_973 0 3.8329546824379270e+00
GS_973_10 0 NS_973 NA_10 0 4.7428518688027549e-01
*
* Real pole n. 974
CS_974 NS_974 0 9.9999999999999998e-13
RS_974 NS_974 0 1.0843846705160875e+04
GS_974_10 0 NS_974 NA_10 0 4.7428518688027549e-01
*
* Real pole n. 975
CS_975 NS_975 0 9.9999999999999998e-13
RS_975 NS_975 0 3.3457029134706481e+03
GS_975_10 0 NS_975 NA_10 0 4.7428518688027549e-01
*
* Real pole n. 976
CS_976 NS_976 0 9.9999999999999998e-13
RS_976 NS_976 0 5.4313394337993634e+02
GS_976_10 0 NS_976 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 977/978
CS_977 NS_977 0 9.9999999999999998e-13
CS_978 NS_978 0 9.9999999999999998e-13
RS_977 NS_977 0 2.0342898045173075e+02
RS_978 NS_978 0 2.0342898045173075e+02
GL_977 0 NS_977 NS_978 0 2.5883098202682536e-01
GL_978 0 NS_978 NS_977 0 -2.5883098202682536e-01
GS_977_10 0 NS_977 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 979/980
CS_979 NS_979 0 9.9999999999999998e-13
CS_980 NS_980 0 9.9999999999999998e-13
RS_979 NS_979 0 1.2739936959261519e+02
RS_980 NS_980 0 1.2739936959261519e+02
GL_979 0 NS_979 NS_980 0 2.5122204303896745e-01
GL_980 0 NS_980 NS_979 0 -2.5122204303896745e-01
GS_979_10 0 NS_979 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 981/982
CS_981 NS_981 0 9.9999999999999998e-13
CS_982 NS_982 0 9.9999999999999998e-13
RS_981 NS_981 0 1.1105129555360161e+02
RS_982 NS_982 0 1.1105129555360161e+02
GL_981 0 NS_981 NS_982 0 2.4643422119526687e-01
GL_982 0 NS_982 NS_981 0 -2.4643422119526687e-01
GS_981_10 0 NS_981 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 983/984
CS_983 NS_983 0 9.9999999999999998e-13
CS_984 NS_984 0 9.9999999999999998e-13
RS_983 NS_983 0 1.0856580972218713e+02
RS_984 NS_984 0 1.0856580972218713e+02
GL_983 0 NS_983 NS_984 0 2.4007148694878275e-01
GL_984 0 NS_984 NS_983 0 -2.4007148694878275e-01
GS_983_10 0 NS_983 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 985/986
CS_985 NS_985 0 9.9999999999999998e-13
CS_986 NS_986 0 9.9999999999999998e-13
RS_985 NS_985 0 1.0135860176893434e+02
RS_986 NS_986 0 1.0135860176893435e+02
GL_985 0 NS_985 NS_986 0 2.3570758371916220e-01
GL_986 0 NS_986 NS_985 0 -2.3570758371916220e-01
GS_985_10 0 NS_985 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 987/988
CS_987 NS_987 0 9.9999999999999998e-13
CS_988 NS_988 0 9.9999999999999998e-13
RS_987 NS_987 0 1.2858526276753685e+02
RS_988 NS_988 0 1.2858526276753685e+02
GL_987 0 NS_987 NS_988 0 2.2966634995600790e-01
GL_988 0 NS_988 NS_987 0 -2.2966634995600790e-01
GS_987_10 0 NS_987 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 989/990
CS_989 NS_989 0 9.9999999999999998e-13
CS_990 NS_990 0 9.9999999999999998e-13
RS_989 NS_989 0 1.1773437593549667e+02
RS_990 NS_990 0 1.1773437593549667e+02
GL_989 0 NS_989 NS_990 0 2.2732609444056490e-01
GL_990 0 NS_990 NS_989 0 -2.2732609444056490e-01
GS_989_10 0 NS_989 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 991/992
CS_991 NS_991 0 9.9999999999999998e-13
CS_992 NS_992 0 9.9999999999999998e-13
RS_991 NS_991 0 9.8170265044265946e+01
RS_992 NS_992 0 9.8170265044265932e+01
GL_991 0 NS_991 NS_992 0 2.2031598117475365e-01
GL_992 0 NS_992 NS_991 0 -2.2031598117475365e-01
GS_991_10 0 NS_991 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 993/994
CS_993 NS_993 0 9.9999999999999998e-13
CS_994 NS_994 0 9.9999999999999998e-13
RS_993 NS_993 0 9.5355901421613709e+01
RS_994 NS_994 0 9.5355901421613694e+01
GL_993 0 NS_993 NS_994 0 2.1739680820836188e-01
GL_994 0 NS_994 NS_993 0 -2.1739680820836188e-01
GS_993_10 0 NS_993 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 995/996
CS_995 NS_995 0 9.9999999999999998e-13
CS_996 NS_996 0 9.9999999999999998e-13
RS_995 NS_995 0 1.0859722031634941e+02
RS_996 NS_996 0 1.0859722031634941e+02
GL_995 0 NS_995 NS_996 0 2.0887403840929383e-01
GL_996 0 NS_996 NS_995 0 -2.0887403840929383e-01
GS_995_10 0 NS_995 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 997/998
CS_997 NS_997 0 9.9999999999999998e-13
CS_998 NS_998 0 9.9999999999999998e-13
RS_997 NS_997 0 7.7959989808728068e+01
RS_998 NS_998 0 7.7959989808728054e+01
GL_997 0 NS_997 NS_998 0 2.0447808896343445e-01
GL_998 0 NS_998 NS_997 0 -2.0447808896343445e-01
GS_997_10 0 NS_997 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 999/1000
CS_999 NS_999 0 9.9999999999999998e-13
CS_1000 NS_1000 0 9.9999999999999998e-13
RS_999 NS_999 0 1.1088851678406323e+02
RS_1000 NS_1000 0 1.1088851678406321e+02
GL_999 0 NS_999 NS_1000 0 1.9843399276071924e-01
GL_1000 0 NS_1000 NS_999 0 -1.9843399276071924e-01
GS_999_10 0 NS_999 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1001/1002
CS_1001 NS_1001 0 9.9999999999999998e-13
CS_1002 NS_1002 0 9.9999999999999998e-13
RS_1001 NS_1001 0 8.1179760966262847e+01
RS_1002 NS_1002 0 8.1179760966262847e+01
GL_1001 0 NS_1001 NS_1002 0 1.8978022990658949e-01
GL_1002 0 NS_1002 NS_1001 0 -1.8978022990658949e-01
GS_1001_10 0 NS_1001 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1003/1004
CS_1003 NS_1003 0 9.9999999999999998e-13
CS_1004 NS_1004 0 9.9999999999999998e-13
RS_1003 NS_1003 0 1.0523970815054612e+02
RS_1004 NS_1004 0 1.0523970815054612e+02
GL_1003 0 NS_1003 NS_1004 0 1.8836779078363333e-01
GL_1004 0 NS_1004 NS_1003 0 -1.8836779078363333e-01
GS_1003_10 0 NS_1003 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1005/1006
CS_1005 NS_1005 0 9.9999999999999998e-13
CS_1006 NS_1006 0 9.9999999999999998e-13
RS_1005 NS_1005 0 1.1208834663822537e+02
RS_1006 NS_1006 0 1.1208834663822537e+02
GL_1005 0 NS_1005 NS_1006 0 1.7925451755127267e-01
GL_1006 0 NS_1006 NS_1005 0 -1.7925451755127267e-01
GS_1005_10 0 NS_1005 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1007/1008
CS_1007 NS_1007 0 9.9999999999999998e-13
CS_1008 NS_1008 0 9.9999999999999998e-13
RS_1007 NS_1007 0 9.2475617668062213e+01
RS_1008 NS_1008 0 9.2475617668062199e+01
GL_1007 0 NS_1007 NS_1008 0 1.7507216970358189e-01
GL_1008 0 NS_1008 NS_1007 0 -1.7507216970358189e-01
GS_1007_10 0 NS_1007 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1009/1010
CS_1009 NS_1009 0 9.9999999999999998e-13
CS_1010 NS_1010 0 9.9999999999999998e-13
RS_1009 NS_1009 0 1.1555782965375326e+02
RS_1010 NS_1010 0 1.1555782965375326e+02
GL_1009 0 NS_1009 NS_1010 0 1.6918904340923188e-01
GL_1010 0 NS_1010 NS_1009 0 -1.6918904340923188e-01
GS_1009_10 0 NS_1009 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1011/1012
CS_1011 NS_1011 0 9.9999999999999998e-13
CS_1012 NS_1012 0 9.9999999999999998e-13
RS_1011 NS_1011 0 9.6856782813111039e+01
RS_1012 NS_1012 0 9.6856782813111039e+01
GL_1011 0 NS_1011 NS_1012 0 1.6488898173469207e-01
GL_1012 0 NS_1012 NS_1011 0 -1.6488898173469207e-01
GS_1011_10 0 NS_1011 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1013/1014
CS_1013 NS_1013 0 9.9999999999999998e-13
CS_1014 NS_1014 0 9.9999999999999998e-13
RS_1013 NS_1013 0 1.1717534841017003e+02
RS_1014 NS_1014 0 1.1717534841017003e+02
GL_1013 0 NS_1013 NS_1014 0 1.5866517390841936e-01
GL_1014 0 NS_1014 NS_1013 0 -1.5866517390841936e-01
GS_1013_10 0 NS_1013 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1015/1016
CS_1015 NS_1015 0 9.9999999999999998e-13
CS_1016 NS_1016 0 9.9999999999999998e-13
RS_1015 NS_1015 0 8.8607873746940697e+01
RS_1016 NS_1016 0 8.8607873746940697e+01
GL_1015 0 NS_1015 NS_1016 0 1.5214737618207635e-01
GL_1016 0 NS_1016 NS_1015 0 -1.5214737618207635e-01
GS_1015_10 0 NS_1015 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1017/1018
CS_1017 NS_1017 0 9.9999999999999998e-13
CS_1018 NS_1018 0 9.9999999999999998e-13
RS_1017 NS_1017 0 1.1741456484283673e+02
RS_1018 NS_1018 0 1.1741456484283673e+02
GL_1017 0 NS_1017 NS_1018 0 1.4829748860889613e-01
GL_1018 0 NS_1018 NS_1017 0 -1.4829748860889613e-01
GS_1017_10 0 NS_1017 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1019/1020
CS_1019 NS_1019 0 9.9999999999999998e-13
CS_1020 NS_1020 0 9.9999999999999998e-13
RS_1019 NS_1019 0 1.3292289814180702e+02
RS_1020 NS_1020 0 1.3292289814180702e+02
GL_1019 0 NS_1019 NS_1020 0 1.4243056778188259e-01
GL_1020 0 NS_1020 NS_1019 0 -1.4243056778188259e-01
GS_1019_10 0 NS_1019 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1021/1022
CS_1021 NS_1021 0 9.9999999999999998e-13
CS_1022 NS_1022 0 9.9999999999999998e-13
RS_1021 NS_1021 0 1.2325134819531741e+02
RS_1022 NS_1022 0 1.2325134819531739e+02
GL_1021 0 NS_1021 NS_1022 0 1.3890785074828846e-01
GL_1022 0 NS_1022 NS_1021 0 -1.3890785074828846e-01
GS_1021_10 0 NS_1021 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1023/1024
CS_1023 NS_1023 0 9.9999999999999998e-13
CS_1024 NS_1024 0 9.9999999999999998e-13
RS_1023 NS_1023 0 9.1909059882883227e+01
RS_1024 NS_1024 0 9.1909059882883227e+01
GL_1023 0 NS_1023 NS_1024 0 1.3373879533989103e-01
GL_1024 0 NS_1024 NS_1023 0 -1.3373879533989103e-01
GS_1023_10 0 NS_1023 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1025/1026
CS_1025 NS_1025 0 9.9999999999999998e-13
CS_1026 NS_1026 0 9.9999999999999998e-13
RS_1025 NS_1025 0 1.2276824880349510e+02
RS_1026 NS_1026 0 1.2276824880349510e+02
GL_1025 0 NS_1025 NS_1026 0 1.2885409674522977e-01
GL_1026 0 NS_1026 NS_1025 0 -1.2885409674522977e-01
GS_1025_10 0 NS_1025 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1027/1028
CS_1027 NS_1027 0 9.9999999999999998e-13
CS_1028 NS_1028 0 9.9999999999999998e-13
RS_1027 NS_1027 0 1.1612442076026501e+02
RS_1028 NS_1028 0 1.1612442076026501e+02
GL_1027 0 NS_1027 NS_1028 0 1.2417838026896348e-01
GL_1028 0 NS_1028 NS_1027 0 -1.2417838026896348e-01
GS_1027_10 0 NS_1027 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1029/1030
CS_1029 NS_1029 0 9.9999999999999998e-13
CS_1030 NS_1030 0 9.9999999999999998e-13
RS_1029 NS_1029 0 1.2130204223875414e+02
RS_1030 NS_1030 0 1.2130204223875414e+02
GL_1029 0 NS_1029 NS_1030 0 1.1919240021970828e-01
GL_1030 0 NS_1030 NS_1029 0 -1.1919240021970828e-01
GS_1029_10 0 NS_1029 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1031/1032
CS_1031 NS_1031 0 9.9999999999999998e-13
CS_1032 NS_1032 0 9.9999999999999998e-13
RS_1031 NS_1031 0 9.3083309227260045e+01
RS_1032 NS_1032 0 9.3083309227260045e+01
GL_1031 0 NS_1031 NS_1032 0 1.1485268189050464e-01
GL_1032 0 NS_1032 NS_1031 0 -1.1485268189050464e-01
GS_1031_10 0 NS_1031 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1033/1034
CS_1033 NS_1033 0 9.9999999999999998e-13
CS_1034 NS_1034 0 9.9999999999999998e-13
RS_1033 NS_1033 0 1.2387094149263906e+02
RS_1034 NS_1034 0 1.2387094149263908e+02
GL_1033 0 NS_1033 NS_1034 0 1.0935451806229070e-01
GL_1034 0 NS_1034 NS_1033 0 -1.0935451806229070e-01
GS_1033_10 0 NS_1033 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1035/1036
CS_1035 NS_1035 0 9.9999999999999998e-13
CS_1036 NS_1036 0 9.9999999999999998e-13
RS_1035 NS_1035 0 1.1186020221520803e+02
RS_1036 NS_1036 0 1.1186020221520802e+02
GL_1035 0 NS_1035 NS_1036 0 1.0538242730807947e-01
GL_1036 0 NS_1036 NS_1035 0 -1.0538242730807947e-01
GS_1035_10 0 NS_1035 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1037/1038
CS_1037 NS_1037 0 9.9999999999999998e-13
CS_1038 NS_1038 0 9.9999999999999998e-13
RS_1037 NS_1037 0 1.2031265815570148e+02
RS_1038 NS_1038 0 1.2031265815570150e+02
GL_1037 0 NS_1037 NS_1038 0 9.9497602364102364e-02
GL_1038 0 NS_1038 NS_1037 0 -9.9497602364102364e-02
GS_1037_10 0 NS_1037 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1039/1040
CS_1039 NS_1039 0 9.9999999999999998e-13
CS_1040 NS_1040 0 9.9999999999999998e-13
RS_1039 NS_1039 0 9.6254518048655143e+01
RS_1040 NS_1040 0 9.6254518048655143e+01
GL_1039 0 NS_1039 NS_1040 0 9.5930770757699110e-02
GL_1040 0 NS_1040 NS_1039 0 -9.5930770757699110e-02
GS_1039_10 0 NS_1039 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1041/1042
CS_1041 NS_1041 0 9.9999999999999998e-13
CS_1042 NS_1042 0 9.9999999999999998e-13
RS_1041 NS_1041 0 1.2318640771018909e+02
RS_1042 NS_1042 0 1.2318640771018909e+02
GL_1041 0 NS_1041 NS_1042 0 8.9880619653662355e-02
GL_1042 0 NS_1042 NS_1041 0 -8.9880619653662355e-02
GS_1041_10 0 NS_1041 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1043/1044
CS_1043 NS_1043 0 9.9999999999999998e-13
CS_1044 NS_1044 0 9.9999999999999998e-13
RS_1043 NS_1043 0 1.1312630346155738e+02
RS_1044 NS_1044 0 1.1312630346155738e+02
GL_1043 0 NS_1043 NS_1044 0 8.6534434501560398e-02
GL_1044 0 NS_1044 NS_1043 0 -8.6534434501560398e-02
GS_1043_10 0 NS_1043 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1045/1046
CS_1045 NS_1045 0 9.9999999999999998e-13
CS_1046 NS_1046 0 9.9999999999999998e-13
RS_1045 NS_1045 0 1.1831504703984019e+02
RS_1046 NS_1046 0 1.1831504703984019e+02
GL_1045 0 NS_1045 NS_1046 0 7.9864296724202116e-02
GL_1046 0 NS_1046 NS_1045 0 -7.9864296724202116e-02
GS_1045_10 0 NS_1045 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1047/1048
CS_1047 NS_1047 0 9.9999999999999998e-13
CS_1048 NS_1048 0 9.9999999999999998e-13
RS_1047 NS_1047 0 1.0281987486447559e+02
RS_1048 NS_1048 0 1.0281987486447559e+02
GL_1047 0 NS_1047 NS_1048 0 7.6950339194481784e-02
GL_1048 0 NS_1048 NS_1047 0 -7.6950339194481784e-02
GS_1047_10 0 NS_1047 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1049/1050
CS_1049 NS_1049 0 9.9999999999999998e-13
CS_1050 NS_1050 0 9.9999999999999998e-13
RS_1049 NS_1049 0 1.2230186914382300e+02
RS_1050 NS_1050 0 1.2230186914382300e+02
GL_1049 0 NS_1049 NS_1050 0 7.0709298709435750e-02
GL_1050 0 NS_1050 NS_1049 0 -7.0709298709435750e-02
GS_1049_10 0 NS_1049 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1051/1052
CS_1051 NS_1051 0 9.9999999999999998e-13
CS_1052 NS_1052 0 9.9999999999999998e-13
RS_1051 NS_1051 0 1.2215699953322022e+02
RS_1052 NS_1052 0 1.2215699953322020e+02
GL_1051 0 NS_1051 NS_1052 0 6.7518227185671367e-02
GL_1052 0 NS_1052 NS_1051 0 -6.7518227185671367e-02
GS_1051_10 0 NS_1051 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1053/1054
CS_1053 NS_1053 0 9.9999999999999998e-13
CS_1054 NS_1054 0 9.9999999999999998e-13
RS_1053 NS_1053 0 3.4305564408226764e+03
RS_1054 NS_1054 0 3.4305564408226769e+03
GL_1053 0 NS_1053 NS_1054 0 5.4396471187208063e-02
GL_1054 0 NS_1054 NS_1053 0 -5.4396471187208063e-02
GS_1053_10 0 NS_1053 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1055/1056
CS_1055 NS_1055 0 9.9999999999999998e-13
CS_1056 NS_1056 0 9.9999999999999998e-13
RS_1055 NS_1055 0 1.1894859826238778e+02
RS_1056 NS_1056 0 1.1894859826238779e+02
GL_1055 0 NS_1055 NS_1056 0 6.0591569497719031e-02
GL_1056 0 NS_1056 NS_1055 0 -6.0591569497719031e-02
GS_1055_10 0 NS_1055 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1057/1058
CS_1057 NS_1057 0 9.9999999999999998e-13
CS_1058 NS_1058 0 9.9999999999999998e-13
RS_1057 NS_1057 0 1.3537641711503298e+02
RS_1058 NS_1058 0 1.3537641711503298e+02
GL_1057 0 NS_1057 NS_1058 0 5.1190778164089609e-02
GL_1058 0 NS_1058 NS_1057 0 -5.1190778164089609e-02
GS_1057_10 0 NS_1057 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1059/1060
CS_1059 NS_1059 0 9.9999999999999998e-13
CS_1060 NS_1060 0 9.9999999999999998e-13
RS_1059 NS_1059 0 1.3105452427659637e+02
RS_1060 NS_1060 0 1.3105452427659637e+02
GL_1059 0 NS_1059 NS_1060 0 4.7418984574880592e-02
GL_1060 0 NS_1060 NS_1059 0 -4.7418984574880592e-02
GS_1059_10 0 NS_1059 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1061/1062
CS_1061 NS_1061 0 9.9999999999999998e-13
CS_1062 NS_1062 0 9.9999999999999998e-13
RS_1061 NS_1061 0 1.2170234397098790e+02
RS_1062 NS_1062 0 1.2170234397098790e+02
GL_1061 0 NS_1061 NS_1062 0 4.0778813929127578e-02
GL_1062 0 NS_1062 NS_1061 0 -4.0778813929127578e-02
GS_1061_10 0 NS_1061 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1063/1064
CS_1063 NS_1063 0 9.9999999999999998e-13
CS_1064 NS_1064 0 9.9999999999999998e-13
RS_1063 NS_1063 0 1.1550510326517782e+02
RS_1064 NS_1064 0 1.1550510326517782e+02
GL_1063 0 NS_1063 NS_1064 0 5.7236026076957713e-02
GL_1064 0 NS_1064 NS_1063 0 -5.7236026076957713e-02
GS_1063_10 0 NS_1063 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1065/1066
CS_1065 NS_1065 0 9.9999999999999998e-13
CS_1066 NS_1066 0 9.9999999999999998e-13
RS_1065 NS_1065 0 6.2039157456337159e+02
RS_1066 NS_1066 0 6.2039157456337159e+02
GL_1065 0 NS_1065 NS_1066 0 1.9354364738401211e-02
GL_1066 0 NS_1066 NS_1065 0 -1.9354364738401211e-02
GS_1065_10 0 NS_1065 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1067/1068
CS_1067 NS_1067 0 9.9999999999999998e-13
CS_1068 NS_1068 0 9.9999999999999998e-13
RS_1067 NS_1067 0 1.1050313240441588e+02
RS_1068 NS_1068 0 1.1050313240441587e+02
GL_1067 0 NS_1067 NS_1068 0 1.6472588786558075e-02
GL_1068 0 NS_1068 NS_1067 0 -1.6472588786558075e-02
GS_1067_10 0 NS_1067 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1069/1070
CS_1069 NS_1069 0 9.9999999999999998e-13
CS_1070 NS_1070 0 9.9999999999999998e-13
RS_1069 NS_1069 0 1.2869119986945731e+02
RS_1070 NS_1070 0 1.2869119986945731e+02
GL_1069 0 NS_1069 NS_1070 0 2.0888592987579706e-02
GL_1070 0 NS_1070 NS_1069 0 -2.0888592987579706e-02
GS_1069_10 0 NS_1069 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1071/1072
CS_1071 NS_1071 0 9.9999999999999998e-13
CS_1072 NS_1072 0 9.9999999999999998e-13
RS_1071 NS_1071 0 1.4314560950270646e+02
RS_1072 NS_1072 0 1.4314560950270646e+02
GL_1071 0 NS_1071 NS_1072 0 9.7871236580563716e-03
GL_1072 0 NS_1072 NS_1071 0 -9.7871236580563716e-03
GS_1071_10 0 NS_1071 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1073/1074
CS_1073 NS_1073 0 9.9999999999999998e-13
CS_1074 NS_1074 0 9.9999999999999998e-13
RS_1073 NS_1073 0 1.1863004336811436e+02
RS_1074 NS_1074 0 1.1863004336811436e+02
GL_1073 0 NS_1073 NS_1074 0 3.7627463994326378e-02
GL_1074 0 NS_1074 NS_1073 0 -3.7627463994326378e-02
GS_1073_10 0 NS_1073 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1075/1076
CS_1075 NS_1075 0 9.9999999999999998e-13
CS_1076 NS_1076 0 9.9999999999999998e-13
RS_1075 NS_1075 0 1.2686172273444870e+02
RS_1076 NS_1076 0 1.2686172273444869e+02
GL_1075 0 NS_1075 NS_1076 0 3.1975218188091938e-02
GL_1076 0 NS_1076 NS_1075 0 -3.1975218188091938e-02
GS_1075_10 0 NS_1075 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1077/1078
CS_1077 NS_1077 0 9.9999999999999998e-13
CS_1078 NS_1078 0 9.9999999999999998e-13
RS_1077 NS_1077 0 1.3141621772977734e+02
RS_1078 NS_1078 0 1.3141621772977737e+02
GL_1077 0 NS_1077 NS_1078 0 2.8228381102665165e-02
GL_1078 0 NS_1078 NS_1077 0 -2.8228381102665165e-02
GS_1077_10 0 NS_1077 NA_10 0 4.7428518688027549e-01
*
* Complex pair n. 1079/1080
CS_1079 NS_1079 0 9.9999999999999998e-13
CS_1080 NS_1080 0 9.9999999999999998e-13
RS_1079 NS_1079 0 1.2452833644614726e+02
RS_1080 NS_1080 0 1.2452833644614726e+02
GL_1079 0 NS_1079 NS_1080 0 2.1457325426059259e-03
GL_1080 0 NS_1080 NS_1079 0 -2.1457325426059259e-03
GS_1079_10 0 NS_1079 NA_10 0 4.7428518688027549e-01
*
* Real pole n. 1081
CS_1081 NS_1081 0 9.9999999999999998e-13
RS_1081 NS_1081 0 3.8329546824379270e+00
GS_1081_11 0 NS_1081 NA_11 0 4.7428518688027549e-01
*
* Real pole n. 1082
CS_1082 NS_1082 0 9.9999999999999998e-13
RS_1082 NS_1082 0 1.0843846705160875e+04
GS_1082_11 0 NS_1082 NA_11 0 4.7428518688027549e-01
*
* Real pole n. 1083
CS_1083 NS_1083 0 9.9999999999999998e-13
RS_1083 NS_1083 0 3.3457029134706481e+03
GS_1083_11 0 NS_1083 NA_11 0 4.7428518688027549e-01
*
* Real pole n. 1084
CS_1084 NS_1084 0 9.9999999999999998e-13
RS_1084 NS_1084 0 5.4313394337993634e+02
GS_1084_11 0 NS_1084 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1085/1086
CS_1085 NS_1085 0 9.9999999999999998e-13
CS_1086 NS_1086 0 9.9999999999999998e-13
RS_1085 NS_1085 0 2.0342898045173075e+02
RS_1086 NS_1086 0 2.0342898045173075e+02
GL_1085 0 NS_1085 NS_1086 0 2.5883098202682536e-01
GL_1086 0 NS_1086 NS_1085 0 -2.5883098202682536e-01
GS_1085_11 0 NS_1085 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1087/1088
CS_1087 NS_1087 0 9.9999999999999998e-13
CS_1088 NS_1088 0 9.9999999999999998e-13
RS_1087 NS_1087 0 1.2739936959261519e+02
RS_1088 NS_1088 0 1.2739936959261519e+02
GL_1087 0 NS_1087 NS_1088 0 2.5122204303896745e-01
GL_1088 0 NS_1088 NS_1087 0 -2.5122204303896745e-01
GS_1087_11 0 NS_1087 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1089/1090
CS_1089 NS_1089 0 9.9999999999999998e-13
CS_1090 NS_1090 0 9.9999999999999998e-13
RS_1089 NS_1089 0 1.1105129555360161e+02
RS_1090 NS_1090 0 1.1105129555360161e+02
GL_1089 0 NS_1089 NS_1090 0 2.4643422119526687e-01
GL_1090 0 NS_1090 NS_1089 0 -2.4643422119526687e-01
GS_1089_11 0 NS_1089 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1091/1092
CS_1091 NS_1091 0 9.9999999999999998e-13
CS_1092 NS_1092 0 9.9999999999999998e-13
RS_1091 NS_1091 0 1.0856580972218713e+02
RS_1092 NS_1092 0 1.0856580972218713e+02
GL_1091 0 NS_1091 NS_1092 0 2.4007148694878275e-01
GL_1092 0 NS_1092 NS_1091 0 -2.4007148694878275e-01
GS_1091_11 0 NS_1091 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1093/1094
CS_1093 NS_1093 0 9.9999999999999998e-13
CS_1094 NS_1094 0 9.9999999999999998e-13
RS_1093 NS_1093 0 1.0135860176893434e+02
RS_1094 NS_1094 0 1.0135860176893435e+02
GL_1093 0 NS_1093 NS_1094 0 2.3570758371916220e-01
GL_1094 0 NS_1094 NS_1093 0 -2.3570758371916220e-01
GS_1093_11 0 NS_1093 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1095/1096
CS_1095 NS_1095 0 9.9999999999999998e-13
CS_1096 NS_1096 0 9.9999999999999998e-13
RS_1095 NS_1095 0 1.2858526276753685e+02
RS_1096 NS_1096 0 1.2858526276753685e+02
GL_1095 0 NS_1095 NS_1096 0 2.2966634995600790e-01
GL_1096 0 NS_1096 NS_1095 0 -2.2966634995600790e-01
GS_1095_11 0 NS_1095 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1097/1098
CS_1097 NS_1097 0 9.9999999999999998e-13
CS_1098 NS_1098 0 9.9999999999999998e-13
RS_1097 NS_1097 0 1.1773437593549667e+02
RS_1098 NS_1098 0 1.1773437593549667e+02
GL_1097 0 NS_1097 NS_1098 0 2.2732609444056490e-01
GL_1098 0 NS_1098 NS_1097 0 -2.2732609444056490e-01
GS_1097_11 0 NS_1097 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1099/1100
CS_1099 NS_1099 0 9.9999999999999998e-13
CS_1100 NS_1100 0 9.9999999999999998e-13
RS_1099 NS_1099 0 9.8170265044265946e+01
RS_1100 NS_1100 0 9.8170265044265932e+01
GL_1099 0 NS_1099 NS_1100 0 2.2031598117475365e-01
GL_1100 0 NS_1100 NS_1099 0 -2.2031598117475365e-01
GS_1099_11 0 NS_1099 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1101/1102
CS_1101 NS_1101 0 9.9999999999999998e-13
CS_1102 NS_1102 0 9.9999999999999998e-13
RS_1101 NS_1101 0 9.5355901421613709e+01
RS_1102 NS_1102 0 9.5355901421613694e+01
GL_1101 0 NS_1101 NS_1102 0 2.1739680820836188e-01
GL_1102 0 NS_1102 NS_1101 0 -2.1739680820836188e-01
GS_1101_11 0 NS_1101 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1103/1104
CS_1103 NS_1103 0 9.9999999999999998e-13
CS_1104 NS_1104 0 9.9999999999999998e-13
RS_1103 NS_1103 0 1.0859722031634941e+02
RS_1104 NS_1104 0 1.0859722031634941e+02
GL_1103 0 NS_1103 NS_1104 0 2.0887403840929383e-01
GL_1104 0 NS_1104 NS_1103 0 -2.0887403840929383e-01
GS_1103_11 0 NS_1103 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1105/1106
CS_1105 NS_1105 0 9.9999999999999998e-13
CS_1106 NS_1106 0 9.9999999999999998e-13
RS_1105 NS_1105 0 7.7959989808728068e+01
RS_1106 NS_1106 0 7.7959989808728054e+01
GL_1105 0 NS_1105 NS_1106 0 2.0447808896343445e-01
GL_1106 0 NS_1106 NS_1105 0 -2.0447808896343445e-01
GS_1105_11 0 NS_1105 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1107/1108
CS_1107 NS_1107 0 9.9999999999999998e-13
CS_1108 NS_1108 0 9.9999999999999998e-13
RS_1107 NS_1107 0 1.1088851678406323e+02
RS_1108 NS_1108 0 1.1088851678406321e+02
GL_1107 0 NS_1107 NS_1108 0 1.9843399276071924e-01
GL_1108 0 NS_1108 NS_1107 0 -1.9843399276071924e-01
GS_1107_11 0 NS_1107 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1109/1110
CS_1109 NS_1109 0 9.9999999999999998e-13
CS_1110 NS_1110 0 9.9999999999999998e-13
RS_1109 NS_1109 0 8.1179760966262847e+01
RS_1110 NS_1110 0 8.1179760966262847e+01
GL_1109 0 NS_1109 NS_1110 0 1.8978022990658949e-01
GL_1110 0 NS_1110 NS_1109 0 -1.8978022990658949e-01
GS_1109_11 0 NS_1109 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1111/1112
CS_1111 NS_1111 0 9.9999999999999998e-13
CS_1112 NS_1112 0 9.9999999999999998e-13
RS_1111 NS_1111 0 1.0523970815054612e+02
RS_1112 NS_1112 0 1.0523970815054612e+02
GL_1111 0 NS_1111 NS_1112 0 1.8836779078363333e-01
GL_1112 0 NS_1112 NS_1111 0 -1.8836779078363333e-01
GS_1111_11 0 NS_1111 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1113/1114
CS_1113 NS_1113 0 9.9999999999999998e-13
CS_1114 NS_1114 0 9.9999999999999998e-13
RS_1113 NS_1113 0 1.1208834663822537e+02
RS_1114 NS_1114 0 1.1208834663822537e+02
GL_1113 0 NS_1113 NS_1114 0 1.7925451755127267e-01
GL_1114 0 NS_1114 NS_1113 0 -1.7925451755127267e-01
GS_1113_11 0 NS_1113 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1115/1116
CS_1115 NS_1115 0 9.9999999999999998e-13
CS_1116 NS_1116 0 9.9999999999999998e-13
RS_1115 NS_1115 0 9.2475617668062213e+01
RS_1116 NS_1116 0 9.2475617668062199e+01
GL_1115 0 NS_1115 NS_1116 0 1.7507216970358189e-01
GL_1116 0 NS_1116 NS_1115 0 -1.7507216970358189e-01
GS_1115_11 0 NS_1115 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1117/1118
CS_1117 NS_1117 0 9.9999999999999998e-13
CS_1118 NS_1118 0 9.9999999999999998e-13
RS_1117 NS_1117 0 1.1555782965375326e+02
RS_1118 NS_1118 0 1.1555782965375326e+02
GL_1117 0 NS_1117 NS_1118 0 1.6918904340923188e-01
GL_1118 0 NS_1118 NS_1117 0 -1.6918904340923188e-01
GS_1117_11 0 NS_1117 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1119/1120
CS_1119 NS_1119 0 9.9999999999999998e-13
CS_1120 NS_1120 0 9.9999999999999998e-13
RS_1119 NS_1119 0 9.6856782813111039e+01
RS_1120 NS_1120 0 9.6856782813111039e+01
GL_1119 0 NS_1119 NS_1120 0 1.6488898173469207e-01
GL_1120 0 NS_1120 NS_1119 0 -1.6488898173469207e-01
GS_1119_11 0 NS_1119 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1121/1122
CS_1121 NS_1121 0 9.9999999999999998e-13
CS_1122 NS_1122 0 9.9999999999999998e-13
RS_1121 NS_1121 0 1.1717534841017003e+02
RS_1122 NS_1122 0 1.1717534841017003e+02
GL_1121 0 NS_1121 NS_1122 0 1.5866517390841936e-01
GL_1122 0 NS_1122 NS_1121 0 -1.5866517390841936e-01
GS_1121_11 0 NS_1121 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1123/1124
CS_1123 NS_1123 0 9.9999999999999998e-13
CS_1124 NS_1124 0 9.9999999999999998e-13
RS_1123 NS_1123 0 8.8607873746940697e+01
RS_1124 NS_1124 0 8.8607873746940697e+01
GL_1123 0 NS_1123 NS_1124 0 1.5214737618207635e-01
GL_1124 0 NS_1124 NS_1123 0 -1.5214737618207635e-01
GS_1123_11 0 NS_1123 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1125/1126
CS_1125 NS_1125 0 9.9999999999999998e-13
CS_1126 NS_1126 0 9.9999999999999998e-13
RS_1125 NS_1125 0 1.1741456484283673e+02
RS_1126 NS_1126 0 1.1741456484283673e+02
GL_1125 0 NS_1125 NS_1126 0 1.4829748860889613e-01
GL_1126 0 NS_1126 NS_1125 0 -1.4829748860889613e-01
GS_1125_11 0 NS_1125 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1127/1128
CS_1127 NS_1127 0 9.9999999999999998e-13
CS_1128 NS_1128 0 9.9999999999999998e-13
RS_1127 NS_1127 0 1.3292289814180702e+02
RS_1128 NS_1128 0 1.3292289814180702e+02
GL_1127 0 NS_1127 NS_1128 0 1.4243056778188259e-01
GL_1128 0 NS_1128 NS_1127 0 -1.4243056778188259e-01
GS_1127_11 0 NS_1127 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1129/1130
CS_1129 NS_1129 0 9.9999999999999998e-13
CS_1130 NS_1130 0 9.9999999999999998e-13
RS_1129 NS_1129 0 1.2325134819531741e+02
RS_1130 NS_1130 0 1.2325134819531739e+02
GL_1129 0 NS_1129 NS_1130 0 1.3890785074828846e-01
GL_1130 0 NS_1130 NS_1129 0 -1.3890785074828846e-01
GS_1129_11 0 NS_1129 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1131/1132
CS_1131 NS_1131 0 9.9999999999999998e-13
CS_1132 NS_1132 0 9.9999999999999998e-13
RS_1131 NS_1131 0 9.1909059882883227e+01
RS_1132 NS_1132 0 9.1909059882883227e+01
GL_1131 0 NS_1131 NS_1132 0 1.3373879533989103e-01
GL_1132 0 NS_1132 NS_1131 0 -1.3373879533989103e-01
GS_1131_11 0 NS_1131 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1133/1134
CS_1133 NS_1133 0 9.9999999999999998e-13
CS_1134 NS_1134 0 9.9999999999999998e-13
RS_1133 NS_1133 0 1.2276824880349510e+02
RS_1134 NS_1134 0 1.2276824880349510e+02
GL_1133 0 NS_1133 NS_1134 0 1.2885409674522977e-01
GL_1134 0 NS_1134 NS_1133 0 -1.2885409674522977e-01
GS_1133_11 0 NS_1133 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1135/1136
CS_1135 NS_1135 0 9.9999999999999998e-13
CS_1136 NS_1136 0 9.9999999999999998e-13
RS_1135 NS_1135 0 1.1612442076026501e+02
RS_1136 NS_1136 0 1.1612442076026501e+02
GL_1135 0 NS_1135 NS_1136 0 1.2417838026896348e-01
GL_1136 0 NS_1136 NS_1135 0 -1.2417838026896348e-01
GS_1135_11 0 NS_1135 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1137/1138
CS_1137 NS_1137 0 9.9999999999999998e-13
CS_1138 NS_1138 0 9.9999999999999998e-13
RS_1137 NS_1137 0 1.2130204223875414e+02
RS_1138 NS_1138 0 1.2130204223875414e+02
GL_1137 0 NS_1137 NS_1138 0 1.1919240021970828e-01
GL_1138 0 NS_1138 NS_1137 0 -1.1919240021970828e-01
GS_1137_11 0 NS_1137 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1139/1140
CS_1139 NS_1139 0 9.9999999999999998e-13
CS_1140 NS_1140 0 9.9999999999999998e-13
RS_1139 NS_1139 0 9.3083309227260045e+01
RS_1140 NS_1140 0 9.3083309227260045e+01
GL_1139 0 NS_1139 NS_1140 0 1.1485268189050464e-01
GL_1140 0 NS_1140 NS_1139 0 -1.1485268189050464e-01
GS_1139_11 0 NS_1139 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1141/1142
CS_1141 NS_1141 0 9.9999999999999998e-13
CS_1142 NS_1142 0 9.9999999999999998e-13
RS_1141 NS_1141 0 1.2387094149263906e+02
RS_1142 NS_1142 0 1.2387094149263908e+02
GL_1141 0 NS_1141 NS_1142 0 1.0935451806229070e-01
GL_1142 0 NS_1142 NS_1141 0 -1.0935451806229070e-01
GS_1141_11 0 NS_1141 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1143/1144
CS_1143 NS_1143 0 9.9999999999999998e-13
CS_1144 NS_1144 0 9.9999999999999998e-13
RS_1143 NS_1143 0 1.1186020221520803e+02
RS_1144 NS_1144 0 1.1186020221520802e+02
GL_1143 0 NS_1143 NS_1144 0 1.0538242730807947e-01
GL_1144 0 NS_1144 NS_1143 0 -1.0538242730807947e-01
GS_1143_11 0 NS_1143 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1145/1146
CS_1145 NS_1145 0 9.9999999999999998e-13
CS_1146 NS_1146 0 9.9999999999999998e-13
RS_1145 NS_1145 0 1.2031265815570148e+02
RS_1146 NS_1146 0 1.2031265815570150e+02
GL_1145 0 NS_1145 NS_1146 0 9.9497602364102364e-02
GL_1146 0 NS_1146 NS_1145 0 -9.9497602364102364e-02
GS_1145_11 0 NS_1145 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1147/1148
CS_1147 NS_1147 0 9.9999999999999998e-13
CS_1148 NS_1148 0 9.9999999999999998e-13
RS_1147 NS_1147 0 9.6254518048655143e+01
RS_1148 NS_1148 0 9.6254518048655143e+01
GL_1147 0 NS_1147 NS_1148 0 9.5930770757699110e-02
GL_1148 0 NS_1148 NS_1147 0 -9.5930770757699110e-02
GS_1147_11 0 NS_1147 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1149/1150
CS_1149 NS_1149 0 9.9999999999999998e-13
CS_1150 NS_1150 0 9.9999999999999998e-13
RS_1149 NS_1149 0 1.2318640771018909e+02
RS_1150 NS_1150 0 1.2318640771018909e+02
GL_1149 0 NS_1149 NS_1150 0 8.9880619653662355e-02
GL_1150 0 NS_1150 NS_1149 0 -8.9880619653662355e-02
GS_1149_11 0 NS_1149 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1151/1152
CS_1151 NS_1151 0 9.9999999999999998e-13
CS_1152 NS_1152 0 9.9999999999999998e-13
RS_1151 NS_1151 0 1.1312630346155738e+02
RS_1152 NS_1152 0 1.1312630346155738e+02
GL_1151 0 NS_1151 NS_1152 0 8.6534434501560398e-02
GL_1152 0 NS_1152 NS_1151 0 -8.6534434501560398e-02
GS_1151_11 0 NS_1151 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1153/1154
CS_1153 NS_1153 0 9.9999999999999998e-13
CS_1154 NS_1154 0 9.9999999999999998e-13
RS_1153 NS_1153 0 1.1831504703984019e+02
RS_1154 NS_1154 0 1.1831504703984019e+02
GL_1153 0 NS_1153 NS_1154 0 7.9864296724202116e-02
GL_1154 0 NS_1154 NS_1153 0 -7.9864296724202116e-02
GS_1153_11 0 NS_1153 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1155/1156
CS_1155 NS_1155 0 9.9999999999999998e-13
CS_1156 NS_1156 0 9.9999999999999998e-13
RS_1155 NS_1155 0 1.0281987486447559e+02
RS_1156 NS_1156 0 1.0281987486447559e+02
GL_1155 0 NS_1155 NS_1156 0 7.6950339194481784e-02
GL_1156 0 NS_1156 NS_1155 0 -7.6950339194481784e-02
GS_1155_11 0 NS_1155 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1157/1158
CS_1157 NS_1157 0 9.9999999999999998e-13
CS_1158 NS_1158 0 9.9999999999999998e-13
RS_1157 NS_1157 0 1.2230186914382300e+02
RS_1158 NS_1158 0 1.2230186914382300e+02
GL_1157 0 NS_1157 NS_1158 0 7.0709298709435750e-02
GL_1158 0 NS_1158 NS_1157 0 -7.0709298709435750e-02
GS_1157_11 0 NS_1157 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1159/1160
CS_1159 NS_1159 0 9.9999999999999998e-13
CS_1160 NS_1160 0 9.9999999999999998e-13
RS_1159 NS_1159 0 1.2215699953322022e+02
RS_1160 NS_1160 0 1.2215699953322020e+02
GL_1159 0 NS_1159 NS_1160 0 6.7518227185671367e-02
GL_1160 0 NS_1160 NS_1159 0 -6.7518227185671367e-02
GS_1159_11 0 NS_1159 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1161/1162
CS_1161 NS_1161 0 9.9999999999999998e-13
CS_1162 NS_1162 0 9.9999999999999998e-13
RS_1161 NS_1161 0 3.4305564408226764e+03
RS_1162 NS_1162 0 3.4305564408226769e+03
GL_1161 0 NS_1161 NS_1162 0 5.4396471187208063e-02
GL_1162 0 NS_1162 NS_1161 0 -5.4396471187208063e-02
GS_1161_11 0 NS_1161 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1163/1164
CS_1163 NS_1163 0 9.9999999999999998e-13
CS_1164 NS_1164 0 9.9999999999999998e-13
RS_1163 NS_1163 0 1.1894859826238778e+02
RS_1164 NS_1164 0 1.1894859826238779e+02
GL_1163 0 NS_1163 NS_1164 0 6.0591569497719031e-02
GL_1164 0 NS_1164 NS_1163 0 -6.0591569497719031e-02
GS_1163_11 0 NS_1163 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1165/1166
CS_1165 NS_1165 0 9.9999999999999998e-13
CS_1166 NS_1166 0 9.9999999999999998e-13
RS_1165 NS_1165 0 1.3537641711503298e+02
RS_1166 NS_1166 0 1.3537641711503298e+02
GL_1165 0 NS_1165 NS_1166 0 5.1190778164089609e-02
GL_1166 0 NS_1166 NS_1165 0 -5.1190778164089609e-02
GS_1165_11 0 NS_1165 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1167/1168
CS_1167 NS_1167 0 9.9999999999999998e-13
CS_1168 NS_1168 0 9.9999999999999998e-13
RS_1167 NS_1167 0 1.3105452427659637e+02
RS_1168 NS_1168 0 1.3105452427659637e+02
GL_1167 0 NS_1167 NS_1168 0 4.7418984574880592e-02
GL_1168 0 NS_1168 NS_1167 0 -4.7418984574880592e-02
GS_1167_11 0 NS_1167 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1169/1170
CS_1169 NS_1169 0 9.9999999999999998e-13
CS_1170 NS_1170 0 9.9999999999999998e-13
RS_1169 NS_1169 0 1.2170234397098790e+02
RS_1170 NS_1170 0 1.2170234397098790e+02
GL_1169 0 NS_1169 NS_1170 0 4.0778813929127578e-02
GL_1170 0 NS_1170 NS_1169 0 -4.0778813929127578e-02
GS_1169_11 0 NS_1169 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1171/1172
CS_1171 NS_1171 0 9.9999999999999998e-13
CS_1172 NS_1172 0 9.9999999999999998e-13
RS_1171 NS_1171 0 1.1550510326517782e+02
RS_1172 NS_1172 0 1.1550510326517782e+02
GL_1171 0 NS_1171 NS_1172 0 5.7236026076957713e-02
GL_1172 0 NS_1172 NS_1171 0 -5.7236026076957713e-02
GS_1171_11 0 NS_1171 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1173/1174
CS_1173 NS_1173 0 9.9999999999999998e-13
CS_1174 NS_1174 0 9.9999999999999998e-13
RS_1173 NS_1173 0 6.2039157456337159e+02
RS_1174 NS_1174 0 6.2039157456337159e+02
GL_1173 0 NS_1173 NS_1174 0 1.9354364738401211e-02
GL_1174 0 NS_1174 NS_1173 0 -1.9354364738401211e-02
GS_1173_11 0 NS_1173 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1175/1176
CS_1175 NS_1175 0 9.9999999999999998e-13
CS_1176 NS_1176 0 9.9999999999999998e-13
RS_1175 NS_1175 0 1.1050313240441588e+02
RS_1176 NS_1176 0 1.1050313240441587e+02
GL_1175 0 NS_1175 NS_1176 0 1.6472588786558075e-02
GL_1176 0 NS_1176 NS_1175 0 -1.6472588786558075e-02
GS_1175_11 0 NS_1175 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1177/1178
CS_1177 NS_1177 0 9.9999999999999998e-13
CS_1178 NS_1178 0 9.9999999999999998e-13
RS_1177 NS_1177 0 1.2869119986945731e+02
RS_1178 NS_1178 0 1.2869119986945731e+02
GL_1177 0 NS_1177 NS_1178 0 2.0888592987579706e-02
GL_1178 0 NS_1178 NS_1177 0 -2.0888592987579706e-02
GS_1177_11 0 NS_1177 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1179/1180
CS_1179 NS_1179 0 9.9999999999999998e-13
CS_1180 NS_1180 0 9.9999999999999998e-13
RS_1179 NS_1179 0 1.4314560950270646e+02
RS_1180 NS_1180 0 1.4314560950270646e+02
GL_1179 0 NS_1179 NS_1180 0 9.7871236580563716e-03
GL_1180 0 NS_1180 NS_1179 0 -9.7871236580563716e-03
GS_1179_11 0 NS_1179 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1181/1182
CS_1181 NS_1181 0 9.9999999999999998e-13
CS_1182 NS_1182 0 9.9999999999999998e-13
RS_1181 NS_1181 0 1.1863004336811436e+02
RS_1182 NS_1182 0 1.1863004336811436e+02
GL_1181 0 NS_1181 NS_1182 0 3.7627463994326378e-02
GL_1182 0 NS_1182 NS_1181 0 -3.7627463994326378e-02
GS_1181_11 0 NS_1181 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1183/1184
CS_1183 NS_1183 0 9.9999999999999998e-13
CS_1184 NS_1184 0 9.9999999999999998e-13
RS_1183 NS_1183 0 1.2686172273444870e+02
RS_1184 NS_1184 0 1.2686172273444869e+02
GL_1183 0 NS_1183 NS_1184 0 3.1975218188091938e-02
GL_1184 0 NS_1184 NS_1183 0 -3.1975218188091938e-02
GS_1183_11 0 NS_1183 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1185/1186
CS_1185 NS_1185 0 9.9999999999999998e-13
CS_1186 NS_1186 0 9.9999999999999998e-13
RS_1185 NS_1185 0 1.3141621772977734e+02
RS_1186 NS_1186 0 1.3141621772977737e+02
GL_1185 0 NS_1185 NS_1186 0 2.8228381102665165e-02
GL_1186 0 NS_1186 NS_1185 0 -2.8228381102665165e-02
GS_1185_11 0 NS_1185 NA_11 0 4.7428518688027549e-01
*
* Complex pair n. 1187/1188
CS_1187 NS_1187 0 9.9999999999999998e-13
CS_1188 NS_1188 0 9.9999999999999998e-13
RS_1187 NS_1187 0 1.2452833644614726e+02
RS_1188 NS_1188 0 1.2452833644614726e+02
GL_1187 0 NS_1187 NS_1188 0 2.1457325426059259e-03
GL_1188 0 NS_1188 NS_1187 0 -2.1457325426059259e-03
GS_1187_11 0 NS_1187 NA_11 0 4.7428518688027549e-01
*
* Real pole n. 1189
CS_1189 NS_1189 0 9.9999999999999998e-13
RS_1189 NS_1189 0 3.8329546824379270e+00
GS_1189_12 0 NS_1189 NA_12 0 4.7428518688027549e-01
*
* Real pole n. 1190
CS_1190 NS_1190 0 9.9999999999999998e-13
RS_1190 NS_1190 0 1.0843846705160875e+04
GS_1190_12 0 NS_1190 NA_12 0 4.7428518688027549e-01
*
* Real pole n. 1191
CS_1191 NS_1191 0 9.9999999999999998e-13
RS_1191 NS_1191 0 3.3457029134706481e+03
GS_1191_12 0 NS_1191 NA_12 0 4.7428518688027549e-01
*
* Real pole n. 1192
CS_1192 NS_1192 0 9.9999999999999998e-13
RS_1192 NS_1192 0 5.4313394337993634e+02
GS_1192_12 0 NS_1192 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1193/1194
CS_1193 NS_1193 0 9.9999999999999998e-13
CS_1194 NS_1194 0 9.9999999999999998e-13
RS_1193 NS_1193 0 2.0342898045173075e+02
RS_1194 NS_1194 0 2.0342898045173075e+02
GL_1193 0 NS_1193 NS_1194 0 2.5883098202682536e-01
GL_1194 0 NS_1194 NS_1193 0 -2.5883098202682536e-01
GS_1193_12 0 NS_1193 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1195/1196
CS_1195 NS_1195 0 9.9999999999999998e-13
CS_1196 NS_1196 0 9.9999999999999998e-13
RS_1195 NS_1195 0 1.2739936959261519e+02
RS_1196 NS_1196 0 1.2739936959261519e+02
GL_1195 0 NS_1195 NS_1196 0 2.5122204303896745e-01
GL_1196 0 NS_1196 NS_1195 0 -2.5122204303896745e-01
GS_1195_12 0 NS_1195 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1197/1198
CS_1197 NS_1197 0 9.9999999999999998e-13
CS_1198 NS_1198 0 9.9999999999999998e-13
RS_1197 NS_1197 0 1.1105129555360161e+02
RS_1198 NS_1198 0 1.1105129555360161e+02
GL_1197 0 NS_1197 NS_1198 0 2.4643422119526687e-01
GL_1198 0 NS_1198 NS_1197 0 -2.4643422119526687e-01
GS_1197_12 0 NS_1197 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1199/1200
CS_1199 NS_1199 0 9.9999999999999998e-13
CS_1200 NS_1200 0 9.9999999999999998e-13
RS_1199 NS_1199 0 1.0856580972218713e+02
RS_1200 NS_1200 0 1.0856580972218713e+02
GL_1199 0 NS_1199 NS_1200 0 2.4007148694878275e-01
GL_1200 0 NS_1200 NS_1199 0 -2.4007148694878275e-01
GS_1199_12 0 NS_1199 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1201/1202
CS_1201 NS_1201 0 9.9999999999999998e-13
CS_1202 NS_1202 0 9.9999999999999998e-13
RS_1201 NS_1201 0 1.0135860176893434e+02
RS_1202 NS_1202 0 1.0135860176893435e+02
GL_1201 0 NS_1201 NS_1202 0 2.3570758371916220e-01
GL_1202 0 NS_1202 NS_1201 0 -2.3570758371916220e-01
GS_1201_12 0 NS_1201 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1203/1204
CS_1203 NS_1203 0 9.9999999999999998e-13
CS_1204 NS_1204 0 9.9999999999999998e-13
RS_1203 NS_1203 0 1.2858526276753685e+02
RS_1204 NS_1204 0 1.2858526276753685e+02
GL_1203 0 NS_1203 NS_1204 0 2.2966634995600790e-01
GL_1204 0 NS_1204 NS_1203 0 -2.2966634995600790e-01
GS_1203_12 0 NS_1203 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1205/1206
CS_1205 NS_1205 0 9.9999999999999998e-13
CS_1206 NS_1206 0 9.9999999999999998e-13
RS_1205 NS_1205 0 1.1773437593549667e+02
RS_1206 NS_1206 0 1.1773437593549667e+02
GL_1205 0 NS_1205 NS_1206 0 2.2732609444056490e-01
GL_1206 0 NS_1206 NS_1205 0 -2.2732609444056490e-01
GS_1205_12 0 NS_1205 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1207/1208
CS_1207 NS_1207 0 9.9999999999999998e-13
CS_1208 NS_1208 0 9.9999999999999998e-13
RS_1207 NS_1207 0 9.8170265044265946e+01
RS_1208 NS_1208 0 9.8170265044265932e+01
GL_1207 0 NS_1207 NS_1208 0 2.2031598117475365e-01
GL_1208 0 NS_1208 NS_1207 0 -2.2031598117475365e-01
GS_1207_12 0 NS_1207 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1209/1210
CS_1209 NS_1209 0 9.9999999999999998e-13
CS_1210 NS_1210 0 9.9999999999999998e-13
RS_1209 NS_1209 0 9.5355901421613709e+01
RS_1210 NS_1210 0 9.5355901421613694e+01
GL_1209 0 NS_1209 NS_1210 0 2.1739680820836188e-01
GL_1210 0 NS_1210 NS_1209 0 -2.1739680820836188e-01
GS_1209_12 0 NS_1209 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1211/1212
CS_1211 NS_1211 0 9.9999999999999998e-13
CS_1212 NS_1212 0 9.9999999999999998e-13
RS_1211 NS_1211 0 1.0859722031634941e+02
RS_1212 NS_1212 0 1.0859722031634941e+02
GL_1211 0 NS_1211 NS_1212 0 2.0887403840929383e-01
GL_1212 0 NS_1212 NS_1211 0 -2.0887403840929383e-01
GS_1211_12 0 NS_1211 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1213/1214
CS_1213 NS_1213 0 9.9999999999999998e-13
CS_1214 NS_1214 0 9.9999999999999998e-13
RS_1213 NS_1213 0 7.7959989808728068e+01
RS_1214 NS_1214 0 7.7959989808728054e+01
GL_1213 0 NS_1213 NS_1214 0 2.0447808896343445e-01
GL_1214 0 NS_1214 NS_1213 0 -2.0447808896343445e-01
GS_1213_12 0 NS_1213 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1215/1216
CS_1215 NS_1215 0 9.9999999999999998e-13
CS_1216 NS_1216 0 9.9999999999999998e-13
RS_1215 NS_1215 0 1.1088851678406323e+02
RS_1216 NS_1216 0 1.1088851678406321e+02
GL_1215 0 NS_1215 NS_1216 0 1.9843399276071924e-01
GL_1216 0 NS_1216 NS_1215 0 -1.9843399276071924e-01
GS_1215_12 0 NS_1215 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1217/1218
CS_1217 NS_1217 0 9.9999999999999998e-13
CS_1218 NS_1218 0 9.9999999999999998e-13
RS_1217 NS_1217 0 8.1179760966262847e+01
RS_1218 NS_1218 0 8.1179760966262847e+01
GL_1217 0 NS_1217 NS_1218 0 1.8978022990658949e-01
GL_1218 0 NS_1218 NS_1217 0 -1.8978022990658949e-01
GS_1217_12 0 NS_1217 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1219/1220
CS_1219 NS_1219 0 9.9999999999999998e-13
CS_1220 NS_1220 0 9.9999999999999998e-13
RS_1219 NS_1219 0 1.0523970815054612e+02
RS_1220 NS_1220 0 1.0523970815054612e+02
GL_1219 0 NS_1219 NS_1220 0 1.8836779078363333e-01
GL_1220 0 NS_1220 NS_1219 0 -1.8836779078363333e-01
GS_1219_12 0 NS_1219 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1221/1222
CS_1221 NS_1221 0 9.9999999999999998e-13
CS_1222 NS_1222 0 9.9999999999999998e-13
RS_1221 NS_1221 0 1.1208834663822537e+02
RS_1222 NS_1222 0 1.1208834663822537e+02
GL_1221 0 NS_1221 NS_1222 0 1.7925451755127267e-01
GL_1222 0 NS_1222 NS_1221 0 -1.7925451755127267e-01
GS_1221_12 0 NS_1221 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1223/1224
CS_1223 NS_1223 0 9.9999999999999998e-13
CS_1224 NS_1224 0 9.9999999999999998e-13
RS_1223 NS_1223 0 9.2475617668062213e+01
RS_1224 NS_1224 0 9.2475617668062199e+01
GL_1223 0 NS_1223 NS_1224 0 1.7507216970358189e-01
GL_1224 0 NS_1224 NS_1223 0 -1.7507216970358189e-01
GS_1223_12 0 NS_1223 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1225/1226
CS_1225 NS_1225 0 9.9999999999999998e-13
CS_1226 NS_1226 0 9.9999999999999998e-13
RS_1225 NS_1225 0 1.1555782965375326e+02
RS_1226 NS_1226 0 1.1555782965375326e+02
GL_1225 0 NS_1225 NS_1226 0 1.6918904340923188e-01
GL_1226 0 NS_1226 NS_1225 0 -1.6918904340923188e-01
GS_1225_12 0 NS_1225 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1227/1228
CS_1227 NS_1227 0 9.9999999999999998e-13
CS_1228 NS_1228 0 9.9999999999999998e-13
RS_1227 NS_1227 0 9.6856782813111039e+01
RS_1228 NS_1228 0 9.6856782813111039e+01
GL_1227 0 NS_1227 NS_1228 0 1.6488898173469207e-01
GL_1228 0 NS_1228 NS_1227 0 -1.6488898173469207e-01
GS_1227_12 0 NS_1227 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1229/1230
CS_1229 NS_1229 0 9.9999999999999998e-13
CS_1230 NS_1230 0 9.9999999999999998e-13
RS_1229 NS_1229 0 1.1717534841017003e+02
RS_1230 NS_1230 0 1.1717534841017003e+02
GL_1229 0 NS_1229 NS_1230 0 1.5866517390841936e-01
GL_1230 0 NS_1230 NS_1229 0 -1.5866517390841936e-01
GS_1229_12 0 NS_1229 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1231/1232
CS_1231 NS_1231 0 9.9999999999999998e-13
CS_1232 NS_1232 0 9.9999999999999998e-13
RS_1231 NS_1231 0 8.8607873746940697e+01
RS_1232 NS_1232 0 8.8607873746940697e+01
GL_1231 0 NS_1231 NS_1232 0 1.5214737618207635e-01
GL_1232 0 NS_1232 NS_1231 0 -1.5214737618207635e-01
GS_1231_12 0 NS_1231 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1233/1234
CS_1233 NS_1233 0 9.9999999999999998e-13
CS_1234 NS_1234 0 9.9999999999999998e-13
RS_1233 NS_1233 0 1.1741456484283673e+02
RS_1234 NS_1234 0 1.1741456484283673e+02
GL_1233 0 NS_1233 NS_1234 0 1.4829748860889613e-01
GL_1234 0 NS_1234 NS_1233 0 -1.4829748860889613e-01
GS_1233_12 0 NS_1233 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1235/1236
CS_1235 NS_1235 0 9.9999999999999998e-13
CS_1236 NS_1236 0 9.9999999999999998e-13
RS_1235 NS_1235 0 1.3292289814180702e+02
RS_1236 NS_1236 0 1.3292289814180702e+02
GL_1235 0 NS_1235 NS_1236 0 1.4243056778188259e-01
GL_1236 0 NS_1236 NS_1235 0 -1.4243056778188259e-01
GS_1235_12 0 NS_1235 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1237/1238
CS_1237 NS_1237 0 9.9999999999999998e-13
CS_1238 NS_1238 0 9.9999999999999998e-13
RS_1237 NS_1237 0 1.2325134819531741e+02
RS_1238 NS_1238 0 1.2325134819531739e+02
GL_1237 0 NS_1237 NS_1238 0 1.3890785074828846e-01
GL_1238 0 NS_1238 NS_1237 0 -1.3890785074828846e-01
GS_1237_12 0 NS_1237 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1239/1240
CS_1239 NS_1239 0 9.9999999999999998e-13
CS_1240 NS_1240 0 9.9999999999999998e-13
RS_1239 NS_1239 0 9.1909059882883227e+01
RS_1240 NS_1240 0 9.1909059882883227e+01
GL_1239 0 NS_1239 NS_1240 0 1.3373879533989103e-01
GL_1240 0 NS_1240 NS_1239 0 -1.3373879533989103e-01
GS_1239_12 0 NS_1239 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1241/1242
CS_1241 NS_1241 0 9.9999999999999998e-13
CS_1242 NS_1242 0 9.9999999999999998e-13
RS_1241 NS_1241 0 1.2276824880349510e+02
RS_1242 NS_1242 0 1.2276824880349510e+02
GL_1241 0 NS_1241 NS_1242 0 1.2885409674522977e-01
GL_1242 0 NS_1242 NS_1241 0 -1.2885409674522977e-01
GS_1241_12 0 NS_1241 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1243/1244
CS_1243 NS_1243 0 9.9999999999999998e-13
CS_1244 NS_1244 0 9.9999999999999998e-13
RS_1243 NS_1243 0 1.1612442076026501e+02
RS_1244 NS_1244 0 1.1612442076026501e+02
GL_1243 0 NS_1243 NS_1244 0 1.2417838026896348e-01
GL_1244 0 NS_1244 NS_1243 0 -1.2417838026896348e-01
GS_1243_12 0 NS_1243 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1245/1246
CS_1245 NS_1245 0 9.9999999999999998e-13
CS_1246 NS_1246 0 9.9999999999999998e-13
RS_1245 NS_1245 0 1.2130204223875414e+02
RS_1246 NS_1246 0 1.2130204223875414e+02
GL_1245 0 NS_1245 NS_1246 0 1.1919240021970828e-01
GL_1246 0 NS_1246 NS_1245 0 -1.1919240021970828e-01
GS_1245_12 0 NS_1245 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1247/1248
CS_1247 NS_1247 0 9.9999999999999998e-13
CS_1248 NS_1248 0 9.9999999999999998e-13
RS_1247 NS_1247 0 9.3083309227260045e+01
RS_1248 NS_1248 0 9.3083309227260045e+01
GL_1247 0 NS_1247 NS_1248 0 1.1485268189050464e-01
GL_1248 0 NS_1248 NS_1247 0 -1.1485268189050464e-01
GS_1247_12 0 NS_1247 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1249/1250
CS_1249 NS_1249 0 9.9999999999999998e-13
CS_1250 NS_1250 0 9.9999999999999998e-13
RS_1249 NS_1249 0 1.2387094149263906e+02
RS_1250 NS_1250 0 1.2387094149263908e+02
GL_1249 0 NS_1249 NS_1250 0 1.0935451806229070e-01
GL_1250 0 NS_1250 NS_1249 0 -1.0935451806229070e-01
GS_1249_12 0 NS_1249 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1251/1252
CS_1251 NS_1251 0 9.9999999999999998e-13
CS_1252 NS_1252 0 9.9999999999999998e-13
RS_1251 NS_1251 0 1.1186020221520803e+02
RS_1252 NS_1252 0 1.1186020221520802e+02
GL_1251 0 NS_1251 NS_1252 0 1.0538242730807947e-01
GL_1252 0 NS_1252 NS_1251 0 -1.0538242730807947e-01
GS_1251_12 0 NS_1251 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1253/1254
CS_1253 NS_1253 0 9.9999999999999998e-13
CS_1254 NS_1254 0 9.9999999999999998e-13
RS_1253 NS_1253 0 1.2031265815570148e+02
RS_1254 NS_1254 0 1.2031265815570150e+02
GL_1253 0 NS_1253 NS_1254 0 9.9497602364102364e-02
GL_1254 0 NS_1254 NS_1253 0 -9.9497602364102364e-02
GS_1253_12 0 NS_1253 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1255/1256
CS_1255 NS_1255 0 9.9999999999999998e-13
CS_1256 NS_1256 0 9.9999999999999998e-13
RS_1255 NS_1255 0 9.6254518048655143e+01
RS_1256 NS_1256 0 9.6254518048655143e+01
GL_1255 0 NS_1255 NS_1256 0 9.5930770757699110e-02
GL_1256 0 NS_1256 NS_1255 0 -9.5930770757699110e-02
GS_1255_12 0 NS_1255 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1257/1258
CS_1257 NS_1257 0 9.9999999999999998e-13
CS_1258 NS_1258 0 9.9999999999999998e-13
RS_1257 NS_1257 0 1.2318640771018909e+02
RS_1258 NS_1258 0 1.2318640771018909e+02
GL_1257 0 NS_1257 NS_1258 0 8.9880619653662355e-02
GL_1258 0 NS_1258 NS_1257 0 -8.9880619653662355e-02
GS_1257_12 0 NS_1257 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1259/1260
CS_1259 NS_1259 0 9.9999999999999998e-13
CS_1260 NS_1260 0 9.9999999999999998e-13
RS_1259 NS_1259 0 1.1312630346155738e+02
RS_1260 NS_1260 0 1.1312630346155738e+02
GL_1259 0 NS_1259 NS_1260 0 8.6534434501560398e-02
GL_1260 0 NS_1260 NS_1259 0 -8.6534434501560398e-02
GS_1259_12 0 NS_1259 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1261/1262
CS_1261 NS_1261 0 9.9999999999999998e-13
CS_1262 NS_1262 0 9.9999999999999998e-13
RS_1261 NS_1261 0 1.1831504703984019e+02
RS_1262 NS_1262 0 1.1831504703984019e+02
GL_1261 0 NS_1261 NS_1262 0 7.9864296724202116e-02
GL_1262 0 NS_1262 NS_1261 0 -7.9864296724202116e-02
GS_1261_12 0 NS_1261 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1263/1264
CS_1263 NS_1263 0 9.9999999999999998e-13
CS_1264 NS_1264 0 9.9999999999999998e-13
RS_1263 NS_1263 0 1.0281987486447559e+02
RS_1264 NS_1264 0 1.0281987486447559e+02
GL_1263 0 NS_1263 NS_1264 0 7.6950339194481784e-02
GL_1264 0 NS_1264 NS_1263 0 -7.6950339194481784e-02
GS_1263_12 0 NS_1263 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1265/1266
CS_1265 NS_1265 0 9.9999999999999998e-13
CS_1266 NS_1266 0 9.9999999999999998e-13
RS_1265 NS_1265 0 1.2230186914382300e+02
RS_1266 NS_1266 0 1.2230186914382300e+02
GL_1265 0 NS_1265 NS_1266 0 7.0709298709435750e-02
GL_1266 0 NS_1266 NS_1265 0 -7.0709298709435750e-02
GS_1265_12 0 NS_1265 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1267/1268
CS_1267 NS_1267 0 9.9999999999999998e-13
CS_1268 NS_1268 0 9.9999999999999998e-13
RS_1267 NS_1267 0 1.2215699953322022e+02
RS_1268 NS_1268 0 1.2215699953322020e+02
GL_1267 0 NS_1267 NS_1268 0 6.7518227185671367e-02
GL_1268 0 NS_1268 NS_1267 0 -6.7518227185671367e-02
GS_1267_12 0 NS_1267 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1269/1270
CS_1269 NS_1269 0 9.9999999999999998e-13
CS_1270 NS_1270 0 9.9999999999999998e-13
RS_1269 NS_1269 0 3.4305564408226764e+03
RS_1270 NS_1270 0 3.4305564408226769e+03
GL_1269 0 NS_1269 NS_1270 0 5.4396471187208063e-02
GL_1270 0 NS_1270 NS_1269 0 -5.4396471187208063e-02
GS_1269_12 0 NS_1269 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1271/1272
CS_1271 NS_1271 0 9.9999999999999998e-13
CS_1272 NS_1272 0 9.9999999999999998e-13
RS_1271 NS_1271 0 1.1894859826238778e+02
RS_1272 NS_1272 0 1.1894859826238779e+02
GL_1271 0 NS_1271 NS_1272 0 6.0591569497719031e-02
GL_1272 0 NS_1272 NS_1271 0 -6.0591569497719031e-02
GS_1271_12 0 NS_1271 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1273/1274
CS_1273 NS_1273 0 9.9999999999999998e-13
CS_1274 NS_1274 0 9.9999999999999998e-13
RS_1273 NS_1273 0 1.3537641711503298e+02
RS_1274 NS_1274 0 1.3537641711503298e+02
GL_1273 0 NS_1273 NS_1274 0 5.1190778164089609e-02
GL_1274 0 NS_1274 NS_1273 0 -5.1190778164089609e-02
GS_1273_12 0 NS_1273 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1275/1276
CS_1275 NS_1275 0 9.9999999999999998e-13
CS_1276 NS_1276 0 9.9999999999999998e-13
RS_1275 NS_1275 0 1.3105452427659637e+02
RS_1276 NS_1276 0 1.3105452427659637e+02
GL_1275 0 NS_1275 NS_1276 0 4.7418984574880592e-02
GL_1276 0 NS_1276 NS_1275 0 -4.7418984574880592e-02
GS_1275_12 0 NS_1275 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1277/1278
CS_1277 NS_1277 0 9.9999999999999998e-13
CS_1278 NS_1278 0 9.9999999999999998e-13
RS_1277 NS_1277 0 1.2170234397098790e+02
RS_1278 NS_1278 0 1.2170234397098790e+02
GL_1277 0 NS_1277 NS_1278 0 4.0778813929127578e-02
GL_1278 0 NS_1278 NS_1277 0 -4.0778813929127578e-02
GS_1277_12 0 NS_1277 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1279/1280
CS_1279 NS_1279 0 9.9999999999999998e-13
CS_1280 NS_1280 0 9.9999999999999998e-13
RS_1279 NS_1279 0 1.1550510326517782e+02
RS_1280 NS_1280 0 1.1550510326517782e+02
GL_1279 0 NS_1279 NS_1280 0 5.7236026076957713e-02
GL_1280 0 NS_1280 NS_1279 0 -5.7236026076957713e-02
GS_1279_12 0 NS_1279 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1281/1282
CS_1281 NS_1281 0 9.9999999999999998e-13
CS_1282 NS_1282 0 9.9999999999999998e-13
RS_1281 NS_1281 0 6.2039157456337159e+02
RS_1282 NS_1282 0 6.2039157456337159e+02
GL_1281 0 NS_1281 NS_1282 0 1.9354364738401211e-02
GL_1282 0 NS_1282 NS_1281 0 -1.9354364738401211e-02
GS_1281_12 0 NS_1281 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1283/1284
CS_1283 NS_1283 0 9.9999999999999998e-13
CS_1284 NS_1284 0 9.9999999999999998e-13
RS_1283 NS_1283 0 1.1050313240441588e+02
RS_1284 NS_1284 0 1.1050313240441587e+02
GL_1283 0 NS_1283 NS_1284 0 1.6472588786558075e-02
GL_1284 0 NS_1284 NS_1283 0 -1.6472588786558075e-02
GS_1283_12 0 NS_1283 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1285/1286
CS_1285 NS_1285 0 9.9999999999999998e-13
CS_1286 NS_1286 0 9.9999999999999998e-13
RS_1285 NS_1285 0 1.2869119986945731e+02
RS_1286 NS_1286 0 1.2869119986945731e+02
GL_1285 0 NS_1285 NS_1286 0 2.0888592987579706e-02
GL_1286 0 NS_1286 NS_1285 0 -2.0888592987579706e-02
GS_1285_12 0 NS_1285 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1287/1288
CS_1287 NS_1287 0 9.9999999999999998e-13
CS_1288 NS_1288 0 9.9999999999999998e-13
RS_1287 NS_1287 0 1.4314560950270646e+02
RS_1288 NS_1288 0 1.4314560950270646e+02
GL_1287 0 NS_1287 NS_1288 0 9.7871236580563716e-03
GL_1288 0 NS_1288 NS_1287 0 -9.7871236580563716e-03
GS_1287_12 0 NS_1287 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1289/1290
CS_1289 NS_1289 0 9.9999999999999998e-13
CS_1290 NS_1290 0 9.9999999999999998e-13
RS_1289 NS_1289 0 1.1863004336811436e+02
RS_1290 NS_1290 0 1.1863004336811436e+02
GL_1289 0 NS_1289 NS_1290 0 3.7627463994326378e-02
GL_1290 0 NS_1290 NS_1289 0 -3.7627463994326378e-02
GS_1289_12 0 NS_1289 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1291/1292
CS_1291 NS_1291 0 9.9999999999999998e-13
CS_1292 NS_1292 0 9.9999999999999998e-13
RS_1291 NS_1291 0 1.2686172273444870e+02
RS_1292 NS_1292 0 1.2686172273444869e+02
GL_1291 0 NS_1291 NS_1292 0 3.1975218188091938e-02
GL_1292 0 NS_1292 NS_1291 0 -3.1975218188091938e-02
GS_1291_12 0 NS_1291 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1293/1294
CS_1293 NS_1293 0 9.9999999999999998e-13
CS_1294 NS_1294 0 9.9999999999999998e-13
RS_1293 NS_1293 0 1.3141621772977734e+02
RS_1294 NS_1294 0 1.3141621772977737e+02
GL_1293 0 NS_1293 NS_1294 0 2.8228381102665165e-02
GL_1294 0 NS_1294 NS_1293 0 -2.8228381102665165e-02
GS_1293_12 0 NS_1293 NA_12 0 4.7428518688027549e-01
*
* Complex pair n. 1295/1296
CS_1295 NS_1295 0 9.9999999999999998e-13
CS_1296 NS_1296 0 9.9999999999999998e-13
RS_1295 NS_1295 0 1.2452833644614726e+02
RS_1296 NS_1296 0 1.2452833644614726e+02
GL_1295 0 NS_1295 NS_1296 0 2.1457325426059259e-03
GL_1296 0 NS_1296 NS_1295 0 -2.1457325426059259e-03
GS_1295_12 0 NS_1295 NA_12 0 4.7428518688027549e-01
*
******************************


.ends
*******************
* End of subcircuit
*******************
