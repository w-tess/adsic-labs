**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [4 2 18] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_10_Module_wire_5mm_highloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 6.0205251484948263e-02
GC_1_2 b_1 NI_1 NS_2 0 7.0943153626971264e-06
GC_1_3 b_1 NI_1 NS_3 0 -1.1476371582700626e-12
GC_1_4 b_1 NI_1 NS_4 0 -2.4577438379349798e-06
GC_1_5 b_1 NI_1 NS_5 0 2.1424806003270924e-05
GC_1_6 b_1 NI_1 NS_6 0 -3.0072781652674183e-06
GC_1_7 b_1 NI_1 NS_7 0 -1.5768793472550066e-03
GC_1_8 b_1 NI_1 NS_8 0 6.8779715886366291e-03
GC_1_9 b_1 NI_1 NS_9 0 1.7132713273899956e-02
GC_1_10 b_1 NI_1 NS_10 0 -5.5821258612093940e-03
GC_1_11 b_1 NI_1 NS_11 0 -2.5778390981369328e-02
GC_1_12 b_1 NI_1 NS_12 0 -3.1260446955133490e-02
GC_1_13 b_1 NI_1 NS_13 0 7.1572695533649684e-03
GC_1_14 b_1 NI_1 NS_14 0 2.9562125843075088e-03
GC_1_15 b_1 NI_1 NS_15 0 -3.0968372041693840e-02
GC_1_16 b_1 NI_1 NS_16 0 -3.3276400518464221e-02
GC_1_17 b_1 NI_1 NS_17 0 1.9531977786943561e-01
GC_1_18 b_1 NI_1 NS_18 0 1.1092557322625719e-04
GC_1_19 b_1 NI_1 NS_19 0 1.5682675589712093e-12
GC_1_20 b_1 NI_1 NS_20 0 4.4032541271731149e-06
GC_1_21 b_1 NI_1 NS_21 0 1.1663255304785503e-04
GC_1_22 b_1 NI_1 NS_22 0 4.6013536732782820e-05
GC_1_23 b_1 NI_1 NS_23 0 -6.1176641058101063e-02
GC_1_24 b_1 NI_1 NS_24 0 -4.4021400941638665e-02
GC_1_25 b_1 NI_1 NS_25 0 3.9561848843105069e-02
GC_1_26 b_1 NI_1 NS_26 0 -1.8838335315735286e-02
GC_1_27 b_1 NI_1 NS_27 0 -1.2336119995522446e-01
GC_1_28 b_1 NI_1 NS_28 0 7.0714523433327334e-02
GC_1_29 b_1 NI_1 NS_29 0 -2.2401392583017082e-02
GC_1_30 b_1 NI_1 NS_30 0 1.2250576766664073e-02
GC_1_31 b_1 NI_1 NS_31 0 2.6304263603534425e-02
GC_1_32 b_1 NI_1 NS_32 0 -6.4426935154424603e-02
GC_1_33 b_1 NI_1 NS_33 0 9.3916310000033334e-03
GC_1_34 b_1 NI_1 NS_34 0 1.2890509398882415e-05
GC_1_35 b_1 NI_1 NS_35 0 2.5386651324276448e-13
GC_1_36 b_1 NI_1 NS_36 0 -3.4312185280572385e-07
GC_1_37 b_1 NI_1 NS_37 0 -2.1090937152936802e-05
GC_1_38 b_1 NI_1 NS_38 0 -3.9310816326749106e-06
GC_1_39 b_1 NI_1 NS_39 0 -1.8572943129050818e-03
GC_1_40 b_1 NI_1 NS_40 0 -1.1603165995088826e-02
GC_1_41 b_1 NI_1 NS_41 0 -2.7111006744116692e-02
GC_1_42 b_1 NI_1 NS_42 0 4.1602552746640778e-03
GC_1_43 b_1 NI_1 NS_43 0 1.3734246053024686e-02
GC_1_44 b_1 NI_1 NS_44 0 3.3872451327831038e-02
GC_1_45 b_1 NI_1 NS_45 0 -1.0082683243490417e-02
GC_1_46 b_1 NI_1 NS_46 0 -1.0952382006085655e-03
GC_1_47 b_1 NI_1 NS_47 0 2.5364175891973300e-02
GC_1_48 b_1 NI_1 NS_48 0 3.4556235553199040e-02
GC_1_49 b_1 NI_1 NS_49 0 -3.8114674624403137e-03
GC_1_50 b_1 NI_1 NS_50 0 4.0468601017153458e-06
GC_1_51 b_1 NI_1 NS_51 0 2.6117693463007082e-13
GC_1_52 b_1 NI_1 NS_52 0 -1.2929380642448919e-08
GC_1_53 b_1 NI_1 NS_53 0 -5.0426015755861583e-05
GC_1_54 b_1 NI_1 NS_54 0 1.1717363001461861e-05
GC_1_55 b_1 NI_1 NS_55 0 -2.9195291497743120e-03
GC_1_56 b_1 NI_1 NS_56 0 -2.2869863001898499e-03
GC_1_57 b_1 NI_1 NS_57 0 -6.9814384794004165e-03
GC_1_58 b_1 NI_1 NS_58 0 1.0662378453447955e-03
GC_1_59 b_1 NI_1 NS_59 0 -8.3763004742843736e-03
GC_1_60 b_1 NI_1 NS_60 0 3.0424302078871524e-02
GC_1_61 b_1 NI_1 NS_61 0 1.0638687100251419e-02
GC_1_62 b_1 NI_1 NS_62 0 -3.4452978654049636e-04
GC_1_63 b_1 NI_1 NS_63 0 1.6778994941729068e-02
GC_1_64 b_1 NI_1 NS_64 0 7.7219988180529412e-03
GC_1_65 b_1 NI_1 NS_65 0 -4.1523818208867988e-03
GC_1_66 b_1 NI_1 NS_66 0 1.7210140330758331e-06
GC_1_67 b_1 NI_1 NS_67 0 -1.6982581254736722e-13
GC_1_68 b_1 NI_1 NS_68 0 4.6462986767592645e-08
GC_1_69 b_1 NI_1 NS_69 0 1.3501259769394363e-05
GC_1_70 b_1 NI_1 NS_70 0 -3.8169465291475171e-06
GC_1_71 b_1 NI_1 NS_71 0 2.5164729664481561e-05
GC_1_72 b_1 NI_1 NS_72 0 2.5210476271255016e-05
GC_1_73 b_1 NI_1 NS_73 0 -3.8970066131061010e-04
GC_1_74 b_1 NI_1 NS_74 0 3.7440407553661863e-04
GC_1_75 b_1 NI_1 NS_75 0 1.1968567668834878e-03
GC_1_76 b_1 NI_1 NS_76 0 1.9813017237245681e-03
GC_1_77 b_1 NI_1 NS_77 0 1.9708689931203743e-04
GC_1_78 b_1 NI_1 NS_78 0 -2.0917018607214435e-04
GC_1_79 b_1 NI_1 NS_79 0 1.7545258902549605e-03
GC_1_80 b_1 NI_1 NS_80 0 1.3468062126914093e-03
GC_1_81 b_1 NI_1 NS_81 0 -5.1038232413588901e-04
GC_1_82 b_1 NI_1 NS_82 0 -1.3759943973706266e-06
GC_1_83 b_1 NI_1 NS_83 0 -1.7070376138007358e-13
GC_1_84 b_1 NI_1 NS_84 0 2.8016737456310675e-08
GC_1_85 b_1 NI_1 NS_85 0 7.0315257051580351e-06
GC_1_86 b_1 NI_1 NS_86 0 -1.3983676095631051e-06
GC_1_87 b_1 NI_1 NS_87 0 6.7658885068303844e-04
GC_1_88 b_1 NI_1 NS_88 0 5.6603060806773790e-04
GC_1_89 b_1 NI_1 NS_89 0 1.6569619427860946e-03
GC_1_90 b_1 NI_1 NS_90 0 -1.3045817546181629e-04
GC_1_91 b_1 NI_1 NS_91 0 2.1462925826014499e-03
GC_1_92 b_1 NI_1 NS_92 0 -6.5332367834813080e-03
GC_1_93 b_1 NI_1 NS_93 0 -2.2964828318146812e-03
GC_1_94 b_1 NI_1 NS_94 0 2.6291046654986247e-05
GC_1_95 b_1 NI_1 NS_95 0 -3.4079523501683549e-03
GC_1_96 b_1 NI_1 NS_96 0 -1.5814693509543160e-03
GC_1_97 b_1 NI_1 NS_97 0 1.4735125392038942e-03
GC_1_98 b_1 NI_1 NS_98 0 -3.7426276886598965e-07
GC_1_99 b_1 NI_1 NS_99 0 2.0729541104523740e-14
GC_1_100 b_1 NI_1 NS_100 0 -1.6072318035552761e-08
GC_1_101 b_1 NI_1 NS_101 0 -3.8273514999394242e-06
GC_1_102 b_1 NI_1 NS_102 0 1.0175438209487778e-06
GC_1_103 b_1 NI_1 NS_103 0 -1.9610747217130337e-05
GC_1_104 b_1 NI_1 NS_104 0 -8.8856162824760339e-05
GC_1_105 b_1 NI_1 NS_105 0 -5.5034649401411377e-05
GC_1_106 b_1 NI_1 NS_106 0 -1.0544989336485160e-04
GC_1_107 b_1 NI_1 NS_107 0 -3.3160039456642980e-04
GC_1_108 b_1 NI_1 NS_108 0 -4.2825946799977192e-04
GC_1_109 b_1 NI_1 NS_109 0 -1.2974747386928175e-04
GC_1_110 b_1 NI_1 NS_110 0 6.5863739714910137e-05
GC_1_111 b_1 NI_1 NS_111 0 -4.1022481359596230e-04
GC_1_112 b_1 NI_1 NS_112 0 -2.0280474986638175e-04
GC_1_113 b_1 NI_1 NS_113 0 -1.1925201589246396e-04
GC_1_114 b_1 NI_1 NS_114 0 -4.5752297865929250e-08
GC_1_115 b_1 NI_1 NS_115 0 2.0535967851557122e-14
GC_1_116 b_1 NI_1 NS_116 0 5.1316971228641972e-09
GC_1_117 b_1 NI_1 NS_117 0 7.9241182304107510e-07
GC_1_118 b_1 NI_1 NS_118 0 -2.5092058318194577e-07
GC_1_119 b_1 NI_1 NS_119 0 6.1190009795600653e-05
GC_1_120 b_1 NI_1 NS_120 0 6.1410070503378915e-05
GC_1_121 b_1 NI_1 NS_121 0 1.6107733292740979e-04
GC_1_122 b_1 NI_1 NS_122 0 -4.5879646151363672e-06
GC_1_123 b_1 NI_1 NS_123 0 2.3879194704770008e-04
GC_1_124 b_1 NI_1 NS_124 0 -6.0017895586455324e-04
GC_1_125 b_1 NI_1 NS_125 0 -2.1677325015477877e-04
GC_1_126 b_1 NI_1 NS_126 0 -4.6054267695783660e-06
GC_1_127 b_1 NI_1 NS_127 0 -3.1210421769126308e-04
GC_1_128 b_1 NI_1 NS_128 0 -1.5288177643754601e-04
GC_1_129 b_1 NI_1 NS_129 0 8.1331867742518530e-05
GC_1_130 b_1 NI_1 NS_130 0 -2.2323934629457193e-08
GC_1_131 b_1 NI_1 NS_131 0 3.4392760855977476e-15
GC_1_132 b_1 NI_1 NS_132 0 -9.4734547744753566e-10
GC_1_133 b_1 NI_1 NS_133 0 -2.1747855548315541e-07
GC_1_134 b_1 NI_1 NS_134 0 6.3855388949437116e-08
GC_1_135 b_1 NI_1 NS_135 0 -1.4295318310883328e-06
GC_1_136 b_1 NI_1 NS_136 0 -5.8091550752597977e-06
GC_1_137 b_1 NI_1 NS_137 0 -4.4249397507260294e-06
GC_1_138 b_1 NI_1 NS_138 0 -4.8386380127304990e-06
GC_1_139 b_1 NI_1 NS_139 0 -1.6839083414878980e-05
GC_1_140 b_1 NI_1 NS_140 0 -2.3392374160341896e-05
GC_1_141 b_1 NI_1 NS_141 0 -8.2689930482527607e-06
GC_1_142 b_1 NI_1 NS_142 0 4.0287093675067526e-06
GC_1_143 b_1 NI_1 NS_143 0 -2.1378508858784737e-05
GC_1_144 b_1 NI_1 NS_144 0 -9.0316774874675093e-06
GC_1_145 b_1 NI_1 NS_145 0 2.2238544040041871e-05
GC_1_146 b_1 NI_1 NS_146 0 -1.0064756417884591e-08
GC_1_147 b_1 NI_1 NS_147 0 3.4193648198259035e-15
GC_1_148 b_1 NI_1 NS_148 0 -3.8807162185424266e-10
GC_1_149 b_1 NI_1 NS_149 0 -4.7675817524582017e-08
GC_1_150 b_1 NI_1 NS_150 0 1.6907816836000958e-08
GC_1_151 b_1 NI_1 NS_151 0 -2.6188596420402065e-06
GC_1_152 b_1 NI_1 NS_152 0 3.2026081629342382e-06
GC_1_153 b_1 NI_1 NS_153 0 3.1866851604520283e-06
GC_1_154 b_1 NI_1 NS_154 0 -1.9347471468756970e-06
GC_1_155 b_1 NI_1 NS_155 0 1.2380035347421740e-06
GC_1_156 b_1 NI_1 NS_156 0 -9.9238805675602338e-06
GC_1_157 b_1 NI_1 NS_157 0 -4.6631466233878171e-06
GC_1_158 b_1 NI_1 NS_158 0 7.8397538049522044e-07
GC_1_159 b_1 NI_1 NS_159 0 -8.5401411630734192e-06
GC_1_160 b_1 NI_1 NS_160 0 -5.6351988201231859e-06
GC_1_161 b_1 NI_1 NS_161 0 9.1074232800494396e-06
GC_1_162 b_1 NI_1 NS_162 0 -5.4503963224388379e-11
GC_1_163 b_1 NI_1 NS_163 0 -9.9062282116010417e-16
GC_1_164 b_1 NI_1 NS_164 0 -1.5773102594273834e-10
GC_1_165 b_1 NI_1 NS_165 0 -4.3660385537143305e-08
GC_1_166 b_1 NI_1 NS_166 0 1.7498227374859664e-08
GC_1_167 b_1 NI_1 NS_167 0 -5.6993811517828405e-07
GC_1_168 b_1 NI_1 NS_168 0 -1.6159752970188905e-06
GC_1_169 b_1 NI_1 NS_169 0 -3.1702340747716266e-06
GC_1_170 b_1 NI_1 NS_170 0 6.9399366047867965e-08
GC_1_171 b_1 NI_1 NS_171 0 2.6919058784478408e-07
GC_1_172 b_1 NI_1 NS_172 0 2.5899185610949878e-06
GC_1_173 b_1 NI_1 NS_173 0 -1.1424458225853375e-06
GC_1_174 b_1 NI_1 NS_174 0 -5.5947059733083705e-07
GC_1_175 b_1 NI_1 NS_175 0 -2.6420655613151241e-07
GC_1_176 b_1 NI_1 NS_176 0 1.0913704237379017e-06
GC_1_177 b_1 NI_1 NS_177 0 8.6589498205072128e-06
GC_1_178 b_1 NI_1 NS_178 0 -8.8451219184059332e-09
GC_1_179 b_1 NI_1 NS_179 0 -9.7886257306803411e-16
GC_1_180 b_1 NI_1 NS_180 0 9.8400245278620121e-11
GC_1_181 b_1 NI_1 NS_181 0 3.1547636649705533e-08
GC_1_182 b_1 NI_1 NS_182 0 -1.3740621488858409e-08
GC_1_183 b_1 NI_1 NS_183 0 -2.8506208960087747e-06
GC_1_184 b_1 NI_1 NS_184 0 2.4730779676767068e-06
GC_1_185 b_1 NI_1 NS_185 0 4.8737771176466801e-07
GC_1_186 b_1 NI_1 NS_186 0 -2.0951091626761403e-06
GC_1_187 b_1 NI_1 NS_187 0 1.2467753480529139e-06
GC_1_188 b_1 NI_1 NS_188 0 2.4328941997773351e-06
GC_1_189 b_1 NI_1 NS_189 0 -1.5009743426458823e-06
GC_1_190 b_1 NI_1 NS_190 0 3.6509715056413818e-07
GC_1_191 b_1 NI_1 NS_191 0 -3.2123308243524511e-07
GC_1_192 b_1 NI_1 NS_192 0 -7.4418315056212979e-07
GD_1_1 b_1 NI_1 NA_1 0 -3.5123744329580028e-02
GD_1_2 b_1 NI_1 NA_2 0 -1.7153451787590202e-02
GD_1_3 b_1 NI_1 NA_3 0 4.8388543200682020e-03
GD_1_4 b_1 NI_1 NA_4 0 -5.0311812670005406e-03
GD_1_5 b_1 NI_1 NA_5 0 1.2298218510396056e-03
GD_1_6 b_1 NI_1 NA_6 0 1.5591662048489708e-03
GD_1_7 b_1 NI_1 NA_7 0 -3.8457943015824867e-04
GD_1_8 b_1 NI_1 NA_8 0 1.6472672024082363e-04
GD_1_9 b_1 NI_1 NA_9 0 -2.0122332077995539e-05
GD_1_10 b_1 NI_1 NA_10 0 -9.6481903477474770e-06
GD_1_11 b_1 NI_1 NA_11 0 -2.1459822762373873e-06
GD_1_12 b_1 NI_1 NA_12 0 -3.8758184969025149e-06
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 1.9531221624773548e-01
GC_2_2 b_2 NI_2 NS_2 0 1.1189589590028651e-04
GC_2_3 b_2 NI_2 NS_3 0 1.5688841708078404e-12
GC_2_4 b_2 NI_2 NS_4 0 4.4028400933338810e-06
GC_2_5 b_2 NI_2 NS_5 0 1.1651318673976967e-04
GC_2_6 b_2 NI_2 NS_6 0 4.6043817438571577e-05
GC_2_7 b_2 NI_2 NS_7 0 -6.1176723629265836e-02
GC_2_8 b_2 NI_2 NS_8 0 -4.4021179628839814e-02
GC_2_9 b_2 NI_2 NS_9 0 3.9561519469657407e-02
GC_2_10 b_2 NI_2 NS_10 0 -1.8837952621568965e-02
GC_2_11 b_2 NI_2 NS_11 0 -1.2336191078236922e-01
GC_2_12 b_2 NI_2 NS_12 0 7.0718552014968225e-02
GC_2_13 b_2 NI_2 NS_13 0 -2.2400230684599731e-02
GC_2_14 b_2 NI_2 NS_14 0 1.2251150923926944e-02
GC_2_15 b_2 NI_2 NS_15 0 2.6308854793943827e-02
GC_2_16 b_2 NI_2 NS_16 0 -6.4419789753437748e-02
GC_2_17 b_2 NI_2 NS_17 0 6.0202694648056665e-02
GC_2_18 b_2 NI_2 NS_18 0 7.2133734969322096e-06
GC_2_19 b_2 NI_2 NS_19 0 -1.1474146835443118e-12
GC_2_20 b_2 NI_2 NS_20 0 -2.4577953025727553e-06
GC_2_21 b_2 NI_2 NS_21 0 2.1410866020874879e-05
GC_2_22 b_2 NI_2 NS_22 0 -3.0036759060418889e-06
GC_2_23 b_2 NI_2 NS_23 0 -1.5768214010540254e-03
GC_2_24 b_2 NI_2 NS_24 0 6.8780787869054776e-03
GC_2_25 b_2 NI_2 NS_25 0 1.7132776895214800e-02
GC_2_26 b_2 NI_2 NS_26 0 -5.5819918018604813e-03
GC_2_27 b_2 NI_2 NS_27 0 -2.5778005600070420e-02
GC_2_28 b_2 NI_2 NS_28 0 -3.1259784573285661e-02
GC_2_29 b_2 NI_2 NS_29 0 7.1574409802910594e-03
GC_2_30 b_2 NI_2 NS_30 0 2.9561865760672347e-03
GC_2_31 b_2 NI_2 NS_31 0 -3.0967585260882453e-02
GC_2_32 b_2 NI_2 NS_32 0 -3.3275470486149782e-02
GC_2_33 b_2 NI_2 NS_33 0 -3.8129459114389060e-03
GC_2_34 b_2 NI_2 NS_34 0 3.9682012335500167e-06
GC_2_35 b_2 NI_2 NS_35 0 2.6115721637012573e-13
GC_2_36 b_2 NI_2 NS_36 0 -1.2839410848137323e-08
GC_2_37 b_2 NI_2 NS_37 0 -5.0410561971092315e-05
GC_2_38 b_2 NI_2 NS_38 0 1.1712775258369226e-05
GC_2_39 b_2 NI_2 NS_39 0 -2.9194636137048965e-03
GC_2_40 b_2 NI_2 NS_40 0 -2.2869230859194215e-03
GC_2_41 b_2 NI_2 NS_41 0 -6.9813407396203953e-03
GC_2_42 b_2 NI_2 NS_42 0 1.0663047402449529e-03
GC_2_43 b_2 NI_2 NS_43 0 -8.3757868098408867e-03
GC_2_44 b_2 NI_2 NS_44 0 3.0424462684715985e-02
GC_2_45 b_2 NI_2 NS_45 0 1.0638726707728138e-02
GC_2_46 b_2 NI_2 NS_46 0 -3.4467506203403905e-04
GC_2_47 b_2 NI_2 NS_47 0 1.6779104441262252e-02
GC_2_48 b_2 NI_2 NS_48 0 7.7216498807375642e-03
GC_2_49 b_2 NI_2 NS_49 0 9.3962866360425539e-03
GC_2_50 b_2 NI_2 NS_50 0 1.2543646447372356e-05
GC_2_51 b_2 NI_2 NS_51 0 2.5386400355012452e-13
GC_2_52 b_2 NI_2 NS_52 0 -3.4297135842972635e-07
GC_2_53 b_2 NI_2 NS_53 0 -2.1050390637433167e-05
GC_2_54 b_2 NI_2 NS_54 0 -3.9414549377976160e-06
GC_2_55 b_2 NI_2 NS_55 0 -1.8572619933614194e-03
GC_2_56 b_2 NI_2 NS_56 0 -1.1603257292804229e-02
GC_2_57 b_2 NI_2 NS_57 0 -2.7110876863627942e-02
GC_2_58 b_2 NI_2 NS_58 0 4.1598959735016129e-03
GC_2_59 b_2 NI_2 NS_59 0 1.3733899176534458e-02
GC_2_60 b_2 NI_2 NS_60 0 3.3870468214837808e-02
GC_2_61 b_2 NI_2 NS_61 0 -1.0083207807807866e-02
GC_2_62 b_2 NI_2 NS_62 0 -1.0953347942565840e-03
GC_2_63 b_2 NI_2 NS_63 0 2.5362048132551659e-02
GC_2_64 b_2 NI_2 NS_64 0 3.4553475500296367e-02
GC_2_65 b_2 NI_2 NS_65 0 -5.1016542699475979e-04
GC_2_66 b_2 NI_2 NS_66 0 -1.3847441641100505e-06
GC_2_67 b_2 NI_2 NS_67 0 -1.7070172125237504e-13
GC_2_68 b_2 NI_2 NS_68 0 2.8016090892267160e-08
GC_2_69 b_2 NI_2 NS_69 0 7.0321259366114545e-06
GC_2_70 b_2 NI_2 NS_70 0 -1.3984659037151064e-06
GC_2_71 b_2 NI_2 NS_71 0 6.7658582717854382e-04
GC_2_72 b_2 NI_2 NS_72 0 5.6602652915084225e-04
GC_2_73 b_2 NI_2 NS_73 0 1.6569514891551713e-03
GC_2_74 b_2 NI_2 NS_74 0 -1.3047091056567591e-04
GC_2_75 b_2 NI_2 NS_75 0 2.1462694601077814e-03
GC_2_76 b_2 NI_2 NS_76 0 -6.5332777343236996e-03
GC_2_77 b_2 NI_2 NS_77 0 -2.2964950720986456e-03
GC_2_78 b_2 NI_2 NS_78 0 2.6288041466637070e-05
GC_2_79 b_2 NI_2 NS_79 0 -3.4080189717581944e-03
GC_2_80 b_2 NI_2 NS_80 0 -1.5815496500284681e-03
GC_2_81 b_2 NI_2 NS_81 0 -4.1559289121792086e-03
GC_2_82 b_2 NI_2 NS_82 0 1.7148659646315351e-06
GC_2_83 b_2 NI_2 NS_83 0 -1.6982644434867122e-13
GC_2_84 b_2 NI_2 NS_84 0 4.6466589063766691e-08
GC_2_85 b_2 NI_2 NS_85 0 1.3502673977502525e-05
GC_2_86 b_2 NI_2 NS_86 0 -3.8175819395826150e-06
GC_2_87 b_2 NI_2 NS_87 0 2.5147125304792348e-05
GC_2_88 b_2 NI_2 NS_88 0 2.5429669357183938e-05
GC_2_89 b_2 NI_2 NS_89 0 -3.8931038067688782e-04
GC_2_90 b_2 NI_2 NS_90 0 3.7479474459714307e-04
GC_2_91 b_2 NI_2 NS_91 0 1.1977166881841058e-03
GC_2_92 b_2 NI_2 NS_92 0 1.9814995404555179e-03
GC_2_93 b_2 NI_2 NS_93 0 1.9727524003284474e-04
GC_2_94 b_2 NI_2 NS_94 0 -2.0918073983072386e-04
GC_2_95 b_2 NI_2 NS_95 0 1.7551917920504800e-03
GC_2_96 b_2 NI_2 NS_96 0 1.3469374017120797e-03
GC_2_97 b_2 NI_2 NS_97 0 -1.1780902937185073e-04
GC_2_98 b_2 NI_2 NS_98 0 -4.6617047246599102e-08
GC_2_99 b_2 NI_2 NS_99 0 2.0534206683678893e-14
GC_2_100 b_2 NI_2 NS_100 0 5.1305075087553212e-09
GC_2_101 b_2 NI_2 NS_101 0 7.9260834831309317e-07
GC_2_102 b_2 NI_2 NS_102 0 -2.5091915014234904e-07
GC_2_103 b_2 NI_2 NS_103 0 6.1088039954247954e-05
GC_2_104 b_2 NI_2 NS_104 0 6.1302953788152560e-05
GC_2_105 b_2 NI_2 NS_105 0 1.6097836972919419e-04
GC_2_106 b_2 NI_2 NS_106 0 -4.7204065192345606e-06
GC_2_107 b_2 NI_2 NS_107 0 2.3816405462596040e-04
GC_2_108 b_2 NI_2 NS_108 0 -6.0017432746003216e-04
GC_2_109 b_2 NI_2 NS_109 0 -2.1673614429876215e-04
GC_2_110 b_2 NI_2 NS_110 0 -4.4693097859784501e-06
GC_2_111 b_2 NI_2 NS_111 0 -3.1215588369055020e-04
GC_2_112 b_2 NI_2 NS_112 0 -1.5281005796470413e-04
GC_2_113 b_2 NI_2 NS_113 0 1.4734830752969193e-03
GC_2_114 b_2 NI_2 NS_114 0 -3.7229162567592411e-07
GC_2_115 b_2 NI_2 NS_115 0 2.0731286953677260e-14
GC_2_116 b_2 NI_2 NS_116 0 -1.6072870802073592e-08
GC_2_117 b_2 NI_2 NS_117 0 -3.8275568722240477e-06
GC_2_118 b_2 NI_2 NS_118 0 1.0175896824919994e-06
GC_2_119 b_2 NI_2 NS_119 0 -1.9607386229125299e-05
GC_2_120 b_2 NI_2 NS_120 0 -8.8854137851485232e-05
GC_2_121 b_2 NI_2 NS_121 0 -5.5031303938276242e-05
GC_2_122 b_2 NI_2 NS_122 0 -1.0545527563378640e-04
GC_2_123 b_2 NI_2 NS_123 0 -3.3160884380628320e-04
GC_2_124 b_2 NI_2 NS_124 0 -4.2825521697793096e-04
GC_2_125 b_2 NI_2 NS_125 0 -1.2974371497085217e-04
GC_2_126 b_2 NI_2 NS_126 0 6.5865118114970719e-05
GC_2_127 b_2 NI_2 NS_127 0 -4.1021672280259792e-04
GC_2_128 b_2 NI_2 NS_128 0 -2.0279105793133707e-04
GC_2_129 b_2 NI_2 NS_129 0 2.2230444195250080e-05
GC_2_130 b_2 NI_2 NS_130 0 -9.9611077646007977e-09
GC_2_131 b_2 NI_2 NS_131 0 3.4193023796842006e-15
GC_2_132 b_2 NI_2 NS_132 0 -3.8794237148410095e-10
GC_2_133 b_2 NI_2 NS_133 0 -4.7665277003022454e-08
GC_2_134 b_2 NI_2 NS_134 0 1.6902941931476875e-08
GC_2_135 b_2 NI_2 NS_135 0 -2.6190329609738968e-06
GC_2_136 b_2 NI_2 NS_136 0 3.2035948758236593e-06
GC_2_137 b_2 NI_2 NS_137 0 3.1867006582806097e-06
GC_2_138 b_2 NI_2 NS_138 0 -1.9336503047898789e-06
GC_2_139 b_2 NI_2 NS_139 0 1.2409565244588597e-06
GC_2_140 b_2 NI_2 NS_140 0 -9.9200548634325310e-06
GC_2_141 b_2 NI_2 NS_141 0 -4.6622930961573895e-06
GC_2_142 b_2 NI_2 NS_142 0 7.8335401702980057e-07
GC_2_143 b_2 NI_2 NS_143 0 -8.5371677390938091e-06
GC_2_144 b_2 NI_2 NS_144 0 -5.6333786489929951e-06
GC_2_145 b_2 NI_2 NS_145 0 8.1142020592817914e-05
GC_2_146 b_2 NI_2 NS_146 0 -2.2162478194587910e-08
GC_2_147 b_2 NI_2 NS_147 0 3.4401096205135251e-15
GC_2_148 b_2 NI_2 NS_148 0 -9.4507065244011945e-10
GC_2_149 b_2 NI_2 NS_149 0 -2.1714846895328482e-07
GC_2_150 b_2 NI_2 NS_150 0 6.3742076745142216e-08
GC_2_151 b_2 NI_2 NS_151 0 -1.4238572160722327e-06
GC_2_152 b_2 NI_2 NS_152 0 -5.8118032770926077e-06
GC_2_153 b_2 NI_2 NS_153 0 -4.4293109027193606e-06
GC_2_154 b_2 NI_2 NS_154 0 -4.8292084423012305e-06
GC_2_155 b_2 NI_2 NS_155 0 -1.6795450240274911e-05
GC_2_156 b_2 NI_2 NS_156 0 -2.3341120537570009e-05
GC_2_157 b_2 NI_2 NS_157 0 -8.2574386714923778e-06
GC_2_158 b_2 NI_2 NS_158 0 4.0167068053552016e-06
GC_2_159 b_2 NI_2 NS_159 0 -2.1338511244282370e-05
GC_2_160 b_2 NI_2 NS_160 0 -9.0143072077242359e-06
GC_2_161 b_2 NI_2 NS_161 0 8.6710802233630906e-06
GC_2_162 b_2 NI_2 NS_162 0 -8.8697614285966126e-09
GC_2_163 b_2 NI_2 NS_163 0 -9.7872188059390193e-16
GC_2_164 b_2 NI_2 NS_164 0 9.8050395946346011e-11
GC_2_165 b_2 NI_2 NS_165 0 3.1496441142266480e-08
GC_2_166 b_2 NI_2 NS_166 0 -1.3723179339223559e-08
GC_2_167 b_2 NI_2 NS_167 0 -2.8503081472244566e-06
GC_2_168 b_2 NI_2 NS_168 0 2.4728469614727527e-06
GC_2_169 b_2 NI_2 NS_169 0 4.8801964048922158e-07
GC_2_170 b_2 NI_2 NS_170 0 -2.0960568676196661e-06
GC_2_171 b_2 NI_2 NS_171 0 1.2450034717764232e-06
GC_2_172 b_2 NI_2 NS_172 0 2.4243907716261938e-06
GC_2_173 b_2 NI_2 NS_173 0 -1.5033993225750322e-06
GC_2_174 b_2 NI_2 NS_174 0 3.6646642951993422e-07
GC_2_175 b_2 NI_2 NS_175 0 -3.2644927029052930e-07
GC_2_176 b_2 NI_2 NS_176 0 -7.4696992301315618e-07
GC_2_177 b_2 NI_2 NS_177 0 9.1085069509395807e-06
GC_2_178 b_2 NI_2 NS_178 0 -1.2930804902054696e-10
GC_2_179 b_2 NI_2 NS_179 0 -9.9059831111710994e-16
GC_2_180 b_2 NI_2 NS_180 0 -1.5771847274366732e-10
GC_2_181 b_2 NI_2 NS_181 0 -4.3653087683898768e-08
GC_2_182 b_2 NI_2 NS_182 0 1.7496626983089938e-08
GC_2_183 b_2 NI_2 NS_183 0 -5.6993398672714282e-07
GC_2_184 b_2 NI_2 NS_184 0 -1.6160235178511357e-06
GC_2_185 b_2 NI_2 NS_185 0 -3.1702273622463025e-06
GC_2_186 b_2 NI_2 NS_186 0 6.9325560710329175e-08
GC_2_187 b_2 NI_2 NS_187 0 2.6911099171007857e-07
GC_2_188 b_2 NI_2 NS_188 0 2.5894647212169075e-06
GC_2_189 b_2 NI_2 NS_189 0 -1.1425720951859781e-06
GC_2_190 b_2 NI_2 NS_190 0 -5.5948721066490814e-07
GC_2_191 b_2 NI_2 NS_191 0 -2.6469510324046541e-07
GC_2_192 b_2 NI_2 NS_192 0 1.0907518541197983e-06
GD_2_1 b_2 NI_2 NA_1 0 -1.7151973382174550e-02
GD_2_2 b_2 NI_2 NA_2 0 -3.5122949055498169e-02
GD_2_3 b_2 NI_2 NA_3 0 -5.0305487497640279e-03
GD_2_4 b_2 NI_2 NA_4 0 4.8377374149174467e-03
GD_2_5 b_2 NI_2 NA_5 0 1.5590866541016807e-03
GD_2_6 b_2 NI_2 NA_6 0 1.2308906516978906e-03
GD_2_7 b_2 NI_2 NA_7 0 1.6428450167124597e-04
GD_2_8 b_2 NI_2 NA_8 0 -3.8455892236264884e-04
GD_2_9 b_2 NI_2 NA_9 0 -9.6479955325940167e-06
GD_2_10 b_2 NI_2 NA_10 0 -2.0032116883942280e-05
GD_2_11 b_2 NI_2 NA_11 0 -3.8789059700978260e-06
GD_2_12 b_2 NI_2 NA_12 0 -2.1462240895311929e-06
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 9.7648374106914810e-03
GC_3_2 b_3 NI_3 NS_2 0 -1.3950169916413264e-05
GC_3_3 b_3 NI_3 NS_3 0 2.4707715800740526e-13
GC_3_4 b_3 NI_3 NS_4 0 -3.3612386530048193e-07
GC_3_5 b_3 NI_3 NS_5 0 -1.8185721987205023e-05
GC_3_6 b_3 NI_3 NS_6 0 -4.6198703785336514e-06
GC_3_7 b_3 NI_3 NS_7 0 -1.8582402292284172e-03
GC_3_8 b_3 NI_3 NS_8 0 -1.1618216948709263e-02
GC_3_9 b_3 NI_3 NS_9 0 -2.7110118518508895e-02
GC_3_10 b_3 NI_3 NS_10 0 4.1370426045139038e-03
GC_3_11 b_3 NI_3 NS_11 0 1.3707060537696499e-02
GC_3_12 b_3 NI_3 NS_12 0 3.3729430709231428e-02
GC_3_13 b_3 NI_3 NS_13 0 -1.0121852461970485e-02
GC_3_14 b_3 NI_3 NS_14 0 -1.1019367249036202e-03
GC_3_15 b_3 NI_3 NS_15 0 2.5203472327585030e-02
GC_3_16 b_3 NI_3 NS_16 0 3.4344052433764392e-02
GC_3_17 b_3 NI_3 NS_17 0 -3.7864505499347664e-03
GC_3_18 b_3 NI_3 NS_18 0 -6.7154362288669465e-06
GC_3_19 b_3 NI_3 NS_19 0 2.4804596412669953e-13
GC_3_20 b_3 NI_3 NS_20 0 -1.1920273251330325e-08
GC_3_21 b_3 NI_3 NS_21 0 -4.9382661485630224e-05
GC_3_22 b_3 NI_3 NS_22 0 1.1500073529994178e-05
GC_3_23 b_3 NI_3 NS_23 0 -2.9134861575221215e-03
GC_3_24 b_3 NI_3 NS_24 0 -2.2858689913082680e-03
GC_3_25 b_3 NI_3 NS_25 0 -6.9716553073172292e-03
GC_3_26 b_3 NI_3 NS_26 0 1.0620032540262251e-03
GC_3_27 b_3 NI_3 NS_27 0 -8.3521765523088595e-03
GC_3_28 b_3 NI_3 NS_28 0 3.0378081745053284e-02
GC_3_29 b_3 NI_3 NS_29 0 1.0625811814701919e-02
GC_3_30 b_3 NI_3 NS_30 0 -3.5509049939222589e-04
GC_3_31 b_3 NI_3 NS_31 0 1.6729237124743664e-02
GC_3_32 b_3 NI_3 NS_32 0 7.6374124497311478e-03
GC_3_33 b_3 NI_3 NS_33 0 5.8323406691399717e-02
GC_3_34 b_3 NI_3 NS_34 0 -7.5808535431962536e-06
GC_3_35 b_3 NI_3 NS_35 0 -1.1651066620791375e-12
GC_3_36 b_3 NI_3 NS_36 0 -2.4303493179658623e-06
GC_3_37 b_3 NI_3 NS_37 0 2.8223257415720176e-05
GC_3_38 b_3 NI_3 NS_38 0 -4.6816240376115138e-06
GC_3_39 b_3 NI_3 NS_39 0 -1.5286018201570162e-03
GC_3_40 b_3 NI_3 NS_40 0 7.1114048340669804e-03
GC_3_41 b_3 NI_3 NS_41 0 1.7510183636992454e-02
GC_3_42 b_3 NI_3 NS_42 0 -5.4961710302043210e-03
GC_3_43 b_3 NI_3 NS_43 0 -2.5486250547244849e-02
GC_3_44 b_3 NI_3 NS_44 0 -3.1173404438581194e-02
GC_3_45 b_3 NI_3 NS_45 0 7.4101516417435795e-03
GC_3_46 b_3 NI_3 NS_46 0 2.8759430408195788e-03
GC_3_47 b_3 NI_3 NS_47 0 -3.0809743596175478e-02
GC_3_48 b_3 NI_3 NS_48 0 -3.3522784897376944e-02
GC_3_49 b_3 NI_3 NS_49 0 1.9562356084125260e-01
GC_3_50 b_3 NI_3 NS_50 0 6.0180004206569856e-05
GC_3_51 b_3 NI_3 NS_51 0 3.3868707594450949e-12
GC_3_52 b_3 NI_3 NS_52 0 4.1877026576175170e-06
GC_3_53 b_3 NI_3 NS_53 0 1.2049826642041033e-04
GC_3_54 b_3 NI_3 NS_54 0 4.6653373315862200e-05
GC_3_55 b_3 NI_3 NS_55 0 -6.0782607548995740e-02
GC_3_56 b_3 NI_3 NS_56 0 -4.3809428940219310e-02
GC_3_57 b_3 NI_3 NS_57 0 4.0382961016770469e-02
GC_3_58 b_3 NI_3 NS_58 0 -1.8956105151677057e-02
GC_3_59 b_3 NI_3 NS_59 0 -1.2229035418822104e-01
GC_3_60 b_3 NI_3 NS_60 0 6.7052042723702243e-02
GC_3_61 b_3 NI_3 NS_61 0 -2.3662109318065946e-02
GC_3_62 b_3 NI_3 NS_62 0 1.2239186680645582e-02
GC_3_63 b_3 NI_3 NS_63 0 2.4212271244987888e-02
GC_3_64 b_3 NI_3 NS_64 0 -6.5693184445951153e-02
GC_3_65 b_3 NI_3 NS_65 0 5.5059728758926974e-03
GC_3_66 b_3 NI_3 NS_66 0 7.7003056763413412e-06
GC_3_67 b_3 NI_3 NS_67 0 1.3788105682611864e-13
GC_3_68 b_3 NI_3 NS_68 0 -1.9135926148597598e-07
GC_3_69 b_3 NI_3 NS_69 0 -1.3183572978950604e-05
GC_3_70 b_3 NI_3 NS_70 0 -5.0851346803883278e-07
GC_3_71 b_3 NI_3 NS_71 0 -7.6462493276486664e-04
GC_3_72 b_3 NI_3 NS_72 0 -4.6323643526796415e-03
GC_3_73 b_3 NI_3 NS_73 0 -1.0665727447876918e-02
GC_3_74 b_3 NI_3 NS_74 0 1.5152621532826308e-03
GC_3_75 b_3 NI_3 NS_75 0 4.9161630929859647e-03
GC_3_76 b_3 NI_3 NS_76 0 1.2766052024697019e-02
GC_3_77 b_3 NI_3 NS_77 0 -4.0675830911787846e-03
GC_3_78 b_3 NI_3 NS_78 0 -3.1206461945180607e-04
GC_3_79 b_3 NI_3 NS_79 0 9.4892185162516619e-03
GC_3_80 b_3 NI_3 NS_80 0 1.3304745763606693e-02
GC_3_81 b_3 NI_3 NS_81 0 -1.7394750282459170e-03
GC_3_82 b_3 NI_3 NS_82 0 3.3820024108218562e-06
GC_3_83 b_3 NI_3 NS_83 0 1.4221561786377336e-13
GC_3_84 b_3 NI_3 NS_84 0 3.7243404558652382e-08
GC_3_85 b_3 NI_3 NS_85 0 -1.9140857678055432e-05
GC_3_86 b_3 NI_3 NS_86 0 4.6723282474439848e-06
GC_3_87 b_3 NI_3 NS_87 0 -1.0767884142939338e-03
GC_3_88 b_3 NI_3 NS_88 0 -7.5112565595436510e-04
GC_3_89 b_3 NI_3 NS_89 0 -2.6165140462386690e-03
GC_3_90 b_3 NI_3 NS_90 0 3.9711045629092393e-04
GC_3_91 b_3 NI_3 NS_91 0 -2.9079867602893293e-03
GC_3_92 b_3 NI_3 NS_92 0 1.1463070923586720e-02
GC_3_93 b_3 NI_3 NS_93 0 4.0077366663204437e-03
GC_3_94 b_3 NI_3 NS_94 0 -1.5797382565522114e-04
GC_3_95 b_3 NI_3 NS_95 0 6.2766039080807690e-03
GC_3_96 b_3 NI_3 NS_96 0 2.8067155412053843e-03
GC_3_97 b_3 NI_3 NS_97 0 -4.1487400121279000e-03
GC_3_98 b_3 NI_3 NS_98 0 1.7193164978677300e-06
GC_3_99 b_3 NI_3 NS_99 0 -1.6578376608954608e-13
GC_3_100 b_3 NI_3 NS_100 0 4.6844363960503253e-08
GC_3_101 b_3 NI_3 NS_101 0 1.3494062986328132e-05
GC_3_102 b_3 NI_3 NS_102 0 -3.8201570218822264e-06
GC_3_103 b_3 NI_3 NS_103 0 2.5302390330118924e-05
GC_3_104 b_3 NI_3 NS_104 0 2.4917238882060585e-05
GC_3_105 b_3 NI_3 NS_105 0 -3.8900143121875118e-04
GC_3_106 b_3 NI_3 NS_106 0 3.7410547426011649e-04
GC_3_107 b_3 NI_3 NS_107 0 1.1958345082756299e-03
GC_3_108 b_3 NI_3 NS_108 0 1.9767281416892004e-03
GC_3_109 b_3 NI_3 NS_109 0 1.9599636162518939e-04
GC_3_110 b_3 NI_3 NS_110 0 -2.0844188134892526e-04
GC_3_111 b_3 NI_3 NS_111 0 1.7521895588501427e-03
GC_3_112 b_3 NI_3 NS_112 0 1.3456704349227328e-03
GC_3_113 b_3 NI_3 NS_113 0 -5.1146931124119879e-04
GC_3_114 b_3 NI_3 NS_114 0 -1.3713202396191042e-06
GC_3_115 b_3 NI_3 NS_115 0 -1.6665611673953767e-13
GC_3_116 b_3 NI_3 NS_116 0 2.7367517017034586e-08
GC_3_117 b_3 NI_3 NS_117 0 7.0045548688286295e-06
GC_3_118 b_3 NI_3 NS_118 0 -1.3820748026847916e-06
GC_3_119 b_3 NI_3 NS_119 0 6.7524390376718074e-04
GC_3_120 b_3 NI_3 NS_120 0 5.6582047691683564e-04
GC_3_121 b_3 NI_3 NS_121 0 1.6548660508495900e-03
GC_3_122 b_3 NI_3 NS_122 0 -1.2957952188087502e-04
GC_3_123 b_3 NI_3 NS_123 0 2.1436138342153855e-03
GC_3_124 b_3 NI_3 NS_124 0 -6.5221941112967316e-03
GC_3_125 b_3 NI_3 NS_125 0 -2.2923218245112782e-03
GC_3_126 b_3 NI_3 NS_126 0 2.6317463645827435e-05
GC_3_127 b_3 NI_3 NS_127 0 -3.4016067588201605e-03
GC_3_128 b_3 NI_3 NS_128 0 -1.5787266878925722e-03
GC_3_129 b_3 NI_3 NS_129 0 5.7604004346915882e-04
GC_3_130 b_3 NI_3 NS_130 0 -1.4813960777110783e-07
GC_3_131 b_3 NI_3 NS_131 0 9.3192768226830682e-15
GC_3_132 b_3 NI_3 NS_132 0 -6.6835137527696250e-09
GC_3_133 b_3 NI_3 NS_133 0 -1.5525074440322830e-06
GC_3_134 b_3 NI_3 NS_134 0 4.2140789914091379e-07
GC_3_135 b_3 NI_3 NS_135 0 -7.8445214876517162e-06
GC_3_136 b_3 NI_3 NS_136 0 -3.5375189575536793e-05
GC_3_137 b_3 NI_3 NS_137 0 -2.2999737127103013e-05
GC_3_138 b_3 NI_3 NS_138 0 -4.0669703635933393e-05
GC_3_139 b_3 NI_3 NS_139 0 -1.2953840631552182e-04
GC_3_140 b_3 NI_3 NS_140 0 -1.6494248533207911e-04
GC_3_141 b_3 NI_3 NS_141 0 -5.0630151524382378e-05
GC_3_142 b_3 NI_3 NS_142 0 2.6196934387625631e-05
GC_3_143 b_3 NI_3 NS_143 0 -1.5795927698733793e-04
GC_3_144 b_3 NI_3 NS_144 0 -7.7191734923896398e-05
GC_3_145 b_3 NI_3 NS_145 0 2.1057591362607593e-05
GC_3_146 b_3 NI_3 NS_146 0 -2.2145156693521190e-08
GC_3_147 b_3 NI_3 NS_147 0 9.1433725595179615e-15
GC_3_148 b_3 NI_3 NS_148 0 2.4623325993161368e-09
GC_3_149 b_3 NI_3 NS_149 0 3.6442228414735785e-07
GC_3_150 b_3 NI_3 NS_150 0 -1.2259894704509073e-07
GC_3_151 b_3 NI_3 NS_151 0 1.8634968993929097e-05
GC_3_152 b_3 NI_3 NS_152 0 2.3649325670251776e-05
GC_3_153 b_3 NI_3 NS_153 0 6.0261935646315597e-05
GC_3_154 b_3 NI_3 NS_154 0 -7.0207497398116698e-06
GC_3_155 b_3 NI_3 NS_155 0 7.3285738291032477e-05
GC_3_156 b_3 NI_3 NS_156 0 -2.3641844525980799e-04
GC_3_157 b_3 NI_3 NS_157 0 -8.4900878009855173e-05
GC_3_158 b_3 NI_3 NS_158 0 2.4596682345648682e-06
GC_3_159 b_3 NI_3 NS_159 0 -1.2825114207399451e-04
GC_3_160 b_3 NI_3 NS_160 0 -6.0502595295269267e-05
GC_3_161 b_3 NI_3 NS_161 0 7.9731454759314257e-05
GC_3_162 b_3 NI_3 NS_162 0 5.1635953379931819e-08
GC_3_163 b_3 NI_3 NS_163 0 3.3841296656100783e-15
GC_3_164 b_3 NI_3 NS_164 0 -9.6266628125485731e-10
GC_3_165 b_3 NI_3 NS_165 0 -2.2495943304261879e-07
GC_3_166 b_3 NI_3 NS_166 0 6.5571060238417756e-08
GC_3_167 b_3 NI_3 NS_167 0 -1.4046001763869008e-06
GC_3_168 b_3 NI_3 NS_168 0 -5.7431794053935748e-06
GC_3_169 b_3 NI_3 NS_169 0 -4.3977422177590732e-06
GC_3_170 b_3 NI_3 NS_170 0 -4.7436534555704998e-06
GC_3_171 b_3 NI_3 NS_171 0 -1.6602977539735581e-05
GC_3_172 b_3 NI_3 NS_172 0 -2.2921752740648777e-05
GC_3_173 b_3 NI_3 NS_173 0 -8.1457190079283208e-06
GC_3_174 b_3 NI_3 NS_174 0 4.0119411988132264e-06
GC_3_175 b_3 NI_3 NS_175 0 -2.0849766424135457e-05
GC_3_176 b_3 NI_3 NS_176 0 -8.4226493276852331e-06
GC_3_177 b_3 NI_3 NS_177 0 2.2128193272185825e-05
GC_3_178 b_3 NI_3 NS_178 0 4.4282602397235972e-09
GC_3_179 b_3 NI_3 NS_179 0 3.4030957418704208e-15
GC_3_180 b_3 NI_3 NS_180 0 -3.8797449845179778e-10
GC_3_181 b_3 NI_3 NS_181 0 -4.9135740382524924e-08
GC_3_182 b_3 NI_3 NS_182 0 1.7206599023173059e-08
GC_3_183 b_3 NI_3 NS_183 0 -2.6246965352124099e-06
GC_3_184 b_3 NI_3 NS_184 0 3.2073568575173013e-06
GC_3_185 b_3 NI_3 NS_185 0 3.1794460626145525e-06
GC_3_186 b_3 NI_3 NS_186 0 -1.9239380754105531e-06
GC_3_187 b_3 NI_3 NS_187 0 1.2297205778567671e-06
GC_3_188 b_3 NI_3 NS_188 0 -9.8482058370228647e-06
GC_3_189 b_3 NI_3 NS_189 0 -4.6421411507197074e-06
GC_3_190 b_3 NI_3 NS_190 0 7.9201514683229954e-07
GC_3_191 b_3 NI_3 NS_191 0 -8.4615037617238716e-06
GC_3_192 b_3 NI_3 NS_192 0 -5.5208428344637894e-06
GD_3_1 b_3 NI_3 NA_1 0 4.7466476246351332e-03
GD_3_2 b_3 NI_3 NA_2 0 -5.0216176986334704e-03
GD_3_3 b_3 NI_3 NA_3 0 -3.4686988187583895e-02
GD_3_4 b_3 NI_3 NA_4 0 -1.6361102882565488e-02
GD_3_5 b_3 NI_3 NA_5 0 1.2913596352773402e-03
GD_3_6 b_3 NI_3 NA_6 0 -1.8761857901835087e-03
GD_3_7 b_3 NI_3 NA_7 0 1.2302668352031500e-03
GD_3_8 b_3 NI_3 NA_8 0 1.5551974776624969e-03
GD_3_9 b_3 NI_3 NA_9 0 -1.5086930907280978e-04
GD_3_10 b_3 NI_3 NA_10 0 3.5971411678865617e-05
GD_3_11 b_3 NI_3 NA_11 0 -1.9646822608078837e-05
GD_3_12 b_3 NI_3 NA_12 0 -9.6398942237135826e-06
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 -3.7839449390852996e-03
GC_4_2 b_4 NI_4 NS_2 0 -6.9186104980433934e-06
GC_4_3 b_4 NI_4 NS_3 0 2.4799834514037500e-13
GC_4_4 b_4 NI_4 NS_4 0 -1.1844274244843595e-08
GC_4_5 b_4 NI_4 NS_5 0 -4.9359480046566557e-05
GC_4_6 b_4 NI_4 NS_6 0 1.1494362693597963e-05
GC_4_7 b_4 NI_4 NS_7 0 -2.9134817810958663e-03
GC_4_8 b_4 NI_4 NS_8 0 -2.2859935695321871e-03
GC_4_9 b_4 NI_4 NS_9 0 -6.9716491733392187e-03
GC_4_10 b_4 NI_4 NS_10 0 1.0618189604751857e-03
GC_4_11 b_4 NI_4 NS_11 0 -8.3523650381807004e-03
GC_4_12 b_4 NI_4 NS_12 0 3.0377086952640037e-02
GC_4_13 b_4 NI_4 NS_13 0 1.0625543400098421e-02
GC_4_14 b_4 NI_4 NS_14 0 -3.5514756508324923e-04
GC_4_15 b_4 NI_4 NS_15 0 1.6728102825701925e-02
GC_4_16 b_4 NI_4 NS_16 0 7.6358527932007137e-03
GC_4_17 b_4 NI_4 NS_17 0 9.7641735457100857e-03
GC_4_18 b_4 NI_4 NS_18 0 -1.4036588939224553e-05
GC_4_19 b_4 NI_4 NS_19 0 2.4706433099998979e-13
GC_4_20 b_4 NI_4 NS_20 0 -3.3606478600510438e-07
GC_4_21 b_4 NI_4 NS_21 0 -1.8171421889376461e-05
GC_4_22 b_4 NI_4 NS_22 0 -4.6237964954558327e-06
GC_4_23 b_4 NI_4 NS_23 0 -1.8582493783796225e-03
GC_4_24 b_4 NI_4 NS_24 0 -1.1618241723925509e-02
GC_4_25 b_4 NI_4 NS_25 0 -2.7110129132865500e-02
GC_4_26 b_4 NI_4 NS_26 0 4.1371782480121152e-03
GC_4_27 b_4 NI_4 NS_27 0 1.3707497528372265e-02
GC_4_28 b_4 NI_4 NS_28 0 3.3729532921113595e-02
GC_4_29 b_4 NI_4 NS_29 0 -1.0121852483197882e-02
GC_4_30 b_4 NI_4 NS_30 0 -1.1020398062306675e-03
GC_4_31 b_4 NI_4 NS_31 0 2.5203488101687179e-02
GC_4_32 b_4 NI_4 NS_32 0 3.4343640131753346e-02
GC_4_33 b_4 NI_4 NS_33 0 1.9562848155653287e-01
GC_4_34 b_4 NI_4 NS_34 0 6.1077387469443030e-05
GC_4_35 b_4 NI_4 NS_35 0 3.3873448378780538e-12
GC_4_36 b_4 NI_4 NS_36 0 4.1871623896896527e-06
GC_4_37 b_4 NI_4 NS_37 0 1.2036015569026501e-04
GC_4_38 b_4 NI_4 NS_38 0 4.6690649755276047e-05
GC_4_39 b_4 NI_4 NS_39 0 -6.0783005033423924e-02
GC_4_40 b_4 NI_4 NS_40 0 -4.3809742031978759e-02
GC_4_41 b_4 NI_4 NS_41 0 4.0382339856218495e-02
GC_4_42 b_4 NI_4 NS_42 0 -1.8956381303373671e-02
GC_4_43 b_4 NI_4 NS_43 0 -1.2229370779430254e-01
GC_4_44 b_4 NI_4 NS_44 0 6.7052677818967996e-02
GC_4_45 b_4 NI_4 NS_45 0 -2.3661904996400168e-02
GC_4_46 b_4 NI_4 NS_46 0 1.2240332608872345e-02
GC_4_47 b_4 NI_4 NS_47 0 2.4213659354669289e-02
GC_4_48 b_4 NI_4 NS_48 0 -6.5687878006775474e-02
GC_4_49 b_4 NI_4 NS_49 0 5.8301374366242123e-02
GC_4_50 b_4 NI_4 NS_50 0 -6.5958938437840116e-06
GC_4_51 b_4 NI_4 NS_51 0 -1.1644014447420192e-12
GC_4_52 b_4 NI_4 NS_52 0 -2.4306421993838770e-06
GC_4_53 b_4 NI_4 NS_53 0 2.8124740392901536e-05
GC_4_54 b_4 NI_4 NS_54 0 -4.6581756604053501e-06
GC_4_55 b_4 NI_4 NS_55 0 -1.5282875182670206e-03
GC_4_56 b_4 NI_4 NS_56 0 7.1124137668110510e-03
GC_4_57 b_4 NI_4 NS_57 0 1.7510598110326726e-02
GC_4_58 b_4 NI_4 NS_58 0 -5.4948477996833427e-03
GC_4_59 b_4 NI_4 NS_59 0 -2.5483050190210115e-02
GC_4_60 b_4 NI_4 NS_60 0 -3.1166674146773383e-02
GC_4_61 b_4 NI_4 NS_61 0 7.4119733534026818e-03
GC_4_62 b_4 NI_4 NS_62 0 2.8757205050070826e-03
GC_4_63 b_4 NI_4 NS_63 0 -3.0802277646636841e-02
GC_4_64 b_4 NI_4 NS_64 0 -3.3514439655673370e-02
GC_4_65 b_4 NI_4 NS_65 0 -1.7415731162775110e-03
GC_4_66 b_4 NI_4 NS_66 0 3.4125207230293427e-06
GC_4_67 b_4 NI_4 NS_67 0 1.4221756291631056e-13
GC_4_68 b_4 NI_4 NS_68 0 3.7246154407933652e-08
GC_4_69 b_4 NI_4 NS_69 0 -1.9143093102448636e-05
GC_4_70 b_4 NI_4 NS_70 0 4.6726567242714727e-06
GC_4_71 b_4 NI_4 NS_71 0 -1.0766818057180124e-03
GC_4_72 b_4 NI_4 NS_72 0 -7.5098971709168624e-04
GC_4_73 b_4 NI_4 NS_73 0 -2.6164094661926219e-03
GC_4_74 b_4 NI_4 NS_74 0 3.9728476501588839e-04
GC_4_75 b_4 NI_4 NS_75 0 -2.9072823397682814e-03
GC_4_76 b_4 NI_4 NS_76 0 1.1463294202518738e-02
GC_4_77 b_4 NI_4 NS_77 0 4.0077636705391374e-03
GC_4_78 b_4 NI_4 NS_78 0 -1.5810813680553563e-04
GC_4_79 b_4 NI_4 NS_79 0 6.2769086409219270e-03
GC_4_80 b_4 NI_4 NS_80 0 2.8069235838086926e-03
GC_4_81 b_4 NI_4 NS_81 0 5.5067189090808174e-03
GC_4_82 b_4 NI_4 NS_82 0 7.6561825918766932e-06
GC_4_83 b_4 NI_4 NS_83 0 1.3787682193519536e-13
GC_4_84 b_4 NI_4 NS_84 0 -1.9134190066206083e-07
GC_4_85 b_4 NI_4 NS_85 0 -1.3178647785741413e-05
GC_4_86 b_4 NI_4 NS_86 0 -5.0973861631122062e-07
GC_4_87 b_4 NI_4 NS_87 0 -7.6463907046557967e-04
GC_4_88 b_4 NI_4 NS_88 0 -4.6323923072515878e-03
GC_4_89 b_4 NI_4 NS_89 0 -1.0665738778188804e-02
GC_4_90 b_4 NI_4 NS_90 0 1.5152279248733340e-03
GC_4_91 b_4 NI_4 NS_91 0 4.9160973390964292e-03
GC_4_92 b_4 NI_4 NS_92 0 1.2765826803691161e-02
GC_4_93 b_4 NI_4 NS_93 0 -4.0676473044819377e-03
GC_4_94 b_4 NI_4 NS_94 0 -3.1207217996283315e-04
GC_4_95 b_4 NI_4 NS_95 0 9.4889474925835115e-03
GC_4_96 b_4 NI_4 NS_96 0 1.3304398350845703e-02
GC_4_97 b_4 NI_4 NS_97 0 -5.1130033161060813e-04
GC_4_98 b_4 NI_4 NS_98 0 -1.3817734386130558e-06
GC_4_99 b_4 NI_4 NS_99 0 -1.6665226682355320e-13
GC_4_100 b_4 NI_4 NS_100 0 2.7367877789340959e-08
GC_4_101 b_4 NI_4 NS_101 0 7.0054341237526634e-06
GC_4_102 b_4 NI_4 NS_102 0 -1.3822465654313400e-06
GC_4_103 b_4 NI_4 NS_103 0 6.7524359401272959e-04
GC_4_104 b_4 NI_4 NS_104 0 5.6581489835402787e-04
GC_4_105 b_4 NI_4 NS_105 0 1.6548687999783534e-03
GC_4_106 b_4 NI_4 NS_106 0 -1.2959045235977817e-04
GC_4_107 b_4 NI_4 NS_107 0 2.1435995658111253e-03
GC_4_108 b_4 NI_4 NS_108 0 -6.5222616441435420e-03
GC_4_109 b_4 NI_4 NS_109 0 -2.2923399350525541e-03
GC_4_110 b_4 NI_4 NS_110 0 2.6315054871072358e-05
GC_4_111 b_4 NI_4 NS_111 0 -3.4016800405182596e-03
GC_4_112 b_4 NI_4 NS_112 0 -1.5788172225786213e-03
GC_4_113 b_4 NI_4 NS_113 0 -4.1449869393719819e-03
GC_4_114 b_4 NI_4 NS_114 0 1.7129473952854222e-06
GC_4_115 b_4 NI_4 NS_115 0 -1.6578973815827577e-13
GC_4_116 b_4 NI_4 NS_116 0 4.6844404576536320e-08
GC_4_117 b_4 NI_4 NS_117 0 1.3493702792594351e-05
GC_4_118 b_4 NI_4 NS_118 0 -3.8197835679869641e-06
GC_4_119 b_4 NI_4 NS_119 0 2.5324160430214994e-05
GC_4_120 b_4 NI_4 NS_120 0 2.4694711206584471e-05
GC_4_121 b_4 NI_4 NS_121 0 -3.8938141989306385e-04
GC_4_122 b_4 NI_4 NS_122 0 3.7369321207316575e-04
GC_4_123 b_4 NI_4 NS_123 0 1.1949620601775246e-03
GC_4_124 b_4 NI_4 NS_124 0 1.9764273175164738e-03
GC_4_125 b_4 NI_4 NS_125 0 1.9577966325587759e-04
GC_4_126 b_4 NI_4 NS_126 0 -2.0844091053023761e-04
GC_4_127 b_4 NI_4 NS_127 0 1.7514099721900123e-03
GC_4_128 b_4 NI_4 NS_128 0 1.3454106403367279e-03
GC_4_129 b_4 NI_4 NS_129 0 2.0505590416518784e-05
GC_4_130 b_4 NI_4 NS_130 0 -2.0995411298014870e-08
GC_4_131 b_4 NI_4 NS_131 0 9.1431534381177255e-15
GC_4_132 b_4 NI_4 NS_132 0 2.4616152276017388e-09
GC_4_133 b_4 NI_4 NS_133 0 3.6420323929760343e-07
GC_4_134 b_4 NI_4 NS_134 0 -1.2255232547837352e-07
GC_4_135 b_4 NI_4 NS_135 0 1.8673845006042564e-05
GC_4_136 b_4 NI_4 NS_136 0 2.3690764657373399e-05
GC_4_137 b_4 NI_4 NS_137 0 6.0298818611801796e-05
GC_4_138 b_4 NI_4 NS_138 0 -6.9694932227159132e-06
GC_4_139 b_4 NI_4 NS_139 0 7.3526077034604255e-05
GC_4_140 b_4 NI_4 NS_140 0 -2.3641638520319999e-04
GC_4_141 b_4 NI_4 NS_141 0 -8.4914372069057564e-05
GC_4_142 b_4 NI_4 NS_142 0 2.4070699087038991e-06
GC_4_143 b_4 NI_4 NS_143 0 -1.2822934121510096e-04
GC_4_144 b_4 NI_4 NS_144 0 -6.0525465876309705e-05
GC_4_145 b_4 NI_4 NS_145 0 5.7608712299926851e-04
GC_4_146 b_4 NI_4 NS_146 0 -1.4657538720113676e-07
GC_4_147 b_4 NI_4 NS_147 0 9.3244362446375220e-15
GC_4_148 b_4 NI_4 NS_148 0 -6.6854069528009988e-09
GC_4_149 b_4 NI_4 NS_149 0 -1.5528541112199680e-06
GC_4_150 b_4 NI_4 NS_150 0 4.2151146449172151e-07
GC_4_151 b_4 NI_4 NS_151 0 -7.8459628816333895e-06
GC_4_152 b_4 NI_4 NS_152 0 -3.5377871385670933e-05
GC_4_153 b_4 NI_4 NS_153 0 -2.3002222777271746e-05
GC_4_154 b_4 NI_4 NS_154 0 -4.0672787697076253e-05
GC_4_155 b_4 NI_4 NS_155 0 -1.2955363374967768e-04
GC_4_156 b_4 NI_4 NS_156 0 -1.6495171741352115e-04
GC_4_157 b_4 NI_4 NS_157 0 -5.0632677337053659e-05
GC_4_158 b_4 NI_4 NS_158 0 2.6201006790635310e-05
GC_4_159 b_4 NI_4 NS_159 0 -1.5796651522502229e-04
GC_4_160 b_4 NI_4 NS_160 0 -7.7186979217268526e-05
GC_4_161 b_4 NI_4 NS_161 0 2.2123342510184360e-05
GC_4_162 b_4 NI_4 NS_162 0 4.5798284355211391e-09
GC_4_163 b_4 NI_4 NS_163 0 3.4031120514767904e-15
GC_4_164 b_4 NI_4 NS_164 0 -3.8801598803157943e-10
GC_4_165 b_4 NI_4 NS_165 0 -4.9149252049742241e-08
GC_4_166 b_4 NI_4 NS_166 0 1.7209891608498449e-08
GC_4_167 b_4 NI_4 NS_167 0 -2.6247850986847272e-06
GC_4_168 b_4 NI_4 NS_168 0 3.2078194035874536e-06
GC_4_169 b_4 NI_4 NS_169 0 3.1791708570043097e-06
GC_4_170 b_4 NI_4 NS_170 0 -1.9233723916164756e-06
GC_4_171 b_4 NI_4 NS_171 0 1.2312401531925058e-06
GC_4_172 b_4 NI_4 NS_172 0 -9.8454312541074350e-06
GC_4_173 b_4 NI_4 NS_173 0 -4.6415017676663326e-06
GC_4_174 b_4 NI_4 NS_174 0 7.9166977049050842e-07
GC_4_175 b_4 NI_4 NS_175 0 -8.4595003534193872e-06
GC_4_176 b_4 NI_4 NS_176 0 -5.5193058162914367e-06
GC_4_177 b_4 NI_4 NS_177 0 7.9942180770709573e-05
GC_4_178 b_4 NI_4 NS_178 0 5.1329186929910524e-08
GC_4_179 b_4 NI_4 NS_179 0 3.3842062651454814e-15
GC_4_180 b_4 NI_4 NS_180 0 -9.6515314277463762e-10
GC_4_181 b_4 NI_4 NS_181 0 -2.2531359926897031e-07
GC_4_182 b_4 NI_4 NS_182 0 6.5694107642715574e-08
GC_4_183 b_4 NI_4 NS_183 0 -1.4109178017705114e-06
GC_4_184 b_4 NI_4 NS_184 0 -5.7415831530954746e-06
GC_4_185 b_4 NI_4 NS_185 0 -4.3942322326458739e-06
GC_4_186 b_4 NI_4 NS_186 0 -4.7541768635328064e-06
GC_4_187 b_4 NI_4 NS_187 0 -1.6651202343755399e-05
GC_4_188 b_4 NI_4 NS_188 0 -2.2977720073906725e-05
GC_4_189 b_4 NI_4 NS_189 0 -8.1586047637357114e-06
GC_4_190 b_4 NI_4 NS_190 0 4.0248482463921888e-06
GC_4_191 b_4 NI_4 NS_191 0 -2.0894706630262764e-05
GC_4_192 b_4 NI_4 NS_192 0 -8.4429540324143901e-06
GD_4_1 b_4 NI_4 NA_1 0 -5.0221336123062897e-03
GD_4_2 b_4 NI_4 NA_2 0 4.7468664793699775e-03
GD_4_3 b_4 NI_4 NA_3 0 -1.6363767158787068e-02
GD_4_4 b_4 NI_4 NA_4 0 -3.4680812992563266e-02
GD_4_5 b_4 NI_4 NA_5 0 -1.8755725648373820e-03
GD_4_6 b_4 NI_4 NA_6 0 1.2911314556672557e-03
GD_4_7 b_4 NI_4 NA_7 0 1.5551535630883248e-03
GD_4_8 b_4 NI_4 NA_8 0 1.2291687754269996e-03
GD_4_9 b_4 NI_4 NA_9 0 3.6137654352235634e-05
GD_4_10 b_4 NI_4 NA_10 0 -1.5088503699056530e-04
GD_4_11 b_4 NI_4 NA_11 0 -9.6395207944564733e-06
GD_4_12 b_4 NI_4 NA_12 0 -1.9743730400752342e-05
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 -4.0763653387725649e-03
GC_5_2 b_5 NI_5 NS_2 0 -3.5139348332274457e-06
GC_5_3 b_5 NI_5 NS_3 0 -1.6899825251860125e-13
GC_5_4 b_5 NI_5 NS_4 0 4.8319702941714611e-08
GC_5_5 b_5 NI_5 NS_5 0 1.4111631685868131e-05
GC_5_6 b_5 NI_5 NS_6 0 -3.9679104081922691e-06
GC_5_7 b_5 NI_5 NS_7 0 2.4210966477969433e-05
GC_5_8 b_5 NI_5 NS_8 0 2.1746593940544978e-05
GC_5_9 b_5 NI_5 NS_9 0 -3.9069639079732067e-04
GC_5_10 b_5 NI_5 NS_10 0 3.7012317478493629e-04
GC_5_11 b_5 NI_5 NS_11 0 1.1892433534129369e-03
GC_5_12 b_5 NI_5 NS_12 0 1.9567873156449284e-03
GC_5_13 b_5 NI_5 NS_13 0 1.9071182493844073e-04
GC_5_14 b_5 NI_5 NS_14 0 -2.0993332542062923e-04
GC_5_15 b_5 NI_5 NS_15 0 1.7254227799217326e-03
GC_5_16 b_5 NI_5 NS_16 0 1.3072469071806700e-03
GC_5_17 b_5 NI_5 NS_17 0 -5.4094483352683524e-04
GC_5_18 b_5 NI_5 NS_18 0 3.1248433582921028e-06
GC_5_19 b_5 NI_5 NS_19 0 -1.6762035653362286e-13
GC_5_20 b_5 NI_5 NS_20 0 2.8394452945125541e-08
GC_5_21 b_5 NI_5 NS_21 0 6.6558991447301758e-06
GC_5_22 b_5 NI_5 NS_22 0 -1.3310382425310942e-06
GC_5_23 b_5 NI_5 NS_23 0 6.7451075762788742e-04
GC_5_24 b_5 NI_5 NS_24 0 5.6659219251695158e-04
GC_5_25 b_5 NI_5 NS_25 0 1.6536844107728401e-03
GC_5_26 b_5 NI_5 NS_26 0 -1.2725809781370049e-04
GC_5_27 b_5 NI_5 NS_27 0 2.1416290515703170e-03
GC_5_28 b_5 NI_5 NS_28 0 -6.5096279269541797e-03
GC_5_29 b_5 NI_5 NS_29 0 -2.2901168124610204e-03
GC_5_30 b_5 NI_5 NS_30 0 2.9660962847864953e-05
GC_5_31 b_5 NI_5 NS_31 0 -3.3826735446881081e-03
GC_5_32 b_5 NI_5 NS_32 0 -1.5439577966785813e-03
GC_5_33 b_5 NI_5 NS_33 0 5.5385161382722359e-03
GC_5_34 b_5 NI_5 NS_34 0 4.5230412917922440e-06
GC_5_35 b_5 NI_5 NS_35 0 1.3658682821442897e-13
GC_5_36 b_5 NI_5 NS_36 0 -1.9080451634611999e-07
GC_5_37 b_5 NI_5 NS_37 0 -1.2843237619562489e-05
GC_5_38 b_5 NI_5 NS_38 0 -5.8655436963370832e-07
GC_5_39 b_5 NI_5 NS_39 0 -7.6459481479012562e-04
GC_5_40 b_5 NI_5 NS_40 0 -4.6329858120412017e-03
GC_5_41 b_5 NI_5 NS_41 0 -1.0664636556693974e-02
GC_5_42 b_5 NI_5 NS_42 0 1.5135464030223223e-03
GC_5_43 b_5 NI_5 NS_43 0 4.9164642827145347e-03
GC_5_44 b_5 NI_5 NS_44 0 1.2751636673708181e-02
GC_5_45 b_5 NI_5 NS_45 0 -4.0714540431925532e-03
GC_5_46 b_5 NI_5 NS_46 0 -3.1361281887545080e-04
GC_5_47 b_5 NI_5 NS_47 0 9.4726823165253177e-03
GC_5_48 b_5 NI_5 NS_48 0 1.3280331546763278e-02
GC_5_49 b_5 NI_5 NS_49 0 -1.7172133359548980e-03
GC_5_50 b_5 NI_5 NS_50 0 1.5931896308230462e-06
GC_5_51 b_5 NI_5 NS_51 0 1.3969585181210695e-13
GC_5_52 b_5 NI_5 NS_52 0 3.6465151148243075e-08
GC_5_53 b_5 NI_5 NS_53 0 -1.9056237856352661e-05
GC_5_54 b_5 NI_5 NS_54 0 4.6709530091138251e-06
GC_5_55 b_5 NI_5 NS_55 0 -1.0758999196700762e-03
GC_5_56 b_5 NI_5 NS_56 0 -7.5179350170314848e-04
GC_5_57 b_5 NI_5 NS_57 0 -2.6152298657685477e-03
GC_5_58 b_5 NI_5 NS_58 0 3.9480670084080682e-04
GC_5_59 b_5 NI_5 NS_59 0 -2.9090022692853561e-03
GC_5_60 b_5 NI_5 NS_60 0 1.1450220710031891e-02
GC_5_61 b_5 NI_5 NS_61 0 4.0044822663212083e-03
GC_5_62 b_5 NI_5 NS_62 0 -1.5873432955014659e-04
GC_5_63 b_5 NI_5 NS_63 0 6.2634728085072030e-03
GC_5_64 b_5 NI_5 NS_64 0 2.7899590994231241e-03
GC_5_65 b_5 NI_5 NS_65 0 5.8537658927887065e-02
GC_5_66 b_5 NI_5 NS_66 0 -2.0388009772182726e-05
GC_5_67 b_5 NI_5 NS_67 0 -1.1567285171598091e-12
GC_5_68 b_5 NI_5 NS_68 0 -2.4256583334623104e-06
GC_5_69 b_5 NI_5 NS_69 0 2.9536350536354070e-05
GC_5_70 b_5 NI_5 NS_70 0 -5.0078894898160047e-06
GC_5_71 b_5 NI_5 NS_71 0 -1.5267425713731059e-03
GC_5_72 b_5 NI_5 NS_72 0 7.1024057181454173e-03
GC_5_73 b_5 NI_5 NS_73 0 1.7512566485903790e-02
GC_5_74 b_5 NI_5 NS_74 0 -5.5132440246384480e-03
GC_5_75 b_5 NI_5 NS_75 0 -2.5510613500844239e-02
GC_5_76 b_5 NI_5 NS_76 0 -3.1264056589822863e-02
GC_5_77 b_5 NI_5 NS_77 0 7.3860029435363905e-03
GC_5_78 b_5 NI_5 NS_78 0 2.8755768030010614e-03
GC_5_79 b_5 NI_5 NS_79 0 -3.0902425657618058e-02
GC_5_80 b_5 NI_5 NS_80 0 -3.3632074607379311e-02
GC_5_81 b_5 NI_5 NS_81 0 1.9575295540411958e-01
GC_5_82 b_5 NI_5 NS_82 0 7.3939749184435461e-05
GC_5_83 b_5 NI_5 NS_83 0 3.8301347563717560e-12
GC_5_84 b_5 NI_5 NS_84 0 4.1282406258349754e-06
GC_5_85 b_5 NI_5 NS_85 0 1.1732974204500372e-04
GC_5_86 b_5 NI_5 NS_86 0 4.7766712965404776e-05
GC_5_87 b_5 NI_5 NS_87 0 -6.0787496810176464e-02
GC_5_88 b_5 NI_5 NS_88 0 -4.3818095864065605e-02
GC_5_89 b_5 NI_5 NS_89 0 4.0371785527266071e-02
GC_5_90 b_5 NI_5 NS_90 0 -1.8968571932595903e-02
GC_5_91 b_5 NI_5 NS_91 0 -1.2235626855643199e-01
GC_5_92 b_5 NI_5 NS_92 0 6.7044071632756039e-02
GC_5_93 b_5 NI_5 NS_93 0 -2.3662993117698979e-02
GC_5_94 b_5 NI_5 NS_94 0 1.2258422602092907e-02
GC_5_95 b_5 NI_5 NS_95 0 2.4212693164183036e-02
GC_5_96 b_5 NI_5 NS_96 0 -6.5629641125533031e-02
GC_5_97 b_5 NI_5 NS_97 0 1.0071526244156493e-02
GC_5_98 b_5 NI_5 NS_98 0 2.1084150628403430e-05
GC_5_99 b_5 NI_5 NS_99 0 2.4087196885088366e-13
GC_5_100 b_5 NI_5 NS_100 0 -3.5278817335385110e-07
GC_5_101 b_5 NI_5 NS_101 0 -2.4087861053678260e-05
GC_5_102 b_5 NI_5 NS_102 0 -3.1646292520566965e-06
GC_5_103 b_5 NI_5 NS_103 0 -1.8595033358923571e-03
GC_5_104 b_5 NI_5 NS_104 0 -1.1634093339683762e-02
GC_5_105 b_5 NI_5 NS_105 0 -2.7106536489944585e-02
GC_5_106 b_5 NI_5 NS_106 0 4.0963638759228078e-03
GC_5_107 b_5 NI_5 NS_107 0 1.3532831207454415e-02
GC_5_108 b_5 NI_5 NS_108 0 3.3625063031517070e-02
GC_5_109 b_5 NI_5 NS_109 0 -1.0133837700454989e-02
GC_5_110 b_5 NI_5 NS_110 0 -1.0505317877471236e-03
GC_5_111 b_5 NI_5 NS_111 0 2.5156734089856313e-02
GC_5_112 b_5 NI_5 NS_112 0 3.4474351496079421e-02
GC_5_113 b_5 NI_5 NS_113 0 -3.7912039552583333e-03
GC_5_114 b_5 NI_5 NS_114 0 3.2656133834399968e-06
GC_5_115 b_5 NI_5 NS_115 0 2.5082678200111126e-13
GC_5_116 b_5 NI_5 NS_116 0 -8.2146112456222347e-09
GC_5_117 b_5 NI_5 NS_117 0 -4.9981286442089525e-05
GC_5_118 b_5 NI_5 NS_118 0 1.1524744131101951e-05
GC_5_119 b_5 NI_5 NS_119 0 -2.9275852730946093e-03
GC_5_120 b_5 NI_5 NS_120 0 -2.2944158380212277e-03
GC_5_121 b_5 NI_5 NS_121 0 -7.0008796323093037e-03
GC_5_122 b_5 NI_5 NS_122 0 1.0673522722546185e-03
GC_5_123 b_5 NI_5 NS_123 0 -8.4047449712130323e-03
GC_5_124 b_5 NI_5 NS_124 0 3.0494357310913295e-02
GC_5_125 b_5 NI_5 NS_125 0 1.0663377904983239e-02
GC_5_126 b_5 NI_5 NS_126 0 -3.4370441218192603e-04
GC_5_127 b_5 NI_5 NS_127 0 1.6815967372478730e-02
GC_5_128 b_5 NI_5 NS_128 0 7.7403477933141685e-03
GC_5_129 b_5 NI_5 NS_129 0 -4.1500710408769823e-03
GC_5_130 b_5 NI_5 NS_130 0 1.7940325096409642e-06
GC_5_131 b_5 NI_5 NS_131 0 -1.6635552629891633e-13
GC_5_132 b_5 NI_5 NS_132 0 4.6897986149808275e-08
GC_5_133 b_5 NI_5 NS_133 0 1.3507565373324364e-05
GC_5_134 b_5 NI_5 NS_134 0 -3.8248277683899741e-06
GC_5_135 b_5 NI_5 NS_135 0 2.5129768200461989e-05
GC_5_136 b_5 NI_5 NS_136 0 2.4986208653677653e-05
GC_5_137 b_5 NI_5 NS_137 0 -3.8959401642085209e-04
GC_5_138 b_5 NI_5 NS_138 0 3.7424071971237300e-04
GC_5_139 b_5 NI_5 NS_139 0 1.1957864592344921e-03
GC_5_140 b_5 NI_5 NS_140 0 1.9797515887772029e-03
GC_5_141 b_5 NI_5 NS_141 0 1.9676164885307554e-04
GC_5_142 b_5 NI_5 NS_142 0 -2.0869747082758377e-04
GC_5_143 b_5 NI_5 NS_143 0 1.7539303692297207e-03
GC_5_144 b_5 NI_5 NS_144 0 1.3471568970169951e-03
GC_5_145 b_5 NI_5 NS_145 0 -5.1277254593000031e-04
GC_5_146 b_5 NI_5 NS_146 0 -1.3843023661016740e-06
GC_5_147 b_5 NI_5 NS_147 0 -1.6603134503163032e-13
GC_5_148 b_5 NI_5 NS_148 0 2.8234118983723228e-08
GC_5_149 b_5 NI_5 NS_149 0 7.0653671823848493e-06
GC_5_150 b_5 NI_5 NS_150 0 -1.4078477155185409e-06
GC_5_151 b_5 NI_5 NS_151 0 6.7492468846949791e-04
GC_5_152 b_5 NI_5 NS_152 0 5.6564968133218218e-04
GC_5_153 b_5 NI_5 NS_153 0 1.6543010065692304e-03
GC_5_154 b_5 NI_5 NS_154 0 -1.2917071477193303e-04
GC_5_155 b_5 NI_5 NS_155 0 2.1438548170665517e-03
GC_5_156 b_5 NI_5 NS_156 0 -6.5202425607100130e-03
GC_5_157 b_5 NI_5 NS_157 0 -2.2919645667916870e-03
GC_5_158 b_5 NI_5 NS_158 0 2.6323740064751714e-05
GC_5_159 b_5 NI_5 NS_159 0 -3.4000915494027894e-03
GC_5_160 b_5 NI_5 NS_160 0 -1.5774047270223977e-03
GC_5_161 b_5 NI_5 NS_161 0 1.4525536737689786e-03
GC_5_162 b_5 NI_5 NS_162 0 8.9304084995018697e-07
GC_5_163 b_5 NI_5 NS_163 0 2.0219508824777049e-14
GC_5_164 b_5 NI_5 NS_164 0 -1.6569490931906633e-08
GC_5_165 b_5 NI_5 NS_165 0 -3.9771659840526025e-06
GC_5_166 b_5 NI_5 NS_166 0 1.0552127314452128e-06
GC_5_167 b_5 NI_5 NS_167 0 -1.9285722373561981e-05
GC_5_168 b_5 NI_5 NS_168 0 -8.7861953718919571e-05
GC_5_169 b_5 NI_5 NS_169 0 -5.4556889046112666e-05
GC_5_170 b_5 NI_5 NS_170 0 -1.0426357691411932e-04
GC_5_171 b_5 NI_5 NS_171 0 -3.2908308903828015e-04
GC_5_172 b_5 NI_5 NS_172 0 -4.2217089376874275e-04
GC_5_173 b_5 NI_5 NS_173 0 -1.2813169600824382e-04
GC_5_174 b_5 NI_5 NS_174 0 6.5944966670752970e-05
GC_5_175 b_5 NI_5 NS_175 0 -4.0283639525851765e-04
GC_5_176 b_5 NI_5 NS_176 0 -1.9319047502036491e-04
GC_5_177 b_5 NI_5 NS_177 0 -1.1963877726773978e-04
GC_5_178 b_5 NI_5 NS_178 0 1.2452241486579756e-07
GC_5_179 b_5 NI_5 NS_179 0 2.0815846885684131e-14
GC_5_180 b_5 NI_5 NS_180 0 5.2285548279704039e-09
GC_5_181 b_5 NI_5 NS_181 0 7.8192406376958070e-07
GC_5_182 b_5 NI_5 NS_182 0 -2.5030431122986106e-07
GC_5_183 b_5 NI_5 NS_183 0 6.1048697813348624e-05
GC_5_184 b_5 NI_5 NS_184 0 6.1343120614884141e-05
GC_5_185 b_5 NI_5 NS_185 0 1.6080265319562705e-04
GC_5_186 b_5 NI_5 NS_186 0 -4.4905725710010854e-06
GC_5_187 b_5 NI_5 NS_187 0 2.3841019574454456e-04
GC_5_188 b_5 NI_5 NS_188 0 -5.9913596968895792e-04
GC_5_189 b_5 NI_5 NS_189 0 -2.1651523940410662e-04
GC_5_190 b_5 NI_5 NS_190 0 -4.4588826360912313e-06
GC_5_191 b_5 NI_5 NS_191 0 -3.1116195383081935e-04
GC_5_192 b_5 NI_5 NS_192 0 -1.5141376997596952e-04
GD_5_1 b_5 NI_5 NA_1 0 1.2095415203192497e-03
GD_5_2 b_5 NI_5 NA_2 0 1.5614565093467253e-03
GD_5_3 b_5 NI_5 NA_3 0 1.2828177330910370e-03
GD_5_4 b_5 NI_5 NA_4 0 -1.8797067338259944e-03
GD_5_5 b_5 NI_5 NA_5 0 -3.4735129975975103e-02
GD_5_6 b_5 NI_5 NA_6 0 -1.6409284326495032e-02
GD_5_7 b_5 NI_5 NA_7 0 4.6641448803460221e-03
GD_5_8 b_5 NI_5 NA_8 0 -5.0537222907538256e-03
GD_5_9 b_5 NI_5 NA_9 0 1.2297204792298996e-03
GD_5_10 b_5 NI_5 NA_10 0 1.5552933131317236e-03
GD_5_11 b_5 NI_5 NA_11 0 -3.7876040402757736e-04
GD_5_12 b_5 NI_5 NA_12 0 1.6455497398053259e-04
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 -5.4146559672623286e-04
GC_6_2 b_6 NI_6 NS_2 0 3.1760437237749666e-06
GC_6_3 b_6 NI_6 NS_3 0 -1.6761063423177138e-13
GC_6_4 b_6 NI_6 NS_4 0 2.8375037368408354e-08
GC_6_5 b_6 NI_6 NS_5 0 6.6499091738928987e-06
GC_6_6 b_6 NI_6 NS_6 0 -1.3295516086108136e-06
GC_6_7 b_6 NI_6 NS_7 0 6.7450496769566679e-04
GC_6_8 b_6 NI_6 NS_8 0 5.6662005922094834e-04
GC_6_9 b_6 NI_6 NS_9 0 1.6536696433882472e-03
GC_6_10 b_6 NI_6 NS_10 0 -1.2722222905281523e-04
GC_6_11 b_6 NI_6 NS_11 0 2.1416409525165099e-03
GC_6_12 b_6 NI_6 NS_12 0 -6.5093649826568224e-03
GC_6_13 b_6 NI_6 NS_13 0 -2.2900445465715374e-03
GC_6_14 b_6 NI_6 NS_14 0 2.9679822683144175e-05
GC_6_15 b_6 NI_6 NS_15 0 -3.3823944254563589e-03
GC_6_16 b_6 NI_6 NS_16 0 -1.5435667976631366e-03
GC_6_17 b_6 NI_6 NS_17 0 -4.0732060081252359e-03
GC_6_18 b_6 NI_6 NS_18 0 -3.4916088182687536e-06
GC_6_19 b_6 NI_6 NS_19 0 -1.6900737396596312e-13
GC_6_20 b_6 NI_6 NS_20 0 4.8312923900474634e-08
GC_6_21 b_6 NI_6 NS_21 0 1.4108786442895083e-05
GC_6_22 b_6 NI_6 NS_22 0 -3.9669647795047416e-06
GC_6_23 b_6 NI_6 NS_23 0 2.4230833846656203e-05
GC_6_24 b_6 NI_6 NS_24 0 2.1547153020919787e-05
GC_6_25 b_6 NI_6 NS_25 0 -3.9108099861043884e-04
GC_6_26 b_6 NI_6 NS_26 0 3.6975939016540296e-04
GC_6_27 b_6 NI_6 NS_27 0 1.1884428190581454e-03
GC_6_28 b_6 NI_6 NS_28 0 1.9567241004904692e-03
GC_6_29 b_6 NI_6 NS_29 0 1.9056063253560722e-04
GC_6_30 b_6 NI_6 NS_30 0 -2.0992903504981041e-04
GC_6_31 b_6 NI_6 NS_31 0 1.7248954903859852e-03
GC_6_32 b_6 NI_6 NS_32 0 1.3072609843563247e-03
GC_6_33 b_6 NI_6 NS_33 0 -1.7197237980441339e-03
GC_6_34 b_6 NI_6 NS_34 0 1.5791064733495147e-06
GC_6_35 b_6 NI_6 NS_35 0 1.3970246862903815e-13
GC_6_36 b_6 NI_6 NS_36 0 3.6508556705444068e-08
GC_6_37 b_6 NI_6 NS_37 0 -1.9050792093320600e-05
GC_6_38 b_6 NI_6 NS_38 0 4.6690697078006420e-06
GC_6_39 b_6 NI_6 NS_39 0 -1.0757685111630316e-03
GC_6_40 b_6 NI_6 NS_40 0 -7.5163352165709429e-04
GC_6_41 b_6 NI_6 NS_41 0 -2.6150853641977285e-03
GC_6_42 b_6 NI_6 NS_42 0 3.9500820009947521e-04
GC_6_43 b_6 NI_6 NS_43 0 -2.9080754848283415e-03
GC_6_44 b_6 NI_6 NS_44 0 1.1450433894163439e-02
GC_6_45 b_6 NI_6 NS_45 0 4.0044997410041390e-03
GC_6_46 b_6 NI_6 NS_46 0 -1.5893614687911110e-04
GC_6_47 b_6 NI_6 NS_47 0 6.2637366615422869e-03
GC_6_48 b_6 NI_6 NS_48 0 2.7899181266351912e-03
GC_6_49 b_6 NI_6 NS_49 0 5.5395688735192803e-03
GC_6_50 b_6 NI_6 NS_50 0 4.3928091167434147e-06
GC_6_51 b_6 NI_6 NS_51 0 1.3659183257768064e-13
GC_6_52 b_6 NI_6 NS_52 0 -1.9073604098284677e-07
GC_6_53 b_6 NI_6 NS_53 0 -1.2826196814400369e-05
GC_6_54 b_6 NI_6 NS_54 0 -5.9106962017271866e-07
GC_6_55 b_6 NI_6 NS_55 0 -7.6457529430407024e-04
GC_6_56 b_6 NI_6 NS_56 0 -4.6330169791555884e-03
GC_6_57 b_6 NI_6 NS_57 0 -1.0664585761645686e-02
GC_6_58 b_6 NI_6 NS_58 0 1.5134775310145991e-03
GC_6_59 b_6 NI_6 NS_59 0 4.9165148992001686e-03
GC_6_60 b_6 NI_6 NS_60 0 1.2751053167238327e-02
GC_6_61 b_6 NI_6 NS_61 0 -4.0716158696530655e-03
GC_6_62 b_6 NI_6 NS_62 0 -3.1367226351607038e-04
GC_6_63 b_6 NI_6 NS_63 0 9.4720602982644887e-03
GC_6_64 b_6 NI_6 NS_64 0 1.3279388589707541e-02
GC_6_65 b_6 NI_6 NS_65 0 1.9575395696798198e-01
GC_6_66 b_6 NI_6 NS_66 0 7.4166032220168192e-05
GC_6_67 b_6 NI_6 NS_67 0 3.8299419875466449e-12
GC_6_68 b_6 NI_6 NS_68 0 4.1281014925933240e-06
GC_6_69 b_6 NI_6 NS_69 0 1.1729456148166728e-04
GC_6_70 b_6 NI_6 NS_70 0 4.7776279431484439e-05
GC_6_71 b_6 NI_6 NS_71 0 -6.0787587721326752e-02
GC_6_72 b_6 NI_6 NS_72 0 -4.3818170835032130e-02
GC_6_73 b_6 NI_6 NS_73 0 4.0371632540314374e-02
GC_6_74 b_6 NI_6 NS_74 0 -1.8968636353113282e-02
GC_6_75 b_6 NI_6 NS_75 0 -1.2235705452545932e-01
GC_6_76 b_6 NI_6 NS_76 0 6.7044273234643820e-02
GC_6_77 b_6 NI_6 NS_77 0 -2.3662931128732426e-02
GC_6_78 b_6 NI_6 NS_78 0 1.2258694307250698e-02
GC_6_79 b_6 NI_6 NS_79 0 2.4213073418292090e-02
GC_6_80 b_6 NI_6 NS_80 0 -6.5628303396243690e-02
GC_6_81 b_6 NI_6 NS_81 0 5.8532742773130454e-02
GC_6_82 b_6 NI_6 NS_82 0 -2.0119458561819157e-05
GC_6_83 b_6 NI_6 NS_83 0 -1.1567031082383423e-12
GC_6_84 b_6 NI_6 NS_84 0 -2.4257595172674199e-06
GC_6_85 b_6 NI_6 NS_85 0 2.9507210027870855e-05
GC_6_86 b_6 NI_6 NS_86 0 -5.0006615694717762e-06
GC_6_87 b_6 NI_6 NS_87 0 -1.5266966554140784e-03
GC_6_88 b_6 NI_6 NS_88 0 7.1026253952755922e-03
GC_6_89 b_6 NI_6 NS_89 0 1.7512621183351670e-02
GC_6_90 b_6 NI_6 NS_90 0 -5.5129412213007203e-03
GC_6_91 b_6 NI_6 NS_91 0 -2.5510020506769926e-02
GC_6_92 b_6 NI_6 NS_92 0 -3.1262396399761687e-02
GC_6_93 b_6 NI_6 NS_93 0 7.3864564354098718e-03
GC_6_94 b_6 NI_6 NS_94 0 2.8755704951028515e-03
GC_6_95 b_6 NI_6 NS_95 0 -3.0900595347686327e-02
GC_6_96 b_6 NI_6 NS_96 0 -3.3629886042504241e-02
GC_6_97 b_6 NI_6 NS_97 0 -3.7913520091602164e-03
GC_6_98 b_6 NI_6 NS_98 0 3.3233149503298840e-06
GC_6_99 b_6 NI_6 NS_99 0 2.5083441167323432e-13
GC_6_100 b_6 NI_6 NS_100 0 -8.2147712466770783e-09
GC_6_101 b_6 NI_6 NS_101 0 -4.9985665160069748e-05
GC_6_102 b_6 NI_6 NS_102 0 1.1525537953983220e-05
GC_6_103 b_6 NI_6 NS_103 0 -2.9276238381579136e-03
GC_6_104 b_6 NI_6 NS_104 0 -2.2944413750390401e-03
GC_6_105 b_6 NI_6 NS_105 0 -7.0009378472657554e-03
GC_6_106 b_6 NI_6 NS_106 0 1.0673288390555967e-03
GC_6_107 b_6 NI_6 NS_107 0 -8.4050409000749459e-03
GC_6_108 b_6 NI_6 NS_108 0 3.0494693220933771e-02
GC_6_109 b_6 NI_6 NS_109 0 1.0663499124809938e-02
GC_6_110 b_6 NI_6 NS_110 0 -3.4360435677023067e-04
GC_6_111 b_6 NI_6 NS_111 0 1.6816338560419350e-02
GC_6_112 b_6 NI_6 NS_112 0 7.7408941989288334e-03
GC_6_113 b_6 NI_6 NS_113 0 1.0072816321015931e-02
GC_6_114 b_6 NI_6 NS_114 0 2.0970404497041843e-05
GC_6_115 b_6 NI_6 NS_115 0 2.4085958215106238e-13
GC_6_116 b_6 NI_6 NS_116 0 -3.5273811096849074e-07
GC_6_117 b_6 NI_6 NS_117 0 -2.4073954652708381e-05
GC_6_118 b_6 NI_6 NS_118 0 -3.1682009090150003e-06
GC_6_119 b_6 NI_6 NS_119 0 -1.8595028682194901e-03
GC_6_120 b_6 NI_6 NS_120 0 -1.1634140396617225e-02
GC_6_121 b_6 NI_6 NS_121 0 -2.7106519416890743e-02
GC_6_122 b_6 NI_6 NS_122 0 4.0962883160134142e-03
GC_6_123 b_6 NI_6 NS_123 0 1.3532789778050853e-02
GC_6_124 b_6 NI_6 NS_124 0 3.3624518934004137e-02
GC_6_125 b_6 NI_6 NS_125 0 -1.0133989089814017e-02
GC_6_126 b_6 NI_6 NS_126 0 -1.0505708550928138e-03
GC_6_127 b_6 NI_6 NS_127 0 2.5156127338384283e-02
GC_6_128 b_6 NI_6 NS_128 0 3.4473497085125149e-02
GC_6_129 b_6 NI_6 NS_129 0 -5.1252127182538896e-04
GC_6_130 b_6 NI_6 NS_130 0 -1.3427328803198571e-06
GC_6_131 b_6 NI_6 NS_131 0 -1.6602276245863333e-13
GC_6_132 b_6 NI_6 NS_132 0 2.8202933506247177e-08
GC_6_133 b_6 NI_6 NS_133 0 7.0587523171020503e-06
GC_6_134 b_6 NI_6 NS_134 0 -1.4060017667636877e-06
GC_6_135 b_6 NI_6 NS_135 0 6.7490313306143744e-04
GC_6_136 b_6 NI_6 NS_136 0 5.6563343429419984e-04
GC_6_137 b_6 NI_6 NS_137 0 1.6542673284142980e-03
GC_6_138 b_6 NI_6 NS_138 0 -1.2918567096974109e-04
GC_6_139 b_6 NI_6 NS_139 0 2.1436814047246116e-03
GC_6_140 b_6 NI_6 NS_140 0 -6.5201950222599581e-03
GC_6_141 b_6 NI_6 NS_141 0 -2.2919461022020064e-03
GC_6_142 b_6 NI_6 NS_142 0 2.6379128309586032e-05
GC_6_143 b_6 NI_6 NS_143 0 -3.4000186248513437e-03
GC_6_144 b_6 NI_6 NS_144 0 -1.5771548334244927e-03
GC_6_145 b_6 NI_6 NS_145 0 -4.1542515688878920e-03
GC_6_146 b_6 NI_6 NS_146 0 1.7845927280279916e-06
GC_6_147 b_6 NI_6 NS_147 0 -1.6637498190128177e-13
GC_6_148 b_6 NI_6 NS_148 0 4.6912660040297892e-08
GC_6_149 b_6 NI_6 NS_149 0 1.3511196468844381e-05
GC_6_150 b_6 NI_6 NS_150 0 -3.8261379519195227e-06
GC_6_151 b_6 NI_6 NS_151 0 2.5123759731639439e-05
GC_6_152 b_6 NI_6 NS_152 0 2.5233955050616002e-05
GC_6_153 b_6 NI_6 NS_153 0 -3.8918595434675484e-04
GC_6_154 b_6 NI_6 NS_154 0 3.7467879440021594e-04
GC_6_155 b_6 NI_6 NS_155 0 1.1967986417549927e-03
GC_6_156 b_6 NI_6 NS_156 0 1.9801166379177712e-03
GC_6_157 b_6 NI_6 NS_157 0 1.9699694104930398e-04
GC_6_158 b_6 NI_6 NS_158 0 -2.0873490594940674e-04
GC_6_159 b_6 NI_6 NS_159 0 1.7547643193868952e-03
GC_6_160 b_6 NI_6 NS_160 0 1.3473597355883266e-03
GC_6_161 b_6 NI_6 NS_161 0 -1.1829039458612943e-04
GC_6_162 b_6 NI_6 NS_162 0 1.2953080107911514e-07
GC_6_163 b_6 NI_6 NS_163 0 2.0814811157491536e-14
GC_6_164 b_6 NI_6 NS_164 0 5.2259452401831932e-09
GC_6_165 b_6 NI_6 NS_165 0 7.8147385668177182e-07
GC_6_166 b_6 NI_6 NS_166 0 -2.5015462934925478e-07
GC_6_167 b_6 NI_6 NS_167 0 6.0947529746893363e-05
GC_6_168 b_6 NI_6 NS_168 0 6.1240344394195240e-05
GC_6_169 b_6 NI_6 NS_169 0 1.6070446822273813e-04
GC_6_170 b_6 NI_6 NS_170 0 -4.6172872028432151e-06
GC_6_171 b_6 NI_6 NS_171 0 2.3779234183976140e-04
GC_6_172 b_6 NI_6 NS_172 0 -5.9909776838191185e-04
GC_6_173 b_6 NI_6 NS_173 0 -2.1646890142746104e-04
GC_6_174 b_6 NI_6 NS_174 0 -4.3225076062364064e-06
GC_6_175 b_6 NI_6 NS_175 0 -3.1117682937502046e-04
GC_6_176 b_6 NI_6 NS_176 0 -1.5129599845809406e-04
GC_6_177 b_6 NI_6 NS_177 0 1.4526940385347262e-03
GC_6_178 b_6 NI_6 NS_178 0 8.8654393993482139e-07
GC_6_179 b_6 NI_6 NS_179 0 2.0222904792021602e-14
GC_6_180 b_6 NI_6 NS_180 0 -1.6567983043345655e-08
GC_6_181 b_6 NI_6 NS_181 0 -3.9765621741093888e-06
GC_6_182 b_6 NI_6 NS_182 0 1.0550775344938051e-06
GC_6_183 b_6 NI_6 NS_183 0 -1.9289550089934166e-05
GC_6_184 b_6 NI_6 NS_184 0 -8.7869552439668794e-05
GC_6_185 b_6 NI_6 NS_185 0 -5.4561607281090210e-05
GC_6_186 b_6 NI_6 NS_186 0 -1.0426629475924924e-04
GC_6_187 b_6 NI_6 NS_187 0 -3.2909249767186928e-04
GC_6_188 b_6 NI_6 NS_188 0 -4.2221402681638773e-04
GC_6_189 b_6 NI_6 NS_189 0 -1.2814597589446401e-04
GC_6_190 b_6 NI_6 NS_190 0 6.5945552144793990e-05
GC_6_191 b_6 NI_6 NS_191 0 -4.0288419783190515e-04
GC_6_192 b_6 NI_6 NS_192 0 -1.9324532558699932e-04
GD_6_1 b_6 NI_6 NA_1 0 1.5615410863399782e-03
GD_6_2 b_6 NI_6 NA_2 0 1.2085697753098073e-03
GD_6_3 b_6 NI_6 NA_3 0 -1.8789078562656816e-03
GD_6_4 b_6 NI_6 NA_4 0 1.2826317495752003e-03
GD_6_5 b_6 NI_6 NA_5 0 -1.6409828077647678e-02
GD_6_6 b_6 NI_6 NA_6 0 -3.4733827510654125e-02
GD_6_7 b_6 NI_6 NA_7 0 -5.0537149341527126e-03
GD_6_8 b_6 NI_6 NA_8 0 4.6638403504647699e-03
GD_6_9 b_6 NI_6 NA_9 0 1.5551585240874033e-03
GD_6_10 b_6 NI_6 NA_10 0 1.2309698494739529e-03
GD_6_11 b_6 NI_6 NA_11 0 1.6413650805274075e-04
GD_6_12 b_6 NI_6 NA_12 0 -3.7880820614663807e-04
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 1.4525550304644406e-03
GC_7_2 b_7 NI_7 NS_2 0 8.9320795594831684e-07
GC_7_3 b_7 NI_7 NS_3 0 2.0243117087603147e-14
GC_7_4 b_7 NI_7 NS_4 0 -1.6542790222841445e-08
GC_7_5 b_7 NI_7 NS_5 0 -3.9776676681961983e-06
GC_7_6 b_7 NI_7 NS_6 0 1.0550364674805596e-06
GC_7_7 b_7 NI_7 NS_7 0 -1.9272782576668799e-05
GC_7_8 b_7 NI_7 NS_8 0 -8.7864866221149020e-05
GC_7_9 b_7 NI_7 NS_9 0 -5.4543314197839332e-05
GC_7_10 b_7 NI_7 NS_10 0 -1.0427792071338744e-04
GC_7_11 b_7 NI_7 NS_11 0 -3.2909116330830720e-04
GC_7_12 b_7 NI_7 NS_12 0 -4.2223511723840553e-04
GC_7_13 b_7 NI_7 NS_13 0 -1.2814499784206775e-04
GC_7_14 b_7 NI_7 NS_14 0 6.5948307840502722e-05
GC_7_15 b_7 NI_7 NS_15 0 -4.0287701967473791e-04
GC_7_16 b_7 NI_7 NS_16 0 -1.9322306167043792e-04
GC_7_17 b_7 NI_7 NS_17 0 -1.1956004235086652e-04
GC_7_18 b_7 NI_7 NS_18 0 1.2461892963662818e-07
GC_7_19 b_7 NI_7 NS_19 0 2.0838976310672610e-14
GC_7_20 b_7 NI_7 NS_20 0 5.2020223830953827e-09
GC_7_21 b_7 NI_7 NS_21 0 7.8261275759862014e-07
GC_7_22 b_7 NI_7 NS_22 0 -2.5019221126997335e-07
GC_7_23 b_7 NI_7 NS_23 0 6.1034005267519038e-05
GC_7_24 b_7 NI_7 NS_24 0 6.1343184943904604e-05
GC_7_25 b_7 NI_7 NS_25 0 1.6078981258284806e-04
GC_7_26 b_7 NI_7 NS_26 0 -4.4828663694905500e-06
GC_7_27 b_7 NI_7 NS_27 0 2.3834670197377952e-04
GC_7_28 b_7 NI_7 NS_28 0 -5.9906339537530112e-04
GC_7_29 b_7 NI_7 NS_29 0 -2.1647827747570025e-04
GC_7_30 b_7 NI_7 NS_30 0 -4.4467766056148156e-06
GC_7_31 b_7 NI_7 NS_31 0 -3.1110709216854214e-04
GC_7_32 b_7 NI_7 NS_32 0 -1.5136595156965059e-04
GC_7_33 b_7 NI_7 NS_33 0 -4.1496944625303792e-03
GC_7_34 b_7 NI_7 NS_34 0 1.7889797583251162e-06
GC_7_35 b_7 NI_7 NS_35 0 -1.6629751034918411e-13
GC_7_36 b_7 NI_7 NS_36 0 4.6962265347497353e-08
GC_7_37 b_7 NI_7 NS_37 0 1.3504682400302401e-05
GC_7_38 b_7 NI_7 NS_38 0 -3.8247383800027045e-06
GC_7_39 b_7 NI_7 NS_39 0 2.5160467772932266e-05
GC_7_40 b_7 NI_7 NS_40 0 2.4965169326812597e-05
GC_7_41 b_7 NI_7 NS_41 0 -3.8954655195375478e-04
GC_7_42 b_7 NI_7 NS_42 0 3.7419071448387050e-04
GC_7_43 b_7 NI_7 NS_43 0 1.1957380195202463e-03
GC_7_44 b_7 NI_7 NS_44 0 1.9793719813866253e-03
GC_7_45 b_7 NI_7 NS_45 0 1.9665944839622313e-04
GC_7_46 b_7 NI_7 NS_46 0 -2.0867241352673220e-04
GC_7_47 b_7 NI_7 NS_47 0 1.7536612684049332e-03
GC_7_48 b_7 NI_7 NS_48 0 1.3469524522395559e-03
GC_7_49 b_7 NI_7 NS_49 0 -5.1289256316103271e-04
GC_7_50 b_7 NI_7 NS_50 0 -1.3814662162981889e-06
GC_7_51 b_7 NI_7 NS_51 0 -1.6597419566774534e-13
GC_7_52 b_7 NI_7 NS_52 0 2.8168878838095287e-08
GC_7_53 b_7 NI_7 NS_53 0 7.0689847503229368e-06
GC_7_54 b_7 NI_7 NS_54 0 -1.4081085767231621e-06
GC_7_55 b_7 NI_7 NS_55 0 6.7488516464603299e-04
GC_7_56 b_7 NI_7 NS_56 0 5.6566698052270702e-04
GC_7_57 b_7 NI_7 NS_57 0 1.6542699723055918e-03
GC_7_58 b_7 NI_7 NS_58 0 -1.2912190911573091e-04
GC_7_59 b_7 NI_7 NS_59 0 2.1437558514718568e-03
GC_7_60 b_7 NI_7 NS_60 0 -6.5199286033341183e-03
GC_7_61 b_7 NI_7 NS_61 0 -2.2918351118807597e-03
GC_7_62 b_7 NI_7 NS_62 0 2.6343710990616843e-05
GC_7_63 b_7 NI_7 NS_63 0 -3.3998302500884048e-03
GC_7_64 b_7 NI_7 NS_64 0 -1.5771925455869446e-03
GC_7_65 b_7 NI_7 NS_65 0 1.0071458613534059e-02
GC_7_66 b_7 NI_7 NS_66 0 2.1089779751821401e-05
GC_7_67 b_7 NI_7 NS_67 0 2.4087388370931397e-13
GC_7_68 b_7 NI_7 NS_68 0 -3.5278884794838507e-07
GC_7_69 b_7 NI_7 NS_69 0 -2.4088408153548713e-05
GC_7_70 b_7 NI_7 NS_70 0 -3.1645135643416673e-06
GC_7_71 b_7 NI_7 NS_71 0 -1.8595038874960087e-03
GC_7_72 b_7 NI_7 NS_72 0 -1.1634090908633285e-02
GC_7_73 b_7 NI_7 NS_73 0 -2.7106537493746068e-02
GC_7_74 b_7 NI_7 NS_74 0 4.0963687875291786e-03
GC_7_75 b_7 NI_7 NS_75 0 1.3532835071946275e-02
GC_7_76 b_7 NI_7 NS_76 0 3.3625090879308386e-02
GC_7_77 b_7 NI_7 NS_77 0 -1.0133830551329999e-02
GC_7_78 b_7 NI_7 NS_78 0 -1.0505296930473939e-03
GC_7_79 b_7 NI_7 NS_79 0 2.5156766128630135e-02
GC_7_80 b_7 NI_7 NS_80 0 3.4474396303092035e-02
GC_7_81 b_7 NI_7 NS_81 0 -3.7910272282965017e-03
GC_7_82 b_7 NI_7 NS_82 0 3.2582514341532384e-06
GC_7_83 b_7 NI_7 NS_83 0 2.5082972008364319e-13
GC_7_84 b_7 NI_7 NS_84 0 -8.2120939761904146e-09
GC_7_85 b_7 NI_7 NS_85 0 -4.9980525067126489e-05
GC_7_86 b_7 NI_7 NS_86 0 1.1524559092498230e-05
GC_7_87 b_7 NI_7 NS_87 0 -2.9275878841658067e-03
GC_7_88 b_7 NI_7 NS_88 0 -2.2944246176950342e-03
GC_7_89 b_7 NI_7 NS_89 0 -7.0008839020514208e-03
GC_7_90 b_7 NI_7 NS_90 0 1.0673413321337631e-03
GC_7_91 b_7 NI_7 NS_91 0 -8.4047733682694817e-03
GC_7_92 b_7 NI_7 NS_92 0 3.0494305139086113e-02
GC_7_93 b_7 NI_7 NS_93 0 1.0663363839693700e-02
GC_7_94 b_7 NI_7 NS_94 0 -3.4370158891565503e-04
GC_7_95 b_7 NI_7 NS_95 0 1.6815910047908993e-02
GC_7_96 b_7 NI_7 NS_96 0 7.7402857264779468e-03
GC_7_97 b_7 NI_7 NS_97 0 5.8538696780432456e-02
GC_7_98 b_7 NI_7 NS_98 0 -2.0399782868520616e-05
GC_7_99 b_7 NI_7 NS_99 0 -1.1566557631734898e-12
GC_7_100 b_7 NI_7 NS_100 0 -2.4256618467947484e-06
GC_7_101 b_7 NI_7 NS_101 0 2.9536171348242052e-05
GC_7_102 b_7 NI_7 NS_102 0 -5.0077393182397205e-06
GC_7_103 b_7 NI_7 NS_103 0 -1.5267499712084834e-03
GC_7_104 b_7 NI_7 NS_104 0 7.1023439171835658e-03
GC_7_105 b_7 NI_7 NS_105 0 1.7512534622240509e-02
GC_7_106 b_7 NI_7 NS_106 0 -5.5133355808700737e-03
GC_7_107 b_7 NI_7 NS_107 0 -2.5510898639119005e-02
GC_7_108 b_7 NI_7 NS_108 0 -3.1264350183263907e-02
GC_7_109 b_7 NI_7 NS_109 0 7.3859331936045134e-03
GC_7_110 b_7 NI_7 NS_110 0 2.8756350237446960e-03
GC_7_111 b_7 NI_7 NS_111 0 -3.0902697276635454e-02
GC_7_112 b_7 NI_7 NS_112 0 -3.3632245136793928e-02
GC_7_113 b_7 NI_7 NS_113 0 1.9575321213387820e-01
GC_7_114 b_7 NI_7 NS_114 0 7.3981178954757123e-05
GC_7_115 b_7 NI_7 NS_115 0 3.8306312114534922e-12
GC_7_116 b_7 NI_7 NS_116 0 4.1281588496749995e-06
GC_7_117 b_7 NI_7 NS_117 0 1.1732266287771489e-04
GC_7_118 b_7 NI_7 NS_118 0 4.7768879959761769e-05
GC_7_119 b_7 NI_7 NS_119 0 -6.0787519151737177e-02
GC_7_120 b_7 NI_7 NS_120 0 -4.3818113064925342e-02
GC_7_121 b_7 NI_7 NS_121 0 4.0371750066582279e-02
GC_7_122 b_7 NI_7 NS_122 0 -1.8968584129851623e-02
GC_7_123 b_7 NI_7 NS_123 0 -1.2235642861607081e-01
GC_7_124 b_7 NI_7 NS_124 0 6.7044113150843077e-02
GC_7_125 b_7 NI_7 NS_125 0 -2.3662980586042614e-02
GC_7_126 b_7 NI_7 NS_126 0 1.2258474430122127e-02
GC_7_127 b_7 NI_7 NS_127 0 2.4212756898685340e-02
GC_7_128 b_7 NI_7 NS_128 0 -6.5629399757968582e-02
GC_7_129 b_7 NI_7 NS_129 0 5.5369735976815646e-03
GC_7_130 b_7 NI_7 NS_130 0 4.5137120600802977e-06
GC_7_131 b_7 NI_7 NS_131 0 1.3678567669485528e-13
GC_7_132 b_7 NI_7 NS_132 0 -1.9083496233259916e-07
GC_7_133 b_7 NI_7 NS_133 0 -1.2837238728502372e-05
GC_7_134 b_7 NI_7 NS_134 0 -5.8769714474655993e-07
GC_7_135 b_7 NI_7 NS_135 0 -7.6448539826566683e-04
GC_7_136 b_7 NI_7 NS_136 0 -4.6329222004263945e-03
GC_7_137 b_7 NI_7 NS_137 0 -1.0664494380214067e-02
GC_7_138 b_7 NI_7 NS_138 0 1.5135503785583815e-03
GC_7_139 b_7 NI_7 NS_139 0 4.9166001687895190e-03
GC_7_140 b_7 NI_7 NS_140 0 1.2751659952078864e-02
GC_7_141 b_7 NI_7 NS_141 0 -4.0713865945526959e-03
GC_7_142 b_7 NI_7 NS_142 0 -3.1357012522918525e-04
GC_7_143 b_7 NI_7 NS_143 0 9.4730023039845609e-03
GC_7_144 b_7 NI_7 NS_144 0 1.3280516256656249e-02
GC_7_145 b_7 NI_7 NS_145 0 -1.7164818059571276e-03
GC_7_146 b_7 NI_7 NS_146 0 1.5984841058252338e-06
GC_7_147 b_7 NI_7 NS_147 0 1.3989482050353263e-13
GC_7_148 b_7 NI_7 NS_148 0 3.6496230043400008e-08
GC_7_149 b_7 NI_7 NS_149 0 -1.9059938687261552e-05
GC_7_150 b_7 NI_7 NS_150 0 4.6715613853917005e-06
GC_7_151 b_7 NI_7 NS_151 0 -1.0759447243572124e-03
GC_7_152 b_7 NI_7 NS_152 0 -7.5181020463978656e-04
GC_7_153 b_7 NI_7 NS_153 0 -2.6152412235010817e-03
GC_7_154 b_7 NI_7 NS_154 0 3.9480799273044153e-04
GC_7_155 b_7 NI_7 NS_155 0 -2.9093021630866639e-03
GC_7_156 b_7 NI_7 NS_156 0 1.1450280482787607e-02
GC_7_157 b_7 NI_7 NS_157 0 4.0045967404318998e-03
GC_7_158 b_7 NI_7 NS_158 0 -1.5872579283479144e-04
GC_7_159 b_7 NI_7 NS_159 0 6.2634041496411521e-03
GC_7_160 b_7 NI_7 NS_160 0 2.7898901284060321e-03
GC_7_161 b_7 NI_7 NS_161 0 -4.0765159827529989e-03
GC_7_162 b_7 NI_7 NS_162 0 -3.5138295180783669e-06
GC_7_163 b_7 NI_7 NS_163 0 -1.6897008450471441e-13
GC_7_164 b_7 NI_7 NS_164 0 4.8311842590533813e-08
GC_7_165 b_7 NI_7 NS_165 0 1.4111559008709911e-05
GC_7_166 b_7 NI_7 NS_166 0 -3.9678298878925915e-06
GC_7_167 b_7 NI_7 NS_167 0 2.4220413372981267e-05
GC_7_168 b_7 NI_7 NS_168 0 2.1750335377029242e-05
GC_7_169 b_7 NI_7 NS_169 0 -3.9069537038919884e-04
GC_7_170 b_7 NI_7 NS_170 0 3.7011700220639999e-04
GC_7_171 b_7 NI_7 NS_171 0 1.1892348770402266e-03
GC_7_172 b_7 NI_7 NS_172 0 1.9568551340291783e-03
GC_7_173 b_7 NI_7 NS_173 0 1.9074277462601544e-04
GC_7_174 b_7 NI_7 NS_174 0 -2.0993602354837660e-04
GC_7_175 b_7 NI_7 NS_175 0 1.7254780417946692e-03
GC_7_176 b_7 NI_7 NS_176 0 1.3072723030466682e-03
GC_7_177 b_7 NI_7 NS_177 0 -5.4059345253431852e-04
GC_7_178 b_7 NI_7 NS_178 0 3.1245540002233907e-06
GC_7_179 b_7 NI_7 NS_179 0 -1.6759121911652797e-13
GC_7_180 b_7 NI_7 NS_180 0 2.8401367050436681e-08
GC_7_181 b_7 NI_7 NS_181 0 6.6560576805152073e-06
GC_7_182 b_7 NI_7 NS_182 0 -1.3310751127914655e-06
GC_7_183 b_7 NI_7 NS_183 0 6.7449136055829995e-04
GC_7_184 b_7 NI_7 NS_184 0 5.6657305491242054e-04
GC_7_185 b_7 NI_7 NS_185 0 1.6536587738663431e-03
GC_7_186 b_7 NI_7 NS_186 0 -1.2727187835772603e-04
GC_7_187 b_7 NI_7 NS_187 0 2.1414850898987181e-03
GC_7_188 b_7 NI_7 NS_188 0 -6.5096130758924052e-03
GC_7_189 b_7 NI_7 NS_189 0 -2.2900887365418254e-03
GC_7_190 b_7 NI_7 NS_190 0 2.9685183786094275e-05
GC_7_191 b_7 NI_7 NS_191 0 -3.3826865265310594e-03
GC_7_192 b_7 NI_7 NS_192 0 -1.5439520871963330e-03
GD_7_1 b_7 NI_7 NA_1 0 -3.7872044310361633e-04
GD_7_2 b_7 NI_7 NA_2 0 1.6446240016533044e-04
GD_7_3 b_7 NI_7 NA_3 0 1.2297369783168029e-03
GD_7_4 b_7 NI_7 NA_4 0 1.5551245006189586e-03
GD_7_5 b_7 NI_7 NA_5 0 4.6641607519285581e-03
GD_7_6 b_7 NI_7 NA_6 0 -5.0537712260213278e-03
GD_7_7 b_7 NI_7 NA_7 0 -3.4735394940648742e-02
GD_7_8 b_7 NI_7 NA_8 0 -1.6409419395124563e-02
GD_7_9 b_7 NI_7 NA_9 0 1.2834812694113341e-03
GD_7_10 b_7 NI_7 NA_10 0 -1.8801625901142857e-03
GD_7_11 b_7 NI_7 NA_11 0 1.2095900535538616e-03
GD_7_12 b_7 NI_7 NA_12 0 1.5612930327666070e-03
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 -1.1818043212203119e-04
GC_8_2 b_8 NI_8 NS_2 0 1.2960814643120497e-07
GC_8_3 b_8 NI_8 NS_3 0 2.0837930888212294e-14
GC_8_4 b_8 NI_8 NS_4 0 5.1985450928847352e-09
GC_8_5 b_8 NI_8 NS_5 0 7.8211516840947877e-07
GC_8_6 b_8 NI_8 NS_6 0 -2.5001735943922154e-07
GC_8_7 b_8 NI_8 NS_7 0 6.0931819262253080e-05
GC_8_8 b_8 NI_8 NS_8 0 6.1238778646171993e-05
GC_8_9 b_8 NI_8 NS_9 0 1.6069019582800963e-04
GC_8_10 b_8 NI_8 NS_10 0 -4.6114147191267874e-06
GC_8_11 b_8 NI_8 NS_11 0 2.3772034875282503e-04
GC_8_12 b_8 NI_8 NS_12 0 -5.9903153618839802e-04
GC_8_13 b_8 NI_8 NS_13 0 -2.1643358128548156e-04
GC_8_14 b_8 NI_8 NS_14 0 -4.3083973348967309e-06
GC_8_15 b_8 NI_8 NS_15 0 -3.1112785471685753e-04
GC_8_16 b_8 NI_8 NS_16 0 -1.5125006197992983e-04
GC_8_17 b_8 NI_8 NS_17 0 1.4526966463267370e-03
GC_8_18 b_8 NI_8 NS_18 0 8.8678960040264558e-07
GC_8_19 b_8 NI_8 NS_19 0 2.0246299489917372e-14
GC_8_20 b_8 NI_8 NS_20 0 -1.6541606054093953e-08
GC_8_21 b_8 NI_8 NS_21 0 -3.9770943145461541e-06
GC_8_22 b_8 NI_8 NS_22 0 1.0549140573831258e-06
GC_8_23 b_8 NI_8 NS_23 0 -1.9277044930996798e-05
GC_8_24 b_8 NI_8 NS_24 0 -8.7872301236694783e-05
GC_8_25 b_8 NI_8 NS_25 0 -5.4548240939756875e-05
GC_8_26 b_8 NI_8 NS_26 0 -1.0428003027022217e-04
GC_8_27 b_8 NI_8 NS_27 0 -3.2909982788775874e-04
GC_8_28 b_8 NI_8 NS_28 0 -4.2227744245706896e-04
GC_8_29 b_8 NI_8 NS_29 0 -1.2815926186437112e-04
GC_8_30 b_8 NI_8 NS_30 0 6.5948721608380972e-05
GC_8_31 b_8 NI_8 NS_31 0 -4.0292459546696239e-04
GC_8_32 b_8 NI_8 NS_32 0 -1.9327761837643407e-04
GC_8_33 b_8 NI_8 NS_33 0 -5.1270224514996356e-04
GC_8_34 b_8 NI_8 NS_34 0 -1.3433188797750988e-06
GC_8_35 b_8 NI_8 NS_35 0 -1.6596546955004489e-13
GC_8_36 b_8 NI_8 NS_36 0 2.8139945027161549e-08
GC_8_37 b_8 NI_8 NS_37 0 7.0628769044140770e-06
GC_8_38 b_8 NI_8 NS_38 0 -1.4064003410147747e-06
GC_8_39 b_8 NI_8 NS_39 0 6.7486708343457175e-04
GC_8_40 b_8 NI_8 NS_40 0 5.6565662026762849e-04
GC_8_41 b_8 NI_8 NS_41 0 1.6542448440713836e-03
GC_8_42 b_8 NI_8 NS_42 0 -1.2913297045469928e-04
GC_8_43 b_8 NI_8 NS_43 0 2.1436117355035705e-03
GC_8_44 b_8 NI_8 NS_44 0 -6.5198862447081209e-03
GC_8_45 b_8 NI_8 NS_45 0 -2.2918190471801808e-03
GC_8_46 b_8 NI_8 NS_46 0 2.6391626927568119e-05
GC_8_47 b_8 NI_8 NS_47 0 -3.3997609985337972e-03
GC_8_48 b_8 NI_8 NS_48 0 -1.5769646316875008e-03
GC_8_49 b_8 NI_8 NS_49 0 -4.1538626304280174e-03
GC_8_50 b_8 NI_8 NS_50 0 1.7863836479552726e-06
GC_8_51 b_8 NI_8 NS_51 0 -1.6631811770939300e-13
GC_8_52 b_8 NI_8 NS_52 0 4.6974226815161665e-08
GC_8_53 b_8 NI_8 NS_53 0 1.3507243237525997e-05
GC_8_54 b_8 NI_8 NS_54 0 -3.8257808993782732e-06
GC_8_55 b_8 NI_8 NS_55 0 2.5148873614381760e-05
GC_8_56 b_8 NI_8 NS_56 0 2.5213091397404070e-05
GC_8_57 b_8 NI_8 NS_57 0 -3.8914601115010259e-04
GC_8_58 b_8 NI_8 NS_58 0 3.7463204214209668e-04
GC_8_59 b_8 NI_8 NS_59 0 1.1967381782213159e-03
GC_8_60 b_8 NI_8 NS_60 0 1.9797670558469342e-03
GC_8_61 b_8 NI_8 NS_61 0 1.9690211036927925e-04
GC_8_62 b_8 NI_8 NS_62 0 -2.0870694219841552e-04
GC_8_63 b_8 NI_8 NS_63 0 1.7545167769352805e-03
GC_8_64 b_8 NI_8 NS_64 0 1.3471972816375909e-03
GC_8_65 b_8 NI_8 NS_65 0 -3.7911324504302985e-03
GC_8_66 b_8 NI_8 NS_66 0 3.3099086685226320e-06
GC_8_67 b_8 NI_8 NS_67 0 2.5083682703274456e-13
GC_8_68 b_8 NI_8 NS_68 0 -8.2091197946472607e-09
GC_8_69 b_8 NI_8 NS_69 0 -4.9984117964933023e-05
GC_8_70 b_8 NI_8 NS_70 0 1.1525146900595748e-05
GC_8_71 b_8 NI_8 NS_71 0 -2.9276254881893558e-03
GC_8_72 b_8 NI_8 NS_72 0 -2.2944519720334566e-03
GC_8_73 b_8 NI_8 NS_73 0 -7.0009407450788248e-03
GC_8_74 b_8 NI_8 NS_74 0 1.0673150190266135e-03
GC_8_75 b_8 NI_8 NS_75 0 -8.4050653484825585e-03
GC_8_76 b_8 NI_8 NS_76 0 3.0494618221964649e-02
GC_8_77 b_8 NI_8 NS_77 0 1.0663478557402264e-02
GC_8_78 b_8 NI_8 NS_78 0 -3.4360520732214375e-04
GC_8_79 b_8 NI_8 NS_79 0 1.6816254216786741e-02
GC_8_80 b_8 NI_8 NS_80 0 7.7407887401041726e-03
GC_8_81 b_8 NI_8 NS_81 0 1.0072824230317102e-02
GC_8_82 b_8 NI_8 NS_82 0 2.0968717314406485e-05
GC_8_83 b_8 NI_8 NS_83 0 2.4086070545144305e-13
GC_8_84 b_8 NI_8 NS_84 0 -3.5273573896819875e-07
GC_8_85 b_8 NI_8 NS_85 0 -2.4073613695951795e-05
GC_8_86 b_8 NI_8 NS_86 0 -3.1683110804644012e-06
GC_8_87 b_8 NI_8 NS_87 0 -1.8595031913329341e-03
GC_8_88 b_8 NI_8 NS_88 0 -1.1634140492335016e-02
GC_8_89 b_8 NI_8 NS_89 0 -2.7106518916204990e-02
GC_8_90 b_8 NI_8 NS_90 0 4.0962888516327019e-03
GC_8_91 b_8 NI_8 NS_91 0 1.3532793116182152e-02
GC_8_92 b_8 NI_8 NS_92 0 3.3624513487218004e-02
GC_8_93 b_8 NI_8 NS_93 0 -1.0133991199008806e-02
GC_8_94 b_8 NI_8 NS_94 0 -1.0505718373664101e-03
GC_8_95 b_8 NI_8 NS_95 0 2.5156121748030343e-02
GC_8_96 b_8 NI_8 NS_96 0 3.4473487201456723e-02
GC_8_97 b_8 NI_8 NS_97 0 1.9575430004552299e-01
GC_8_98 b_8 NI_8 NS_98 0 7.4182051879380758e-05
GC_8_99 b_8 NI_8 NS_99 0 3.8304395990106077e-12
GC_8_100 b_8 NI_8 NS_100 0 4.1280321874192179e-06
GC_8_101 b_8 NI_8 NS_101 0 1.1729086518814670e-04
GC_8_102 b_8 NI_8 NS_102 0 4.7777564635107211e-05
GC_8_103 b_8 NI_8 NS_103 0 -6.0787602773528820e-02
GC_8_104 b_8 NI_8 NS_104 0 -4.3818189996638501e-02
GC_8_105 b_8 NI_8 NS_105 0 4.0371608705668131e-02
GC_8_106 b_8 NI_8 NS_106 0 -1.8968655432443460e-02
GC_8_107 b_8 NI_8 NS_107 0 -1.2235717387680711e-01
GC_8_108 b_8 NI_8 NS_108 0 6.7044234116371740e-02
GC_8_109 b_8 NI_8 NS_109 0 -2.3662941617966678e-02
GC_8_110 b_8 NI_8 NS_110 0 1.2258725958369753e-02
GC_8_111 b_8 NI_8 NS_111 0 2.4213041326742062e-02
GC_8_112 b_8 NI_8 NS_112 0 -6.5628237957012586e-02
GC_8_113 b_8 NI_8 NS_113 0 5.8534059871912777e-02
GC_8_114 b_8 NI_8 NS_114 0 -2.0146024384932370e-05
GC_8_115 b_8 NI_8 NS_115 0 -1.1566350921487712e-12
GC_8_116 b_8 NI_8 NS_116 0 -2.4257573680195847e-06
GC_8_117 b_8 NI_8 NS_117 0 2.9508661821527766e-05
GC_8_118 b_8 NI_8 NS_118 0 -5.0009182195944519e-06
GC_8_119 b_8 NI_8 NS_119 0 -1.5267076491579368e-03
GC_8_120 b_8 NI_8 NS_120 0 7.1025512519599888e-03
GC_8_121 b_8 NI_8 NS_121 0 1.7512585109870728e-02
GC_8_122 b_8 NI_8 NS_122 0 -5.5130492856973372e-03
GC_8_123 b_8 NI_8 NS_123 0 -2.5510341289859823e-02
GC_8_124 b_8 NI_8 NS_124 0 -3.1262778315834967e-02
GC_8_125 b_8 NI_8 NS_125 0 7.3863628416985117e-03
GC_8_126 b_8 NI_8 NS_126 0 2.8756295636967071e-03
GC_8_127 b_8 NI_8 NS_127 0 -3.0900966373280780e-02
GC_8_128 b_8 NI_8 NS_128 0 -3.3630175725056000e-02
GC_8_129 b_8 NI_8 NS_129 0 -1.7186591299489687e-03
GC_8_130 b_8 NI_8 NS_130 0 1.5761284829600282e-06
GC_8_131 b_8 NI_8 NS_131 0 1.3990438323117892e-13
GC_8_132 b_8 NI_8 NS_132 0 3.6542220375740614e-08
GC_8_133 b_8 NI_8 NS_133 0 -1.9053724657341371e-05
GC_8_134 b_8 NI_8 NS_134 0 4.6694878883848410e-06
GC_8_135 b_8 NI_8 NS_135 0 -1.0758251926550784e-03
GC_8_136 b_8 NI_8 NS_136 0 -7.5166726942623699e-04
GC_8_137 b_8 NI_8 NS_137 0 -2.6151130095226436e-03
GC_8_138 b_8 NI_8 NS_138 0 3.9499533836876951e-04
GC_8_139 b_8 NI_8 NS_139 0 -2.9084346479425847e-03
GC_8_140 b_8 NI_8 NS_140 0 1.1450430965305148e-02
GC_8_141 b_8 NI_8 NS_141 0 4.0045961644253891e-03
GC_8_142 b_8 NI_8 NS_142 0 -1.5892156744752359e-04
GC_8_143 b_8 NI_8 NS_143 0 6.2635844611555556e-03
GC_8_144 b_8 NI_8 NS_144 0 2.7897718929863306e-03
GC_8_145 b_8 NI_8 NS_145 0 5.5381479522115425e-03
GC_8_146 b_8 NI_8 NS_146 0 4.3906472253344768e-06
GC_8_147 b_8 NI_8 NS_147 0 1.3679101754990040e-13
GC_8_148 b_8 NI_8 NS_148 0 -1.9077038742651429e-07
GC_8_149 b_8 NI_8 NS_149 0 -1.2821326772958605e-05
GC_8_150 b_8 NI_8 NS_150 0 -5.9190358620126031e-07
GC_8_151 b_8 NI_8 NS_151 0 -7.6447612391830383e-04
GC_8_152 b_8 NI_8 NS_152 0 -4.6329567195340753e-03
GC_8_153 b_8 NI_8 NS_153 0 -1.0664457823350347e-02
GC_8_154 b_8 NI_8 NS_154 0 1.5134791067726459e-03
GC_8_155 b_8 NI_8 NS_155 0 4.9166059217149935e-03
GC_8_156 b_8 NI_8 NS_156 0 1.2751100042545779e-02
GC_8_157 b_8 NI_8 NS_157 0 -4.0715418511358499e-03
GC_8_158 b_8 NI_8 NS_158 0 -3.1361944372414961e-04
GC_8_159 b_8 NI_8 NS_159 0 9.4723921574752044e-03
GC_8_160 b_8 NI_8 NS_160 0 1.3279617879870448e-02
GC_8_161 b_8 NI_8 NS_161 0 -5.4123096911943137e-04
GC_8_162 b_8 NI_8 NS_162 0 3.1761667123083244e-06
GC_8_163 b_8 NI_8 NS_163 0 -1.6758164942892160e-13
GC_8_164 b_8 NI_8 NS_164 0 2.8381789799728809e-08
GC_8_165 b_8 NI_8 NS_165 0 6.6500621279930602e-06
GC_8_166 b_8 NI_8 NS_166 0 -1.3295866957996542e-06
GC_8_167 b_8 NI_8 NS_167 0 6.7449017895573004e-04
GC_8_168 b_8 NI_8 NS_168 0 5.6660901861900568e-04
GC_8_169 b_8 NI_8 NS_169 0 1.6536550571717849e-03
GC_8_170 b_8 NI_8 NS_170 0 -1.2722879938291268e-04
GC_8_171 b_8 NI_8 NS_171 0 2.1415322470503578e-03
GC_8_172 b_8 NI_8 NS_172 0 -6.5093451478056936e-03
GC_8_173 b_8 NI_8 NS_173 0 -2.2900161124990433e-03
GC_8_174 b_8 NI_8 NS_174 0 2.9697963141291443e-05
GC_8_175 b_8 NI_8 NS_175 0 -3.3823932605495976e-03
GC_8_176 b_8 NI_8 NS_176 0 -1.5435562035715029e-03
GC_8_177 b_8 NI_8 NS_177 0 -4.0733154397862110e-03
GC_8_178 b_8 NI_8 NS_178 0 -3.4913050327228537e-06
GC_8_179 b_8 NI_8 NS_179 0 -1.6897956913188288e-13
GC_8_180 b_8 NI_8 NS_180 0 4.8300790577477420e-08
GC_8_181 b_8 NI_8 NS_181 0 1.4108330694597187e-05
GC_8_182 b_8 NI_8 NS_182 0 -3.9667327864229318e-06
GC_8_183 b_8 NI_8 NS_183 0 2.4234187978849323e-05
GC_8_184 b_8 NI_8 NS_184 0 2.1551035726504546e-05
GC_8_185 b_8 NI_8 NS_185 0 -3.9108293831849875e-04
GC_8_186 b_8 NI_8 NS_186 0 3.6975918303477489e-04
GC_8_187 b_8 NI_8 NS_187 0 1.1884464777538713e-03
GC_8_188 b_8 NI_8 NS_188 0 1.9567884878511329e-03
GC_8_189 b_8 NI_8 NS_189 0 1.9058562238076569e-04
GC_8_190 b_8 NI_8 NS_190 0 -2.0993638439585917e-04
GC_8_191 b_8 NI_8 NS_191 0 1.7249371133049635e-03
GC_8_192 b_8 NI_8 NS_192 0 1.3072757404810149e-03
GD_8_1 b_8 NI_8 NA_1 0 1.6403382721092474e-04
GD_8_2 b_8 NI_8 NA_2 0 -3.7877021787587414e-04
GD_8_3 b_8 NI_8 NA_3 0 1.5550127932137275e-03
GD_8_4 b_8 NI_8 NA_4 0 1.2309618840217723e-03
GD_8_5 b_8 NI_8 NA_5 0 -5.0537701899001789e-03
GD_8_6 b_8 NI_8 NA_6 0 4.6638387670759592e-03
GD_8_7 b_8 NI_8 NA_7 0 -1.6409959146417120e-02
GD_8_8 b_8 NI_8 NA_8 0 -3.4734169699674029e-02
GD_8_9 b_8 NI_8 NA_9 0 -1.8794748989783539e-03
GD_8_10 b_8 NI_8 NA_10 0 1.2832202137095807e-03
GD_8_11 b_8 NI_8 NA_11 0 1.5614191375289690e-03
GD_8_12 b_8 NI_8 NA_12 0 1.2085963414491495e-03
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 7.9729132707908338e-05
GC_9_2 b_9 NI_9 NS_2 0 5.1636672043567738e-08
GC_9_3 b_9 NI_9 NS_3 0 3.3837852918713668e-15
GC_9_4 b_9 NI_9 NS_4 0 -9.6172977313997591e-10
GC_9_5 b_9 NI_9 NS_5 0 -2.2497095335863727e-07
GC_9_6 b_9 NI_9 NS_6 0 6.5563669191066010e-08
GC_9_7 b_9 NI_9 NS_7 0 -1.4041362968472972e-06
GC_9_8 b_9 NI_9 NS_8 0 -5.7433681830341865e-06
GC_9_9 b_9 NI_9 NS_9 0 -4.3977598948638347e-06
GC_9_10 b_9 NI_9 NS_10 0 -4.7443079509572674e-06
GC_9_11 b_9 NI_9 NS_11 0 -1.6603336889262479e-05
GC_9_12 b_9 NI_9 NS_12 0 -2.2920992117448651e-05
GC_9_13 b_9 NI_9 NS_13 0 -8.1452252378693382e-06
GC_9_14 b_9 NI_9 NS_14 0 4.0115373657215039e-06
GC_9_15 b_9 NI_9 NS_15 0 -2.0849955817307341e-05
GC_9_16 b_9 NI_9 NS_16 0 -8.4234399955201994e-06
GC_9_17 b_9 NI_9 NS_17 0 2.2130007559608558e-05
GC_9_18 b_9 NI_9 NS_18 0 4.4307063437605187e-09
GC_9_19 b_9 NI_9 NS_19 0 3.4027026843600403e-15
GC_9_20 b_9 NI_9 NS_20 0 -3.8847966425358328e-10
GC_9_21 b_9 NI_9 NS_21 0 -4.9110031264124792e-08
GC_9_22 b_9 NI_9 NS_22 0 1.7205438762414635e-08
GC_9_23 b_9 NI_9 NS_23 0 -2.6246932385873067e-06
GC_9_24 b_9 NI_9 NS_24 0 3.2070908120339062e-06
GC_9_25 b_9 NI_9 NS_25 0 3.1790053565598192e-06
GC_9_26 b_9 NI_9 NS_26 0 -1.9242413607100858e-06
GC_9_27 b_9 NI_9 NS_27 0 1.2276278141746326e-06
GC_9_28 b_9 NI_9 NS_28 0 -9.8471842198924135e-06
GC_9_29 b_9 NI_9 NS_29 0 -4.6415167670853241e-06
GC_9_30 b_9 NI_9 NS_30 0 7.9253667799682214e-07
GC_9_31 b_9 NI_9 NS_31 0 -8.4603968214495455e-06
GC_9_32 b_9 NI_9 NS_32 0 -5.5195221494228634e-06
GC_9_33 b_9 NI_9 NS_33 0 5.7603505161798313e-04
GC_9_34 b_9 NI_9 NS_34 0 -1.4756363727965888e-07
GC_9_35 b_9 NI_9 NS_35 0 9.3191389389217790e-15
GC_9_36 b_9 NI_9 NS_36 0 -6.6837578000553088e-09
GC_9_37 b_9 NI_9 NS_37 0 -1.5525788265280804e-06
GC_9_38 b_9 NI_9 NS_38 0 4.2142631765015138e-07
GC_9_39 b_9 NI_9 NS_39 0 -7.8446283624960195e-06
GC_9_40 b_9 NI_9 NS_40 0 -3.5374955071437467e-05
GC_9_41 b_9 NI_9 NS_41 0 -2.2999860568797556e-05
GC_9_42 b_9 NI_9 NS_42 0 -4.0669305936103050e-05
GC_9_43 b_9 NI_9 NS_43 0 -1.2953846505628450e-04
GC_9_44 b_9 NI_9 NS_44 0 -1.6493997450079794e-04
GC_9_45 b_9 NI_9 NS_45 0 -5.0629463687716417e-05
GC_9_46 b_9 NI_9 NS_46 0 2.6197222608035887e-05
GC_9_47 b_9 NI_9 NS_47 0 -1.5795641519509624e-04
GC_9_48 b_9 NI_9 NS_48 0 -7.7187448906239903e-05
GC_9_49 b_9 NI_9 NS_49 0 2.1055651961545268e-05
GC_9_50 b_9 NI_9 NS_50 0 -2.1990012416083612e-08
GC_9_51 b_9 NI_9 NS_51 0 9.1433408777434356e-15
GC_9_52 b_9 NI_9 NS_52 0 2.4622781285223573e-09
GC_9_53 b_9 NI_9 NS_53 0 3.6440447048755706e-07
GC_9_54 b_9 NI_9 NS_54 0 -1.2259458310014687e-07
GC_9_55 b_9 NI_9 NS_55 0 1.8634961362702463e-05
GC_9_56 b_9 NI_9 NS_56 0 2.3649417973142744e-05
GC_9_57 b_9 NI_9 NS_57 0 6.0261932730260830e-05
GC_9_58 b_9 NI_9 NS_58 0 -7.0206161819254694e-06
GC_9_59 b_9 NI_9 NS_59 0 7.3285864378129783e-05
GC_9_60 b_9 NI_9 NS_60 0 -2.3641765760594802e-04
GC_9_61 b_9 NI_9 NS_61 0 -8.4900661281850720e-05
GC_9_62 b_9 NI_9 NS_62 0 2.4597121758836029e-06
GC_9_63 b_9 NI_9 NS_63 0 -1.2825025916511585e-04
GC_9_64 b_9 NI_9 NS_64 0 -6.0501398447498949e-05
GC_9_65 b_9 NI_9 NS_65 0 -4.1491667735925322e-03
GC_9_66 b_9 NI_9 NS_66 0 1.7202681294618845e-06
GC_9_67 b_9 NI_9 NS_67 0 -1.6584146661305731e-13
GC_9_68 b_9 NI_9 NS_68 0 4.6782603407993323e-08
GC_9_69 b_9 NI_9 NS_69 0 1.3497745599171589e-05
GC_9_70 b_9 NI_9 NS_70 0 -3.8204583480288324e-06
GC_9_71 b_9 NI_9 NS_71 0 2.5277391043072440e-05
GC_9_72 b_9 NI_9 NS_72 0 2.4939849430714670e-05
GC_9_73 b_9 NI_9 NS_73 0 -3.8904116638520235e-04
GC_9_74 b_9 NI_9 NS_74 0 3.7415462490745735e-04
GC_9_75 b_9 NI_9 NS_75 0 1.1958978967532032e-03
GC_9_76 b_9 NI_9 NS_76 0 1.9770916077404971e-03
GC_9_77 b_9 NI_9 NS_77 0 1.9609496300642686e-04
GC_9_78 b_9 NI_9 NS_78 0 -2.0846911797504813e-04
GC_9_79 b_9 NI_9 NS_79 0 1.7524532349889300e-03
GC_9_80 b_9 NI_9 NS_80 0 1.3458545823809990e-03
GC_9_81 b_9 NI_9 NS_81 0 -5.1140365856038310e-04
GC_9_82 b_9 NI_9 NS_82 0 -1.3710984653101326e-06
GC_9_83 b_9 NI_9 NS_83 0 -1.6671366967752733e-13
GC_9_84 b_9 NI_9 NS_84 0 2.7430453208852173e-08
GC_9_85 b_9 NI_9 NS_85 0 7.0005230574573777e-06
GC_9_86 b_9 NI_9 NS_86 0 -1.3816970114662862e-06
GC_9_87 b_9 NI_9 NS_87 0 6.7528414486517081e-04
GC_9_88 b_9 NI_9 NS_88 0 5.6580598145526153e-04
GC_9_89 b_9 NI_9 NS_89 0 1.6548984129641990e-03
GC_9_90 b_9 NI_9 NS_90 0 -1.2962499530809156e-04
GC_9_91 b_9 NI_9 NS_91 0 2.1437203864783567e-03
GC_9_92 b_9 NI_9 NS_92 0 -6.5224917061969361e-03
GC_9_93 b_9 NI_9 NS_93 0 -2.2924468615532247e-03
GC_9_94 b_9 NI_9 NS_94 0 2.6297145848818051e-05
GC_9_95 b_9 NI_9 NS_95 0 -3.4018494608953767e-03
GC_9_96 b_9 NI_9 NS_96 0 -1.5789160492377990e-03
GC_9_97 b_9 NI_9 NS_97 0 5.5045567813056962e-03
GC_9_98 b_9 NI_9 NS_98 0 7.6977561774955634e-06
GC_9_99 b_9 NI_9 NS_99 0 1.3807973118511282e-13
GC_9_100 b_9 NI_9 NS_100 0 -1.9139372408702200e-07
GC_9_101 b_9 NI_9 NS_101 0 -1.3178669960466075e-05
GC_9_102 b_9 NI_9 NS_102 0 -5.0935260922807535e-07
GC_9_103 b_9 NI_9 NS_103 0 -7.6452587903454324e-04
GC_9_104 b_9 NI_9 NS_104 0 -4.6323042837315125e-03
GC_9_105 b_9 NI_9 NS_105 0 -1.0665599758027430e-02
GC_9_106 b_9 NI_9 NS_106 0 1.5152634121783010e-03
GC_9_107 b_9 NI_9 NS_107 0 4.9162533738198863e-03
GC_9_108 b_9 NI_9 NS_108 0 1.2766098599891074e-02
GC_9_109 b_9 NI_9 NS_109 0 -4.0675089609761338e-03
GC_9_110 b_9 NI_9 NS_110 0 -3.1201201100893125e-04
GC_9_111 b_9 NI_9 NS_111 0 9.4895489437278723e-03
GC_9_112 b_9 NI_9 NS_112 0 1.3304972279059277e-02
GC_9_113 b_9 NI_9 NS_113 0 -1.7387472536427593e-03
GC_9_114 b_9 NI_9 NS_114 0 3.3844914856621857e-06
GC_9_115 b_9 NI_9 NS_115 0 1.4241557227615289e-13
GC_9_116 b_9 NI_9 NS_116 0 3.7276047993039472e-08
GC_9_117 b_9 NI_9 NS_117 0 -1.9144152108445355e-05
GC_9_118 b_9 NI_9 NS_118 0 4.6728287629064467e-06
GC_9_119 b_9 NI_9 NS_119 0 -1.0768323520573377e-03
GC_9_120 b_9 NI_9 NS_120 0 -7.5114209148142812e-04
GC_9_121 b_9 NI_9 NS_121 0 -2.6165243318033351e-03
GC_9_122 b_9 NI_9 NS_122 0 3.9711204900221659e-04
GC_9_123 b_9 NI_9 NS_123 0 -2.9082785714389710e-03
GC_9_124 b_9 NI_9 NS_124 0 1.1463127336805478e-02
GC_9_125 b_9 NI_9 NS_125 0 4.0078499766629198e-03
GC_9_126 b_9 NI_9 NS_126 0 -1.5796865237660080e-04
GC_9_127 b_9 NI_9 NS_127 0 6.2765284990584699e-03
GC_9_128 b_9 NI_9 NS_128 0 2.8066287709139766e-03
GC_9_129 b_9 NI_9 NS_129 0 5.8324393288564681e-02
GC_9_130 b_9 NI_9 NS_130 0 -7.5750912873790252e-06
GC_9_131 b_9 NI_9 NS_131 0 -1.1650579143916058e-12
GC_9_132 b_9 NI_9 NS_132 0 -2.4303778669764744e-06
GC_9_133 b_9 NI_9 NS_133 0 2.8219664172341523e-05
GC_9_134 b_9 NI_9 NS_134 0 -4.6803798276501536e-06
GC_9_135 b_9 NI_9 NS_135 0 -1.5286252505367752e-03
GC_9_136 b_9 NI_9 NS_136 0 7.1113443934310199e-03
GC_9_137 b_9 NI_9 NS_137 0 1.7510122821835519e-02
GC_9_138 b_9 NI_9 NS_138 0 -5.4962426125809288e-03
GC_9_139 b_9 NI_9 NS_139 0 -2.5486524590942427e-02
GC_9_140 b_9 NI_9 NS_140 0 -3.1173567313001471e-02
GC_9_141 b_9 NI_9 NS_141 0 7.4101108952942260e-03
GC_9_142 b_9 NI_9 NS_142 0 2.8759912083722522e-03
GC_9_143 b_9 NI_9 NS_143 0 -3.0809941490717783e-02
GC_9_144 b_9 NI_9 NS_144 0 -3.3522851500927875e-02
GC_9_145 b_9 NI_9 NS_145 0 1.9562354555801867e-01
GC_9_146 b_9 NI_9 NS_146 0 6.0207255326817782e-05
GC_9_147 b_9 NI_9 NS_147 0 3.3891413275533787e-12
GC_9_148 b_9 NI_9 NS_148 0 4.1874328525749313e-06
GC_9_149 b_9 NI_9 NS_149 0 1.2048998865789507e-04
GC_9_150 b_9 NI_9 NS_150 0 4.6656840671793248e-05
GC_9_151 b_9 NI_9 NS_151 0 -6.0782605418120465e-02
GC_9_152 b_9 NI_9 NS_152 0 -4.3809427881697588e-02
GC_9_153 b_9 NI_9 NS_153 0 4.0382961365952319e-02
GC_9_154 b_9 NI_9 NS_154 0 -1.8956109124575876e-02
GC_9_155 b_9 NI_9 NS_155 0 -1.2229038087963495e-01
GC_9_156 b_9 NI_9 NS_156 0 6.7052044479621722e-02
GC_9_157 b_9 NI_9 NS_157 0 -2.3662110864315716e-02
GC_9_158 b_9 NI_9 NS_158 0 1.2239199059846839e-02
GC_9_159 b_9 NI_9 NS_159 0 2.4212290113314019e-02
GC_9_160 b_9 NI_9 NS_160 0 -6.5693075875292134e-02
GC_9_161 b_9 NI_9 NS_161 0 9.7646980274384339e-03
GC_9_162 b_9 NI_9 NS_162 0 -1.3948793479294420e-05
GC_9_163 b_9 NI_9 NS_163 0 2.4707412377460436e-13
GC_9_164 b_9 NI_9 NS_164 0 -3.3612310995843697e-07
GC_9_165 b_9 NI_9 NS_165 0 -1.8185656468472924e-05
GC_9_166 b_9 NI_9 NS_166 0 -4.6199027518140825e-06
GC_9_167 b_9 NI_9 NS_167 0 -1.8582383122872255e-03
GC_9_168 b_9 NI_9 NS_168 0 -1.1618210813343336e-02
GC_9_169 b_9 NI_9 NS_169 0 -2.7110116349494343e-02
GC_9_170 b_9 NI_9 NS_170 0 4.1370517465618732e-03
GC_9_171 b_9 NI_9 NS_171 0 1.3707091961262435e-02
GC_9_172 b_9 NI_9 NS_172 0 3.3729475712676420e-02
GC_9_173 b_9 NI_9 NS_173 0 -1.0121840316874192e-02
GC_9_174 b_9 NI_9 NS_174 0 -1.1019446233926510e-03
GC_9_175 b_9 NI_9 NS_175 0 2.5203510468226692e-02
GC_9_176 b_9 NI_9 NS_176 0 3.4344075355729337e-02
GC_9_177 b_9 NI_9 NS_177 0 -3.7864915734637816e-03
GC_9_178 b_9 NI_9 NS_178 0 -6.7149129460149070e-06
GC_9_179 b_9 NI_9 NS_179 0 2.4804447355673485e-13
GC_9_180 b_9 NI_9 NS_180 0 -1.1920879156714809e-08
GC_9_181 b_9 NI_9 NS_181 0 -4.9382742309299040e-05
GC_9_182 b_9 NI_9 NS_182 0 1.1500099475696079e-05
GC_9_183 b_9 NI_9 NS_183 0 -2.9134859513938183e-03
GC_9_184 b_9 NI_9 NS_184 0 -2.2858663501166680e-03
GC_9_185 b_9 NI_9 NS_185 0 -6.9716540015497585e-03
GC_9_186 b_9 NI_9 NS_186 0 1.0620071524246638e-03
GC_9_187 b_9 NI_9 NS_187 0 -8.3521619052031506e-03
GC_9_188 b_9 NI_9 NS_188 0 3.0378092842247885e-02
GC_9_189 b_9 NI_9 NS_189 0 1.0625813540673211e-02
GC_9_190 b_9 NI_9 NS_190 0 -3.5509426634026394e-04
GC_9_191 b_9 NI_9 NS_191 0 1.6729245384958086e-02
GC_9_192 b_9 NI_9 NS_192 0 7.6374167087320073e-03
GD_9_1 b_9 NI_9 NA_1 0 -1.9644716021815505e-05
GD_9_2 b_9 NI_9 NA_2 0 -9.6408825624290336e-06
GD_9_3 b_9 NI_9 NA_3 0 -1.5086858373049078e-04
GD_9_4 b_9 NI_9 NA_4 0 3.5971827455118786e-05
GD_9_5 b_9 NI_9 NA_5 0 1.2302838217287811e-03
GD_9_6 b_9 NI_9 NA_6 0 1.5553807253317785e-03
GD_9_7 b_9 NI_9 NA_7 0 1.2919463503727163e-03
GD_9_8 b_9 NI_9 NA_8 0 -1.8766376825671608e-03
GD_9_9 b_9 NI_9 NA_9 0 -3.4687299564332780e-02
GD_9_10 b_9 NI_9 NA_10 0 -1.6361108648325323e-02
GD_9_11 b_9 NI_9 NA_11 0 4.7466897934198308e-03
GD_9_12 b_9 NI_9 NA_12 0 -5.0216068559711747e-03
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 2.2119275238874653e-05
GC_10_2 b_10 NI_10 NS_2 0 4.5743982783698239e-09
GC_10_3 b_10 NI_10 NS_3 0 3.4028111137934281e-15
GC_10_4 b_10 NI_10 NS_4 0 -3.8840872464666749e-10
GC_10_5 b_10 NI_10 NS_5 0 -4.9107612433468920e-08
GC_10_6 b_10 NI_10 NS_6 0 1.7203227307015861e-08
GC_10_7 b_10 NI_10 NS_7 0 -2.6247205088846106e-06
GC_10_8 b_10 NI_10 NS_8 0 3.2081765725003273e-06
GC_10_9 b_10 NI_10 NS_9 0 3.1791851171494243e-06
GC_10_10 b_10 NI_10 NS_10 0 -1.9230748856245417e-06
GC_10_11 b_10 NI_10 NS_11 0 1.2311696336766057e-06
GC_10_12 b_10 NI_10 NS_12 0 -9.8431512474164809e-06
GC_10_13 b_10 NI_10 NS_13 0 -4.6406134249574798e-06
GC_10_14 b_10 NI_10 NS_14 0 7.9180975595243106e-07
GC_10_15 b_10 NI_10 NS_15 0 -8.4570546264112864e-06
GC_10_16 b_10 NI_10 NS_16 0 -5.5174435340256207e-06
GC_10_17 b_10 NI_10 NS_17 0 7.9935434163174067e-05
GC_10_18 b_10 NI_10 NS_18 0 5.1336417679910985e-08
GC_10_19 b_10 NI_10 NS_19 0 3.3838984317328122e-15
GC_10_20 b_10 NI_10 NS_20 0 -9.6421093678841851e-10
GC_10_21 b_10 NI_10 NS_21 0 -2.2531669109669770e-07
GC_10_22 b_10 NI_10 NS_22 0 6.5684082024459943e-08
GC_10_23 b_10 NI_10 NS_23 0 -1.4101659912621390e-06
GC_10_24 b_10 NI_10 NS_24 0 -5.7416068915966753e-06
GC_10_25 b_10 NI_10 NS_25 0 -4.3940176236486289e-06
GC_10_26 b_10 NI_10 NS_26 0 -4.7547917578019262e-06
GC_10_27 b_10 NI_10 NS_27 0 -1.6650797496614348e-05
GC_10_28 b_10 NI_10 NS_28 0 -2.2976339808895000e-05
GC_10_29 b_10 NI_10 NS_29 0 -8.1578925097982126e-06
GC_10_30 b_10 NI_10 NS_30 0 4.0242996222732091e-06
GC_10_31 b_10 NI_10 NS_31 0 -2.0894058480400915e-05
GC_10_32 b_10 NI_10 NS_32 0 -8.4433143944921164e-06
GC_10_33 b_10 NI_10 NS_33 0 2.0506449024154850e-05
GC_10_34 b_10 NI_10 NS_34 0 -2.1073735103997632e-08
GC_10_35 b_10 NI_10 NS_35 0 9.1432053600592069e-15
GC_10_36 b_10 NI_10 NS_36 0 2.4616232464354995e-09
GC_10_37 b_10 NI_10 NS_37 0 3.6421134340316709e-07
GC_10_38 b_10 NI_10 NS_38 0 -1.2255406235181875e-07
GC_10_39 b_10 NI_10 NS_39 0 1.8673851763436220e-05
GC_10_40 b_10 NI_10 NS_40 0 2.3690733120679359e-05
GC_10_41 b_10 NI_10 NS_41 0 6.0298835622667033e-05
GC_10_42 b_10 NI_10 NS_42 0 -6.9695482450759352e-06
GC_10_43 b_10 NI_10 NS_43 0 7.3526062299136797e-05
GC_10_44 b_10 NI_10 NS_44 0 -2.3641677516930630e-04
GC_10_45 b_10 NI_10 NS_45 0 -8.4914480481993297e-05
GC_10_46 b_10 NI_10 NS_46 0 2.4070386583053099e-06
GC_10_47 b_10 NI_10 NS_47 0 -1.2822977345579011e-04
GC_10_48 b_10 NI_10 NS_48 0 -6.0526075408350885e-05
GC_10_49 b_10 NI_10 NS_49 0 5.7608703120219640e-04
GC_10_50 b_10 NI_10 NS_50 0 -1.4674213268625771e-07
GC_10_51 b_10 NI_10 NS_51 0 9.3244608687296483e-15
GC_10_52 b_10 NI_10 NS_52 0 -6.6853099623153366e-09
GC_10_53 b_10 NI_10 NS_53 0 -1.5528296031781904e-06
GC_10_54 b_10 NI_10 NS_54 0 4.2150462090923766e-07
GC_10_55 b_10 NI_10 NS_55 0 -7.8458753732288548e-06
GC_10_56 b_10 NI_10 NS_56 0 -3.5377891600324235e-05
GC_10_57 b_10 NI_10 NS_57 0 -2.3002141108941712e-05
GC_10_58 b_10 NI_10 NS_58 0 -4.0672851599620635e-05
GC_10_59 b_10 NI_10 NS_59 0 -1.2955330818076121e-04
GC_10_60 b_10 NI_10 NS_60 0 -1.6495209250749694e-04
GC_10_61 b_10 NI_10 NS_61 0 -5.0632770468033536e-05
GC_10_62 b_10 NI_10 NS_62 0 2.6200842237287966e-05
GC_10_63 b_10 NI_10 NS_63 0 -1.5796701995976403e-04
GC_10_64 b_10 NI_10 NS_64 0 -7.7188083936040607e-05
GC_10_65 b_10 NI_10 NS_65 0 -5.1116312075418001e-04
GC_10_66 b_10 NI_10 NS_66 0 -1.3799927796967660e-06
GC_10_67 b_10 NI_10 NS_67 0 -1.6670923713567873e-13
GC_10_68 b_10 NI_10 NS_68 0 2.7429811729503983e-08
GC_10_69 b_10 NI_10 NS_69 0 7.0011632520808519e-06
GC_10_70 b_10 NI_10 NS_70 0 -1.3818045572078834e-06
GC_10_71 b_10 NI_10 NS_71 0 6.7528070246365116e-04
GC_10_72 b_10 NI_10 NS_72 0 5.6579423363677713e-04
GC_10_73 b_10 NI_10 NS_73 0 1.6548932565212204e-03
GC_10_74 b_10 NI_10 NS_74 0 -1.2964057674855290e-04
GC_10_75 b_10 NI_10 NS_75 0 2.1436781001842940e-03
GC_10_76 b_10 NI_10 NS_76 0 -6.5225603349048124e-03
GC_10_77 b_10 NI_10 NS_77 0 -2.2924642221656337e-03
GC_10_78 b_10 NI_10 NS_78 0 2.6301233158090834e-05
GC_10_79 b_10 NI_10 NS_79 0 -3.4019261938776513e-03
GC_10_80 b_10 NI_10 NS_80 0 -1.5789970563499674e-03
GC_10_81 b_10 NI_10 NS_81 0 -4.1453292933238380e-03
GC_10_82 b_10 NI_10 NS_82 0 1.7140717507762649e-06
GC_10_83 b_10 NI_10 NS_83 0 -1.6584678855222335e-13
GC_10_84 b_10 NI_10 NS_84 0 4.6782114194276408e-08
GC_10_85 b_10 NI_10 NS_85 0 1.3497091602594379e-05
GC_10_86 b_10 NI_10 NS_86 0 -3.8200055657187723e-06
GC_10_87 b_10 NI_10 NS_87 0 2.5293961013092601e-05
GC_10_88 b_10 NI_10 NS_88 0 2.4714433675054382e-05
GC_10_89 b_10 NI_10 NS_89 0 -3.8942798527382522e-04
GC_10_90 b_10 NI_10 NS_90 0 3.7374090831979504e-04
GC_10_91 b_10 NI_10 NS_91 0 1.1950111179570254e-03
GC_10_92 b_10 NI_10 NS_92 0 1.9767902425477223e-03
GC_10_93 b_10 NI_10 NS_93 0 1.9587725746407264e-04
GC_10_94 b_10 NI_10 NS_94 0 -2.0846776367463944e-04
GC_10_95 b_10 NI_10 NS_95 0 1.7516603043650359e-03
GC_10_96 b_10 NI_10 NS_96 0 1.3455865934461539e-03
GC_10_97 b_10 NI_10 NS_97 0 -1.7406020937752119e-03
GC_10_98 b_10 NI_10 NS_98 0 3.4170973616688832e-06
GC_10_99 b_10 NI_10 NS_99 0 1.4241742415600740e-13
GC_10_100 b_10 NI_10 NS_100 0 3.7276426027941863e-08
GC_10_101 b_10 NI_10 NS_101 0 -1.9146949361082609e-05
GC_10_102 b_10 NI_10 NS_102 0 4.6733118881730892e-06
GC_10_103 b_10 NI_10 NS_103 0 -1.0767387253174938e-03
GC_10_104 b_10 NI_10 NS_104 0 -7.5101949934678594e-04
GC_10_105 b_10 NI_10 NS_105 0 -2.6164378777632229e-03
GC_10_106 b_10 NI_10 NS_106 0 3.9727808904181482e-04
GC_10_107 b_10 NI_10 NS_107 0 -2.9076351418987401e-03
GC_10_108 b_10 NI_10 NS_108 0 1.1463330291385182e-02
GC_10_109 b_10 NI_10 NS_109 0 4.0078707020276810e-03
GC_10_110 b_10 NI_10 NS_110 0 -1.5809203425368987e-04
GC_10_111 b_10 NI_10 NS_111 0 6.2767984362089831e-03
GC_10_112 b_10 NI_10 NS_112 0 2.8068343156839154e-03
GC_10_113 b_10 NI_10 NS_113 0 5.5050582452250679e-03
GC_10_114 b_10 NI_10 NS_114 0 7.6564799803265457e-06
GC_10_115 b_10 NI_10 NS_115 0 1.3807491178181411e-13
GC_10_116 b_10 NI_10 NS_116 0 -1.9137691576114115e-07
GC_10_117 b_10 NI_10 NS_117 0 -1.3173820579021810e-05
GC_10_118 b_10 NI_10 NS_118 0 -5.1057819598319648e-07
GC_10_119 b_10 NI_10 NS_119 0 -7.6452984536688501e-04
GC_10_120 b_10 NI_10 NS_120 0 -4.6323238769425124e-03
GC_10_121 b_10 NI_10 NS_121 0 -1.0665597687106886e-02
GC_10_122 b_10 NI_10 NS_122 0 1.5152393000641160e-03
GC_10_123 b_10 NI_10 NS_123 0 4.9162392972690681e-03
GC_10_124 b_10 NI_10 NS_124 0 1.2765899736624356e-02
GC_10_125 b_10 NI_10 NS_125 0 -4.0675659715885965e-03
GC_10_126 b_10 NI_10 NS_126 0 -3.1202683755084489e-04
GC_10_127 b_10 NI_10 NS_127 0 9.4893216436898707e-03
GC_10_128 b_10 NI_10 NS_128 0 1.3304656449509799e-02
GC_10_129 b_10 NI_10 NS_129 0 1.9563059077350026e-01
GC_10_130 b_10 NI_10 NS_130 0 6.1042623914342407e-05
GC_10_131 b_10 NI_10 NS_131 0 3.3895647636170156e-12
GC_10_132 b_10 NI_10 NS_132 0 4.1869103389072592e-06
GC_10_133 b_10 NI_10 NS_133 0 1.2035869483929546e-04
GC_10_134 b_10 NI_10 NS_134 0 4.6692498212275532e-05
GC_10_135 b_10 NI_10 NS_135 0 -6.0783095951076310e-02
GC_10_136 b_10 NI_10 NS_136 0 -4.3809843663656430e-02
GC_10_137 b_10 NI_10 NS_137 0 4.0382204922112613e-02
GC_10_138 b_10 NI_10 NS_138 0 -1.8956465905449603e-02
GC_10_139 b_10 NI_10 NS_139 0 -1.2229413549360559e-01
GC_10_140 b_10 NI_10 NS_140 0 6.7052443117781635e-02
GC_10_141 b_10 NI_10 NS_141 0 -2.3661967843010841e-02
GC_10_142 b_10 NI_10 NS_142 0 1.2240381584028456e-02
GC_10_143 b_10 NI_10 NS_143 0 2.4213240263797536e-02
GC_10_144 b_10 NI_10 NS_144 0 -6.5688245067041170e-02
GC_10_145 b_10 NI_10 NS_145 0 5.8302073720192055e-02
GC_10_146 b_10 NI_10 NS_146 0 -6.5905950168083563e-06
GC_10_147 b_10 NI_10 NS_147 0 -1.1643763236597675e-12
GC_10_148 b_10 NI_10 NS_148 0 -2.4306521305599706e-06
GC_10_149 b_10 NI_10 NS_149 0 2.8122693983717822e-05
GC_10_150 b_10 NI_10 NS_150 0 -4.6575585171111395e-06
GC_10_151 b_10 NI_10 NS_151 0 -1.5283049652664697e-03
GC_10_152 b_10 NI_10 NS_152 0 7.1123687452975468e-03
GC_10_153 b_10 NI_10 NS_153 0 1.7510548009446479e-02
GC_10_154 b_10 NI_10 NS_154 0 -5.4949007198397560e-03
GC_10_155 b_10 NI_10 NS_155 0 -2.5483258611382360e-02
GC_10_156 b_10 NI_10 NS_156 0 -3.1166764838095364e-02
GC_10_157 b_10 NI_10 NS_157 0 7.4119524626673206e-03
GC_10_158 b_10 NI_10 NS_158 0 2.8757567457169241e-03
GC_10_159 b_10 NI_10 NS_159 0 -3.0802399971382954e-02
GC_10_160 b_10 NI_10 NS_160 0 -3.3514465395643366e-02
GC_10_161 b_10 NI_10 NS_161 0 -3.7839734259171864e-03
GC_10_162 b_10 NI_10 NS_162 0 -6.9187786676171825e-06
GC_10_163 b_10 NI_10 NS_163 0 2.4799543039044478e-13
GC_10_164 b_10 NI_10 NS_164 0 -1.1843657792129593e-08
GC_10_165 b_10 NI_10 NS_165 0 -4.9359374570938963e-05
GC_10_166 b_10 NI_10 NS_166 0 1.1494328619569558e-05
GC_10_167 b_10 NI_10 NS_167 0 -2.9134804065403127e-03
GC_10_168 b_10 NI_10 NS_168 0 -2.2859929737860211e-03
GC_10_169 b_10 NI_10 NS_169 0 -6.9716484917650848e-03
GC_10_170 b_10 NI_10 NS_170 0 1.0618195442934127e-03
GC_10_171 b_10 NI_10 NS_171 0 -8.3523603835182186e-03
GC_10_172 b_10 NI_10 NS_172 0 3.0377092803694307e-02
GC_10_173 b_10 NI_10 NS_173 0 1.0625545332111630e-02
GC_10_174 b_10 NI_10 NS_174 0 -3.5514832565747116e-04
GC_10_175 b_10 NI_10 NS_175 0 1.6728109393441805e-02
GC_10_176 b_10 NI_10 NS_176 0 7.6358555393304375e-03
GC_10_177 b_10 NI_10 NS_177 0 9.7641343668942015e-03
GC_10_178 b_10 NI_10 NS_178 0 -1.4048250753154480e-05
GC_10_179 b_10 NI_10 NS_179 0 2.4705989938805609e-13
GC_10_180 b_10 NI_10 NS_180 0 -3.3605987151731390e-07
GC_10_181 b_10 NI_10 NS_181 0 -1.8169871426358643e-05
GC_10_182 b_10 NI_10 NS_182 0 -4.6241849715583297e-06
GC_10_183 b_10 NI_10 NS_183 0 -1.8582510064197404e-03
GC_10_184 b_10 NI_10 NS_184 0 -1.1618235131344024e-02
GC_10_185 b_10 NI_10 NS_185 0 -2.7110126205266157e-02
GC_10_186 b_10 NI_10 NS_186 0 4.1371886714540416e-03
GC_10_187 b_10 NI_10 NS_187 0 1.3707549391878938e-02
GC_10_188 b_10 NI_10 NS_188 0 3.3729551535474314e-02
GC_10_189 b_10 NI_10 NS_189 0 -1.0121849139815038e-02
GC_10_190 b_10 NI_10 NS_190 0 -1.1020620058801271e-03
GC_10_191 b_10 NI_10 NS_191 0 2.5203473168714092e-02
GC_10_192 b_10 NI_10 NS_192 0 3.4343566603960998e-02
GD_10_1 b_10 NI_10 NA_1 0 -9.6395497821355686e-06
GD_10_2 b_10 NI_10 NA_2 0 -1.9739871924578357e-05
GD_10_3 b_10 NI_10 NA_3 0 3.6137465638472004e-05
GD_10_4 b_10 NI_10 NA_4 0 -1.5088462180394164e-04
GD_10_5 b_10 NI_10 NA_5 0 1.5553121323494785e-03
GD_10_6 b_10 NI_10 NA_6 0 1.2291457743062663e-03
GD_10_7 b_10 NI_10 NA_7 0 -1.8761184885585480e-03
GD_10_8 b_10 NI_10 NA_8 0 1.2918219760920733e-03
GD_10_9 b_10 NI_10 NA_9 0 -1.6364566438648483e-02
GD_10_10 b_10 NI_10 NA_10 0 -3.4681038826393652e-02
GD_10_11 b_10 NI_10 NA_11 0 -5.0221216256232538e-03
GD_10_12 b_10 NI_10 NA_12 0 4.7468659666572970e-03
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 9.1075113336638307e-06
GC_11_2 b_11 NI_11 NS_2 0 -5.4733794775662118e-11
GC_11_3 b_11 NI_11 NS_3 0 -9.9062283444200456e-16
GC_11_4 b_11 NI_11 NS_4 0 -1.5773193269437166e-10
GC_11_5 b_11 NI_11 NS_5 0 -4.3660507033947705e-08
GC_11_6 b_11 NI_11 NS_6 0 1.7498273091226080e-08
GC_11_7 b_11 NI_11 NS_7 0 -5.6994077731473896e-07
GC_11_8 b_11 NI_11 NS_8 0 -1.6159800278530146e-06
GC_11_9 b_11 NI_11 NS_9 0 -3.1702374656274930e-06
GC_11_10 b_11 NI_11 NS_10 0 6.9394824147322155e-08
GC_11_11 b_11 NI_11 NS_11 0 2.6916827272382062e-07
GC_11_12 b_11 NI_11 NS_12 0 2.5898974285843566e-06
GC_11_13 b_11 NI_11 NS_13 0 -1.1424511483908018e-06
GC_11_14 b_11 NI_11 NS_14 0 -5.5946485768767386e-07
GC_11_15 b_11 NI_11 NS_15 0 -2.6422521455756709e-07
GC_11_16 b_11 NI_11 NS_16 0 1.0913622236508704e-06
GC_11_17 b_11 NI_11 NS_17 0 8.6589945365994225e-06
GC_11_18 b_11 NI_11 NS_18 0 -8.8475152491517554e-09
GC_11_19 b_11 NI_11 NS_19 0 -9.7886161566283663e-16
GC_11_20 b_11 NI_11 NS_20 0 9.8400723054480753e-11
GC_11_21 b_11 NI_11 NS_21 0 3.1547875504542483e-08
GC_11_22 b_11 NI_11 NS_22 0 -1.3740675323490961e-08
GC_11_23 b_11 NI_11 NS_23 0 -2.8506214256307990e-06
GC_11_24 b_11 NI_11 NS_24 0 2.4730760192193413e-06
GC_11_25 b_11 NI_11 NS_25 0 4.8737710062987554e-07
GC_11_26 b_11 NI_11 NS_26 0 -2.0951117520569557e-06
GC_11_27 b_11 NI_11 NS_27 0 1.2467702161520636e-06
GC_11_28 b_11 NI_11 NS_28 0 2.4328796841675783e-06
GC_11_29 b_11 NI_11 NS_29 0 -1.5009783603967409e-06
GC_11_30 b_11 NI_11 NS_30 0 3.6509709477122969e-07
GC_11_31 b_11 NI_11 NS_31 0 -3.2124952843965179e-07
GC_11_32 b_11 NI_11 NS_32 0 -7.4420291499310980e-07
GC_11_33 b_11 NI_11 NS_33 0 8.1337621775396277e-05
GC_11_34 b_11 NI_11 NS_34 0 -2.2240789430556961e-08
GC_11_35 b_11 NI_11 NS_35 0 3.4395523694472227e-15
GC_11_36 b_11 NI_11 NS_36 0 -9.4833201388269050e-10
GC_11_37 b_11 NI_11 NS_37 0 -2.1748681409392924e-07
GC_11_38 b_11 NI_11 NS_38 0 6.3868366091799794e-08
GC_11_39 b_11 NI_11 NS_39 0 -1.4302855266226140e-06
GC_11_40 b_11 NI_11 NS_40 0 -5.8090906397348600e-06
GC_11_41 b_11 NI_11 NS_41 0 -4.4251618895561599e-06
GC_11_42 b_11 NI_11 NS_42 0 -4.8379620016880379e-06
GC_11_43 b_11 NI_11 NS_43 0 -1.6839453713221730e-05
GC_11_44 b_11 NI_11 NS_44 0 -2.3393345560403074e-05
GC_11_45 b_11 NI_11 NS_45 0 -8.2695920600449368e-06
GC_11_46 b_11 NI_11 NS_46 0 4.0292901336456155e-06
GC_11_47 b_11 NI_11 NS_47 0 -2.1378690643079857e-05
GC_11_48 b_11 NI_11 NS_48 0 -9.0306483710774948e-06
GC_11_49 b_11 NI_11 NS_49 0 2.2236622567205171e-05
GC_11_50 b_11 NI_11 NS_50 0 -1.0074078974222791e-08
GC_11_51 b_11 NI_11 NS_51 0 3.4197506027658642e-15
GC_11_52 b_11 NI_11 NS_52 0 -3.8753280891742728e-10
GC_11_53 b_11 NI_11 NS_53 0 -4.7696527551389257e-08
GC_11_54 b_11 NI_11 NS_54 0 1.6907214703236759e-08
GC_11_55 b_11 NI_11 NS_55 0 -2.6188755140442299e-06
GC_11_56 b_11 NI_11 NS_56 0 3.2028839258574255e-06
GC_11_57 b_11 NI_11 NS_57 0 3.1871147672872440e-06
GC_11_58 b_11 NI_11 NS_58 0 -1.9344237001809394e-06
GC_11_59 b_11 NI_11 NS_59 0 1.2401019650132631e-06
GC_11_60 b_11 NI_11 NS_60 0 -9.9247887391870140e-06
GC_11_61 b_11 NI_11 NS_61 0 -4.6637366821434787e-06
GC_11_62 b_11 NI_11 NS_62 0 7.8345590434921858e-07
GC_11_63 b_11 NI_11 NS_63 0 -8.5411477727863900e-06
GC_11_64 b_11 NI_11 NS_64 0 -5.6364578391214139e-06
GC_11_65 b_11 NI_11 NS_65 0 1.4735110530203425e-03
GC_11_66 b_11 NI_11 NS_66 0 -3.7422394291817194e-07
GC_11_67 b_11 NI_11 NS_67 0 2.0706701640243327e-14
GC_11_68 b_11 NI_11 NS_68 0 -1.6099242927263318e-08
GC_11_69 b_11 NI_11 NS_69 0 -3.8268870409445698e-06
GC_11_70 b_11 NI_11 NS_70 0 1.0177298416704687e-06
GC_11_71 b_11 NI_11 NS_71 0 -1.9623230369171674e-05
GC_11_72 b_11 NI_11 NS_72 0 -8.8853535128423830e-05
GC_11_73 b_11 NI_11 NS_73 0 -5.5048080911938993e-05
GC_11_74 b_11 NI_11 NS_74 0 -1.0543635125801715e-04
GC_11_75 b_11 NI_11 NS_75 0 -3.3159387375498734e-04
GC_11_76 b_11 NI_11 NS_76 0 -4.2819645549459516e-04
GC_11_77 b_11 NI_11 NS_77 0 -1.2973430143234399e-04
GC_11_78 b_11 NI_11 NS_78 0 6.5860850261969836e-05
GC_11_79 b_11 NI_11 NS_79 0 -4.1018447718774176e-04
GC_11_80 b_11 NI_11 NS_80 0 -2.0277129409686204e-04
GC_11_81 b_11 NI_11 NS_81 0 -1.1933664602634772e-04
GC_11_82 b_11 NI_11 NS_82 0 -4.5602931743174164e-08
GC_11_83 b_11 NI_11 NS_83 0 2.0512382325376512e-14
GC_11_84 b_11 NI_11 NS_84 0 5.1585743761202189e-09
GC_11_85 b_11 NI_11 NS_85 0 7.9172495162485870e-07
GC_11_86 b_11 NI_11 NS_86 0 -2.5103866945136490e-07
GC_11_87 b_11 NI_11 NS_87 0 6.1204716224100826e-05
GC_11_88 b_11 NI_11 NS_88 0 6.1410287358497250e-05
GC_11_89 b_11 NI_11 NS_89 0 1.6109023006616972e-04
GC_11_90 b_11 NI_11 NS_90 0 -4.5952614577605459e-06
GC_11_91 b_11 NI_11 NS_91 0 2.3885609574643809e-04
GC_11_92 b_11 NI_11 NS_92 0 -6.0024941529810251e-04
GC_11_93 b_11 NI_11 NS_93 0 -2.1680961671000822e-04
GC_11_94 b_11 NI_11 NS_94 0 -4.6174837166720860e-06
GC_11_95 b_11 NI_11 NS_95 0 -3.1215666900048051e-04
GC_11_96 b_11 NI_11 NS_96 0 -1.5292694958830491e-04
GC_11_97 b_11 NI_11 NS_97 0 -4.1524693868362980e-03
GC_11_98 b_11 NI_11 NS_98 0 1.7202739205252622e-06
GC_11_99 b_11 NI_11 NS_99 0 -1.6979668978374798e-13
GC_11_100 b_11 NI_11 NS_100 0 4.6451070295484267e-08
GC_11_101 b_11 NI_11 NS_101 0 1.3500910559535535e-05
GC_11_102 b_11 NI_11 NS_102 0 -3.8167386028507314e-06
GC_11_103 b_11 NI_11 NS_103 0 2.5167833418765002e-05
GC_11_104 b_11 NI_11 NS_104 0 2.5213245630249068e-05
GC_11_105 b_11 NI_11 NS_105 0 -3.8970306868505366e-04
GC_11_106 b_11 NI_11 NS_106 0 3.7440246562122969e-04
GC_11_107 b_11 NI_11 NS_107 0 1.1968571210668273e-03
GC_11_108 b_11 NI_11 NS_108 0 1.9813592973353228e-03
GC_11_109 b_11 NI_11 NS_109 0 1.9711006594005999e-04
GC_11_110 b_11 NI_11 NS_110 0 -2.0917726696089537e-04
GC_11_111 b_11 NI_11 NS_111 0 1.7545600406715137e-03
GC_11_112 b_11 NI_11 NS_112 0 1.3468124232981120e-03
GC_11_113 b_11 NI_11 NS_113 0 -5.1000519814260064e-04
GC_11_114 b_11 NI_11 NS_114 0 -1.3763374944598162e-06
GC_11_115 b_11 NI_11 NS_115 0 -1.7067509949749102e-13
GC_11_116 b_11 NI_11 NS_116 0 2.8023640407365982e-08
GC_11_117 b_11 NI_11 NS_117 0 7.0316617346256222e-06
GC_11_118 b_11 NI_11 NS_118 0 -1.3983975704863844e-06
GC_11_119 b_11 NI_11 NS_119 0 6.7656863455211875e-04
GC_11_120 b_11 NI_11 NS_120 0 5.6601003688081821e-04
GC_11_121 b_11 NI_11 NS_121 0 1.6569348898511492e-03
GC_11_122 b_11 NI_11 NS_122 0 -1.3047347969266830e-04
GC_11_123 b_11 NI_11 NS_123 0 2.1461417789966773e-03
GC_11_124 b_11 NI_11 NS_124 0 -6.5332264070953466e-03
GC_11_125 b_11 NI_11 NS_125 0 -2.2964558845839523e-03
GC_11_126 b_11 NI_11 NS_126 0 2.6316675724386351e-05
GC_11_127 b_11 NI_11 NS_127 0 -3.4079702074384919e-03
GC_11_128 b_11 NI_11 NS_128 0 -1.5814656580351201e-03
GC_11_129 b_11 NI_11 NS_129 0 9.3917094913053955e-03
GC_11_130 b_11 NI_11 NS_130 0 1.2870475247296324e-05
GC_11_131 b_11 NI_11 NS_131 0 2.5386271570619567e-13
GC_11_132 b_11 NI_11 NS_132 0 -3.4311216729063255e-07
GC_11_133 b_11 NI_11 NS_133 0 -2.1088335054396739e-05
GC_11_134 b_11 NI_11 NS_134 0 -3.9317522293036448e-06
GC_11_135 b_11 NI_11 NS_135 0 -1.8572960020416787e-03
GC_11_136 b_11 NI_11 NS_136 0 -1.1603164508792676e-02
GC_11_137 b_11 NI_11 NS_137 0 -2.7111003517445519e-02
GC_11_138 b_11 NI_11 NS_138 0 4.1602579803196576e-03
GC_11_139 b_11 NI_11 NS_139 0 1.3734287535951758e-02
GC_11_140 b_11 NI_11 NS_140 0 3.3872423240372228e-02
GC_11_141 b_11 NI_11 NS_141 0 -1.0082692743939982e-02
GC_11_142 b_11 NI_11 NS_142 0 -1.0952613566719085e-03
GC_11_143 b_11 NI_11 NS_143 0 2.5364111278142341e-02
GC_11_144 b_11 NI_11 NS_144 0 3.4556097974818907e-02
GC_11_145 b_11 NI_11 NS_145 0 -3.8116937809492524e-03
GC_11_146 b_11 NI_11 NS_146 0 4.0624524229200693e-06
GC_11_147 b_11 NI_11 NS_147 0 2.6117212374988533e-13
GC_11_148 b_11 NI_11 NS_148 0 -1.2936475546777570e-08
GC_11_149 b_11 NI_11 NS_149 0 -5.0427908808713245e-05
GC_11_150 b_11 NI_11 NS_150 0 1.1717849140240677e-05
GC_11_151 b_11 NI_11 NS_151 0 -2.9195292853919650e-03
GC_11_152 b_11 NI_11 NS_152 0 -2.2869752431779757e-03
GC_11_153 b_11 NI_11 NS_153 0 -6.9814375227679566e-03
GC_11_154 b_11 NI_11 NS_154 0 1.0662539369709920e-03
GC_11_155 b_11 NI_11 NS_155 0 -8.3762742659540187e-03
GC_11_156 b_11 NI_11 NS_156 0 3.0424387387227424e-02
GC_11_157 b_11 NI_11 NS_157 0 1.0638709248842000e-02
GC_11_158 b_11 NI_11 NS_158 0 -3.4452938558611219e-04
GC_11_159 b_11 NI_11 NS_159 0 1.6779086523598542e-02
GC_11_160 b_11 NI_11 NS_160 0 7.7221173242471696e-03
GC_11_161 b_11 NI_11 NS_161 0 6.0205323372037767e-02
GC_11_162 b_11 NI_11 NS_162 0 7.0901804757799690e-06
GC_11_163 b_11 NI_11 NS_163 0 -1.1476404740054533e-12
GC_11_164 b_11 NI_11 NS_164 0 -2.4577415901833895e-06
GC_11_165 b_11 NI_11 NS_165 0 2.1425300733544325e-05
GC_11_166 b_11 NI_11 NS_166 0 -3.0074083276946602e-06
GC_11_167 b_11 NI_11 NS_167 0 -1.5768800580942355e-03
GC_11_168 b_11 NI_11 NS_168 0 6.8779680937498585e-03
GC_11_169 b_11 NI_11 NS_169 0 1.7132712095719791e-02
GC_11_170 b_11 NI_11 NS_170 0 -5.5821303109003751e-03
GC_11_171 b_11 NI_11 NS_171 0 -2.5778399771245797e-02
GC_11_172 b_11 NI_11 NS_172 0 -3.1260470539679196e-02
GC_11_173 b_11 NI_11 NS_173 0 7.1572631031797951e-03
GC_11_174 b_11 NI_11 NS_174 0 2.9562126288017422e-03
GC_11_175 b_11 NI_11 NS_175 0 -3.0968398510784065e-02
GC_11_176 b_11 NI_11 NS_176 0 -3.3276432946358486e-02
GC_11_177 b_11 NI_11 NS_177 0 1.9531990624724319e-01
GC_11_178 b_11 NI_11 NS_178 0 1.1089949296769764e-04
GC_11_179 b_11 NI_11 NS_179 0 1.5678424309695368e-12
GC_11_180 b_11 NI_11 NS_180 0 4.4033140177286095e-06
GC_11_181 b_11 NI_11 NS_181 0 1.1663679510842817e-04
GC_11_182 b_11 NI_11 NS_182 0 4.6012193235557817e-05
GC_11_183 b_11 NI_11 NS_183 0 -6.1176636152861438e-02
GC_11_184 b_11 NI_11 NS_184 0 -4.4021406027253955e-02
GC_11_185 b_11 NI_11 NS_185 0 3.9561856052839510e-02
GC_11_186 b_11 NI_11 NS_186 0 -1.8838344768229969e-02
GC_11_187 b_11 NI_11 NS_187 0 -1.2336117729326648e-01
GC_11_188 b_11 NI_11 NS_188 0 7.0714443646176739e-02
GC_11_189 b_11 NI_11 NS_189 0 -2.2401414341780682e-02
GC_11_190 b_11 NI_11 NS_190 0 1.2250561272138621e-02
GC_11_191 b_11 NI_11 NS_191 0 2.6304168999551913e-02
GC_11_192 b_11 NI_11 NS_192 0 -6.4427105496198109e-02
GD_11_1 b_11 NI_11 NA_1 0 -2.1460113886217121e-06
GD_11_2 b_11 NI_11 NA_2 0 -3.8758308714656937e-06
GD_11_3 b_11 NI_11 NA_3 0 -2.0125964040036315e-05
GD_11_4 b_11 NI_11 NA_4 0 -9.6472272824813411e-06
GD_11_5 b_11 NI_11 NA_5 0 -3.8461760294061992e-04
GD_11_6 b_11 NI_11 NA_6 0 1.6482072202236820e-04
GD_11_7 b_11 NI_11 NA_7 0 1.2298426472795393e-03
GD_11_8 b_11 NI_11 NA_8 0 1.5589941559713200e-03
GD_11_9 b_11 NI_11 NA_9 0 4.8388259879316216e-03
GD_11_10 b_11 NI_11 NA_10 0 -5.0311289137721059e-03
GD_11_11 b_11 NI_11 NA_11 0 -3.5123762934377932e-02
GD_11_12 b_11 NI_11 NA_12 0 -1.7153463095995213e-02
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 8.6710727068003231e-06
GC_12_2 b_12 NI_12 NS_2 0 -8.8693872083519922e-09
GC_12_3 b_12 NI_12 NS_3 0 -9.7872216948720694e-16
GC_12_4 b_12 NI_12 NS_4 0 9.8050344366897581e-11
GC_12_5 b_12 NI_12 NS_5 0 3.1496406380341183e-08
GC_12_6 b_12 NI_12 NS_6 0 -1.3723171912876780e-08
GC_12_7 b_12 NI_12 NS_7 0 -2.8503080955826167e-06
GC_12_8 b_12 NI_12 NS_8 0 2.4728473286741023e-06
GC_12_9 b_12 NI_12 NS_9 0 4.8801974326467150e-07
GC_12_10 b_12 NI_12 NS_10 0 -2.0960563683232102e-06
GC_12_11 b_12 NI_12 NS_11 0 1.2450044771532780e-06
GC_12_12 b_12 NI_12 NS_12 0 2.4243933334752879e-06
GC_12_13 b_12 NI_12 NS_13 0 -1.5033986241279559e-06
GC_12_14 b_12 NI_12 NS_14 0 3.6646638819379838e-07
GC_12_15 b_12 NI_12 NS_15 0 -3.2644648538806129e-07
GC_12_16 b_12 NI_12 NS_16 0 -7.4696672965475627e-07
GC_12_17 b_12 NI_12 NS_17 0 9.1083800567208458e-06
GC_12_18 b_12 NI_12 NS_18 0 -1.2580628327180148e-10
GC_12_19 b_12 NI_12 NS_19 0 -9.9059911702724387e-16
GC_12_20 b_12 NI_12 NS_20 0 -1.5771801273570259e-10
GC_12_21 b_12 NI_12 NS_21 0 -4.3653312276925353e-08
GC_12_22 b_12 NI_12 NS_22 0 1.7496658727155016e-08
GC_12_23 b_12 NI_12 NS_23 0 -5.6993159274932852e-07
GC_12_24 b_12 NI_12 NS_24 0 -1.6160171643372833e-06
GC_12_25 b_12 NI_12 NS_25 0 -3.1702244488663693e-06
GC_12_26 b_12 NI_12 NS_26 0 6.9332736072078161e-08
GC_12_27 b_12 NI_12 NS_27 0 2.6913490757824911e-07
GC_12_28 b_12 NI_12 NS_28 0 2.5895027487000970e-06
GC_12_29 b_12 NI_12 NS_29 0 -1.1425621007036362e-06
GC_12_30 b_12 NI_12 NS_30 0 -5.5949177506357027e-07
GC_12_31 b_12 NI_12 NS_31 0 -2.6465764737911885e-07
GC_12_32 b_12 NI_12 NS_32 0 1.0907858023125197e-06
GC_12_33 b_12 NI_12 NS_33 0 2.2234082318352182e-05
GC_12_34 b_12 NI_12 NS_34 0 -9.9394728766550696e-09
GC_12_35 b_12 NI_12 NS_35 0 3.4195806139884398e-15
GC_12_36 b_12 NI_12 NS_36 0 -3.8753863413714940e-10
GC_12_37 b_12 NI_12 NS_37 0 -4.7707527319332941e-08
GC_12_38 b_12 NI_12 NS_38 0 1.6909545976828535e-08
GC_12_39 b_12 NI_12 NS_39 0 -2.6190944671917111e-06
GC_12_40 b_12 NI_12 NS_40 0 3.2032594502529045e-06
GC_12_41 b_12 NI_12 NS_41 0 3.1866931716370906e-06
GC_12_42 b_12 NI_12 NS_42 0 -1.9339186511100252e-06
GC_12_43 b_12 NI_12 NS_43 0 1.2410898872770705e-06
GC_12_44 b_12 NI_12 NS_44 0 -9.9221892833316768e-06
GC_12_45 b_12 NI_12 NS_45 0 -4.6631411598478319e-06
GC_12_46 b_12 NI_12 NS_46 0 7.8320959804798861e-07
GC_12_47 b_12 NI_12 NS_47 0 -8.5394570366416382e-06
GC_12_48 b_12 NI_12 NS_48 0 -5.6350786901111697e-06
GC_12_49 b_12 NI_12 NS_49 0 8.1144836023105108e-05
GC_12_50 b_12 NI_12 NS_50 0 -2.2192337915418952e-08
GC_12_51 b_12 NI_12 NS_51 0 3.4405162392990466e-15
GC_12_52 b_12 NI_12 NS_52 0 -9.4602886258277631e-10
GC_12_53 b_12 NI_12 NS_53 0 -2.1713551091239050e-07
GC_12_54 b_12 NI_12 NS_54 0 6.3749501880380676e-08
GC_12_55 b_12 NI_12 NS_55 0 -1.4243171009333198e-06
GC_12_56 b_12 NI_12 NS_56 0 -5.8116387142715012e-06
GC_12_57 b_12 NI_12 NS_57 0 -4.4292909949009299e-06
GC_12_58 b_12 NI_12 NS_58 0 -4.8285913374122823e-06
GC_12_59 b_12 NI_12 NS_59 0 -1.6795134514612659e-05
GC_12_60 b_12 NI_12 NS_60 0 -2.3342091801274903e-05
GC_12_61 b_12 NI_12 NS_61 0 -8.2579908646071908e-06
GC_12_62 b_12 NI_12 NS_62 0 4.0171046786984908e-06
GC_12_63 b_12 NI_12 NS_63 0 -2.1338547258410183e-05
GC_12_64 b_12 NI_12 NS_64 0 -9.0137858668552587e-06
GC_12_65 b_12 NI_12 NS_65 0 -1.1792655209018123e-04
GC_12_66 b_12 NI_12 NS_66 0 -4.6304145402282422e-08
GC_12_67 b_12 NI_12 NS_67 0 2.0510612859688721e-14
GC_12_68 b_12 NI_12 NS_68 0 5.1582160940840051e-09
GC_12_69 b_12 NI_12 NS_69 0 7.9195343620399705e-07
GC_12_70 b_12 NI_12 NS_70 0 -2.5105880658638088e-07
GC_12_71 b_12 NI_12 NS_71 0 6.1103738140544565e-05
GC_12_72 b_12 NI_12 NS_72 0 6.1304875541409143e-05
GC_12_73 b_12 NI_12 NS_73 0 1.6099266752157216e-04
GC_12_74 b_12 NI_12 NS_74 0 -4.7257417745186489e-06
GC_12_75 b_12 NI_12 NS_75 0 2.3823676918369811e-04
GC_12_76 b_12 NI_12 NS_76 0 -6.0023765151425671e-04
GC_12_77 b_12 NI_12 NS_77 0 -2.1677064971494005e-04
GC_12_78 b_12 NI_12 NS_78 0 -4.4833212468429114e-06
GC_12_79 b_12 NI_12 NS_79 0 -3.1220159700124674e-04
GC_12_80 b_12 NI_12 NS_80 0 -1.5285220129125114e-04
GC_12_81 b_12 NI_12 NS_81 0 1.4734876141312089e-03
GC_12_82 b_12 NI_12 NS_82 0 -3.7230525656522257e-07
GC_12_83 b_12 NI_12 NS_83 0 2.0708523306316809e-14
GC_12_84 b_12 NI_12 NS_84 0 -1.6100148381387063e-08
GC_12_85 b_12 NI_12 NS_85 0 -3.8271169441528012e-06
GC_12_86 b_12 NI_12 NS_86 0 1.0177881003238184e-06
GC_12_87 b_12 NI_12 NS_87 0 -1.9620353235270839e-05
GC_12_88 b_12 NI_12 NS_88 0 -8.8851582865977441e-05
GC_12_89 b_12 NI_12 NS_89 0 -5.5045032216004277e-05
GC_12_90 b_12 NI_12 NS_90 0 -1.0544144878040834e-04
GC_12_91 b_12 NI_12 NS_91 0 -3.3160243395201854e-04
GC_12_92 b_12 NI_12 NS_92 0 -4.2819294642989814e-04
GC_12_93 b_12 NI_12 NS_93 0 -1.2973095473704414e-04
GC_12_94 b_12 NI_12 NS_94 0 6.5862187493095608e-05
GC_12_95 b_12 NI_12 NS_95 0 -4.1017771375680031e-04
GC_12_96 b_12 NI_12 NS_96 0 -2.0275870359170751e-04
GC_12_97 b_12 NI_12 NS_97 0 -5.0989191660364037e-04
GC_12_98 b_12 NI_12 NS_98 0 -1.3866566193946168e-06
GC_12_99 b_12 NI_12 NS_99 0 -1.7067332834635853e-13
GC_12_100 b_12 NI_12 NS_100 0 2.8023865743603637e-08
GC_12_101 b_12 NI_12 NS_101 0 7.0325158600676317e-06
GC_12_102 b_12 NI_12 NS_102 0 -1.3985622006970159e-06
GC_12_103 b_12 NI_12 NS_103 0 6.7657052300662004e-04
GC_12_104 b_12 NI_12 NS_104 0 5.6601348794055556e-04
GC_12_105 b_12 NI_12 NS_105 0 1.6569359312314474e-03
GC_12_106 b_12 NI_12 NS_106 0 -1.3047983119293921e-04
GC_12_107 b_12 NI_12 NS_107 0 2.1461555947041785e-03
GC_12_108 b_12 NI_12 NS_108 0 -6.5332695983442808e-03
GC_12_109 b_12 NI_12 NS_109 0 -2.2964698790434957e-03
GC_12_110 b_12 NI_12 NS_110 0 2.6306288294296817e-05
GC_12_111 b_12 NI_12 NS_111 0 -3.4080313647015643e-03
GC_12_112 b_12 NI_12 NS_112 0 -1.5815552385794139e-03
GC_12_113 b_12 NI_12 NS_113 0 -4.1560557775754559e-03
GC_12_114 b_12 NI_12 NS_114 0 1.7139426366545770e-06
GC_12_115 b_12 NI_12 NS_115 0 -1.6979710964731061e-13
GC_12_116 b_12 NI_12 NS_116 0 4.6458948118174903e-08
GC_12_117 b_12 NI_12 NS_117 0 1.3502704931430932e-05
GC_12_118 b_12 NI_12 NS_118 0 -3.8175248859984823e-06
GC_12_119 b_12 NI_12 NS_119 0 2.5156215264516882e-05
GC_12_120 b_12 NI_12 NS_120 0 2.5432195744922051e-05
GC_12_121 b_12 NI_12 NS_121 0 -3.8930998249809195e-04
GC_12_122 b_12 NI_12 NS_122 0 3.7478710002571928e-04
GC_12_123 b_12 NI_12 NS_123 0 1.1977043889985751e-03
GC_12_124 b_12 NI_12 NS_124 0 1.9815604496822019e-03
GC_12_125 b_12 NI_12 NS_125 0 1.9730434187730225e-04
GC_12_126 b_12 NI_12 NS_126 0 -2.0918307062500738e-04
GC_12_127 b_12 NI_12 NS_127 0 1.7552393646532863e-03
GC_12_128 b_12 NI_12 NS_128 0 1.3469542731062200e-03
GC_12_129 b_12 NI_12 NS_129 0 -3.8129262164872863e-03
GC_12_130 b_12 NI_12 NS_130 0 3.9607457613584647e-06
GC_12_131 b_12 NI_12 NS_131 0 2.6115830765524794e-13
GC_12_132 b_12 NI_12 NS_132 0 -1.2835687119094594e-08
GC_12_133 b_12 NI_12 NS_133 0 -5.0409515012063782e-05
GC_12_134 b_12 NI_12 NS_134 0 1.1712501493831180e-05
GC_12_135 b_12 NI_12 NS_135 0 -2.9194609672189534e-03
GC_12_136 b_12 NI_12 NS_136 0 -2.2869238510411986e-03
GC_12_137 b_12 NI_12 NS_137 0 -6.9813375833556813e-03
GC_12_138 b_12 NI_12 NS_138 0 1.0663020174983783e-03
GC_12_139 b_12 NI_12 NS_139 0 -8.3757776230425404e-03
GC_12_140 b_12 NI_12 NS_140 0 3.0424441558210235e-02
GC_12_141 b_12 NI_12 NS_141 0 1.0638721395726412e-02
GC_12_142 b_12 NI_12 NS_142 0 -3.4467976820512752e-04
GC_12_143 b_12 NI_12 NS_143 0 1.6779080246226478e-02
GC_12_144 b_12 NI_12 NS_144 0 7.7216015319844815e-03
GC_12_145 b_12 NI_12 NS_145 0 9.3962459305299492e-03
GC_12_146 b_12 NI_12 NS_146 0 1.2536357178510421e-05
GC_12_147 b_12 NI_12 NS_147 0 2.5386044483703679e-13
GC_12_148 b_12 NI_12 NS_148 0 -3.4296736633209767e-07
GC_12_149 b_12 NI_12 NS_149 0 -2.1049309801311891e-05
GC_12_150 b_12 NI_12 NS_150 0 -3.9417396493263322e-06
GC_12_151 b_12 NI_12 NS_151 0 -1.8572595216007233e-03
GC_12_152 b_12 NI_12 NS_152 0 -1.1603255107540919e-02
GC_12_153 b_12 NI_12 NS_153 0 -2.7110873421980469e-02
GC_12_154 b_12 NI_12 NS_154 0 4.1598986166486883e-03
GC_12_155 b_12 NI_12 NS_155 0 1.3733926726581649e-02
GC_12_156 b_12 NI_12 NS_156 0 3.3870470678028564e-02
GC_12_157 b_12 NI_12 NS_157 0 -1.0083207369031209e-02
GC_12_158 b_12 NI_12 NS_158 0 -1.0953456611492599e-03
GC_12_159 b_12 NI_12 NS_159 0 2.5362038981058568e-02
GC_12_160 b_12 NI_12 NS_160 0 3.4553432362724748e-02
GC_12_161 b_12 NI_12 NS_161 0 1.9531231252107836e-01
GC_12_162 b_12 NI_12 NS_162 0 1.1188404770774734e-04
GC_12_163 b_12 NI_12 NS_163 0 1.5684534954802531e-12
GC_12_164 b_12 NI_12 NS_164 0 4.4028933003423356e-06
GC_12_165 b_12 NI_12 NS_165 0 1.1651552616245988e-04
GC_12_166 b_12 NI_12 NS_166 0 4.6042965410768455e-05
GC_12_167 b_12 NI_12 NS_167 0 -6.1176723006502738e-02
GC_12_168 b_12 NI_12 NS_168 0 -4.4021184493371147e-02
GC_12_169 b_12 NI_12 NS_169 0 3.9561519720181022e-02
GC_12_170 b_12 NI_12 NS_170 0 -1.8837959478211576e-02
GC_12_171 b_12 NI_12 NS_171 0 -1.2336191531711513e-01
GC_12_172 b_12 NI_12 NS_172 0 7.0718512584403148e-02
GC_12_173 b_12 NI_12 NS_173 0 -2.2400240826414768e-02
GC_12_174 b_12 NI_12 NS_174 0 1.2251147807508080e-02
GC_12_175 b_12 NI_12 NS_175 0 2.6308809871746663e-02
GC_12_176 b_12 NI_12 NS_176 0 -6.4419863054978849e-02
GC_12_177 b_12 NI_12 NS_177 0 6.0202494909286121e-02
GC_12_178 b_12 NI_12 NS_178 0 7.2267047623587099e-06
GC_12_179 b_12 NI_12 NS_179 0 -1.1474135829035945e-12
GC_12_180 b_12 NI_12 NS_180 0 -2.4578005332612988e-06
GC_12_181 b_12 NI_12 NS_181 0 2.1409342788713746e-05
GC_12_182 b_12 NI_12 NS_182 0 -3.0032933438254368e-06
GC_12_183 b_12 NI_12 NS_183 0 -1.5768202972111917e-03
GC_12_184 b_12 NI_12 NS_184 0 6.8780872594455386e-03
GC_12_185 b_12 NI_12 NS_185 0 1.7132777784430807e-02
GC_12_186 b_12 NI_12 NS_186 0 -5.5819793690011507e-03
GC_12_187 b_12 NI_12 NS_187 0 -2.5777986817383917e-02
GC_12_188 b_12 NI_12 NS_188 0 -3.1259713043061507e-02
GC_12_189 b_12 NI_12 NS_189 0 7.1574603463663332e-03
GC_12_190 b_12 NI_12 NS_190 0 2.9561886803687342e-03
GC_12_191 b_12 NI_12 NS_191 0 -3.0967504649685024e-02
GC_12_192 b_12 NI_12 NS_192 0 -3.3275366105864540e-02
GD_12_1 b_12 NI_12 NA_1 0 -3.8789040661303740e-06
GD_12_2 b_12 NI_12 NA_2 0 -2.1461866496789893e-06
GD_12_3 b_12 NI_12 NA_3 0 -9.6478587004228178e-06
GD_12_4 b_12 NI_12 NA_4 0 -2.0034324652920251e-05
GD_12_5 b_12 NI_12 NA_5 0 1.6438891897302218e-04
GD_12_6 b_12 NI_12 NA_6 0 -3.8460035209557820e-04
GD_12_7 b_12 NI_12 NA_7 0 1.5589543349922529e-03
GD_12_8 b_12 NI_12 NA_8 0 1.2309326439975655e-03
GD_12_9 b_12 NI_12 NA_9 0 -5.0305449593314542e-03
GD_12_10 b_12 NI_12 NA_10 0 4.8377577611601512e-03
GD_12_11 b_12 NI_12 NA_11 0 -1.7151991519583253e-02
GD_12_12 b_12 NI_12 NA_12 0 -3.5122897929639345e-02
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 2.5672877468519357e+00
GS_1_1 0 NS_1 NA_1 0 1.0122801651643585e+00
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 2.2430162391226233e+01
GS_2_1 0 NS_2 NA_1 0 1.0122801651643585e+00
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 2.7538444474213284e+07
GS_3_1 0 NS_3 NA_1 0 1.0122801651643585e+00
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 4.0001297681631996e+02
GS_4_1 0 NS_4 NA_1 0 1.0122801651643585e+00
*
* Real pole n. 5
CS_5 NS_5 0 9.9999999999999998e-13
RS_5 NS_5 0 5.0368733495324598e+01
GS_5_1 0 NS_5 NA_1 0 1.0122801651643585e+00
*
* Real pole n. 6
CS_6 NS_6 0 9.9999999999999998e-13
RS_6 NS_6 0 7.9588225794903536e+01
GS_6_1 0 NS_6 NA_1 0 1.0122801651643585e+00
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 1.3668579217853052e+01
RS_8 NS_8 0 1.3668579217853051e+01
GL_7 0 NS_7 NS_8 0 2.7584469331003131e-01
GL_8 0 NS_8 NS_7 0 -2.7584469331003131e-01
GS_7_1 0 NS_7 NA_1 0 1.0122801651643585e+00
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 1.2586243420126262e+01
RS_10 NS_10 0 1.2586243420126261e+01
GL_9 0 NS_9 NS_10 0 2.0570892785941347e-01
GL_10 0 NS_10 NS_9 0 -2.0570892785941347e-01
GS_9_1 0 NS_9 NA_1 0 1.0122801651643585e+00
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 1.0104148971761660e+01
RS_12 NS_12 0 1.0104148971761662e+01
GL_11 0 NS_11 NS_12 0 1.3061824103629194e-01
GL_12 0 NS_12 NS_11 0 -1.3061824103629194e-01
GS_11_1 0 NS_11 NA_1 0 1.0122801651643585e+00
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 1.4792959057818901e+01
RS_14 NS_14 0 1.4792959057818901e+01
GL_13 0 NS_13 NS_14 0 1.0109973535635272e-01
GL_14 0 NS_14 NS_13 0 -1.0109973535635272e-01
GS_13_1 0 NS_13 NA_1 0 1.0122801651643585e+00
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 1.2191222956881845e+01
RS_16 NS_16 0 1.2191222956881846e+01
GL_15 0 NS_15 NS_16 0 2.7789121104222367e-02
GL_16 0 NS_16 NS_15 0 -2.7789121104222367e-02
GS_15_1 0 NS_15 NA_1 0 1.0122801651643585e+00
*
* Real pole n. 17
CS_17 NS_17 0 9.9999999999999998e-13
RS_17 NS_17 0 2.5672877468519357e+00
GS_17_2 0 NS_17 NA_2 0 1.0122801651643585e+00
*
* Real pole n. 18
CS_18 NS_18 0 9.9999999999999998e-13
RS_18 NS_18 0 2.2430162391226233e+01
GS_18_2 0 NS_18 NA_2 0 1.0122801651643585e+00
*
* Real pole n. 19
CS_19 NS_19 0 9.9999999999999998e-13
RS_19 NS_19 0 2.7538444474213284e+07
GS_19_2 0 NS_19 NA_2 0 1.0122801651643585e+00
*
* Real pole n. 20
CS_20 NS_20 0 9.9999999999999998e-13
RS_20 NS_20 0 4.0001297681631996e+02
GS_20_2 0 NS_20 NA_2 0 1.0122801651643585e+00
*
* Real pole n. 21
CS_21 NS_21 0 9.9999999999999998e-13
RS_21 NS_21 0 5.0368733495324598e+01
GS_21_2 0 NS_21 NA_2 0 1.0122801651643585e+00
*
* Real pole n. 22
CS_22 NS_22 0 9.9999999999999998e-13
RS_22 NS_22 0 7.9588225794903536e+01
GS_22_2 0 NS_22 NA_2 0 1.0122801651643585e+00
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 1.3668579217853052e+01
RS_24 NS_24 0 1.3668579217853051e+01
GL_23 0 NS_23 NS_24 0 2.7584469331003131e-01
GL_24 0 NS_24 NS_23 0 -2.7584469331003131e-01
GS_23_2 0 NS_23 NA_2 0 1.0122801651643585e+00
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 1.2586243420126262e+01
RS_26 NS_26 0 1.2586243420126261e+01
GL_25 0 NS_25 NS_26 0 2.0570892785941347e-01
GL_26 0 NS_26 NS_25 0 -2.0570892785941347e-01
GS_25_2 0 NS_25 NA_2 0 1.0122801651643585e+00
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 1.0104148971761660e+01
RS_28 NS_28 0 1.0104148971761662e+01
GL_27 0 NS_27 NS_28 0 1.3061824103629194e-01
GL_28 0 NS_28 NS_27 0 -1.3061824103629194e-01
GS_27_2 0 NS_27 NA_2 0 1.0122801651643585e+00
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 1.4792959057818901e+01
RS_30 NS_30 0 1.4792959057818901e+01
GL_29 0 NS_29 NS_30 0 1.0109973535635272e-01
GL_30 0 NS_30 NS_29 0 -1.0109973535635272e-01
GS_29_2 0 NS_29 NA_2 0 1.0122801651643585e+00
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 1.2191222956881845e+01
RS_32 NS_32 0 1.2191222956881846e+01
GL_31 0 NS_31 NS_32 0 2.7789121104222367e-02
GL_32 0 NS_32 NS_31 0 -2.7789121104222367e-02
GS_31_2 0 NS_31 NA_2 0 1.0122801651643585e+00
*
* Real pole n. 33
CS_33 NS_33 0 9.9999999999999998e-13
RS_33 NS_33 0 2.5672877468519357e+00
GS_33_3 0 NS_33 NA_3 0 1.0122801651643585e+00
*
* Real pole n. 34
CS_34 NS_34 0 9.9999999999999998e-13
RS_34 NS_34 0 2.2430162391226233e+01
GS_34_3 0 NS_34 NA_3 0 1.0122801651643585e+00
*
* Real pole n. 35
CS_35 NS_35 0 9.9999999999999998e-13
RS_35 NS_35 0 2.7538444474213284e+07
GS_35_3 0 NS_35 NA_3 0 1.0122801651643585e+00
*
* Real pole n. 36
CS_36 NS_36 0 9.9999999999999998e-13
RS_36 NS_36 0 4.0001297681631996e+02
GS_36_3 0 NS_36 NA_3 0 1.0122801651643585e+00
*
* Real pole n. 37
CS_37 NS_37 0 9.9999999999999998e-13
RS_37 NS_37 0 5.0368733495324598e+01
GS_37_3 0 NS_37 NA_3 0 1.0122801651643585e+00
*
* Real pole n. 38
CS_38 NS_38 0 9.9999999999999998e-13
RS_38 NS_38 0 7.9588225794903536e+01
GS_38_3 0 NS_38 NA_3 0 1.0122801651643585e+00
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 1.3668579217853052e+01
RS_40 NS_40 0 1.3668579217853051e+01
GL_39 0 NS_39 NS_40 0 2.7584469331003131e-01
GL_40 0 NS_40 NS_39 0 -2.7584469331003131e-01
GS_39_3 0 NS_39 NA_3 0 1.0122801651643585e+00
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 1.2586243420126262e+01
RS_42 NS_42 0 1.2586243420126261e+01
GL_41 0 NS_41 NS_42 0 2.0570892785941347e-01
GL_42 0 NS_42 NS_41 0 -2.0570892785941347e-01
GS_41_3 0 NS_41 NA_3 0 1.0122801651643585e+00
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 1.0104148971761660e+01
RS_44 NS_44 0 1.0104148971761662e+01
GL_43 0 NS_43 NS_44 0 1.3061824103629194e-01
GL_44 0 NS_44 NS_43 0 -1.3061824103629194e-01
GS_43_3 0 NS_43 NA_3 0 1.0122801651643585e+00
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 1.4792959057818901e+01
RS_46 NS_46 0 1.4792959057818901e+01
GL_45 0 NS_45 NS_46 0 1.0109973535635272e-01
GL_46 0 NS_46 NS_45 0 -1.0109973535635272e-01
GS_45_3 0 NS_45 NA_3 0 1.0122801651643585e+00
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 1.2191222956881845e+01
RS_48 NS_48 0 1.2191222956881846e+01
GL_47 0 NS_47 NS_48 0 2.7789121104222367e-02
GL_48 0 NS_48 NS_47 0 -2.7789121104222367e-02
GS_47_3 0 NS_47 NA_3 0 1.0122801651643585e+00
*
* Real pole n. 49
CS_49 NS_49 0 9.9999999999999998e-13
RS_49 NS_49 0 2.5672877468519357e+00
GS_49_4 0 NS_49 NA_4 0 1.0122801651643585e+00
*
* Real pole n. 50
CS_50 NS_50 0 9.9999999999999998e-13
RS_50 NS_50 0 2.2430162391226233e+01
GS_50_4 0 NS_50 NA_4 0 1.0122801651643585e+00
*
* Real pole n. 51
CS_51 NS_51 0 9.9999999999999998e-13
RS_51 NS_51 0 2.7538444474213284e+07
GS_51_4 0 NS_51 NA_4 0 1.0122801651643585e+00
*
* Real pole n. 52
CS_52 NS_52 0 9.9999999999999998e-13
RS_52 NS_52 0 4.0001297681631996e+02
GS_52_4 0 NS_52 NA_4 0 1.0122801651643585e+00
*
* Real pole n. 53
CS_53 NS_53 0 9.9999999999999998e-13
RS_53 NS_53 0 5.0368733495324598e+01
GS_53_4 0 NS_53 NA_4 0 1.0122801651643585e+00
*
* Real pole n. 54
CS_54 NS_54 0 9.9999999999999998e-13
RS_54 NS_54 0 7.9588225794903536e+01
GS_54_4 0 NS_54 NA_4 0 1.0122801651643585e+00
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 1.3668579217853052e+01
RS_56 NS_56 0 1.3668579217853051e+01
GL_55 0 NS_55 NS_56 0 2.7584469331003131e-01
GL_56 0 NS_56 NS_55 0 -2.7584469331003131e-01
GS_55_4 0 NS_55 NA_4 0 1.0122801651643585e+00
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 1.2586243420126262e+01
RS_58 NS_58 0 1.2586243420126261e+01
GL_57 0 NS_57 NS_58 0 2.0570892785941347e-01
GL_58 0 NS_58 NS_57 0 -2.0570892785941347e-01
GS_57_4 0 NS_57 NA_4 0 1.0122801651643585e+00
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 1.0104148971761660e+01
RS_60 NS_60 0 1.0104148971761662e+01
GL_59 0 NS_59 NS_60 0 1.3061824103629194e-01
GL_60 0 NS_60 NS_59 0 -1.3061824103629194e-01
GS_59_4 0 NS_59 NA_4 0 1.0122801651643585e+00
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 1.4792959057818901e+01
RS_62 NS_62 0 1.4792959057818901e+01
GL_61 0 NS_61 NS_62 0 1.0109973535635272e-01
GL_62 0 NS_62 NS_61 0 -1.0109973535635272e-01
GS_61_4 0 NS_61 NA_4 0 1.0122801651643585e+00
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 1.2191222956881845e+01
RS_64 NS_64 0 1.2191222956881846e+01
GL_63 0 NS_63 NS_64 0 2.7789121104222367e-02
GL_64 0 NS_64 NS_63 0 -2.7789121104222367e-02
GS_63_4 0 NS_63 NA_4 0 1.0122801651643585e+00
*
* Real pole n. 65
CS_65 NS_65 0 9.9999999999999998e-13
RS_65 NS_65 0 2.5672877468519357e+00
GS_65_5 0 NS_65 NA_5 0 1.0122801651643585e+00
*
* Real pole n. 66
CS_66 NS_66 0 9.9999999999999998e-13
RS_66 NS_66 0 2.2430162391226233e+01
GS_66_5 0 NS_66 NA_5 0 1.0122801651643585e+00
*
* Real pole n. 67
CS_67 NS_67 0 9.9999999999999998e-13
RS_67 NS_67 0 2.7538444474213284e+07
GS_67_5 0 NS_67 NA_5 0 1.0122801651643585e+00
*
* Real pole n. 68
CS_68 NS_68 0 9.9999999999999998e-13
RS_68 NS_68 0 4.0001297681631996e+02
GS_68_5 0 NS_68 NA_5 0 1.0122801651643585e+00
*
* Real pole n. 69
CS_69 NS_69 0 9.9999999999999998e-13
RS_69 NS_69 0 5.0368733495324598e+01
GS_69_5 0 NS_69 NA_5 0 1.0122801651643585e+00
*
* Real pole n. 70
CS_70 NS_70 0 9.9999999999999998e-13
RS_70 NS_70 0 7.9588225794903536e+01
GS_70_5 0 NS_70 NA_5 0 1.0122801651643585e+00
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 1.3668579217853052e+01
RS_72 NS_72 0 1.3668579217853051e+01
GL_71 0 NS_71 NS_72 0 2.7584469331003131e-01
GL_72 0 NS_72 NS_71 0 -2.7584469331003131e-01
GS_71_5 0 NS_71 NA_5 0 1.0122801651643585e+00
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 1.2586243420126262e+01
RS_74 NS_74 0 1.2586243420126261e+01
GL_73 0 NS_73 NS_74 0 2.0570892785941347e-01
GL_74 0 NS_74 NS_73 0 -2.0570892785941347e-01
GS_73_5 0 NS_73 NA_5 0 1.0122801651643585e+00
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 1.0104148971761660e+01
RS_76 NS_76 0 1.0104148971761662e+01
GL_75 0 NS_75 NS_76 0 1.3061824103629194e-01
GL_76 0 NS_76 NS_75 0 -1.3061824103629194e-01
GS_75_5 0 NS_75 NA_5 0 1.0122801651643585e+00
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 1.4792959057818901e+01
RS_78 NS_78 0 1.4792959057818901e+01
GL_77 0 NS_77 NS_78 0 1.0109973535635272e-01
GL_78 0 NS_78 NS_77 0 -1.0109973535635272e-01
GS_77_5 0 NS_77 NA_5 0 1.0122801651643585e+00
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 1.2191222956881845e+01
RS_80 NS_80 0 1.2191222956881846e+01
GL_79 0 NS_79 NS_80 0 2.7789121104222367e-02
GL_80 0 NS_80 NS_79 0 -2.7789121104222367e-02
GS_79_5 0 NS_79 NA_5 0 1.0122801651643585e+00
*
* Real pole n. 81
CS_81 NS_81 0 9.9999999999999998e-13
RS_81 NS_81 0 2.5672877468519357e+00
GS_81_6 0 NS_81 NA_6 0 1.0122801651643585e+00
*
* Real pole n. 82
CS_82 NS_82 0 9.9999999999999998e-13
RS_82 NS_82 0 2.2430162391226233e+01
GS_82_6 0 NS_82 NA_6 0 1.0122801651643585e+00
*
* Real pole n. 83
CS_83 NS_83 0 9.9999999999999998e-13
RS_83 NS_83 0 2.7538444474213284e+07
GS_83_6 0 NS_83 NA_6 0 1.0122801651643585e+00
*
* Real pole n. 84
CS_84 NS_84 0 9.9999999999999998e-13
RS_84 NS_84 0 4.0001297681631996e+02
GS_84_6 0 NS_84 NA_6 0 1.0122801651643585e+00
*
* Real pole n. 85
CS_85 NS_85 0 9.9999999999999998e-13
RS_85 NS_85 0 5.0368733495324598e+01
GS_85_6 0 NS_85 NA_6 0 1.0122801651643585e+00
*
* Real pole n. 86
CS_86 NS_86 0 9.9999999999999998e-13
RS_86 NS_86 0 7.9588225794903536e+01
GS_86_6 0 NS_86 NA_6 0 1.0122801651643585e+00
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 1.3668579217853052e+01
RS_88 NS_88 0 1.3668579217853051e+01
GL_87 0 NS_87 NS_88 0 2.7584469331003131e-01
GL_88 0 NS_88 NS_87 0 -2.7584469331003131e-01
GS_87_6 0 NS_87 NA_6 0 1.0122801651643585e+00
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 1.2586243420126262e+01
RS_90 NS_90 0 1.2586243420126261e+01
GL_89 0 NS_89 NS_90 0 2.0570892785941347e-01
GL_90 0 NS_90 NS_89 0 -2.0570892785941347e-01
GS_89_6 0 NS_89 NA_6 0 1.0122801651643585e+00
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 1.0104148971761660e+01
RS_92 NS_92 0 1.0104148971761662e+01
GL_91 0 NS_91 NS_92 0 1.3061824103629194e-01
GL_92 0 NS_92 NS_91 0 -1.3061824103629194e-01
GS_91_6 0 NS_91 NA_6 0 1.0122801651643585e+00
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 1.4792959057818901e+01
RS_94 NS_94 0 1.4792959057818901e+01
GL_93 0 NS_93 NS_94 0 1.0109973535635272e-01
GL_94 0 NS_94 NS_93 0 -1.0109973535635272e-01
GS_93_6 0 NS_93 NA_6 0 1.0122801651643585e+00
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 1.2191222956881845e+01
RS_96 NS_96 0 1.2191222956881846e+01
GL_95 0 NS_95 NS_96 0 2.7789121104222367e-02
GL_96 0 NS_96 NS_95 0 -2.7789121104222367e-02
GS_95_6 0 NS_95 NA_6 0 1.0122801651643585e+00
*
* Real pole n. 97
CS_97 NS_97 0 9.9999999999999998e-13
RS_97 NS_97 0 2.5672877468519357e+00
GS_97_7 0 NS_97 NA_7 0 1.0122801651643585e+00
*
* Real pole n. 98
CS_98 NS_98 0 9.9999999999999998e-13
RS_98 NS_98 0 2.2430162391226233e+01
GS_98_7 0 NS_98 NA_7 0 1.0122801651643585e+00
*
* Real pole n. 99
CS_99 NS_99 0 9.9999999999999998e-13
RS_99 NS_99 0 2.7538444474213284e+07
GS_99_7 0 NS_99 NA_7 0 1.0122801651643585e+00
*
* Real pole n. 100
CS_100 NS_100 0 9.9999999999999998e-13
RS_100 NS_100 0 4.0001297681631996e+02
GS_100_7 0 NS_100 NA_7 0 1.0122801651643585e+00
*
* Real pole n. 101
CS_101 NS_101 0 9.9999999999999998e-13
RS_101 NS_101 0 5.0368733495324598e+01
GS_101_7 0 NS_101 NA_7 0 1.0122801651643585e+00
*
* Real pole n. 102
CS_102 NS_102 0 9.9999999999999998e-13
RS_102 NS_102 0 7.9588225794903536e+01
GS_102_7 0 NS_102 NA_7 0 1.0122801651643585e+00
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 1.3668579217853052e+01
RS_104 NS_104 0 1.3668579217853051e+01
GL_103 0 NS_103 NS_104 0 2.7584469331003131e-01
GL_104 0 NS_104 NS_103 0 -2.7584469331003131e-01
GS_103_7 0 NS_103 NA_7 0 1.0122801651643585e+00
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 1.2586243420126262e+01
RS_106 NS_106 0 1.2586243420126261e+01
GL_105 0 NS_105 NS_106 0 2.0570892785941347e-01
GL_106 0 NS_106 NS_105 0 -2.0570892785941347e-01
GS_105_7 0 NS_105 NA_7 0 1.0122801651643585e+00
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 1.0104148971761660e+01
RS_108 NS_108 0 1.0104148971761662e+01
GL_107 0 NS_107 NS_108 0 1.3061824103629194e-01
GL_108 0 NS_108 NS_107 0 -1.3061824103629194e-01
GS_107_7 0 NS_107 NA_7 0 1.0122801651643585e+00
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 1.4792959057818901e+01
RS_110 NS_110 0 1.4792959057818901e+01
GL_109 0 NS_109 NS_110 0 1.0109973535635272e-01
GL_110 0 NS_110 NS_109 0 -1.0109973535635272e-01
GS_109_7 0 NS_109 NA_7 0 1.0122801651643585e+00
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 1.2191222956881845e+01
RS_112 NS_112 0 1.2191222956881846e+01
GL_111 0 NS_111 NS_112 0 2.7789121104222367e-02
GL_112 0 NS_112 NS_111 0 -2.7789121104222367e-02
GS_111_7 0 NS_111 NA_7 0 1.0122801651643585e+00
*
* Real pole n. 113
CS_113 NS_113 0 9.9999999999999998e-13
RS_113 NS_113 0 2.5672877468519357e+00
GS_113_8 0 NS_113 NA_8 0 1.0122801651643585e+00
*
* Real pole n. 114
CS_114 NS_114 0 9.9999999999999998e-13
RS_114 NS_114 0 2.2430162391226233e+01
GS_114_8 0 NS_114 NA_8 0 1.0122801651643585e+00
*
* Real pole n. 115
CS_115 NS_115 0 9.9999999999999998e-13
RS_115 NS_115 0 2.7538444474213284e+07
GS_115_8 0 NS_115 NA_8 0 1.0122801651643585e+00
*
* Real pole n. 116
CS_116 NS_116 0 9.9999999999999998e-13
RS_116 NS_116 0 4.0001297681631996e+02
GS_116_8 0 NS_116 NA_8 0 1.0122801651643585e+00
*
* Real pole n. 117
CS_117 NS_117 0 9.9999999999999998e-13
RS_117 NS_117 0 5.0368733495324598e+01
GS_117_8 0 NS_117 NA_8 0 1.0122801651643585e+00
*
* Real pole n. 118
CS_118 NS_118 0 9.9999999999999998e-13
RS_118 NS_118 0 7.9588225794903536e+01
GS_118_8 0 NS_118 NA_8 0 1.0122801651643585e+00
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 1.3668579217853052e+01
RS_120 NS_120 0 1.3668579217853051e+01
GL_119 0 NS_119 NS_120 0 2.7584469331003131e-01
GL_120 0 NS_120 NS_119 0 -2.7584469331003131e-01
GS_119_8 0 NS_119 NA_8 0 1.0122801651643585e+00
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 1.2586243420126262e+01
RS_122 NS_122 0 1.2586243420126261e+01
GL_121 0 NS_121 NS_122 0 2.0570892785941347e-01
GL_122 0 NS_122 NS_121 0 -2.0570892785941347e-01
GS_121_8 0 NS_121 NA_8 0 1.0122801651643585e+00
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 1.0104148971761660e+01
RS_124 NS_124 0 1.0104148971761662e+01
GL_123 0 NS_123 NS_124 0 1.3061824103629194e-01
GL_124 0 NS_124 NS_123 0 -1.3061824103629194e-01
GS_123_8 0 NS_123 NA_8 0 1.0122801651643585e+00
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 1.4792959057818901e+01
RS_126 NS_126 0 1.4792959057818901e+01
GL_125 0 NS_125 NS_126 0 1.0109973535635272e-01
GL_126 0 NS_126 NS_125 0 -1.0109973535635272e-01
GS_125_8 0 NS_125 NA_8 0 1.0122801651643585e+00
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 1.2191222956881845e+01
RS_128 NS_128 0 1.2191222956881846e+01
GL_127 0 NS_127 NS_128 0 2.7789121104222367e-02
GL_128 0 NS_128 NS_127 0 -2.7789121104222367e-02
GS_127_8 0 NS_127 NA_8 0 1.0122801651643585e+00
*
* Real pole n. 129
CS_129 NS_129 0 9.9999999999999998e-13
RS_129 NS_129 0 2.5672877468519357e+00
GS_129_9 0 NS_129 NA_9 0 1.0122801651643585e+00
*
* Real pole n. 130
CS_130 NS_130 0 9.9999999999999998e-13
RS_130 NS_130 0 2.2430162391226233e+01
GS_130_9 0 NS_130 NA_9 0 1.0122801651643585e+00
*
* Real pole n. 131
CS_131 NS_131 0 9.9999999999999998e-13
RS_131 NS_131 0 2.7538444474213284e+07
GS_131_9 0 NS_131 NA_9 0 1.0122801651643585e+00
*
* Real pole n. 132
CS_132 NS_132 0 9.9999999999999998e-13
RS_132 NS_132 0 4.0001297681631996e+02
GS_132_9 0 NS_132 NA_9 0 1.0122801651643585e+00
*
* Real pole n. 133
CS_133 NS_133 0 9.9999999999999998e-13
RS_133 NS_133 0 5.0368733495324598e+01
GS_133_9 0 NS_133 NA_9 0 1.0122801651643585e+00
*
* Real pole n. 134
CS_134 NS_134 0 9.9999999999999998e-13
RS_134 NS_134 0 7.9588225794903536e+01
GS_134_9 0 NS_134 NA_9 0 1.0122801651643585e+00
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 1.3668579217853052e+01
RS_136 NS_136 0 1.3668579217853051e+01
GL_135 0 NS_135 NS_136 0 2.7584469331003131e-01
GL_136 0 NS_136 NS_135 0 -2.7584469331003131e-01
GS_135_9 0 NS_135 NA_9 0 1.0122801651643585e+00
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 1.2586243420126262e+01
RS_138 NS_138 0 1.2586243420126261e+01
GL_137 0 NS_137 NS_138 0 2.0570892785941347e-01
GL_138 0 NS_138 NS_137 0 -2.0570892785941347e-01
GS_137_9 0 NS_137 NA_9 0 1.0122801651643585e+00
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 1.0104148971761660e+01
RS_140 NS_140 0 1.0104148971761662e+01
GL_139 0 NS_139 NS_140 0 1.3061824103629194e-01
GL_140 0 NS_140 NS_139 0 -1.3061824103629194e-01
GS_139_9 0 NS_139 NA_9 0 1.0122801651643585e+00
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 1.4792959057818901e+01
RS_142 NS_142 0 1.4792959057818901e+01
GL_141 0 NS_141 NS_142 0 1.0109973535635272e-01
GL_142 0 NS_142 NS_141 0 -1.0109973535635272e-01
GS_141_9 0 NS_141 NA_9 0 1.0122801651643585e+00
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 1.2191222956881845e+01
RS_144 NS_144 0 1.2191222956881846e+01
GL_143 0 NS_143 NS_144 0 2.7789121104222367e-02
GL_144 0 NS_144 NS_143 0 -2.7789121104222367e-02
GS_143_9 0 NS_143 NA_9 0 1.0122801651643585e+00
*
* Real pole n. 145
CS_145 NS_145 0 9.9999999999999998e-13
RS_145 NS_145 0 2.5672877468519357e+00
GS_145_10 0 NS_145 NA_10 0 1.0122801651643585e+00
*
* Real pole n. 146
CS_146 NS_146 0 9.9999999999999998e-13
RS_146 NS_146 0 2.2430162391226233e+01
GS_146_10 0 NS_146 NA_10 0 1.0122801651643585e+00
*
* Real pole n. 147
CS_147 NS_147 0 9.9999999999999998e-13
RS_147 NS_147 0 2.7538444474213284e+07
GS_147_10 0 NS_147 NA_10 0 1.0122801651643585e+00
*
* Real pole n. 148
CS_148 NS_148 0 9.9999999999999998e-13
RS_148 NS_148 0 4.0001297681631996e+02
GS_148_10 0 NS_148 NA_10 0 1.0122801651643585e+00
*
* Real pole n. 149
CS_149 NS_149 0 9.9999999999999998e-13
RS_149 NS_149 0 5.0368733495324598e+01
GS_149_10 0 NS_149 NA_10 0 1.0122801651643585e+00
*
* Real pole n. 150
CS_150 NS_150 0 9.9999999999999998e-13
RS_150 NS_150 0 7.9588225794903536e+01
GS_150_10 0 NS_150 NA_10 0 1.0122801651643585e+00
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 1.3668579217853052e+01
RS_152 NS_152 0 1.3668579217853051e+01
GL_151 0 NS_151 NS_152 0 2.7584469331003131e-01
GL_152 0 NS_152 NS_151 0 -2.7584469331003131e-01
GS_151_10 0 NS_151 NA_10 0 1.0122801651643585e+00
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 1.2586243420126262e+01
RS_154 NS_154 0 1.2586243420126261e+01
GL_153 0 NS_153 NS_154 0 2.0570892785941347e-01
GL_154 0 NS_154 NS_153 0 -2.0570892785941347e-01
GS_153_10 0 NS_153 NA_10 0 1.0122801651643585e+00
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 1.0104148971761660e+01
RS_156 NS_156 0 1.0104148971761662e+01
GL_155 0 NS_155 NS_156 0 1.3061824103629194e-01
GL_156 0 NS_156 NS_155 0 -1.3061824103629194e-01
GS_155_10 0 NS_155 NA_10 0 1.0122801651643585e+00
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 1.4792959057818901e+01
RS_158 NS_158 0 1.4792959057818901e+01
GL_157 0 NS_157 NS_158 0 1.0109973535635272e-01
GL_158 0 NS_158 NS_157 0 -1.0109973535635272e-01
GS_157_10 0 NS_157 NA_10 0 1.0122801651643585e+00
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 1.2191222956881845e+01
RS_160 NS_160 0 1.2191222956881846e+01
GL_159 0 NS_159 NS_160 0 2.7789121104222367e-02
GL_160 0 NS_160 NS_159 0 -2.7789121104222367e-02
GS_159_10 0 NS_159 NA_10 0 1.0122801651643585e+00
*
* Real pole n. 161
CS_161 NS_161 0 9.9999999999999998e-13
RS_161 NS_161 0 2.5672877468519357e+00
GS_161_11 0 NS_161 NA_11 0 1.0122801651643585e+00
*
* Real pole n. 162
CS_162 NS_162 0 9.9999999999999998e-13
RS_162 NS_162 0 2.2430162391226233e+01
GS_162_11 0 NS_162 NA_11 0 1.0122801651643585e+00
*
* Real pole n. 163
CS_163 NS_163 0 9.9999999999999998e-13
RS_163 NS_163 0 2.7538444474213284e+07
GS_163_11 0 NS_163 NA_11 0 1.0122801651643585e+00
*
* Real pole n. 164
CS_164 NS_164 0 9.9999999999999998e-13
RS_164 NS_164 0 4.0001297681631996e+02
GS_164_11 0 NS_164 NA_11 0 1.0122801651643585e+00
*
* Real pole n. 165
CS_165 NS_165 0 9.9999999999999998e-13
RS_165 NS_165 0 5.0368733495324598e+01
GS_165_11 0 NS_165 NA_11 0 1.0122801651643585e+00
*
* Real pole n. 166
CS_166 NS_166 0 9.9999999999999998e-13
RS_166 NS_166 0 7.9588225794903536e+01
GS_166_11 0 NS_166 NA_11 0 1.0122801651643585e+00
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 1.3668579217853052e+01
RS_168 NS_168 0 1.3668579217853051e+01
GL_167 0 NS_167 NS_168 0 2.7584469331003131e-01
GL_168 0 NS_168 NS_167 0 -2.7584469331003131e-01
GS_167_11 0 NS_167 NA_11 0 1.0122801651643585e+00
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 1.2586243420126262e+01
RS_170 NS_170 0 1.2586243420126261e+01
GL_169 0 NS_169 NS_170 0 2.0570892785941347e-01
GL_170 0 NS_170 NS_169 0 -2.0570892785941347e-01
GS_169_11 0 NS_169 NA_11 0 1.0122801651643585e+00
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 1.0104148971761660e+01
RS_172 NS_172 0 1.0104148971761662e+01
GL_171 0 NS_171 NS_172 0 1.3061824103629194e-01
GL_172 0 NS_172 NS_171 0 -1.3061824103629194e-01
GS_171_11 0 NS_171 NA_11 0 1.0122801651643585e+00
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 1.4792959057818901e+01
RS_174 NS_174 0 1.4792959057818901e+01
GL_173 0 NS_173 NS_174 0 1.0109973535635272e-01
GL_174 0 NS_174 NS_173 0 -1.0109973535635272e-01
GS_173_11 0 NS_173 NA_11 0 1.0122801651643585e+00
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 1.2191222956881845e+01
RS_176 NS_176 0 1.2191222956881846e+01
GL_175 0 NS_175 NS_176 0 2.7789121104222367e-02
GL_176 0 NS_176 NS_175 0 -2.7789121104222367e-02
GS_175_11 0 NS_175 NA_11 0 1.0122801651643585e+00
*
* Real pole n. 177
CS_177 NS_177 0 9.9999999999999998e-13
RS_177 NS_177 0 2.5672877468519357e+00
GS_177_12 0 NS_177 NA_12 0 1.0122801651643585e+00
*
* Real pole n. 178
CS_178 NS_178 0 9.9999999999999998e-13
RS_178 NS_178 0 2.2430162391226233e+01
GS_178_12 0 NS_178 NA_12 0 1.0122801651643585e+00
*
* Real pole n. 179
CS_179 NS_179 0 9.9999999999999998e-13
RS_179 NS_179 0 2.7538444474213284e+07
GS_179_12 0 NS_179 NA_12 0 1.0122801651643585e+00
*
* Real pole n. 180
CS_180 NS_180 0 9.9999999999999998e-13
RS_180 NS_180 0 4.0001297681631996e+02
GS_180_12 0 NS_180 NA_12 0 1.0122801651643585e+00
*
* Real pole n. 181
CS_181 NS_181 0 9.9999999999999998e-13
RS_181 NS_181 0 5.0368733495324598e+01
GS_181_12 0 NS_181 NA_12 0 1.0122801651643585e+00
*
* Real pole n. 182
CS_182 NS_182 0 9.9999999999999998e-13
RS_182 NS_182 0 7.9588225794903536e+01
GS_182_12 0 NS_182 NA_12 0 1.0122801651643585e+00
*
* Complex pair n. 183/184
CS_183 NS_183 0 9.9999999999999998e-13
CS_184 NS_184 0 9.9999999999999998e-13
RS_183 NS_183 0 1.3668579217853052e+01
RS_184 NS_184 0 1.3668579217853051e+01
GL_183 0 NS_183 NS_184 0 2.7584469331003131e-01
GL_184 0 NS_184 NS_183 0 -2.7584469331003131e-01
GS_183_12 0 NS_183 NA_12 0 1.0122801651643585e+00
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 1.2586243420126262e+01
RS_186 NS_186 0 1.2586243420126261e+01
GL_185 0 NS_185 NS_186 0 2.0570892785941347e-01
GL_186 0 NS_186 NS_185 0 -2.0570892785941347e-01
GS_185_12 0 NS_185 NA_12 0 1.0122801651643585e+00
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 1.0104148971761660e+01
RS_188 NS_188 0 1.0104148971761662e+01
GL_187 0 NS_187 NS_188 0 1.3061824103629194e-01
GL_188 0 NS_188 NS_187 0 -1.3061824103629194e-01
GS_187_12 0 NS_187 NA_12 0 1.0122801651643585e+00
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 1.4792959057818901e+01
RS_190 NS_190 0 1.4792959057818901e+01
GL_189 0 NS_189 NS_190 0 1.0109973535635272e-01
GL_190 0 NS_190 NS_189 0 -1.0109973535635272e-01
GS_189_12 0 NS_189 NA_12 0 1.0122801651643585e+00
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 1.2191222956881845e+01
RS_192 NS_192 0 1.2191222956881846e+01
GL_191 0 NS_191 NS_192 0 2.7789121104222367e-02
GL_192 0 NS_192 NS_191 0 -2.7789121104222367e-02
GS_191_12 0 NS_191 NA_12 0 1.0122801651643585e+00
*
******************************


.ends
*******************
* End of subcircuit
*******************
