**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [6 4 28] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** n/a - passivity was not enforced
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_12_PCB_wire_0p25inch_highloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 -1.0222189382686536e-03
GC_1_2 b_1 NI_1 NS_2 0 -1.7322668026375918e-02
GC_1_3 b_1 NI_1 NS_3 0 1.1757822387305574e-02
GC_1_4 b_1 NI_1 NS_4 0 2.8947520427771859e-06
GC_1_5 b_1 NI_1 NS_5 0 -5.0926480052766377e-07
GC_1_6 b_1 NI_1 NS_6 0 -2.9660693246163502e-08
GC_1_7 b_1 NI_1 NS_7 0 3.0704128506545028e-03
GC_1_8 b_1 NI_1 NS_8 0 1.2919121928318890e-03
GC_1_9 b_1 NI_1 NS_9 0 -2.9518618707215006e-03
GC_1_10 b_1 NI_1 NS_10 0 -9.9170148249821972e-03
GC_1_11 b_1 NI_1 NS_11 0 5.8893975062115043e-04
GC_1_12 b_1 NI_1 NS_12 0 1.3640194001803980e-02
GC_1_13 b_1 NI_1 NS_13 0 1.7423650650642906e-02
GC_1_14 b_1 NI_1 NS_14 0 -2.3868296008015436e-02
GC_1_15 b_1 NI_1 NS_15 0 -3.3167484266264612e-02
GC_1_16 b_1 NI_1 NS_16 0 2.1401807985247351e-02
GC_1_17 b_1 NI_1 NS_17 0 4.0587922746253592e-03
GC_1_18 b_1 NI_1 NS_18 0 -2.2320128311773386e-03
GC_1_19 b_1 NI_1 NS_19 0 1.5116274598290057e-02
GC_1_20 b_1 NI_1 NS_20 0 5.6072380779884686e-03
GC_1_21 b_1 NI_1 NS_21 0 -2.8699862317699099e-01
GC_1_22 b_1 NI_1 NS_22 0 1.2135733771095281e-01
GC_1_23 b_1 NI_1 NS_23 0 7.0298545669318551e-03
GC_1_24 b_1 NI_1 NS_24 0 5.7777308956970074e-05
GC_1_25 b_1 NI_1 NS_25 0 1.2954678181379544e-06
GC_1_26 b_1 NI_1 NS_26 0 1.4196126589821395e-08
GC_1_27 b_1 NI_1 NS_27 0 3.0514922267685724e-02
GC_1_28 b_1 NI_1 NS_28 0 4.1652932579782607e-03
GC_1_29 b_1 NI_1 NS_29 0 -7.3042421194979314e-03
GC_1_30 b_1 NI_1 NS_30 0 2.2210834258712158e-02
GC_1_31 b_1 NI_1 NS_31 0 -1.6943497309199432e-02
GC_1_32 b_1 NI_1 NS_32 0 -1.8718581187072925e-02
GC_1_33 b_1 NI_1 NS_33 0 4.4820939568194884e-02
GC_1_34 b_1 NI_1 NS_34 0 1.4501642688124481e-02
GC_1_35 b_1 NI_1 NS_35 0 8.2245808728605471e-02
GC_1_36 b_1 NI_1 NS_36 0 3.0932524324755656e-02
GC_1_37 b_1 NI_1 NS_37 0 -1.0134600388785650e-02
GC_1_38 b_1 NI_1 NS_38 0 -4.8138172557028232e-03
GC_1_39 b_1 NI_1 NS_39 0 -2.1451566364332434e-02
GC_1_40 b_1 NI_1 NS_40 0 -4.8857374149900096e-03
GC_1_41 b_1 NI_1 NS_41 0 2.2274176795434541e-02
GC_1_42 b_1 NI_1 NS_42 0 8.9558630542299258e-03
GC_1_43 b_1 NI_1 NS_43 0 -1.1409760099151504e-02
GC_1_44 b_1 NI_1 NS_44 0 -5.3360833874138167e-06
GC_1_45 b_1 NI_1 NS_45 0 -9.5822579627153655e-08
GC_1_46 b_1 NI_1 NS_46 0 -1.2412250849481511e-09
GC_1_47 b_1 NI_1 NS_47 0 -3.3143877241228791e-03
GC_1_48 b_1 NI_1 NS_48 0 -2.3911427672548280e-03
GC_1_49 b_1 NI_1 NS_49 0 2.7261769899454592e-03
GC_1_50 b_1 NI_1 NS_50 0 1.1171778125940076e-02
GC_1_51 b_1 NI_1 NS_51 0 -3.5307706731909776e-04
GC_1_52 b_1 NI_1 NS_52 0 -1.7759590133167649e-02
GC_1_53 b_1 NI_1 NS_53 0 -2.2020926264061297e-02
GC_1_54 b_1 NI_1 NS_54 0 2.1326546211935585e-02
GC_1_55 b_1 NI_1 NS_55 0 2.8908349472181977e-02
GC_1_56 b_1 NI_1 NS_56 0 -1.8397053919704077e-02
GC_1_57 b_1 NI_1 NS_57 0 -2.4507569379336796e-03
GC_1_58 b_1 NI_1 NS_58 0 1.4218494192317892e-03
GC_1_59 b_1 NI_1 NS_59 0 -1.7818879771854996e-02
GC_1_60 b_1 NI_1 NS_60 0 -7.1265648084851618e-03
GC_1_61 b_1 NI_1 NS_61 0 -8.2288461374579264e-02
GC_1_62 b_1 NI_1 NS_62 0 6.5322021849922376e-02
GC_1_63 b_1 NI_1 NS_63 0 -1.0307113987320324e-02
GC_1_64 b_1 NI_1 NS_64 0 -2.3858543740764415e-06
GC_1_65 b_1 NI_1 NS_65 0 1.6335231281682485e-08
GC_1_66 b_1 NI_1 NS_66 0 1.6410073241915433e-09
GC_1_67 b_1 NI_1 NS_67 0 -3.9597044083589306e-04
GC_1_68 b_1 NI_1 NS_68 0 -1.4000567030019084e-03
GC_1_69 b_1 NI_1 NS_69 0 -6.9917491209412919e-03
GC_1_70 b_1 NI_1 NS_70 0 -3.7822426985025200e-03
GC_1_71 b_1 NI_1 NS_71 0 -9.0594503188277595e-03
GC_1_72 b_1 NI_1 NS_72 0 1.3121192278131088e-02
GC_1_73 b_1 NI_1 NS_73 0 -1.5240954434080477e-02
GC_1_74 b_1 NI_1 NS_74 0 2.8718756402281151e-02
GC_1_75 b_1 NI_1 NS_75 0 4.5110991427149472e-02
GC_1_76 b_1 NI_1 NS_76 0 1.6488627627910361e-02
GC_1_77 b_1 NI_1 NS_77 0 -2.2090755317901853e-03
GC_1_78 b_1 NI_1 NS_78 0 -1.3391797800839161e-03
GC_1_79 b_1 NI_1 NS_79 0 1.2863710674879012e-02
GC_1_80 b_1 NI_1 NS_80 0 6.9572426669046996e-03
GC_1_81 b_1 NI_1 NS_81 0 2.7174115821772000e-04
GC_1_82 b_1 NI_1 NS_82 0 -1.1194127112613104e-05
GC_1_83 b_1 NI_1 NS_83 0 -9.5765069074447400e-06
GC_1_84 b_1 NI_1 NS_84 0 6.1170048036647436e-08
GC_1_85 b_1 NI_1 NS_85 0 -3.1755797022978616e-10
GC_1_86 b_1 NI_1 NS_86 0 9.0305714976593636e-12
GC_1_87 b_1 NI_1 NS_87 0 -4.6037800608859903e-07
GC_1_88 b_1 NI_1 NS_88 0 -1.5384218975440852e-05
GC_1_89 b_1 NI_1 NS_89 0 -9.5047719624023158e-06
GC_1_90 b_1 NI_1 NS_90 0 -2.0753489822213513e-05
GC_1_91 b_1 NI_1 NS_91 0 -3.7497052545528499e-05
GC_1_92 b_1 NI_1 NS_92 0 -1.9825266004699476e-05
GC_1_93 b_1 NI_1 NS_93 0 -7.4897115463339327e-05
GC_1_94 b_1 NI_1 NS_94 0 -7.8245278481738734e-05
GC_1_95 b_1 NI_1 NS_95 0 -7.3342906412342430e-05
GC_1_96 b_1 NI_1 NS_96 0 2.1906424126283996e-04
GC_1_97 b_1 NI_1 NS_97 0 1.4840686609615702e-05
GC_1_98 b_1 NI_1 NS_98 0 -5.7290357263067270e-05
GC_1_99 b_1 NI_1 NS_99 0 -4.6091055545733033e-06
GC_1_100 b_1 NI_1 NS_100 0 1.3659348391919208e-05
GC_1_101 b_1 NI_1 NS_101 0 3.0050323718818617e-04
GC_1_102 b_1 NI_1 NS_102 0 -2.6759729181300047e-04
GC_1_103 b_1 NI_1 NS_103 0 4.2937842849253362e-05
GC_1_104 b_1 NI_1 NS_104 0 1.3911739318512860e-08
GC_1_105 b_1 NI_1 NS_105 0 -1.4978353405891414e-10
GC_1_106 b_1 NI_1 NS_106 0 1.4933238226627101e-11
GC_1_107 b_1 NI_1 NS_107 0 2.1659411432353123e-06
GC_1_108 b_1 NI_1 NS_108 0 7.3080135507372240e-06
GC_1_109 b_1 NI_1 NS_109 0 3.3345692068580734e-05
GC_1_110 b_1 NI_1 NS_110 0 2.1778354057868978e-05
GC_1_111 b_1 NI_1 NS_111 0 4.6482455849148190e-05
GC_1_112 b_1 NI_1 NS_112 0 -5.6793318374757557e-05
GC_1_113 b_1 NI_1 NS_113 0 7.4769075185396295e-05
GC_1_114 b_1 NI_1 NS_114 0 -1.2484402667173656e-04
GC_1_115 b_1 NI_1 NS_115 0 -1.8751986130427462e-04
GC_1_116 b_1 NI_1 NS_116 0 -7.7199056108160168e-05
GC_1_117 b_1 NI_1 NS_117 0 8.1439071000455390e-06
GC_1_118 b_1 NI_1 NS_118 0 4.1237466923363233e-06
GC_1_119 b_1 NI_1 NS_119 0 -5.4121468631203835e-05
GC_1_120 b_1 NI_1 NS_120 0 -3.1122573958567608e-05
GC_1_121 b_1 NI_1 NS_121 0 -8.6861198400690117e-05
GC_1_122 b_1 NI_1 NS_122 0 1.4645967683878723e-05
GC_1_123 b_1 NI_1 NS_123 0 -1.4880453955215419e-06
GC_1_124 b_1 NI_1 NS_124 0 -1.2743198722750780e-08
GC_1_125 b_1 NI_1 NS_125 0 2.5843959549143818e-10
GC_1_126 b_1 NI_1 NS_126 0 -1.6682804801532088e-11
GC_1_127 b_1 NI_1 NS_127 0 -1.1230022019952073e-06
GC_1_128 b_1 NI_1 NS_128 0 3.9730700565037270e-06
GC_1_129 b_1 NI_1 NS_129 0 2.2350120861744729e-06
GC_1_130 b_1 NI_1 NS_130 0 9.1477028494247728e-06
GC_1_131 b_1 NI_1 NS_131 0 1.0925656292127522e-05
GC_1_132 b_1 NI_1 NS_132 0 3.7171221365333942e-06
GC_1_133 b_1 NI_1 NS_133 0 1.4672172692365044e-05
GC_1_134 b_1 NI_1 NS_134 0 3.1019472490304148e-05
GC_1_135 b_1 NI_1 NS_135 0 3.7950165705387814e-05
GC_1_136 b_1 NI_1 NS_136 0 -6.4987152579985193e-05
GC_1_137 b_1 NI_1 NS_137 0 -7.1220149208146759e-06
GC_1_138 b_1 NI_1 NS_138 0 1.5944609022413496e-05
GC_1_139 b_1 NI_1 NS_139 0 -1.4986071140652405e-06
GC_1_140 b_1 NI_1 NS_140 0 -5.1723139725574585e-06
GC_1_141 b_1 NI_1 NS_141 0 5.0854222089303821e-05
GC_1_142 b_1 NI_1 NS_142 0 -3.8778256953404159e-05
GC_1_143 b_1 NI_1 NS_143 0 6.8081277313992227e-06
GC_1_144 b_1 NI_1 NS_144 0 -1.4682990708260841e-08
GC_1_145 b_1 NI_1 NS_145 0 -3.5990523365917259e-11
GC_1_146 b_1 NI_1 NS_146 0 8.7893645634310847e-13
GC_1_147 b_1 NI_1 NS_147 0 -3.8162801567230239e-07
GC_1_148 b_1 NI_1 NS_148 0 -1.0212853529113893e-06
GC_1_149 b_1 NI_1 NS_149 0 2.1520818382620026e-06
GC_1_150 b_1 NI_1 NS_150 0 2.5509758361901706e-06
GC_1_151 b_1 NI_1 NS_151 0 3.8434424963564309e-06
GC_1_152 b_1 NI_1 NS_152 0 -4.0510586480238736e-06
GC_1_153 b_1 NI_1 NS_153 0 9.5840558260081111e-06
GC_1_154 b_1 NI_1 NS_154 0 -1.5381445166057243e-05
GC_1_155 b_1 NI_1 NS_155 0 -2.5653773362983723e-05
GC_1_156 b_1 NI_1 NS_156 0 -8.5208277581455236e-06
GC_1_157 b_1 NI_1 NS_157 0 2.3656838935736340e-06
GC_1_158 b_1 NI_1 NS_158 0 2.6330662706018348e-07
GC_1_159 b_1 NI_1 NS_159 0 -6.9147863554886559e-06
GC_1_160 b_1 NI_1 NS_160 0 -3.8167757801324720e-06
GC_1_161 b_1 NI_1 NS_161 0 5.6957078589317183e-06
GC_1_162 b_1 NI_1 NS_162 0 1.3939729309714481e-06
GC_1_163 b_1 NI_1 NS_163 0 -8.6838689453685892e-07
GC_1_164 b_1 NI_1 NS_164 0 3.5299822202200857e-09
GC_1_165 b_1 NI_1 NS_165 0 5.0050039741821726e-11
GC_1_166 b_1 NI_1 NS_166 0 -5.2578434755579337e-13
GC_1_167 b_1 NI_1 NS_167 0 -4.1796103188657673e-07
GC_1_168 b_1 NI_1 NS_168 0 -3.4615031928794605e-07
GC_1_169 b_1 NI_1 NS_169 0 -2.5593579159445760e-07
GC_1_170 b_1 NI_1 NS_170 0 2.1882228006657227e-07
GC_1_171 b_1 NI_1 NS_171 0 -7.9356264370504717e-07
GC_1_172 b_1 NI_1 NS_172 0 -6.7751049490229573e-07
GC_1_173 b_1 NI_1 NS_173 0 -2.5395446892360772e-06
GC_1_174 b_1 NI_1 NS_174 0 -5.4510480920204044e-08
GC_1_175 b_1 NI_1 NS_175 0 3.9405128705713880e-07
GC_1_176 b_1 NI_1 NS_176 0 3.5255764539304816e-06
GC_1_177 b_1 NI_1 NS_177 0 1.6398897929622087e-07
GC_1_178 b_1 NI_1 NS_178 0 -8.5380562625846708e-07
GC_1_179 b_1 NI_1 NS_179 0 -5.5850074062002046e-07
GC_1_180 b_1 NI_1 NS_180 0 2.6967845329241072e-07
GC_1_181 b_1 NI_1 NS_181 0 2.0691347130963628e-05
GC_1_182 b_1 NI_1 NS_182 0 -5.0104189578278726e-06
GC_1_183 b_1 NI_1 NS_183 0 9.9579383426208865e-07
GC_1_184 b_1 NI_1 NS_184 0 -5.5012565982915650e-09
GC_1_185 b_1 NI_1 NS_185 0 -2.5924673896373743e-11
GC_1_186 b_1 NI_1 NS_186 0 -1.2333431834935791e-12
GC_1_187 b_1 NI_1 NS_187 0 -1.3186628476169182e-06
GC_1_188 b_1 NI_1 NS_188 0 -1.6811875391948890e-06
GC_1_189 b_1 NI_1 NS_189 0 -1.8034002166945665e-06
GC_1_190 b_1 NI_1 NS_190 0 1.3685259497731990e-07
GC_1_191 b_1 NI_1 NS_191 0 -2.4181788574415175e-06
GC_1_192 b_1 NI_1 NS_192 0 2.2165264281078320e-06
GC_1_193 b_1 NI_1 NS_193 0 -3.9553369199296092e-06
GC_1_194 b_1 NI_1 NS_194 0 -2.1598084328824272e-06
GC_1_195 b_1 NI_1 NS_195 0 1.2334122830184309e-06
GC_1_196 b_1 NI_1 NS_196 0 8.3243685029840140e-06
GC_1_197 b_1 NI_1 NS_197 0 -3.9465893517720630e-07
GC_1_198 b_1 NI_1 NS_198 0 -1.7930222420454247e-06
GC_1_199 b_1 NI_1 NS_199 0 -3.7110457532973728e-07
GC_1_200 b_1 NI_1 NS_200 0 1.7920447625762634e-07
GC_1_201 b_1 NI_1 NS_201 0 7.3331175758441455e-06
GC_1_202 b_1 NI_1 NS_202 0 -2.5197811676477146e-06
GC_1_203 b_1 NI_1 NS_203 0 1.5310189338446640e-07
GC_1_204 b_1 NI_1 NS_204 0 -4.0111443223945841e-09
GC_1_205 b_1 NI_1 NS_205 0 1.6388490745715528e-10
GC_1_206 b_1 NI_1 NS_206 0 -1.2217803739948424e-11
GC_1_207 b_1 NI_1 NS_207 0 -3.1670348498420010e-07
GC_1_208 b_1 NI_1 NS_208 0 -2.3700963496602472e-07
GC_1_209 b_1 NI_1 NS_209 0 -7.6440599693101310e-08
GC_1_210 b_1 NI_1 NS_210 0 9.2571227597350734e-08
GC_1_211 b_1 NI_1 NS_211 0 -7.8260990262121858e-07
GC_1_212 b_1 NI_1 NS_212 0 -4.1598991822905669e-07
GC_1_213 b_1 NI_1 NS_213 0 -9.7698214886938907e-07
GC_1_214 b_1 NI_1 NS_214 0 4.5608533649495976e-07
GC_1_215 b_1 NI_1 NS_215 0 2.6664085224432563e-07
GC_1_216 b_1 NI_1 NS_216 0 3.1017425434540972e-07
GC_1_217 b_1 NI_1 NS_217 0 -1.5147407088239185e-07
GC_1_218 b_1 NI_1 NS_218 0 -3.1214807552743551e-07
GC_1_219 b_1 NI_1 NS_219 0 -8.8434219582879401e-07
GC_1_220 b_1 NI_1 NS_220 0 -4.0322299204533123e-07
GC_1_221 b_1 NI_1 NS_221 0 -6.3363383158008942e-07
GC_1_222 b_1 NI_1 NS_222 0 -6.2720233513433424e-07
GC_1_223 b_1 NI_1 NS_223 0 -7.3992681743997451e-08
GC_1_224 b_1 NI_1 NS_224 0 4.6611083992340127e-09
GC_1_225 b_1 NI_1 NS_225 0 -1.7625100700396750e-10
GC_1_226 b_1 NI_1 NS_226 0 1.2487328262934047e-11
GC_1_227 b_1 NI_1 NS_227 0 9.0959399721026150e-07
GC_1_228 b_1 NI_1 NS_228 0 -8.4398007282656367e-07
GC_1_229 b_1 NI_1 NS_229 0 1.2588118524643978e-06
GC_1_230 b_1 NI_1 NS_230 0 -1.6665155546594817e-07
GC_1_231 b_1 NI_1 NS_231 0 -1.8644413649230941e-07
GC_1_232 b_1 NI_1 NS_232 0 -1.1990627923211708e-06
GC_1_233 b_1 NI_1 NS_233 0 2.8924859388333922e-06
GC_1_234 b_1 NI_1 NS_234 0 -4.1240301185804683e-06
GC_1_235 b_1 NI_1 NS_235 0 -8.7582632744413000e-06
GC_1_236 b_1 NI_1 NS_236 0 4.8513133872891340e-08
GC_1_237 b_1 NI_1 NS_237 0 2.1514264106252252e-06
GC_1_238 b_1 NI_1 NS_238 0 -3.9711516241141303e-07
GC_1_239 b_1 NI_1 NS_239 0 -8.8852833478672687e-07
GC_1_240 b_1 NI_1 NS_240 0 8.3679149916746122e-07
GD_1_1 b_1 NI_1 NA_1 0 -6.6119424152693285e-03
GD_1_2 b_1 NI_1 NA_2 0 5.7256231429356333e-02
GD_1_3 b_1 NI_1 NA_3 0 6.2239313359402247e-03
GD_1_4 b_1 NI_1 NA_4 0 2.3474509773005838e-03
GD_1_5 b_1 NI_1 NA_5 0 -6.6464568311446059e-05
GD_1_6 b_1 NI_1 NA_6 0 7.8745445807131756e-06
GD_1_7 b_1 NI_1 NA_7 0 1.9756190513807335e-05
GD_1_8 b_1 NI_1 NA_8 0 -3.9272307753418902e-06
GD_1_9 b_1 NI_1 NA_9 0 -2.2799323424937022e-06
GD_1_10 b_1 NI_1 NA_10 0 -1.0364077262790966e-05
GD_1_11 b_1 NI_1 NA_11 0 -2.3878575458006216e-06
GD_1_12 b_1 NI_1 NA_12 0 6.5403346453427850e-06
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 -2.8699894458250119e-01
GC_2_2 b_2 NI_2 NS_2 0 1.2135745353105520e-01
GC_2_3 b_2 NI_2 NS_3 0 7.0298414593019179e-03
GC_2_4 b_2 NI_2 NS_4 0 5.7777328223358546e-05
GC_2_5 b_2 NI_2 NS_5 0 1.2954678440773548e-06
GC_2_6 b_2 NI_2 NS_6 0 1.4196095550236526e-08
GC_2_7 b_2 NI_2 NS_7 0 3.0514954625909849e-02
GC_2_8 b_2 NI_2 NS_8 0 4.1653129350299849e-03
GC_2_9 b_2 NI_2 NS_9 0 -7.3041993281922103e-03
GC_2_10 b_2 NI_2 NS_10 0 2.2210831950473894e-02
GC_2_11 b_2 NI_2 NS_11 0 -1.6943519262066008e-02
GC_2_12 b_2 NI_2 NS_12 0 -1.8718656039767408e-02
GC_2_13 b_2 NI_2 NS_13 0 4.4820829361716961e-02
GC_2_14 b_2 NI_2 NS_14 0 1.4501652354770979e-02
GC_2_15 b_2 NI_2 NS_15 0 8.2246056282419433e-02
GC_2_16 b_2 NI_2 NS_16 0 3.0932605629839460e-02
GC_2_17 b_2 NI_2 NS_17 0 -1.0134686024784798e-02
GC_2_18 b_2 NI_2 NS_18 0 -4.8138241034932031e-03
GC_2_19 b_2 NI_2 NS_19 0 -2.1451541522689219e-02
GC_2_20 b_2 NI_2 NS_20 0 -4.8857424813007590e-03
GC_2_21 b_2 NI_2 NS_21 0 -1.0222189382686536e-03
GC_2_22 b_2 NI_2 NS_22 0 -1.7322668026375908e-02
GC_2_23 b_2 NI_2 NS_23 0 1.1757822387305567e-02
GC_2_24 b_2 NI_2 NS_24 0 2.8947520427772757e-06
GC_2_25 b_2 NI_2 NS_25 0 -5.0926480052767828e-07
GC_2_26 b_2 NI_2 NS_26 0 -2.9660693246163512e-08
GC_2_27 b_2 NI_2 NS_27 0 3.0704128506545063e-03
GC_2_28 b_2 NI_2 NS_28 0 1.2919121928318910e-03
GC_2_29 b_2 NI_2 NS_29 0 -2.9518618707215062e-03
GC_2_30 b_2 NI_2 NS_30 0 -9.9170148249822024e-03
GC_2_31 b_2 NI_2 NS_31 0 5.8893975062115607e-04
GC_2_32 b_2 NI_2 NS_32 0 1.3640194001803980e-02
GC_2_33 b_2 NI_2 NS_33 0 1.7423650650642910e-02
GC_2_34 b_2 NI_2 NS_34 0 -2.3868296008015443e-02
GC_2_35 b_2 NI_2 NS_35 0 -3.3167484266264688e-02
GC_2_36 b_2 NI_2 NS_36 0 2.1401807985247365e-02
GC_2_37 b_2 NI_2 NS_37 0 4.0587922746253930e-03
GC_2_38 b_2 NI_2 NS_38 0 -2.2320128311773412e-03
GC_2_39 b_2 NI_2 NS_39 0 1.5116274598290062e-02
GC_2_40 b_2 NI_2 NS_40 0 5.6072380779884686e-03
GC_2_41 b_2 NI_2 NS_41 0 -8.2288459820620066e-02
GC_2_42 b_2 NI_2 NS_42 0 6.5322021497881744e-02
GC_2_43 b_2 NI_2 NS_43 0 -1.0307113947331676e-02
GC_2_44 b_2 NI_2 NS_44 0 -2.3858545423345970e-06
GC_2_45 b_2 NI_2 NS_45 0 1.6335232744058055e-08
GC_2_46 b_2 NI_2 NS_46 0 1.6410072798340605e-09
GC_2_47 b_2 NI_2 NS_47 0 -3.9597056283257069e-04
GC_2_48 b_2 NI_2 NS_48 0 -1.4000568072940981e-03
GC_2_49 b_2 NI_2 NS_49 0 -6.9917492851545643e-03
GC_2_50 b_2 NI_2 NS_50 0 -3.7822427319941032e-03
GC_2_51 b_2 NI_2 NS_51 0 -9.0594504362458816e-03
GC_2_52 b_2 NI_2 NS_52 0 1.3121192465553386e-02
GC_2_53 b_2 NI_2 NS_53 0 -1.5240954526060871e-02
GC_2_54 b_2 NI_2 NS_54 0 2.8718756330228731e-02
GC_2_55 b_2 NI_2 NS_55 0 4.5110991131374546e-02
GC_2_56 b_2 NI_2 NS_56 0 1.6488627946037705e-02
GC_2_57 b_2 NI_2 NS_57 0 -2.2090754467328131e-03
GC_2_58 b_2 NI_2 NS_58 0 -1.3391798350294770e-03
GC_2_59 b_2 NI_2 NS_59 0 1.2863710635988242e-02
GC_2_60 b_2 NI_2 NS_60 0 6.9572426980069003e-03
GC_2_61 b_2 NI_2 NS_61 0 2.2267884546061077e-02
GC_2_62 b_2 NI_2 NS_62 0 8.9573195774672893e-03
GC_2_63 b_2 NI_2 NS_63 0 -1.1409899388773091e-02
GC_2_64 b_2 NI_2 NS_64 0 -5.3357066118445833e-06
GC_2_65 b_2 NI_2 NS_65 0 -9.5823210023365753e-08
GC_2_66 b_2 NI_2 NS_66 0 -1.2410082342728397e-09
GC_2_67 b_2 NI_2 NS_67 0 -3.3142114616009346e-03
GC_2_68 b_2 NI_2 NS_68 0 -2.3908942851530901e-03
GC_2_69 b_2 NI_2 NS_69 0 2.7265905726581536e-03
GC_2_70 b_2 NI_2 NS_70 0 1.1171998297267328e-02
GC_2_71 b_2 NI_2 NS_71 0 -3.5268616804207239e-04
GC_2_72 b_2 NI_2 NS_72 0 -1.7759691461714484e-02
GC_2_73 b_2 NI_2 NS_73 0 -2.2020324822123571e-02
GC_2_74 b_2 NI_2 NS_74 0 2.1327615899668265e-02
GC_2_75 b_2 NI_2 NS_75 0 2.8910199692313818e-02
GC_2_76 b_2 NI_2 NS_76 0 -1.8399087807940258e-02
GC_2_77 b_2 NI_2 NS_77 0 -2.4511198413732656e-03
GC_2_78 b_2 NI_2 NS_78 0 1.4222320248858224e-03
GC_2_79 b_2 NI_2 NS_79 0 -1.7818694628047235e-02
GC_2_80 b_2 NI_2 NS_80 0 -7.1267647328478977e-03
GC_2_81 b_2 NI_2 NS_81 0 3.0050542053710228e-04
GC_2_82 b_2 NI_2 NS_82 0 -2.6759720550306542e-04
GC_2_83 b_2 NI_2 NS_83 0 4.2937783943979142e-05
GC_2_84 b_2 NI_2 NS_84 0 1.3912054734518844e-08
GC_2_85 b_2 NI_2 NS_85 0 -1.4978819714139652e-10
GC_2_86 b_2 NI_2 NS_86 0 1.4933412186004478e-11
GC_2_87 b_2 NI_2 NS_87 0 2.1661615986515927e-06
GC_2_88 b_2 NI_2 NS_88 0 7.3079536077980415e-06
GC_2_89 b_2 NI_2 NS_89 0 3.3345900348392432e-05
GC_2_90 b_2 NI_2 NS_90 0 2.1777980028651739e-05
GC_2_91 b_2 NI_2 NS_91 0 4.6481490590295578e-05
GC_2_92 b_2 NI_2 NS_92 0 -5.6794136976896553e-05
GC_2_93 b_2 NI_2 NS_93 0 7.4766882138452856e-05
GC_2_94 b_2 NI_2 NS_94 0 -1.2484469947891569e-04
GC_2_95 b_2 NI_2 NS_95 0 -1.8751805292421250e-04
GC_2_96 b_2 NI_2 NS_96 0 -7.7196110248134689e-05
GC_2_97 b_2 NI_2 NS_97 0 8.1430442366634552e-06
GC_2_98 b_2 NI_2 NS_98 0 4.1233497114678235e-06
GC_2_99 b_2 NI_2 NS_99 0 -5.4121375029434786e-05
GC_2_100 b_2 NI_2 NS_100 0 -3.1122467438644958e-05
GC_2_101 b_2 NI_2 NS_101 0 2.7270670865859719e-04
GC_2_102 b_2 NI_2 NS_102 0 -1.1383754918183681e-05
GC_2_103 b_2 NI_2 NS_103 0 -9.5559239890018922e-06
GC_2_104 b_2 NI_2 NS_104 0 6.1073863577110944e-08
GC_2_105 b_2 NI_2 NS_105 0 -3.1719513694265935e-10
GC_2_106 b_2 NI_2 NS_106 0 9.0131926092120304e-12
GC_2_107 b_2 NI_2 NS_107 0 -4.9941248535091549e-07
GC_2_108 b_2 NI_2 NS_108 0 -1.5410044228998580e-05
GC_2_109 b_2 NI_2 NS_109 0 -9.6053241956152017e-06
GC_2_110 b_2 NI_2 NS_110 0 -2.0782388683127278e-05
GC_2_111 b_2 NI_2 NS_111 0 -3.7546626578110078e-05
GC_2_112 b_2 NI_2 NS_112 0 -1.9743152762149715e-05
GC_2_113 b_2 NI_2 NS_113 0 -7.4988912989486836e-05
GC_2_114 b_2 NI_2 NS_114 0 -7.8362507787239563e-05
GC_2_115 b_2 NI_2 NS_115 0 -7.3509913341744849e-05
GC_2_116 b_2 NI_2 NS_116 0 2.1939666113014335e-04
GC_2_117 b_2 NI_2 NS_117 0 1.4867517443734584e-05
GC_2_118 b_2 NI_2 NS_118 0 -5.7361994193714254e-05
GC_2_119 b_2 NI_2 NS_119 0 -4.6235340300279596e-06
GC_2_120 b_2 NI_2 NS_120 0 1.3685042718479841e-05
GC_2_121 b_2 NI_2 NS_121 0 5.0922300318150649e-05
GC_2_122 b_2 NI_2 NS_122 0 -3.8768878137450510e-05
GC_2_123 b_2 NI_2 NS_123 0 6.8058308923623234e-06
GC_2_124 b_2 NI_2 NS_124 0 -1.4678932838006855e-08
GC_2_125 b_2 NI_2 NS_125 0 -3.5984990025810006e-11
GC_2_126 b_2 NI_2 NS_126 0 8.7816991199916913e-13
GC_2_127 b_2 NI_2 NS_127 0 -3.9997179124826264e-07
GC_2_128 b_2 NI_2 NS_128 0 -1.0354839597402132e-06
GC_2_129 b_2 NI_2 NS_129 0 2.1268629798489244e-06
GC_2_130 b_2 NI_2 NS_130 0 2.5480817560958453e-06
GC_2_131 b_2 NI_2 NS_131 0 3.8281434013993134e-06
GC_2_132 b_2 NI_2 NS_132 0 -4.0076899451993602e-06
GC_2_133 b_2 NI_2 NS_133 0 9.5696476413966318e-06
GC_2_134 b_2 NI_2 NS_134 0 -1.5346625777712684e-05
GC_2_135 b_2 NI_2 NS_135 0 -2.5610119870208083e-05
GC_2_136 b_2 NI_2 NS_136 0 -8.5179434818633077e-06
GC_2_137 b_2 NI_2 NS_137 0 2.3607084068265978e-06
GC_2_138 b_2 NI_2 NS_138 0 2.6764576103192390e-07
GC_2_139 b_2 NI_2 NS_139 0 -6.9119888644840941e-06
GC_2_140 b_2 NI_2 NS_140 0 -3.8140226249673423e-06
GC_2_141 b_2 NI_2 NS_141 0 -8.6883715509151753e-05
GC_2_142 b_2 NI_2 NS_142 0 1.4652651970756272e-05
GC_2_143 b_2 NI_2 NS_143 0 -1.4888053428043621e-06
GC_2_144 b_2 NI_2 NS_144 0 -1.2740379588515129e-08
GC_2_145 b_2 NI_2 NS_145 0 2.5839541817869070e-10
GC_2_146 b_2 NI_2 NS_146 0 -1.6679185663090425e-11
GC_2_147 b_2 NI_2 NS_147 0 -1.1229325319838877e-06
GC_2_148 b_2 NI_2 NS_148 0 3.9744249291720533e-06
GC_2_149 b_2 NI_2 NS_149 0 2.2362284542230004e-06
GC_2_150 b_2 NI_2 NS_150 0 9.1490008594632574e-06
GC_2_151 b_2 NI_2 NS_151 0 1.0926853409797484e-05
GC_2_152 b_2 NI_2 NS_152 0 3.7178690530487305e-06
GC_2_153 b_2 NI_2 NS_153 0 1.4674343645948292e-05
GC_2_154 b_2 NI_2 NS_154 0 3.1025615722756359e-05
GC_2_155 b_2 NI_2 NS_155 0 3.7960203886374840e-05
GC_2_156 b_2 NI_2 NS_156 0 -6.4994945843353219e-05
GC_2_157 b_2 NI_2 NS_157 0 -7.1240281916145294e-06
GC_2_158 b_2 NI_2 NS_158 0 1.5945791166708479e-05
GC_2_159 b_2 NI_2 NS_159 0 -1.4978347788730602e-06
GC_2_160 b_2 NI_2 NS_160 0 -5.1730650951062279e-06
GC_2_161 b_2 NI_2 NS_161 0 2.0691198168796381e-05
GC_2_162 b_2 NI_2 NS_162 0 -5.0103740550481953e-06
GC_2_163 b_2 NI_2 NS_163 0 9.9579017701263890e-07
GC_2_164 b_2 NI_2 NS_164 0 -5.5012629444656805e-09
GC_2_165 b_2 NI_2 NS_165 0 -2.5924586063993116e-11
GC_2_166 b_2 NI_2 NS_166 0 -1.2333507835956672e-12
GC_2_167 b_2 NI_2 NS_167 0 -1.3186727749723603e-06
GC_2_168 b_2 NI_2 NS_168 0 -1.6811813959867443e-06
GC_2_169 b_2 NI_2 NS_169 0 -1.8034084224086242e-06
GC_2_170 b_2 NI_2 NS_170 0 1.3686982559270639e-07
GC_2_171 b_2 NI_2 NS_171 0 -2.4181483922279950e-06
GC_2_172 b_2 NI_2 NS_172 0 2.2165533373700290e-06
GC_2_173 b_2 NI_2 NS_173 0 -3.9553010071183763e-06
GC_2_174 b_2 NI_2 NS_174 0 -2.1597716303056818e-06
GC_2_175 b_2 NI_2 NS_175 0 1.2334459301345174e-06
GC_2_176 b_2 NI_2 NS_176 0 8.3243112226966604e-06
GC_2_177 b_2 NI_2 NS_177 0 -3.9465642639280213e-07
GC_2_178 b_2 NI_2 NS_178 0 -1.7930162893825012e-06
GC_2_179 b_2 NI_2 NS_179 0 -3.7109497862337424e-07
GC_2_180 b_2 NI_2 NS_180 0 1.7920059558833948e-07
GC_2_181 b_2 NI_2 NS_181 0 5.7390983489177019e-06
GC_2_182 b_2 NI_2 NS_182 0 1.3787314949332164e-06
GC_2_183 b_2 NI_2 NS_183 0 -8.6637353524023401e-07
GC_2_184 b_2 NI_2 NS_184 0 3.5224550118579967e-09
GC_2_185 b_2 NI_2 NS_185 0 5.0090034504675750e-11
GC_2_186 b_2 NI_2 NS_186 0 -5.2606127766883666e-13
GC_2_187 b_2 NI_2 NS_187 0 -4.1959946098212356e-07
GC_2_188 b_2 NI_2 NS_188 0 -3.4603312569527518e-07
GC_2_189 b_2 NI_2 NS_189 0 -2.5691671794445418e-07
GC_2_190 b_2 NI_2 NS_190 0 2.1863620693730043e-07
GC_2_191 b_2 NI_2 NS_191 0 -7.9604795155344134e-07
GC_2_192 b_2 NI_2 NS_192 0 -6.7621312443822101e-07
GC_2_193 b_2 NI_2 NS_193 0 -2.5375268014869291e-06
GC_2_194 b_2 NI_2 NS_194 0 -5.5017973704381433e-08
GC_2_195 b_2 NI_2 NS_195 0 3.8307261139220780e-07
GC_2_196 b_2 NI_2 NS_196 0 3.5238201770390337e-06
GC_2_197 b_2 NI_2 NS_197 0 1.6617776593318304e-07
GC_2_198 b_2 NI_2 NS_198 0 -8.5364107575662573e-07
GC_2_199 b_2 NI_2 NS_199 0 -5.6158084151636612e-07
GC_2_200 b_2 NI_2 NS_200 0 2.6962865361425876e-07
GC_2_201 b_2 NI_2 NS_201 0 -6.3290792754018104e-07
GC_2_202 b_2 NI_2 NS_202 0 -6.2866891407781015e-07
GC_2_203 b_2 NI_2 NS_203 0 -7.3718811956199496e-08
GC_2_204 b_2 NI_2 NS_204 0 4.6597131236442592e-09
GC_2_205 b_2 NI_2 NS_205 0 -1.7622882774429318e-10
GC_2_206 b_2 NI_2 NS_206 0 1.2485704757046103e-11
GC_2_207 b_2 NI_2 NS_207 0 9.0995539361595203e-07
GC_2_208 b_2 NI_2 NS_208 0 -8.4388376522697450e-07
GC_2_209 b_2 NI_2 NS_209 0 1.2594059030871272e-06
GC_2_210 b_2 NI_2 NS_210 0 -1.6700305830922089e-07
GC_2_211 b_2 NI_2 NS_211 0 -1.8724478297083948e-07
GC_2_212 b_2 NI_2 NS_212 0 -1.1999801573792754e-06
GC_2_213 b_2 NI_2 NS_213 0 2.8912207838340882e-06
GC_2_214 b_2 NI_2 NS_214 0 -4.1236266531124756e-06
GC_2_215 b_2 NI_2 NS_215 0 -8.7556922816342635e-06
GC_2_216 b_2 NI_2 NS_216 0 4.7054618193474399e-08
GC_2_217 b_2 NI_2 NS_217 0 2.1502533922955005e-06
GC_2_218 b_2 NI_2 NS_218 0 -3.9617847804228137e-07
GC_2_219 b_2 NI_2 NS_219 0 -8.8887429927983292e-07
GC_2_220 b_2 NI_2 NS_220 0 8.3645542566945973e-07
GC_2_221 b_2 NI_2 NS_221 0 7.3320647045636195e-06
GC_2_222 b_2 NI_2 NS_222 0 -2.5195979229801521e-06
GC_2_223 b_2 NI_2 NS_223 0 1.5308903242283245e-07
GC_2_224 b_2 NI_2 NS_224 0 -4.0110866472051807e-09
GC_2_225 b_2 NI_2 NS_225 0 1.6388396416454157e-10
GC_2_226 b_2 NI_2 NS_226 0 -1.2217730760225527e-11
GC_2_227 b_2 NI_2 NS_227 0 -3.1665109368060729e-07
GC_2_228 b_2 NI_2 NS_228 0 -2.3698644395225053e-07
GC_2_229 b_2 NI_2 NS_229 0 -7.6390776579433845e-08
GC_2_230 b_2 NI_2 NS_230 0 9.2605485366437068e-08
GC_2_231 b_2 NI_2 NS_231 0 -7.8248638765588618e-07
GC_2_232 b_2 NI_2 NS_232 0 -4.1603029503422030e-07
GC_2_233 b_2 NI_2 NS_233 0 -9.7686400442770293e-07
GC_2_234 b_2 NI_2 NS_234 0 4.5613973112896631e-07
GC_2_235 b_2 NI_2 NS_235 0 2.6679512100947969e-07
GC_2_236 b_2 NI_2 NS_236 0 3.0984695492726131e-07
GC_2_237 b_2 NI_2 NS_237 0 -1.5150711809875050e-07
GC_2_238 b_2 NI_2 NS_238 0 -3.1207026403153876e-07
GC_2_239 b_2 NI_2 NS_239 0 -8.8431500781467000e-07
GC_2_240 b_2 NI_2 NS_240 0 -4.0325455569697637e-07
GD_2_1 b_2 NI_2 NA_1 0 5.7256339596373149e-02
GD_2_2 b_2 NI_2 NA_2 0 -6.6119424152692730e-03
GD_2_3 b_2 NI_2 NA_3 0 2.3474503953194430e-03
GD_2_4 b_2 NI_2 NA_4 0 6.2259683072083327e-03
GD_2_5 b_2 NI_2 NA_5 0 7.8739705187710485e-06
GD_2_6 b_2 NI_2 NA_6 0 -6.6955532859409590e-05
GD_2_7 b_2 NI_2 NA_7 0 -3.9775986893964339e-06
GD_2_8 b_2 NI_2 NA_8 0 1.9757259604378204e-05
GD_2_9 b_2 NI_2 NA_9 0 -1.0364068610811252e-05
GD_2_10 b_2 NI_2 NA_10 0 -2.3046839896073086e-06
GD_2_11 b_2 NI_2 NA_11 0 6.5411158686230532e-06
GD_2_12 b_2 NI_2 NA_12 0 -2.3872964722855127e-06
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 2.2267884546061229e-02
GC_3_2 b_3 NI_3 NS_2 0 8.9573195774672112e-03
GC_3_3 b_3 NI_3 NS_3 0 -1.1409899388773070e-02
GC_3_4 b_3 NI_3 NS_4 0 -5.3357066118453770e-06
GC_3_5 b_3 NI_3 NS_5 0 -9.5823210023361981e-08
GC_3_6 b_3 NI_3 NS_6 0 -1.2410082342723525e-09
GC_3_7 b_3 NI_3 NS_7 0 -3.3142114616009277e-03
GC_3_8 b_3 NI_3 NS_8 0 -2.3908942851530932e-03
GC_3_9 b_3 NI_3 NS_9 0 2.7265905726581289e-03
GC_3_10 b_3 NI_3 NS_10 0 1.1171998297267330e-02
GC_3_11 b_3 NI_3 NS_11 0 -3.5268616804206036e-04
GC_3_12 b_3 NI_3 NS_12 0 -1.7759691461714477e-02
GC_3_13 b_3 NI_3 NS_13 0 -2.2020324822123558e-02
GC_3_14 b_3 NI_3 NS_14 0 2.1327615899668268e-02
GC_3_15 b_3 NI_3 NS_15 0 2.8910199692313749e-02
GC_3_16 b_3 NI_3 NS_16 0 -1.8399087807940289e-02
GC_3_17 b_3 NI_3 NS_17 0 -2.4511198413732418e-03
GC_3_18 b_3 NI_3 NS_18 0 1.4222320248858324e-03
GC_3_19 b_3 NI_3 NS_19 0 -1.7818694628047249e-02
GC_3_20 b_3 NI_3 NS_20 0 -7.1267647328478977e-03
GC_3_21 b_3 NI_3 NS_21 0 -8.2288461357651374e-02
GC_3_22 b_3 NI_3 NS_22 0 6.5322021842723801e-02
GC_3_23 b_3 NI_3 NS_23 0 -1.0307113986153655e-02
GC_3_24 b_3 NI_3 NS_24 0 -2.3858543821315970e-06
GC_3_25 b_3 NI_3 NS_25 0 1.6335231358585063e-08
GC_3_26 b_3 NI_3 NS_26 0 1.6410073214708445e-09
GC_3_27 b_3 NI_3 NS_27 0 -3.9597044109948983e-04
GC_3_28 b_3 NI_3 NS_28 0 -1.4000567034305651e-03
GC_3_29 b_3 NI_3 NS_29 0 -6.9917491213848685e-03
GC_3_30 b_3 NI_3 NS_30 0 -3.7822426989903655e-03
GC_3_31 b_3 NI_3 NS_31 0 -9.0594503196265407e-03
GC_3_32 b_3 NI_3 NS_32 0 1.3121192277925849e-02
GC_3_33 b_3 NI_3 NS_33 0 -1.5240954433953841e-02
GC_3_34 b_3 NI_3 NS_34 0 2.8718756400073122e-02
GC_3_35 b_3 NI_3 NS_35 0 4.5110991420963739e-02
GC_3_36 b_3 NI_3 NS_36 0 1.6488627629001454e-02
GC_3_37 b_3 NI_3 NS_37 0 -2.2090755305097859e-03
GC_3_38 b_3 NI_3 NS_38 0 -1.3391797801787248e-03
GC_3_39 b_3 NI_3 NS_39 0 1.2863710673931708e-02
GC_3_40 b_3 NI_3 NS_40 0 6.9572426668203053e-03
GC_3_41 b_3 NI_3 NS_41 0 -1.4551902072501201e-03
GC_3_42 b_3 NI_3 NS_42 0 -1.7225749581186531e-02
GC_3_43 b_3 NI_3 NS_43 0 1.1743970365723822e-02
GC_3_44 b_3 NI_3 NS_44 0 2.9971096683402701e-06
GC_3_45 b_3 NI_3 NS_45 0 -5.0997795379026973e-07
GC_3_46 b_3 NI_3 NS_46 0 -2.9633812117832443e-08
GC_3_47 b_3 NI_3 NS_47 0 3.0965325001513226e-03
GC_3_48 b_3 NI_3 NS_48 0 1.3051943670992392e-03
GC_3_49 b_3 NI_3 NS_49 0 -2.9261127150177488e-03
GC_3_50 b_3 NI_3 NS_50 0 -9.9123416426922378e-03
GC_3_51 b_3 NI_3 NS_51 0 6.3752755685791160e-04
GC_3_52 b_3 NI_3 NS_52 0 1.3628527547780793e-02
GC_3_53 b_3 NI_3 NS_53 0 1.7509588834278004e-02
GC_3_54 b_3 NI_3 NS_54 0 -2.3852006616147687e-02
GC_3_55 b_3 NI_3 NS_55 0 -3.3177959639940809e-02
GC_3_56 b_3 NI_3 NS_56 0 2.1222695048691346e-02
GC_3_57 b_3 NI_3 NS_57 0 4.0623997774704946e-03
GC_3_58 b_3 NI_3 NS_58 0 -2.1854449406243453e-03
GC_3_59 b_3 NI_3 NS_59 0 1.5119316701147677e-02
GC_3_60 b_3 NI_3 NS_60 0 5.6106547450701112e-03
GC_3_61 b_3 NI_3 NS_61 0 -2.8564000682351648e-01
GC_3_62 b_3 NI_3 NS_62 0 1.2097605663919701e-01
GC_3_63 b_3 NI_3 NS_63 0 7.0824863396637856e-03
GC_3_64 b_3 NI_3 NS_64 0 5.7464553490901451e-05
GC_3_65 b_3 NI_3 NS_65 0 1.3019123350575353e-06
GC_3_66 b_3 NI_3 NS_66 0 1.3695318513044394e-08
GC_3_67 b_3 NI_3 NS_67 0 3.0465780292360575e-02
GC_3_68 b_3 NI_3 NS_68 0 4.1090451362333792e-03
GC_3_69 b_3 NI_3 NS_69 0 -7.3763975158783425e-03
GC_3_70 b_3 NI_3 NS_70 0 2.2180118554762790e-02
GC_3_71 b_3 NI_3 NS_71 0 -1.7056204165724221e-02
GC_3_72 b_3 NI_3 NS_72 0 -1.8685516556591893e-02
GC_3_73 b_3 NI_3 NS_73 0 4.4665639744307116e-02
GC_3_74 b_3 NI_3 NS_74 0 1.4315030871751155e-02
GC_3_75 b_3 NI_3 NS_75 0 8.2000112574895159e-02
GC_3_76 b_3 NI_3 NS_76 0 3.1380076795064660e-02
GC_3_77 b_3 NI_3 NS_77 0 -1.0089097276106938e-02
GC_3_78 b_3 NI_3 NS_78 0 -4.9101507320294729e-03
GC_3_79 b_3 NI_3 NS_79 0 -2.1483626036327204e-02
GC_3_80 b_3 NI_3 NS_80 0 -4.8833393807782644e-03
GC_3_81 b_3 NI_3 NS_81 0 1.2460295911826696e-04
GC_3_82 b_3 NI_3 NS_82 0 8.0357130131917249e-05
GC_3_83 b_3 NI_3 NS_83 0 -9.5148169956568070e-05
GC_3_84 b_3 NI_3 NS_84 0 -1.1560586044515251e-07
GC_3_85 b_3 NI_3 NS_85 0 -4.2556432309500420e-10
GC_3_86 b_3 NI_3 NS_86 0 -1.2107893778945519e-10
GC_3_87 b_3 NI_3 NS_87 0 -2.9524729677071776e-05
GC_3_88 b_3 NI_3 NS_88 0 -1.6598751286767264e-05
GC_3_89 b_3 NI_3 NS_89 0 2.8263593289912682e-05
GC_3_90 b_3 NI_3 NS_90 0 9.8568706608732527e-05
GC_3_91 b_3 NI_3 NS_91 0 -6.2941192305394754e-07
GC_3_92 b_3 NI_3 NS_92 0 -1.4684426129597057e-04
GC_3_93 b_3 NI_3 NS_93 0 -1.7067067314414602e-04
GC_3_94 b_3 NI_3 NS_94 0 2.0939417415112869e-04
GC_3_95 b_3 NI_3 NS_95 0 2.7022139311703406e-04
GC_3_96 b_3 NI_3 NS_96 0 -2.1560536352375351e-04
GC_3_97 b_3 NI_3 NS_97 0 -2.5134850254888577e-05
GC_3_98 b_3 NI_3 NS_98 0 2.6863414416776110e-05
GC_3_99 b_3 NI_3 NS_99 0 -1.5209446859752230e-04
GC_3_100 b_3 NI_3 NS_100 0 -6.3894955659849983e-05
GC_3_101 b_3 NI_3 NS_101 0 -5.3979227016776336e-04
GC_3_102 b_3 NI_3 NS_102 0 4.9388521344228425e-04
GC_3_103 b_3 NI_3 NS_103 0 -7.8319138674097725e-05
GC_3_104 b_3 NI_3 NS_104 0 9.9521379965561606e-09
GC_3_105 b_3 NI_3 NS_105 0 2.8669969292597587e-10
GC_3_106 b_3 NI_3 NS_106 0 8.0713861859436118e-11
GC_3_107 b_3 NI_3 NS_107 0 -1.2925624726765163e-05
GC_3_108 b_3 NI_3 NS_108 0 -9.1377576337082143e-06
GC_3_109 b_3 NI_3 NS_109 0 -6.7846976609626055e-05
GC_3_110 b_3 NI_3 NS_110 0 -3.2036623881078055e-05
GC_3_111 b_3 NI_3 NS_111 0 -7.1365955992728060e-05
GC_3_112 b_3 NI_3 NS_112 0 1.1523613554753181e-04
GC_3_113 b_3 NI_3 NS_113 0 -1.3883879516015209e-04
GC_3_114 b_3 NI_3 NS_114 0 2.2241980674553652e-04
GC_3_115 b_3 NI_3 NS_115 0 3.5584091692507906e-04
GC_3_116 b_3 NI_3 NS_116 0 1.6517825975792652e-04
GC_3_117 b_3 NI_3 NS_117 0 -1.7005467605479965e-05
GC_3_118 b_3 NI_3 NS_118 0 -1.8451588227691447e-05
GC_3_119 b_3 NI_3 NS_119 0 1.0145875857576514e-04
GC_3_120 b_3 NI_3 NS_120 0 5.6315095486523486e-05
GC_3_121 b_3 NI_3 NS_121 0 2.8249440155792764e-04
GC_3_122 b_3 NI_3 NS_122 0 -1.3810042512492373e-05
GC_3_123 b_3 NI_3 NS_123 0 -9.2728558000077270e-06
GC_3_124 b_3 NI_3 NS_124 0 5.9696244996697190e-08
GC_3_125 b_3 NI_3 NS_125 0 -3.0906100824666400e-10
GC_3_126 b_3 NI_3 NS_126 0 9.3204334711095520e-12
GC_3_127 b_3 NI_3 NS_127 0 -7.6635914674945889e-07
GC_3_128 b_3 NI_3 NS_128 0 -1.5748718103283603e-05
GC_3_129 b_3 NI_3 NS_129 0 -1.0078797578414015e-05
GC_3_130 b_3 NI_3 NS_130 0 -2.1107423636476820e-05
GC_3_131 b_3 NI_3 NS_131 0 -3.8248667532999075e-05
GC_3_132 b_3 NI_3 NS_132 0 -1.9774688647789564e-05
GC_3_133 b_3 NI_3 NS_133 0 -7.5998900403247350e-05
GC_3_134 b_3 NI_3 NS_134 0 -7.9943369328120892e-05
GC_3_135 b_3 NI_3 NS_135 0 -7.6445578776235818e-05
GC_3_136 b_3 NI_3 NS_136 0 2.2266396007953668e-04
GC_3_137 b_3 NI_3 NS_137 0 1.5542652459594939e-05
GC_3_138 b_3 NI_3 NS_138 0 -5.8015180970683710e-05
GC_3_139 b_3 NI_3 NS_139 0 -4.8512122609528725e-06
GC_3_140 b_3 NI_3 NS_140 0 1.3939680175418020e-05
GC_3_141 b_3 NI_3 NS_141 0 3.0534411163382126e-04
GC_3_142 b_3 NI_3 NS_142 0 -2.6784573336185931e-04
GC_3_143 b_3 NI_3 NS_143 0 4.2963844114348496e-05
GC_3_144 b_3 NI_3 NS_144 0 1.4101512850513284e-08
GC_3_145 b_3 NI_3 NS_145 0 -1.4707755849198867e-10
GC_3_146 b_3 NI_3 NS_146 0 1.3946692202775977e-11
GC_3_147 b_3 NI_3 NS_147 0 1.6536677828931433e-06
GC_3_148 b_3 NI_3 NS_148 0 7.0334548612297815e-06
GC_3_149 b_3 NI_3 NS_149 0 3.2641712283870301e-05
GC_3_150 b_3 NI_3 NS_150 0 2.1791257091342988e-05
GC_3_151 b_3 NI_3 NS_151 0 4.5840777214586724e-05
GC_3_152 b_3 NI_3 NS_152 0 -5.5994684673124077e-05
GC_3_153 b_3 NI_3 NS_153 0 7.2919506540748295e-05
GC_3_154 b_3 NI_3 NS_154 0 -1.2481997785567358e-04
GC_3_155 b_3 NI_3 NS_155 0 -1.8541625529138291e-04
GC_3_156 b_3 NI_3 NS_156 0 -7.4145716712830092e-05
GC_3_157 b_3 NI_3 NS_157 0 7.6332247874851240e-06
GC_3_158 b_3 NI_3 NS_158 0 3.5082933426251249e-06
GC_3_159 b_3 NI_3 NS_159 0 -5.3960457227613747e-05
GC_3_160 b_3 NI_3 NS_160 0 -3.1131045528218698e-05
GC_3_161 b_3 NI_3 NS_161 0 2.2539396688841493e-05
GC_3_162 b_3 NI_3 NS_162 0 -5.1374412038923287e-06
GC_3_163 b_3 NI_3 NS_163 0 3.6837553602524484e-07
GC_3_164 b_3 NI_3 NS_164 0 -8.1493386787328071e-09
GC_3_165 b_3 NI_3 NS_165 0 1.7606318050915514e-10
GC_3_166 b_3 NI_3 NS_166 0 -9.7889987614895562e-12
GC_3_167 b_3 NI_3 NS_167 0 -1.2142846318321459e-06
GC_3_168 b_3 NI_3 NS_168 0 -9.1145978060417937e-07
GC_3_169 b_3 NI_3 NS_169 0 -1.3989593787513050e-06
GC_3_170 b_3 NI_3 NS_170 0 -4.6250397239763857e-08
GC_3_171 b_3 NI_3 NS_171 0 -2.2030210655732329e-06
GC_3_172 b_3 NI_3 NS_172 0 2.2975035868267901e-08
GC_3_173 b_3 NI_3 NS_173 0 -4.7812862191182529e-06
GC_3_174 b_3 NI_3 NS_174 0 -4.5199496261919391e-07
GC_3_175 b_3 NI_3 NS_175 0 1.0107469669123644e-06
GC_3_176 b_3 NI_3 NS_176 0 7.1426263055338426e-06
GC_3_177 b_3 NI_3 NS_177 0 -3.5884019268405694e-07
GC_3_178 b_3 NI_3 NS_178 0 -1.8237683028864596e-06
GC_3_179 b_3 NI_3 NS_179 0 -1.0678367423979764e-06
GC_3_180 b_3 NI_3 NS_180 0 -3.9178573168513363e-07
GC_3_181 b_3 NI_3 NS_181 0 7.9173691911981434e-06
GC_3_182 b_3 NI_3 NS_182 0 -6.3418641539435330e-06
GC_3_183 b_3 NI_3 NS_183 0 4.7307442140779733e-07
GC_3_184 b_3 NI_3 NS_184 0 6.3738327127577391e-09
GC_3_185 b_3 NI_3 NS_185 0 -1.7569995882885665e-10
GC_3_186 b_3 NI_3 NS_186 0 8.2809630672677681e-12
GC_3_187 b_3 NI_3 NS_187 0 2.1359813963213082e-06
GC_3_188 b_3 NI_3 NS_188 0 -1.0057334268923017e-06
GC_3_189 b_3 NI_3 NS_189 0 2.8515667257536478e-06
GC_3_190 b_3 NI_3 NS_190 0 -1.3365742540816388e-06
GC_3_191 b_3 NI_3 NS_191 0 -2.5442343224583742e-07
GC_3_192 b_3 NI_3 NS_192 0 -3.4600118745845103e-06
GC_3_193 b_3 NI_3 NS_193 0 6.9380334949875354e-06
GC_3_194 b_3 NI_3 NS_194 0 -9.0883171087916401e-06
GC_3_195 b_3 NI_3 NS_195 0 -2.3892364876173340e-05
GC_3_196 b_3 NI_3 NS_196 0 -2.8584542951265020e-06
GC_3_197 b_3 NI_3 NS_197 0 5.9682595493284461e-06
GC_3_198 b_3 NI_3 NS_198 0 3.0695716082239256e-07
GC_3_199 b_3 NI_3 NS_199 0 -2.6280914026732648e-06
GC_3_200 b_3 NI_3 NS_200 0 1.4076505089819106e-06
GC_3_201 b_3 NI_3 NS_201 0 5.6987573133480891e-06
GC_3_202 b_3 NI_3 NS_202 0 1.3907358206525792e-06
GC_3_203 b_3 NI_3 NS_203 0 -8.6920422656663429e-07
GC_3_204 b_3 NI_3 NS_204 0 3.5211619203111102e-09
GC_3_205 b_3 NI_3 NS_205 0 5.0063241198897914e-11
GC_3_206 b_3 NI_3 NS_206 0 -5.2297015395387499e-13
GC_3_207 b_3 NI_3 NS_207 0 -4.1974768465539645e-07
GC_3_208 b_3 NI_3 NS_208 0 -3.4327712457799377e-07
GC_3_209 b_3 NI_3 NS_209 0 -2.5399992355724006e-07
GC_3_210 b_3 NI_3 NS_210 0 2.2159700747607230e-07
GC_3_211 b_3 NI_3 NS_211 0 -7.9481937980927909e-07
GC_3_212 b_3 NI_3 NS_212 0 -6.7506845190095032e-07
GC_3_213 b_3 NI_3 NS_213 0 -2.5308339226384579e-06
GC_3_214 b_3 NI_3 NS_214 0 -3.7212587283318559e-08
GC_3_215 b_3 NI_3 NS_215 0 4.0514420639834170e-07
GC_3_216 b_3 NI_3 NS_216 0 3.4974523945683412e-06
GC_3_217 b_3 NI_3 NS_217 0 1.6145097878951460e-07
GC_3_218 b_3 NI_3 NS_218 0 -8.5014425366163759e-07
GC_3_219 b_3 NI_3 NS_219 0 -5.6427564143747217e-07
GC_3_220 b_3 NI_3 NS_220 0 2.6709321780374799e-07
GC_3_221 b_3 NI_3 NS_221 0 2.0604781474281978e-05
GC_3_222 b_3 NI_3 NS_222 0 -4.9935578795759698e-06
GC_3_223 b_3 NI_3 NS_223 0 9.9303260511228488e-07
GC_3_224 b_3 NI_3 NS_224 0 -5.4984996775530316e-09
GC_3_225 b_3 NI_3 NS_225 0 -2.5967349839975071e-11
GC_3_226 b_3 NI_3 NS_226 0 -1.2308357975414393e-12
GC_3_227 b_3 NI_3 NS_227 0 -1.3115853203401860e-06
GC_3_228 b_3 NI_3 NS_228 0 -1.6746876351685390e-06
GC_3_229 b_3 NI_3 NS_229 0 -1.7990785522565544e-06
GC_3_230 b_3 NI_3 NS_230 0 1.3848541571339683e-07
GC_3_231 b_3 NI_3 NS_231 0 -2.4070255039826695e-06
GC_3_232 b_3 NI_3 NS_232 0 2.2075749138845694e-06
GC_3_233 b_3 NI_3 NS_233 0 -3.9348564810437927e-06
GC_3_234 b_3 NI_3 NS_234 0 -2.1436719780917977e-06
GC_3_235 b_3 NI_3 NS_235 0 1.2291045117435839e-06
GC_3_236 b_3 NI_3 NS_236 0 8.2805525602846495e-06
GC_3_237 b_3 NI_3 NS_237 0 -3.9212386807537402e-07
GC_3_238 b_3 NI_3 NS_238 0 -1.7846276179825112e-06
GC_3_239 b_3 NI_3 NS_239 0 -3.6943313999697318e-07
GC_3_240 b_3 NI_3 NS_240 0 1.7726572638980068e-07
GD_3_1 b_3 NI_3 NA_1 0 6.2259683072082659e-03
GD_3_2 b_3 NI_3 NA_2 0 2.3474509727493182e-03
GD_3_3 b_3 NI_3 NA_3 0 -6.3838899589371504e-03
GD_3_4 b_3 NI_3 NA_4 0 5.6719414776441095e-02
GD_3_5 b_3 NI_3 NA_5 0 7.4682395383388763e-05
GD_3_6 b_3 NI_3 NA_6 0 -5.2020156290454401e-05
GD_3_7 b_3 NI_3 NA_7 0 -7.0349371154274659e-05
GD_3_8 b_3 NI_3 NA_8 0 4.0802501924538473e-06
GD_3_9 b_3 NI_3 NA_9 0 -9.6644135619597490e-06
GD_3_10 b_3 NI_3 NA_10 0 1.1836313198024613e-05
GD_3_11 b_3 NI_3 NA_11 0 -2.2999152041507315e-06
GD_3_12 b_3 NI_3 NA_12 0 -1.0327427477503275e-05
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 -8.2288459819198495e-02
GC_4_2 b_4 NI_4 NS_2 0 6.5322021497353638e-02
GC_4_3 b_4 NI_4 NS_3 0 -1.0307113947270369e-02
GC_4_4 b_4 NI_4 NS_4 0 -2.3858545425141193e-06
GC_4_5 b_4 NI_4 NS_5 0 1.6335232743110106e-08
GC_4_6 b_4 NI_4 NS_6 0 1.6410072799657847e-09
GC_4_7 b_4 NI_4 NS_7 0 -3.9597056283940740e-04
GC_4_8 b_4 NI_4 NS_8 0 -1.4000568073199177e-03
GC_4_9 b_4 NI_4 NS_9 0 -6.9917492851527333e-03
GC_4_10 b_4 NI_4 NS_10 0 -3.7822427320226381e-03
GC_4_11 b_4 NI_4 NS_11 0 -9.0594504362612269e-03
GC_4_12 b_4 NI_4 NS_12 0 1.3121192465484844e-02
GC_4_13 b_4 NI_4 NS_13 0 -1.5240954525849816e-02
GC_4_14 b_4 NI_4 NS_14 0 2.8718756329897805e-02
GC_4_15 b_4 NI_4 NS_15 0 4.5110991130268757e-02
GC_4_16 b_4 NI_4 NS_16 0 1.6488627946115230e-02
GC_4_17 b_4 NI_4 NS_17 0 -2.2090754464435098e-03
GC_4_18 b_4 NI_4 NS_18 0 -1.3391798350514735e-03
GC_4_19 b_4 NI_4 NS_19 0 1.2863710635893625e-02
GC_4_20 b_4 NI_4 NS_20 0 6.9572426980583782e-03
GC_4_21 b_4 NI_4 NS_21 0 2.2274176797544301e-02
GC_4_22 b_4 NI_4 NS_22 0 8.9558630531341530e-03
GC_4_23 b_4 NI_4 NS_23 0 -1.1409760098995594e-02
GC_4_24 b_4 NI_4 NS_24 0 -5.3360833878899856e-06
GC_4_25 b_4 NI_4 NS_25 0 -9.5822579621924338e-08
GC_4_26 b_4 NI_4 NS_26 0 -1.2412250853179486e-09
GC_4_27 b_4 NI_4 NS_27 0 -3.3143877240879287e-03
GC_4_28 b_4 NI_4 NS_28 0 -2.3911427672941663e-03
GC_4_29 b_4 NI_4 NS_29 0 2.7261769899886734e-03
GC_4_30 b_4 NI_4 NS_30 0 1.1171778125851090e-02
GC_4_31 b_4 NI_4 NS_31 0 -3.5307706736995161e-04
GC_4_32 b_4 NI_4 NS_32 0 -1.7759590133315854e-02
GC_4_33 b_4 NI_4 NS_33 0 -2.2020926263780858e-02
GC_4_34 b_4 NI_4 NS_34 0 2.1326546211518693e-02
GC_4_35 b_4 NI_4 NS_35 0 2.8908349470800787e-02
GC_4_36 b_4 NI_4 NS_36 0 -1.8397053919956913e-02
GC_4_37 b_4 NI_4 NS_37 0 -2.4507569376264922e-03
GC_4_38 b_4 NI_4 NS_38 0 1.4218494193147277e-03
GC_4_39 b_4 NI_4 NS_39 0 -1.7818879772058833e-02
GC_4_40 b_4 NI_4 NS_40 0 -7.1265648084886677e-03
GC_4_41 b_4 NI_4 NS_41 0 -2.8564004784537411e-01
GC_4_42 b_4 NI_4 NS_42 0 1.2097604399740693e-01
GC_4_43 b_4 NI_4 NS_43 0 7.0824886025124215e-03
GC_4_44 b_4 NI_4 NS_44 0 5.7464564958274266e-05
GC_4_45 b_4 NI_4 NS_45 0 1.3019118326841696e-06
GC_4_46 b_4 NI_4 NS_46 0 1.3695385533275196e-08
GC_4_47 b_4 NI_4 NS_47 0 3.0465750935702744e-02
GC_4_48 b_4 NI_4 NS_48 0 4.1090315761284791e-03
GC_4_49 b_4 NI_4 NS_49 0 -7.3764419067182136e-03
GC_4_50 b_4 NI_4 NS_50 0 2.2180136525064512e-02
GC_4_51 b_4 NI_4 NS_51 0 -1.7056157523198053e-02
GC_4_52 b_4 NI_4 NS_52 0 -1.8685420136203935e-02
GC_4_53 b_4 NI_4 NS_53 0 4.4665768431487819e-02
GC_4_54 b_4 NI_4 NS_54 0 1.4315106013721631e-02
GC_4_55 b_4 NI_4 NS_55 0 8.2000031398742262e-02
GC_4_56 b_4 NI_4 NS_56 0 3.1379882771994362e-02
GC_4_57 b_4 NI_4 NS_57 0 -1.0089046784998109e-02
GC_4_58 b_4 NI_4 NS_58 0 -4.9101192870033483e-03
GC_4_59 b_4 NI_4 NS_59 0 -2.1483635707441200e-02
GC_4_60 b_4 NI_4 NS_60 0 -4.8833462056285934e-03
GC_4_61 b_4 NI_4 NS_61 0 -1.4551902072501254e-03
GC_4_62 b_4 NI_4 NS_62 0 -1.7225749581186531e-02
GC_4_63 b_4 NI_4 NS_63 0 1.1743970365723817e-02
GC_4_64 b_4 NI_4 NS_64 0 2.9971096683403582e-06
GC_4_65 b_4 NI_4 NS_65 0 -5.0997795379025490e-07
GC_4_66 b_4 NI_4 NS_66 0 -2.9633812117832777e-08
GC_4_67 b_4 NI_4 NS_67 0 3.0965325001513248e-03
GC_4_68 b_4 NI_4 NS_68 0 1.3051943670992355e-03
GC_4_69 b_4 NI_4 NS_69 0 -2.9261127150177436e-03
GC_4_70 b_4 NI_4 NS_70 0 -9.9123416426922430e-03
GC_4_71 b_4 NI_4 NS_71 0 6.3752755685791160e-04
GC_4_72 b_4 NI_4 NS_72 0 1.3628527547780784e-02
GC_4_73 b_4 NI_4 NS_73 0 1.7509588834278004e-02
GC_4_74 b_4 NI_4 NS_74 0 -2.3852006616147715e-02
GC_4_75 b_4 NI_4 NS_75 0 -3.3177959639940829e-02
GC_4_76 b_4 NI_4 NS_76 0 2.1222695048691349e-02
GC_4_77 b_4 NI_4 NS_77 0 4.0623997774704946e-03
GC_4_78 b_4 NI_4 NS_78 0 -2.1854449406243453e-03
GC_4_79 b_4 NI_4 NS_79 0 1.5119316701147672e-02
GC_4_80 b_4 NI_4 NS_80 0 5.6106547450701112e-03
GC_4_81 b_4 NI_4 NS_81 0 -5.3986446414241388e-04
GC_4_82 b_4 NI_4 NS_82 0 4.9387677195845861e-04
GC_4_83 b_4 NI_4 NS_83 0 -7.8316883412608609e-05
GC_4_84 b_4 NI_4 NS_84 0 9.9479530808034863e-09
GC_4_85 b_4 NI_4 NS_85 0 2.8671032482079601e-10
GC_4_86 b_4 NI_4 NS_86 0 8.0714486955357228e-11
GC_4_87 b_4 NI_4 NS_87 0 -1.2907650857387630e-05
GC_4_88 b_4 NI_4 NS_88 0 -9.1233029760387841e-06
GC_4_89 b_4 NI_4 NS_89 0 -6.7822033339019400e-05
GC_4_90 b_4 NI_4 NS_90 0 -3.2033060854955261e-05
GC_4_91 b_4 NI_4 NS_91 0 -7.1350116730616478e-05
GC_4_92 b_4 NI_4 NS_92 0 1.1519365007894424e-04
GC_4_93 b_4 NI_4 NS_93 0 -1.3882393687989465e-04
GC_4_94 b_4 NI_4 NS_94 0 2.2238771977410978e-04
GC_4_95 b_4 NI_4 NS_95 0 3.5580111242229618e-04
GC_4_96 b_4 NI_4 NS_96 0 1.6517132581635090e-04
GC_4_97 b_4 NI_4 NS_97 0 -1.7001250922303337e-05
GC_4_98 b_4 NI_4 NS_98 0 -1.8454775701678902e-05
GC_4_99 b_4 NI_4 NS_99 0 1.0145602736659403e-04
GC_4_100 b_4 NI_4 NS_100 0 5.6312012311391360e-05
GC_4_101 b_4 NI_4 NS_101 0 1.2462394263345019e-04
GC_4_102 b_4 NI_4 NS_102 0 8.0350031538262536e-05
GC_4_103 b_4 NI_4 NS_103 0 -9.5147267598533788e-05
GC_4_104 b_4 NI_4 NS_104 0 -1.1560845657038583e-07
GC_4_105 b_4 NI_4 NS_105 0 -4.2553955078061321e-10
GC_4_106 b_4 NI_4 NS_106 0 -1.2108016696551860e-10
GC_4_107 b_4 NI_4 NS_107 0 -2.9524917232452643e-05
GC_4_108 b_4 NI_4 NS_108 0 -1.6599768361297139e-05
GC_4_109 b_4 NI_4 NS_109 0 2.8262319577069992e-05
GC_4_110 b_4 NI_4 NS_110 0 9.8567738888713147e-05
GC_4_111 b_4 NI_4 NS_111 0 -6.3018385681517033e-07
GC_4_112 b_4 NI_4 NS_112 0 -1.4684437267063806e-04
GC_4_113 b_4 NI_4 NS_113 0 -1.7067166828734688e-04
GC_4_114 b_4 NI_4 NS_114 0 2.0938949285958299e-04
GC_4_115 b_4 NI_4 NS_115 0 2.7021268006723818e-04
GC_4_116 b_4 NI_4 NS_116 0 -2.1560055771258565e-04
GC_4_117 b_4 NI_4 NS_117 0 -2.5133118527089512e-05
GC_4_118 b_4 NI_4 NS_118 0 2.6862783610684094e-05
GC_4_119 b_4 NI_4 NS_119 0 -1.5209539352302147e-04
GC_4_120 b_4 NI_4 NS_120 0 -6.3894565954001215e-05
GC_4_121 b_4 NI_4 NS_121 0 3.0534162039899817e-04
GC_4_122 b_4 NI_4 NS_122 0 -2.6784547221724502e-04
GC_4_123 b_4 NI_4 NS_123 0 4.2963856605225915e-05
GC_4_124 b_4 NI_4 NS_124 0 1.4101248460641856e-08
GC_4_125 b_4 NI_4 NS_125 0 -1.4707385658245227e-10
GC_4_126 b_4 NI_4 NS_126 0 1.3946538426036530e-11
GC_4_127 b_4 NI_4 NS_127 0 1.6535510295020695e-06
GC_4_128 b_4 NI_4 NS_128 0 7.0335453033696513e-06
GC_4_129 b_4 NI_4 NS_129 0 3.2641608526611874e-05
GC_4_130 b_4 NI_4 NS_130 0 2.1791552444166234e-05
GC_4_131 b_4 NI_4 NS_131 0 4.5841507228432952e-05
GC_4_132 b_4 NI_4 NS_132 0 -5.5994157796701879e-05
GC_4_133 b_4 NI_4 NS_133 0 7.2920974373642656e-05
GC_4_134 b_4 NI_4 NS_134 0 -1.2481942306054086e-04
GC_4_135 b_4 NI_4 NS_135 0 -1.8541708860784489e-04
GC_4_136 b_4 NI_4 NS_136 0 -7.4147696132777460e-05
GC_4_137 b_4 NI_4 NS_137 0 7.6337242892666254e-06
GC_4_138 b_4 NI_4 NS_138 0 3.5085201547275717e-06
GC_4_139 b_4 NI_4 NS_139 0 -5.3960441112190942e-05
GC_4_140 b_4 NI_4 NS_140 0 -3.1131141111296012e-05
GC_4_141 b_4 NI_4 NS_141 0 2.8152218833617780e-04
GC_4_142 b_4 NI_4 NS_142 0 -1.3618967167957612e-05
GC_4_143 b_4 NI_4 NS_143 0 -9.2935602813164918e-06
GC_4_144 b_4 NI_4 NS_144 0 5.9792833077865781e-08
GC_4_145 b_4 NI_4 NS_145 0 -3.0942232913762972e-10
GC_4_146 b_4 NI_4 NS_146 0 9.3377840434860162e-12
GC_4_147 b_4 NI_4 NS_147 0 -7.2720607613426332e-07
GC_4_148 b_4 NI_4 NS_148 0 -1.5722571164572560e-05
GC_4_149 b_4 NI_4 NS_149 0 -9.9778774994439601e-06
GC_4_150 b_4 NI_4 NS_150 0 -2.1078181834483482e-05
GC_4_151 b_4 NI_4 NS_151 0 -3.8198546424459136e-05
GC_4_152 b_4 NI_4 NS_152 0 -1.9856757466134410e-05
GC_4_153 b_4 NI_4 NS_153 0 -7.5906332125097770e-05
GC_4_154 b_4 NI_4 NS_154 0 -7.9824772147423935e-05
GC_4_155 b_4 NI_4 NS_155 0 -7.6276335475169941e-05
GC_4_156 b_4 NI_4 NS_156 0 2.2232889416944272e-04
GC_4_157 b_4 NI_4 NS_157 0 1.5515373754012152e-05
GC_4_158 b_4 NI_4 NS_158 0 -5.7943007459913686e-05
GC_4_159 b_4 NI_4 NS_159 0 -4.8366112664142021e-06
GC_4_160 b_4 NI_4 NS_160 0 1.3913723536885291e-05
GC_4_161 b_4 NI_4 NS_161 0 7.9171040270804091e-06
GC_4_162 b_4 NI_4 NS_162 0 -6.3407566851962175e-06
GC_4_163 b_4 NI_4 NS_163 0 4.7284628722710264e-07
GC_4_164 b_4 NI_4 NS_164 0 6.3751300439348563e-09
GC_4_165 b_4 NI_4 NS_165 0 -1.7572033049102582e-10
GC_4_166 b_4 NI_4 NS_166 0 8.2824454187989839e-12
GC_4_167 b_4 NI_4 NS_167 0 2.1357709466034782e-06
GC_4_168 b_4 NI_4 NS_168 0 -1.0057450614457255e-06
GC_4_169 b_4 NI_4 NS_169 0 2.8511711620749625e-06
GC_4_170 b_4 NI_4 NS_170 0 -1.3362567277647321e-06
GC_4_171 b_4 NI_4 NS_171 0 -2.5357602930850181e-07
GC_4_172 b_4 NI_4 NS_172 0 -3.4595027094696057e-06
GC_4_173 b_4 NI_4 NS_173 0 6.9393796039215547e-06
GC_4_174 b_4 NI_4 NS_174 0 -9.0892538008567099e-06
GC_4_175 b_4 NI_4 NS_175 0 -2.3895809073880413e-05
GC_4_176 b_4 NI_4 NS_176 0 -2.8566943333039529e-06
GC_4_177 b_4 NI_4 NS_177 0 5.9695862446222483e-06
GC_4_178 b_4 NI_4 NS_178 0 3.0591205563942899e-07
GC_4_179 b_4 NI_4 NS_179 0 -2.6278122288018788e-06
GC_4_180 b_4 NI_4 NS_180 0 1.4080032472892418e-06
GC_4_181 b_4 NI_4 NS_181 0 2.2540461907508493e-05
GC_4_182 b_4 NI_4 NS_182 0 -5.1376210386454256e-06
GC_4_183 b_4 NI_4 NS_183 0 3.6838722103469533e-07
GC_4_184 b_4 NI_4 NS_184 0 -8.1493943494085690e-09
GC_4_185 b_4 NI_4 NS_185 0 1.7606410101236766e-10
GC_4_186 b_4 NI_4 NS_186 0 -9.7890773739934753e-12
GC_4_187 b_4 NI_4 NS_187 0 -1.2143346807677555e-06
GC_4_188 b_4 NI_4 NS_188 0 -9.1148481821950527e-07
GC_4_189 b_4 NI_4 NS_189 0 -1.3990076159823766e-06
GC_4_190 b_4 NI_4 NS_190 0 -4.6289000983209950e-08
GC_4_191 b_4 NI_4 NS_191 0 -2.2031483356578035e-06
GC_4_192 b_4 NI_4 NS_192 0 2.3009494322055350e-08
GC_4_193 b_4 NI_4 NS_193 0 -4.7814128481049877e-06
GC_4_194 b_4 NI_4 NS_194 0 -4.5206608511116708e-07
GC_4_195 b_4 NI_4 NS_195 0 1.0105771221302708e-06
GC_4_196 b_4 NI_4 NS_196 0 7.1429857578765478e-06
GC_4_197 b_4 NI_4 NS_197 0 -3.5880414665850058e-07
GC_4_198 b_4 NI_4 NS_198 0 -1.8238538831706607e-06
GC_4_199 b_4 NI_4 NS_199 0 -1.0678623429262091e-06
GC_4_200 b_4 NI_4 NS_200 0 -3.9175125824456833e-07
GC_4_201 b_4 NI_4 NS_201 0 2.0605006317673025e-05
GC_4_202 b_4 NI_4 NS_202 0 -4.9936209244266564e-06
GC_4_203 b_4 NI_4 NS_203 0 9.9303788802134085e-07
GC_4_204 b_4 NI_4 NS_204 0 -5.4984961928680149e-09
GC_4_205 b_4 NI_4 NS_205 0 -2.5967424863202019e-11
GC_4_206 b_4 NI_4 NS_206 0 -1.2308295708744959e-12
GC_4_207 b_4 NI_4 NS_207 0 -1.3115723955874906e-06
GC_4_208 b_4 NI_4 NS_208 0 -1.6746979099244771e-06
GC_4_209 b_4 NI_4 NS_209 0 -1.7990698880008700e-06
GC_4_210 b_4 NI_4 NS_210 0 1.3846236586080762e-07
GC_4_211 b_4 NI_4 NS_211 0 -2.4070676291433273e-06
GC_4_212 b_4 NI_4 NS_212 0 2.2075382729982401e-06
GC_4_213 b_4 NI_4 NS_213 0 -3.9349088550230061e-06
GC_4_214 b_4 NI_4 NS_214 0 -2.1437295806718179e-06
GC_4_215 b_4 NI_4 NS_215 0 1.2290490484578453e-06
GC_4_216 b_4 NI_4 NS_216 0 8.2806508099196448e-06
GC_4_217 b_4 NI_4 NS_217 0 -3.9212457016821423e-07
GC_4_218 b_4 NI_4 NS_218 0 -1.7846417168686507e-06
GC_4_219 b_4 NI_4 NS_219 0 -3.6944483678978371e-07
GC_4_220 b_4 NI_4 NS_220 0 1.7727242837473507e-07
GC_4_221 b_4 NI_4 NS_221 0 5.6551608191214848e-06
GC_4_222 b_4 NI_4 NS_222 0 1.4060288392568065e-06
GC_4_223 b_4 NI_4 NS_223 0 -8.7122201817113258e-07
GC_4_224 b_4 NI_4 NS_224 0 3.5286918648699379e-09
GC_4_225 b_4 NI_4 NS_225 0 5.0023230935341653e-11
GC_4_226 b_4 NI_4 NS_226 0 -5.2267582058699089e-13
GC_4_227 b_4 NI_4 NS_227 0 -4.1810709406951872e-07
GC_4_228 b_4 NI_4 NS_228 0 -3.4338252003625659e-07
GC_4_229 b_4 NI_4 NS_229 0 -2.5300981511186497e-07
GC_4_230 b_4 NI_4 NS_230 0 2.2179392706599256e-07
GC_4_231 b_4 NI_4 NS_231 0 -7.9231991693866990e-07
GC_4_232 b_4 NI_4 NS_232 0 -6.7635775969175156e-07
GC_4_233 b_4 NI_4 NS_233 0 -2.5328282705043950e-06
GC_4_234 b_4 NI_4 NS_234 0 -3.6654012901161399e-08
GC_4_235 b_4 NI_4 NS_235 0 4.1620915142346701e-07
GC_4_236 b_4 NI_4 NS_236 0 3.4991362889921496e-06
GC_4_237 b_4 NI_4 NS_237 0 1.5924466670306977e-07
GC_4_238 b_4 NI_4 NS_238 0 -8.5029830196310475e-07
GC_4_239 b_4 NI_4 NS_239 0 -5.6118828701422422e-07
GC_4_240 b_4 NI_4 NS_240 0 2.6713392431131773e-07
GD_4_1 b_4 NI_4 NA_1 0 2.3474503950476457e-03
GD_4_2 b_4 NI_4 NA_2 0 6.2239313357730624e-03
GD_4_3 b_4 NI_4 NA_3 0 5.6719404092723649e-02
GD_4_4 b_4 NI_4 NA_4 0 -6.3838899589371261e-03
GD_4_5 b_4 NI_4 NA_5 0 -5.1970821850192507e-05
GD_4_6 b_4 NI_4 NA_6 0 7.4679720274325122e-05
GD_4_7 b_4 NI_4 NA_7 0 4.0808617673254657e-06
GD_4_8 b_4 NI_4 NA_8 0 -6.9856716547272529e-05
GD_4_9 b_4 NI_4 NA_9 0 1.1835727161843281e-05
GD_4_10 b_4 NI_4 NA_10 0 -9.6649620829937273e-06
GD_4_11 b_4 NI_4 NA_11 0 -1.0327450105039692e-05
GD_4_12 b_4 NI_4 NA_12 0 -2.2751427490797291e-06
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 2.7270670797563005e-04
GC_5_2 b_5 NI_5 NS_2 0 -1.1383754636797318e-05
GC_5_3 b_5 NI_5 NS_3 0 -9.5559240216873046e-06
GC_5_4 b_5 NI_5 NS_4 0 6.1073863591250994e-08
GC_5_5 b_5 NI_5 NS_5 0 -3.1719513787908478e-10
GC_5_6 b_5 NI_5 NS_6 0 9.0131933735920277e-12
GC_5_7 b_5 NI_5 NS_7 0 -4.9941249024049280e-07
GC_5_8 b_5 NI_5 NS_8 0 -1.5410044213610397e-05
GC_5_9 b_5 NI_5 NS_9 0 -9.6053242000127325e-06
GC_5_10 b_5 NI_5 NS_10 0 -2.0782388655193137e-05
GC_5_11 b_5 NI_5 NS_11 0 -3.7546626554692070e-05
GC_5_12 b_5 NI_5 NS_12 0 -1.9743152723514577e-05
GC_5_13 b_5 NI_5 NS_13 0 -7.4988913056754208e-05
GC_5_14 b_5 NI_5 NS_14 0 -7.8362507652211561e-05
GC_5_15 b_5 NI_5 NS_15 0 -7.3509912901264352e-05
GC_5_16 b_5 NI_5 NS_16 0 2.1939666115101093e-04
GC_5_17 b_5 NI_5 NS_17 0 1.4867517341468921e-05
GC_5_18 b_5 NI_5 NS_18 0 -5.7361994209980343e-05
GC_5_19 b_5 NI_5 NS_19 0 -4.6235339718104136e-06
GC_5_20 b_5 NI_5 NS_20 0 1.3685042702583554e-05
GC_5_21 b_5 NI_5 NS_21 0 3.0050323984163129e-04
GC_5_22 b_5 NI_5 NS_22 0 -2.6759729308189974e-04
GC_5_23 b_5 NI_5 NS_23 0 4.2937843047902083e-05
GC_5_24 b_5 NI_5 NS_24 0 1.3911738157861497e-08
GC_5_25 b_5 NI_5 NS_25 0 -1.4978350942303630e-10
GC_5_26 b_5 NI_5 NS_26 0 1.4933236064041154e-11
GC_5_27 b_5 NI_5 NS_27 0 2.1659410937954281e-06
GC_5_28 b_5 NI_5 NS_28 0 7.3080135403415132e-06
GC_5_29 b_5 NI_5 NS_29 0 3.3345692080145356e-05
GC_5_30 b_5 NI_5 NS_30 0 2.1778354058450670e-05
GC_5_31 b_5 NI_5 NS_31 0 4.6482455857450129e-05
GC_5_32 b_5 NI_5 NS_32 0 -5.6793318483704839e-05
GC_5_33 b_5 NI_5 NS_33 0 7.4769075437913107e-05
GC_5_34 b_5 NI_5 NS_34 0 -1.2484402716658920e-04
GC_5_35 b_5 NI_5 NS_35 0 -1.8751986264623464e-04
GC_5_36 b_5 NI_5 NS_36 0 -7.7199056129450416e-05
GC_5_37 b_5 NI_5 NS_37 0 8.1439073697440651e-06
GC_5_38 b_5 NI_5 NS_38 0 4.1237466902171756e-06
GC_5_39 b_5 NI_5 NS_39 0 -5.4121468831604580e-05
GC_5_40 b_5 NI_5 NS_40 0 -3.1122573981807658e-05
GC_5_41 b_5 NI_5 NS_41 0 1.2462394377981597e-04
GC_5_42 b_5 NI_5 NS_42 0 8.0350030928110389e-05
GC_5_43 b_5 NI_5 NS_43 0 -9.5147267512226809e-05
GC_5_44 b_5 NI_5 NS_44 0 -1.1560845695645489e-07
GC_5_45 b_5 NI_5 NS_45 0 -4.2553954713121286e-10
GC_5_46 b_5 NI_5 NS_46 0 -1.2108016707068797e-10
GC_5_47 b_5 NI_5 NS_47 0 -2.9524917172394866e-05
GC_5_48 b_5 NI_5 NS_48 0 -1.6599768381149253e-05
GC_5_49 b_5 NI_5 NS_49 0 2.8262319654891699e-05
GC_5_50 b_5 NI_5 NS_50 0 9.8567738807564287e-05
GC_5_51 b_5 NI_5 NS_51 0 -6.3018388165699189e-07
GC_5_52 b_5 NI_5 NS_52 0 -1.4684437283425363e-04
GC_5_53 b_5 NI_5 NS_53 0 -1.7067166804607314e-04
GC_5_54 b_5 NI_5 NS_54 0 2.0938949243982368e-04
GC_5_55 b_5 NI_5 NS_55 0 2.7021267887976326e-04
GC_5_56 b_5 NI_5 NS_56 0 -2.1560055766604581e-04
GC_5_57 b_5 NI_5 NS_57 0 -2.5133118233423755e-05
GC_5_58 b_5 NI_5 NS_58 0 2.6862783583407884e-05
GC_5_59 b_5 NI_5 NS_59 0 -1.5209539362190773e-04
GC_5_60 b_5 NI_5 NS_60 0 -6.3894565930140406e-05
GC_5_61 b_5 NI_5 NS_61 0 -5.3979227558290826e-04
GC_5_62 b_5 NI_5 NS_62 0 4.9388521508943292e-04
GC_5_63 b_5 NI_5 NS_63 0 -7.8319138852137450e-05
GC_5_64 b_5 NI_5 NS_64 0 9.9521385198953099e-09
GC_5_65 b_5 NI_5 NS_65 0 2.8669965414866935e-10
GC_5_66 b_5 NI_5 NS_66 0 8.0713872771496091e-11
GC_5_67 b_5 NI_5 NS_67 0 -1.2925624692853075e-05
GC_5_68 b_5 NI_5 NS_68 0 -9.1377574942458015e-06
GC_5_69 b_5 NI_5 NS_69 0 -6.7846976568498025e-05
GC_5_70 b_5 NI_5 NS_70 0 -3.2036623696598602e-05
GC_5_71 b_5 NI_5 NS_71 0 -7.1365955774260861e-05
GC_5_72 b_5 NI_5 NS_72 0 1.1523613583160625e-04
GC_5_73 b_5 NI_5 NS_73 0 -1.3883879523976273e-04
GC_5_74 b_5 NI_5 NS_74 0 2.2241980822483486e-04
GC_5_75 b_5 NI_5 NS_75 0 3.5584092009343461e-04
GC_5_76 b_5 NI_5 NS_76 0 1.6517825811149318e-04
GC_5_77 b_5 NI_5 NS_77 0 -1.7005468321778808e-05
GC_5_78 b_5 NI_5 NS_78 0 -1.8451587801420375e-05
GC_5_79 b_5 NI_5 NS_79 0 1.0145875881539049e-04
GC_5_80 b_5 NI_5 NS_80 0 5.6315095297176582e-05
GC_5_81 b_5 NI_5 NS_81 0 -9.3726655116822951e-04
GC_5_82 b_5 NI_5 NS_82 0 -1.7325122753597964e-02
GC_5_83 b_5 NI_5 NS_83 0 1.1756094123794279e-02
GC_5_84 b_5 NI_5 NS_84 0 2.9426102902452176e-06
GC_5_85 b_5 NI_5 NS_85 0 -5.0962286620962446e-07
GC_5_86 b_5 NI_5 NS_86 0 -2.9668205457973490e-08
GC_5_87 b_5 NI_5 NS_87 0 3.0719126848572859e-03
GC_5_88 b_5 NI_5 NS_88 0 1.2847124259509830e-03
GC_5_89 b_5 NI_5 NS_89 0 -2.9639168272317115e-03
GC_5_90 b_5 NI_5 NS_90 0 -9.9278285614478948e-03
GC_5_91 b_5 NI_5 NS_91 0 5.8579924652858413e-04
GC_5_92 b_5 NI_5 NS_92 0 1.3645080551189272e-02
GC_5_93 b_5 NI_5 NS_93 0 1.7411063181380474e-02
GC_5_94 b_5 NI_5 NS_94 0 -2.3905073452168128e-02
GC_5_95 b_5 NI_5 NS_95 0 -3.3221885726839026e-02
GC_5_96 b_5 NI_5 NS_96 0 2.1449490462518022e-02
GC_5_97 b_5 NI_5 NS_97 0 4.0698736023087939e-03
GC_5_98 b_5 NI_5 NS_98 0 -2.2340707647231497e-03
GC_5_99 b_5 NI_5 NS_99 0 1.5117890334129035e-02
GC_5_100 b_5 NI_5 NS_100 0 5.6202762008539953e-03
GC_5_101 b_5 NI_5 NS_101 0 -2.8556594911078675e-01
GC_5_102 b_5 NI_5 NS_102 0 1.2097574679039476e-01
GC_5_103 b_5 NI_5 NS_103 0 7.0770605070180721e-03
GC_5_104 b_5 NI_5 NS_104 0 5.7565193887564934e-05
GC_5_105 b_5 NI_5 NS_105 0 1.2985822547435219e-06
GC_5_106 b_5 NI_5 NS_106 0 1.4018750273668521e-08
GC_5_107 b_5 NI_5 NS_107 0 3.0464941337271473e-02
GC_5_108 b_5 NI_5 NS_108 0 4.1070459849588230e-03
GC_5_109 b_5 NI_5 NS_109 0 -7.3803888565569303e-03
GC_5_110 b_5 NI_5 NS_110 0 2.2172609358355092e-02
GC_5_111 b_5 NI_5 NS_111 0 -1.7062230455883492e-02
GC_5_112 b_5 NI_5 NS_112 0 -1.8682680320462126e-02
GC_5_113 b_5 NI_5 NS_113 0 4.4646617493442432e-02
GC_5_114 b_5 NI_5 NS_114 0 1.4294514024690851e-02
GC_5_115 b_5 NI_5 NS_115 0 8.1981868478833764e-02
GC_5_116 b_5 NI_5 NS_116 0 3.1414612583227232e-02
GC_5_117 b_5 NI_5 NS_117 0 -1.0082921128176686e-02
GC_5_118 b_5 NI_5 NS_118 0 -4.9140409030850162e-03
GC_5_119 b_5 NI_5 NS_119 0 -2.1489484228921996e-02
GC_5_120 b_5 NI_5 NS_120 0 -4.8797257350585181e-03
GC_5_121 b_5 NI_5 NS_121 0 2.2333485084293267e-02
GC_5_122 b_5 NI_5 NS_122 0 8.9184338921983446e-03
GC_5_123 b_5 NI_5 NS_123 0 -1.1401600408274900e-02
GC_5_124 b_5 NI_5 NS_124 0 -5.3823441502445202e-06
GC_5_125 b_5 NI_5 NS_125 0 -9.5308344342130914e-08
GC_5_126 b_5 NI_5 NS_126 0 -1.2685911015156329e-09
GC_5_127 b_5 NI_5 NS_127 0 -3.3183157155340405e-03
GC_5_128 b_5 NI_5 NS_128 0 -2.3921302575102021e-03
GC_5_129 b_5 NI_5 NS_129 0 2.7239195453364132e-03
GC_5_130 b_5 NI_5 NS_130 0 1.1169875325987040e-02
GC_5_131 b_5 NI_5 NS_131 0 -3.6330705414727683e-04
GC_5_132 b_5 NI_5 NS_132 0 -1.7752735332879431e-02
GC_5_133 b_5 NI_5 NS_133 0 -2.2016949437053776e-02
GC_5_134 b_5 NI_5 NS_134 0 2.1338989327258532e-02
GC_5_135 b_5 NI_5 NS_135 0 2.8916848613792966e-02
GC_5_136 b_5 NI_5 NS_136 0 -1.8399470310471837e-02
GC_5_137 b_5 NI_5 NS_137 0 -2.4531764736285761e-03
GC_5_138 b_5 NI_5 NS_138 0 1.4162712460930379e-03
GC_5_139 b_5 NI_5 NS_139 0 -1.7821660735131032e-02
GC_5_140 b_5 NI_5 NS_140 0 -7.1344518915960791e-03
GC_5_141 b_5 NI_5 NS_141 0 -8.2237001688338987e-02
GC_5_142 b_5 NI_5 NS_142 0 6.5305852816874177e-02
GC_5_143 b_5 NI_5 NS_143 0 -1.0305226885530833e-02
GC_5_144 b_5 NI_5 NS_144 0 -2.4029859711971136e-06
GC_5_145 b_5 NI_5 NS_145 0 1.6307886669065151e-08
GC_5_146 b_5 NI_5 NS_146 0 1.6568107851290218e-09
GC_5_147 b_5 NI_5 NS_147 0 -3.9692405239336942e-04
GC_5_148 b_5 NI_5 NS_148 0 -1.4031043331831363e-03
GC_5_149 b_5 NI_5 NS_149 0 -6.9955150578639453e-03
GC_5_150 b_5 NI_5 NS_150 0 -3.7827359493684885e-03
GC_5_151 b_5 NI_5 NS_151 0 -9.0599083973671637e-03
GC_5_152 b_5 NI_5 NS_152 0 1.3124883429509761e-02
GC_5_153 b_5 NI_5 NS_153 0 -1.5228217954426668e-02
GC_5_154 b_5 NI_5 NS_154 0 2.8706591444776785e-02
GC_5_155 b_5 NI_5 NS_155 0 4.5065279289461080e-02
GC_5_156 b_5 NI_5 NS_156 0 1.6496171682930879e-02
GC_5_157 b_5 NI_5 NS_157 0 -2.1949566512916526e-03
GC_5_158 b_5 NI_5 NS_158 0 -1.3428667030015782e-03
GC_5_159 b_5 NI_5 NS_159 0 1.2861366874249044e-02
GC_5_160 b_5 NI_5 NS_160 0 6.9592344555460574e-03
GC_5_161 b_5 NI_5 NS_161 0 2.7705412667916167e-04
GC_5_162 b_5 NI_5 NS_162 0 -1.2387381301197637e-05
GC_5_163 b_5 NI_5 NS_163 0 -9.4633644382173773e-06
GC_5_164 b_5 NI_5 NS_164 0 6.0728928977705360e-08
GC_5_165 b_5 NI_5 NS_165 0 -3.1805478171541015e-10
GC_5_166 b_5 NI_5 NS_166 0 9.7939353399745333e-12
GC_5_167 b_5 NI_5 NS_167 0 -5.8027995776733224e-07
GC_5_168 b_5 NI_5 NS_168 0 -1.5576453642976063e-05
GC_5_169 b_5 NI_5 NS_169 0 -9.7465693579262124e-06
GC_5_170 b_5 NI_5 NS_170 0 -2.0953109029566185e-05
GC_5_171 b_5 NI_5 NS_171 0 -3.7868615402687072e-05
GC_5_172 b_5 NI_5 NS_172 0 -1.9889341243796711e-05
GC_5_173 b_5 NI_5 NS_173 0 -7.5415010402439579e-05
GC_5_174 b_5 NI_5 NS_174 0 -7.9253549225928376e-05
GC_5_175 b_5 NI_5 NS_175 0 -7.5278067513166220e-05
GC_5_176 b_5 NI_5 NS_176 0 2.2097702677586977e-04
GC_5_177 b_5 NI_5 NS_177 0 1.5306009389452864e-05
GC_5_178 b_5 NI_5 NS_178 0 -5.7665549259534716e-05
GC_5_179 b_5 NI_5 NS_179 0 -4.7284458551073584e-06
GC_5_180 b_5 NI_5 NS_180 0 1.3857052575360210e-05
GC_5_181 b_5 NI_5 NS_181 0 3.0487060207122312e-04
GC_5_182 b_5 NI_5 NS_182 0 -2.6795564136938686e-04
GC_5_183 b_5 NI_5 NS_183 0 4.3029677725815956e-05
GC_5_184 b_5 NI_5 NS_184 0 1.3275143603432587e-08
GC_5_185 b_5 NI_5 NS_185 0 -1.3642185380248016e-10
GC_5_186 b_5 NI_5 NS_186 0 1.3413643033037057e-11
GC_5_187 b_5 NI_5 NS_187 0 1.6673087928350513e-06
GC_5_188 b_5 NI_5 NS_188 0 7.0536131999090906e-06
GC_5_189 b_5 NI_5 NS_189 0 3.2663687574631964e-05
GC_5_190 b_5 NI_5 NS_190 0 2.1834068071842076e-05
GC_5_191 b_5 NI_5 NS_191 0 4.5895161509100195e-05
GC_5_192 b_5 NI_5 NS_192 0 -5.6019838278533292e-05
GC_5_193 b_5 NI_5 NS_193 0 7.3005720024375622e-05
GC_5_194 b_5 NI_5 NS_194 0 -1.2465455937387245e-04
GC_5_195 b_5 NI_5 NS_195 0 -1.8515939577169331e-04
GC_5_196 b_5 NI_5 NS_196 0 -7.4482522558536342e-05
GC_5_197 b_5 NI_5 NS_197 0 7.5437637602545312e-06
GC_5_198 b_5 NI_5 NS_198 0 3.5788428385373756e-06
GC_5_199 b_5 NI_5 NS_199 0 -5.3931892107295272e-05
GC_5_200 b_5 NI_5 NS_200 0 -3.1184819980291598e-05
GC_5_201 b_5 NI_5 NS_201 0 -7.8386262692553899e-05
GC_5_202 b_5 NI_5 NS_202 0 1.3378293575870036e-05
GC_5_203 b_5 NI_5 NS_203 0 -1.3936000038697851e-06
GC_5_204 b_5 NI_5 NS_204 0 -1.3100500970503667e-08
GC_5_205 b_5 NI_5 NS_205 0 2.6340787395270520e-10
GC_5_206 b_5 NI_5 NS_206 0 -1.7096275821107206e-11
GC_5_207 b_5 NI_5 NS_207 0 -1.5341826743089738e-06
GC_5_208 b_5 NI_5 NS_208 0 3.6435271319800677e-06
GC_5_209 b_5 NI_5 NS_209 0 1.6179623081688881e-06
GC_5_210 b_5 NI_5 NS_210 0 8.9335050018294747e-06
GC_5_211 b_5 NI_5 NS_211 0 1.0126601569764030e-05
GC_5_212 b_5 NI_5 NS_212 0 3.9283519260325954e-06
GC_5_213 b_5 NI_5 NS_213 0 1.3024106484684229e-05
GC_5_214 b_5 NI_5 NS_214 0 2.9985525556983375e-05
GC_5_215 b_5 NI_5 NS_215 0 3.6902719855553611e-05
GC_5_216 b_5 NI_5 NS_216 0 -6.0917486571398373e-05
GC_5_217 b_5 NI_5 NS_217 0 -6.8806255581356324e-06
GC_5_218 b_5 NI_5 NS_218 0 1.5060253515729353e-05
GC_5_219 b_5 NI_5 NS_219 0 -1.5080846923272749e-06
GC_5_220 b_5 NI_5 NS_220 0 -4.9189622593664072e-06
GC_5_221 b_5 NI_5 NS_221 0 6.1496279003032939e-05
GC_5_222 b_5 NI_5 NS_222 0 -4.0968511513297937e-05
GC_5_223 b_5 NI_5 NS_223 0 7.0419747230294941e-06
GC_5_224 b_5 NI_5 NS_224 0 -1.5383551171581694e-08
GC_5_225 b_5 NI_5 NS_225 0 -2.8243287262267063e-11
GC_5_226 b_5 NI_5 NS_226 0 2.8286463984862836e-13
GC_5_227 b_5 NI_5 NS_227 0 -9.0513692188917243e-07
GC_5_228 b_5 NI_5 NS_228 0 -1.4038336501479816e-06
GC_5_229 b_5 NI_5 NS_229 0 1.3494591296112959e-06
GC_5_230 b_5 NI_5 NS_230 0 2.2662979758648903e-06
GC_5_231 b_5 NI_5 NS_231 0 2.9358435737974158e-06
GC_5_232 b_5 NI_5 NS_232 0 -3.4739240968756017e-06
GC_5_233 b_5 NI_5 NS_233 0 7.8879427214495532e-06
GC_5_234 b_5 NI_5 NS_234 0 -1.6508173944916280e-05
GC_5_235 b_5 NI_5 NS_235 0 -2.6704649221956404e-05
GC_5_236 b_5 NI_5 NS_236 0 -4.5356303941220136e-06
GC_5_237 b_5 NI_5 NS_237 0 2.5910949144379550e-06
GC_5_238 b_5 NI_5 NS_238 0 -5.5008349315717848e-07
GC_5_239 b_5 NI_5 NS_239 0 -7.0849925880063254e-06
GC_5_240 b_5 NI_5 NS_240 0 -3.6888956188645406e-06
GD_5_1 b_5 NI_5 NA_1 0 -6.6955532767880280e-05
GD_5_2 b_5 NI_5 NA_2 0 7.8745438886619517e-06
GD_5_3 b_5 NI_5 NA_3 0 7.4679720387294584e-05
GD_5_4 b_5 NI_5 NA_4 0 -5.2020155077352970e-05
GD_5_5 b_5 NI_5 NA_5 0 -6.6185230473112594e-03
GD_5_6 b_5 NI_5 NA_6 0 5.6693614557915474e-02
GD_5_7 b_5 NI_5 NA_7 0 6.1947474638149600e-03
GD_5_8 b_5 NI_5 NA_8 0 2.3344520445871824e-03
GD_5_9 b_5 NI_5 NA_9 0 -6.8166037211890901e-05
GD_5_10 b_5 NI_5 NA_10 0 4.2508828557616228e-06
GD_5_11 b_5 NI_5 NA_11 0 1.5819161345759031e-05
GD_5_12 b_5 NI_5 NA_12 0 -8.9720782546948026e-06
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 3.0050542332200902e-04
GC_6_2 b_6 NI_6 NS_2 0 -2.6759720626367054e-04
GC_6_3 b_6 NI_6 NS_3 0 4.2937784011652582e-05
GC_6_4 b_6 NI_6 NS_4 0 1.3912054823751590e-08
GC_6_5 b_6 NI_6 NS_5 0 -1.4978819691118667e-10
GC_6_6 b_6 NI_6 NS_6 0 1.4933411280037539e-11
GC_6_7 b_6 NI_6 NS_7 0 2.1661615913595026e-06
GC_6_8 b_6 NI_6 NS_8 0 7.3079535578510260e-06
GC_6_9 b_6 NI_6 NS_9 0 3.3345900355513662e-05
GC_6_10 b_6 NI_6 NS_10 0 2.1777979889757573e-05
GC_6_11 b_6 NI_6 NS_11 0 4.6481490404613095e-05
GC_6_12 b_6 NI_6 NS_12 0 -5.6794137122474107e-05
GC_6_13 b_6 NI_6 NS_13 0 7.4766882143051459e-05
GC_6_14 b_6 NI_6 NS_14 0 -1.2484470014994923e-04
GC_6_15 b_6 NI_6 NS_15 0 -1.8751805452203046e-04
GC_6_16 b_6 NI_6 NS_16 0 -7.7196109448434512e-05
GC_6_17 b_6 NI_6 NS_17 0 8.1430446200182293e-06
GC_6_18 b_6 NI_6 NS_18 0 4.1233495227007976e-06
GC_6_19 b_6 NI_6 NS_19 0 -5.4121375150576740e-05
GC_6_20 b_6 NI_6 NS_20 0 -3.1122467319710209e-05
GC_6_21 b_6 NI_6 NS_21 0 2.7174115870622772e-04
GC_6_22 b_6 NI_6 NS_22 0 -1.1194127265913965e-05
GC_6_23 b_6 NI_6 NS_23 0 -9.5765068857577642e-06
GC_6_24 b_6 NI_6 NS_24 0 6.1170047781967896e-08
GC_6_25 b_6 NI_6 NS_25 0 -3.1755796488761146e-10
GC_6_26 b_6 NI_6 NS_26 0 9.0305706826264186e-12
GC_6_27 b_6 NI_6 NS_27 0 -4.6037800875030610e-07
GC_6_28 b_6 NI_6 NS_28 0 -1.5384218992790987e-05
GC_6_29 b_6 NI_6 NS_29 0 -9.5047719747768658e-06
GC_6_30 b_6 NI_6 NS_30 0 -2.0753489848541591e-05
GC_6_31 b_6 NI_6 NS_31 0 -3.7497052582706334e-05
GC_6_32 b_6 NI_6 NS_32 0 -1.9825266018949670e-05
GC_6_33 b_6 NI_6 NS_33 0 -7.4897115485665462e-05
GC_6_34 b_6 NI_6 NS_34 0 -7.8245278584966016e-05
GC_6_35 b_6 NI_6 NS_35 0 -7.3342906625140620e-05
GC_6_36 b_6 NI_6 NS_36 0 2.1906424141363286e-04
GC_6_37 b_6 NI_6 NS_37 0 1.4840686656832197e-05
GC_6_38 b_6 NI_6 NS_38 0 -5.7290357298156104e-05
GC_6_39 b_6 NI_6 NS_39 0 -4.6091055710131058e-06
GC_6_40 b_6 NI_6 NS_40 0 1.3659348404213419e-05
GC_6_41 b_6 NI_6 NS_41 0 -5.3986446151776956e-04
GC_6_42 b_6 NI_6 NS_42 0 4.9387677187228145e-04
GC_6_43 b_6 NI_6 NS_43 0 -7.8316883411938193e-05
GC_6_44 b_6 NI_6 NS_44 0 9.9479530017795474e-09
GC_6_45 b_6 NI_6 NS_45 0 2.8671033684364877e-10
GC_6_46 b_6 NI_6 NS_46 0 8.0714484690985882e-11
GC_6_47 b_6 NI_6 NS_47 0 -1.2907650969491363e-05
GC_6_48 b_6 NI_6 NS_48 0 -9.1233033379930912e-06
GC_6_49 b_6 NI_6 NS_49 0 -6.7822033930036178e-05
GC_6_50 b_6 NI_6 NS_50 0 -3.2033061170606547e-05
GC_6_51 b_6 NI_6 NS_51 0 -7.1350117376576448e-05
GC_6_52 b_6 NI_6 NS_52 0 1.1519365052430621e-04
GC_6_53 b_6 NI_6 NS_53 0 -1.3882393824788563e-04
GC_6_54 b_6 NI_6 NS_54 0 2.2238771992412164e-04
GC_6_55 b_6 NI_6 NS_55 0 3.5580111399265938e-04
GC_6_56 b_6 NI_6 NS_56 0 1.6517132775501698e-04
GC_6_57 b_6 NI_6 NS_57 0 -1.7001251401868709e-05
GC_6_58 b_6 NI_6 NS_58 0 -1.8454776073749034e-05
GC_6_59 b_6 NI_6 NS_59 0 1.0145602746692786e-04
GC_6_60 b_6 NI_6 NS_60 0 5.6312012330663446e-05
GC_6_61 b_6 NI_6 NS_61 0 1.2460296003865301e-04
GC_6_62 b_6 NI_6 NS_62 0 8.0357129809888821e-05
GC_6_63 b_6 NI_6 NS_63 0 -9.5148169915632431e-05
GC_6_64 b_6 NI_6 NS_64 0 -1.1560586074313003e-07
GC_6_65 b_6 NI_6 NS_65 0 -4.2556430304141940e-10
GC_6_66 b_6 NI_6 NS_66 0 -1.2107894005194887e-10
GC_6_67 b_6 NI_6 NS_67 0 -2.9524729649007298e-05
GC_6_68 b_6 NI_6 NS_68 0 -1.6598751326236156e-05
GC_6_69 b_6 NI_6 NS_69 0 2.8263593289345197e-05
GC_6_70 b_6 NI_6 NS_70 0 9.8568706517968176e-05
GC_6_71 b_6 NI_6 NS_71 0 -6.2941201967303707e-07
GC_6_72 b_6 NI_6 NS_72 0 -1.4684426135867090e-04
GC_6_73 b_6 NI_6 NS_73 0 -1.7067067318769964e-04
GC_6_74 b_6 NI_6 NS_74 0 2.0939417391088882e-04
GC_6_75 b_6 NI_6 NS_75 0 2.7022139264303317e-04
GC_6_76 b_6 NI_6 NS_76 0 -2.1560536323909777e-04
GC_6_77 b_6 NI_6 NS_77 0 -2.5134850157550668e-05
GC_6_78 b_6 NI_6 NS_78 0 2.6863414352312928e-05
GC_6_79 b_6 NI_6 NS_79 0 -1.5209446864317139e-04
GC_6_80 b_6 NI_6 NS_80 0 -6.3894955636233959e-05
GC_6_81 b_6 NI_6 NS_81 0 -2.8556595864610695e-01
GC_6_82 b_6 NI_6 NS_82 0 1.2097574617388222e-01
GC_6_83 b_6 NI_6 NS_83 0 7.0770606811213438e-03
GC_6_84 b_6 NI_6 NS_84 0 5.7565192861024468e-05
GC_6_85 b_6 NI_6 NS_85 0 1.2985822761262931e-06
GC_6_86 b_6 NI_6 NS_86 0 1.4018748554634769e-08
GC_6_87 b_6 NI_6 NS_87 0 3.0464942094306155e-02
GC_6_88 b_6 NI_6 NS_88 0 4.1070473709543592e-03
GC_6_89 b_6 NI_6 NS_89 0 -7.3803861754361821e-03
GC_6_90 b_6 NI_6 NS_90 0 2.2172610619047038e-02
GC_6_91 b_6 NI_6 NS_91 0 -1.7062227553409953e-02
GC_6_92 b_6 NI_6 NS_92 0 -1.8682682946140321e-02
GC_6_93 b_6 NI_6 NS_93 0 4.4646623065784104e-02
GC_6_94 b_6 NI_6 NS_94 0 1.4294511526699841e-02
GC_6_95 b_6 NI_6 NS_95 0 8.1981860142589721e-02
GC_6_96 b_6 NI_6 NS_96 0 3.1414606586404346e-02
GC_6_97 b_6 NI_6 NS_97 0 -1.0082918955962505e-02
GC_6_98 b_6 NI_6 NS_98 0 -4.9140400519538732e-03
GC_6_99 b_6 NI_6 NS_99 0 -2.1489484713166206e-02
GC_6_100 b_6 NI_6 NS_100 0 -4.8797258277443103e-03
GC_6_101 b_6 NI_6 NS_101 0 -9.3726655116826096e-04
GC_6_102 b_6 NI_6 NS_102 0 -1.7325122753597929e-02
GC_6_103 b_6 NI_6 NS_103 0 1.1756094123794256e-02
GC_6_104 b_6 NI_6 NS_104 0 2.9426102902458414e-06
GC_6_105 b_6 NI_6 NS_105 0 -5.0962286620964881e-07
GC_6_106 b_6 NI_6 NS_106 0 -2.9668205457972788e-08
GC_6_107 b_6 NI_6 NS_107 0 3.0719126848572924e-03
GC_6_108 b_6 NI_6 NS_108 0 1.2847124259509793e-03
GC_6_109 b_6 NI_6 NS_109 0 -2.9639168272317042e-03
GC_6_110 b_6 NI_6 NS_110 0 -9.9278285614479017e-03
GC_6_111 b_6 NI_6 NS_111 0 5.8579924652857297e-04
GC_6_112 b_6 NI_6 NS_112 0 1.3645080551189263e-02
GC_6_113 b_6 NI_6 NS_113 0 1.7411063181380471e-02
GC_6_114 b_6 NI_6 NS_114 0 -2.3905073452168128e-02
GC_6_115 b_6 NI_6 NS_115 0 -3.3221885726838991e-02
GC_6_116 b_6 NI_6 NS_116 0 2.1449490462518012e-02
GC_6_117 b_6 NI_6 NS_117 0 4.0698736023087757e-03
GC_6_118 b_6 NI_6 NS_118 0 -2.2340707647231462e-03
GC_6_119 b_6 NI_6 NS_119 0 1.5117890334129028e-02
GC_6_120 b_6 NI_6 NS_120 0 5.6202762008539945e-03
GC_6_121 b_6 NI_6 NS_121 0 -8.2237002142653018e-02
GC_6_122 b_6 NI_6 NS_122 0 6.5305853068506198e-02
GC_6_123 b_6 NI_6 NS_123 0 -1.0305226917751733e-02
GC_6_124 b_6 NI_6 NS_124 0 -2.4029859112384393e-06
GC_6_125 b_6 NI_6 NS_125 0 1.6307886450570868e-08
GC_6_126 b_6 NI_6 NS_126 0 1.6568107762406657e-09
GC_6_127 b_6 NI_6 NS_127 0 -3.9692419139674442e-04
GC_6_128 b_6 NI_6 NS_128 0 -1.4031044037180322e-03
GC_6_129 b_6 NI_6 NS_129 0 -6.9955152485385282e-03
GC_6_130 b_6 NI_6 NS_130 0 -3.7827359195603148e-03
GC_6_131 b_6 NI_6 NS_131 0 -9.0599084283642002e-03
GC_6_132 b_6 NI_6 NS_132 0 1.3124883864152280e-02
GC_6_133 b_6 NI_6 NS_133 0 -1.5228217849689887e-02
GC_6_134 b_6 NI_6 NS_134 0 2.8706592104651863e-02
GC_6_135 b_6 NI_6 NS_135 0 4.5065279965253210e-02
GC_6_136 b_6 NI_6 NS_136 0 1.6496170898854124e-02
GC_6_137 b_6 NI_6 NS_137 0 -2.1949567267126277e-03
GC_6_138 b_6 NI_6 NS_138 0 -1.3428664568818822e-03
GC_6_139 b_6 NI_6 NS_139 0 1.2861366894724339e-02
GC_6_140 b_6 NI_6 NS_140 0 6.9592344379893799e-03
GC_6_141 b_6 NI_6 NS_141 0 2.2333485082340402e-02
GC_6_142 b_6 NI_6 NS_142 0 8.9184338894236527e-03
GC_6_143 b_6 NI_6 NS_143 0 -1.1401600407329293e-02
GC_6_144 b_6 NI_6 NS_144 0 -5.3823441542968173e-06
GC_6_145 b_6 NI_6 NS_145 0 -9.5308344304806182e-08
GC_6_146 b_6 NI_6 NS_146 0 -1.2685910996484772e-09
GC_6_147 b_6 NI_6 NS_147 0 -3.3183157151447829e-03
GC_6_148 b_6 NI_6 NS_148 0 -2.3921302584309300e-03
GC_6_149 b_6 NI_6 NS_149 0 2.7239195437716822e-03
GC_6_150 b_6 NI_6 NS_150 0 1.1169875324060987e-02
GC_6_151 b_6 NI_6 NS_151 0 -3.6330705741110289e-04
GC_6_152 b_6 NI_6 NS_152 0 -1.7752735330577137e-02
GC_6_153 b_6 NI_6 NS_153 0 -2.2016949442888688e-02
GC_6_154 b_6 NI_6 NS_154 0 2.1338989335300450e-02
GC_6_155 b_6 NI_6 NS_155 0 2.8916848633880460e-02
GC_6_156 b_6 NI_6 NS_156 0 -1.8399470316659484e-02
GC_6_157 b_6 NI_6 NS_157 0 -2.4531764794582861e-03
GC_6_158 b_6 NI_6 NS_158 0 1.4162712486315164e-03
GC_6_159 b_6 NI_6 NS_159 0 -1.7821660735425404e-02
GC_6_160 b_6 NI_6 NS_160 0 -7.1344518936834874e-03
GC_6_161 b_6 NI_6 NS_161 0 3.0487036770151100e-04
GC_6_162 b_6 NI_6 NS_162 0 -2.6795571908672241e-04
GC_6_163 b_6 NI_6 NS_163 0 4.3029734422070946e-05
GC_6_164 b_6 NI_6 NS_164 0 1.3274605055770553e-08
GC_6_165 b_6 NI_6 NS_165 0 -1.3641658921538358e-10
GC_6_166 b_6 NI_6 NS_166 0 1.3413397197807212e-11
GC_6_167 b_6 NI_6 NS_167 0 1.6671640463830022e-06
GC_6_168 b_6 NI_6 NS_168 0 7.0535563348925194e-06
GC_6_169 b_6 NI_6 NS_169 0 3.2663510605685353e-05
GC_6_170 b_6 NI_6 NS_170 0 2.1834099265482967e-05
GC_6_171 b_6 NI_6 NS_171 0 4.5895159242491996e-05
GC_6_172 b_6 NI_6 NS_172 0 -5.6019428514834158e-05
GC_6_173 b_6 NI_6 NS_173 0 7.3005783978062356e-05
GC_6_174 b_6 NI_6 NS_174 0 -1.2465398889318724e-04
GC_6_175 b_6 NI_6 NS_175 0 -1.8515862198182923e-04
GC_6_176 b_6 NI_6 NS_176 0 -7.4483192202616410e-05
GC_6_177 b_6 NI_6 NS_177 0 7.5436292806076263e-06
GC_6_178 b_6 NI_6 NS_178 0 3.5790292340666843e-06
GC_6_179 b_6 NI_6 NS_179 0 -5.3931860686000954e-05
GC_6_180 b_6 NI_6 NS_180 0 -3.1184917819956529e-05
GC_6_181 b_6 NI_6 NS_181 0 2.7806787001742069e-04
GC_6_182 b_6 NI_6 NS_182 0 -1.2586345330828274e-05
GC_6_183 b_6 NI_6 NS_183 0 -9.4421655146635851e-06
GC_6_184 b_6 NI_6 NS_184 0 6.0630184616777390e-08
GC_6_185 b_6 NI_6 NS_185 0 -3.1771024454991478e-10
GC_6_186 b_6 NI_6 NS_186 0 9.7760244483526859e-12
GC_6_187 b_6 NI_6 NS_187 0 -6.2007907334757023e-07
GC_6_188 b_6 NI_6 NS_188 0 -1.5605308658945998e-05
GC_6_189 b_6 NI_6 NS_189 0 -9.8498685523339603e-06
GC_6_190 b_6 NI_6 NS_190 0 -2.0984727328939275e-05
GC_6_191 b_6 NI_6 NS_191 0 -3.7922143310376194e-05
GC_6_192 b_6 NI_6 NS_192 0 -1.9808608600866335e-05
GC_6_193 b_6 NI_6 NS_193 0 -7.5514369264105888e-05
GC_6_194 b_6 NI_6 NS_194 0 -7.9383282830217778e-05
GC_6_195 b_6 NI_6 NS_195 0 -7.5463293764268627e-05
GC_6_196 b_6 NI_6 NS_196 0 2.2133252111202644e-04
GC_6_197 b_6 NI_6 NS_197 0 1.5336579749990457e-05
GC_6_198 b_6 NI_6 NS_198 0 -5.7741341319775823e-05
GC_6_199 b_6 NI_6 NS_199 0 -4.7436873600306193e-06
GC_6_200 b_6 NI_6 NS_200 0 1.3885238299127374e-05
GC_6_201 b_6 NI_6 NS_201 0 6.1561232277284540e-05
GC_6_202 b_6 NI_6 NS_202 0 -4.0958851327243106e-05
GC_6_203 b_6 NI_6 NS_203 0 7.0396238552834453e-06
GC_6_204 b_6 NI_6 NS_204 0 -1.5378936863652846e-08
GC_6_205 b_6 NI_6 NS_205 0 -2.8245685399940692e-11
GC_6_206 b_6 NI_6 NS_206 0 2.8279517224295048e-13
GC_6_207 b_6 NI_6 NS_207 0 -9.2347572534945145e-07
GC_6_208 b_6 NI_6 NS_208 0 -1.4177402006611045e-06
GC_6_209 b_6 NI_6 NS_209 0 1.3243137868398770e-06
GC_6_210 b_6 NI_6 NS_210 0 2.2639607768106032e-06
GC_6_211 b_6 NI_6 NS_211 0 2.9219974031308718e-06
GC_6_212 b_6 NI_6 NS_212 0 -3.4302900310771816e-06
GC_6_213 b_6 NI_6 NS_213 0 7.8764337499714824e-06
GC_6_214 b_6 NI_6 NS_214 0 -1.6473451794091647e-05
GC_6_215 b_6 NI_6 NS_215 0 -2.6664824238541586e-05
GC_6_216 b_6 NI_6 NS_216 0 -4.5354760301102486e-06
GC_6_217 b_6 NI_6 NS_217 0 2.5875752919255341e-06
GC_6_218 b_6 NI_6 NS_218 0 -5.4559823784414740e-07
GC_6_219 b_6 NI_6 NS_219 0 -7.0823181496860345e-06
GC_6_220 b_6 NI_6 NS_220 0 -3.6861006324849771e-06
GC_6_221 b_6 NI_6 NS_221 0 -7.8387633646845409e-05
GC_6_222 b_6 NI_6 NS_222 0 1.3376513925100590e-05
GC_6_223 b_6 NI_6 NS_223 0 -1.3932390723009537e-06
GC_6_224 b_6 NI_6 NS_224 0 -1.3101589273503809e-08
GC_6_225 b_6 NI_6 NS_225 0 2.6342333048867608e-10
GC_6_226 b_6 NI_6 NS_226 0 -1.7097214040876024e-11
GC_6_227 b_6 NI_6 NS_227 0 -1.5337478874633816e-06
GC_6_228 b_6 NI_6 NS_228 0 3.6436027986629095e-06
GC_6_229 b_6 NI_6 NS_229 0 1.6182179111486819e-06
GC_6_230 b_6 NI_6 NS_230 0 8.9333690473558351e-06
GC_6_231 b_6 NI_6 NS_231 0 1.0127223109284448e-05
GC_6_232 b_6 NI_6 NS_232 0 3.9280734808743202e-06
GC_6_233 b_6 NI_6 NS_233 0 1.3025656671164421e-05
GC_6_234 b_6 NI_6 NS_234 0 2.9985128935436111e-05
GC_6_235 b_6 NI_6 NS_235 0 3.6900818450398162e-05
GC_6_236 b_6 NI_6 NS_236 0 -6.0920660399038548e-05
GC_6_237 b_6 NI_6 NS_237 0 -6.8802554862126541e-06
GC_6_238 b_6 NI_6 NS_238 0 1.5061063942818654e-05
GC_6_239 b_6 NI_6 NS_239 0 -1.5084569558250485e-06
GC_6_240 b_6 NI_6 NS_240 0 -4.9192660630591973e-06
GD_6_1 b_6 NI_6 NA_1 0 7.8739698181100837e-06
GD_6_2 b_6 NI_6 NA_2 0 -6.6464568425211434e-05
GD_6_3 b_6 NI_6 NA_3 0 -5.1970822980635143e-05
GD_6_4 b_6 NI_6 NA_4 0 7.4682395307145973e-05
GD_6_5 b_6 NI_6 NA_5 0 5.6693619931360156e-02
GD_6_6 b_6 NI_6 NA_6 0 -6.6185230473112732e-03
GD_6_7 b_6 NI_6 NA_7 0 2.3344518749601269e-03
GD_6_8 b_6 NI_6 NA_8 0 6.1947474642983355e-03
GD_6_9 b_6 NI_6 NA_9 0 4.2506850972205058e-06
GD_6_10 b_6 NI_6 NA_10 0 -6.8663486095372169e-05
GD_6_11 b_6 NI_6 NA_11 0 -9.0215006098939255e-06
GD_6_12 b_6 NI_6 NA_12 0 1.5822121407145430e-05
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 -8.6883716774969715e-05
GC_7_2 b_7 NI_7 NS_2 0 1.4652652382011632e-05
GC_7_3 b_7 NI_7 NS_3 0 -1.4888053907279354e-06
GC_7_4 b_7 NI_7 NS_4 0 -1.2740379673556924e-08
GC_7_5 b_7 NI_7 NS_5 0 2.5839542480465907e-10
GC_7_6 b_7 NI_7 NS_6 0 -1.6679185718995595e-11
GC_7_7 b_7 NI_7 NS_7 0 -1.1229325177294131e-06
GC_7_8 b_7 NI_7 NS_8 0 3.9744249654717764e-06
GC_7_9 b_7 NI_7 NS_9 0 2.2362284825400268e-06
GC_7_10 b_7 NI_7 NS_10 0 9.1490009085799282e-06
GC_7_11 b_7 NI_7 NS_11 0 1.0926853483875681e-05
GC_7_12 b_7 NI_7 NS_12 0 3.7178690856904064e-06
GC_7_13 b_7 NI_7 NS_13 0 1.4674343662880763e-05
GC_7_14 b_7 NI_7 NS_14 0 3.1025615956708194e-05
GC_7_15 b_7 NI_7 NS_15 0 3.7960204442695665e-05
GC_7_16 b_7 NI_7 NS_16 0 -6.4994946093387316e-05
GC_7_17 b_7 NI_7 NS_17 0 -7.1240283132317715e-06
GC_7_18 b_7 NI_7 NS_18 0 1.5945791217210999e-05
GC_7_19 b_7 NI_7 NS_19 0 -1.4978347153059889e-06
GC_7_20 b_7 NI_7 NS_20 0 -5.1730651214532987e-06
GC_7_21 b_7 NI_7 NS_21 0 5.0854210557924887e-05
GC_7_22 b_7 NI_7 NS_22 0 -3.8778252944601612e-05
GC_7_23 b_7 NI_7 NS_23 0 6.8081272333724269e-06
GC_7_24 b_7 NI_7 NS_24 0 -1.4682988975439075e-08
GC_7_25 b_7 NI_7 NS_25 0 -3.5990551015752974e-11
GC_7_26 b_7 NI_7 NS_26 0 8.7893841270895063e-13
GC_7_27 b_7 NI_7 NS_27 0 -3.8162795702844354e-07
GC_7_28 b_7 NI_7 NS_28 0 -1.0212850006642958e-06
GC_7_29 b_7 NI_7 NS_29 0 2.1520820639075009e-06
GC_7_30 b_7 NI_7 NS_30 0 2.5509763676785854e-06
GC_7_31 b_7 NI_7 NS_31 0 3.8434432084512335e-06
GC_7_32 b_7 NI_7 NS_32 0 -4.0510583149479809e-06
GC_7_33 b_7 NI_7 NS_33 0 9.5840558311886663e-06
GC_7_34 b_7 NI_7 NS_34 0 -1.5381443089607903e-05
GC_7_35 b_7 NI_7 NS_35 0 -2.5653768039655851e-05
GC_7_36 b_7 NI_7 NS_36 0 -8.5208295233697479e-06
GC_7_37 b_7 NI_7 NS_37 0 2.3656827184604186e-06
GC_7_38 b_7 NI_7 NS_38 0 2.6330692729917449e-07
GC_7_39 b_7 NI_7 NS_39 0 -6.9147857088505088e-06
GC_7_40 b_7 NI_7 NS_40 0 -3.8167760109744729e-06
GC_7_41 b_7 NI_7 NS_41 0 2.8152219020954287e-04
GC_7_42 b_7 NI_7 NS_42 0 -1.3618967873203273e-05
GC_7_43 b_7 NI_7 NS_43 0 -9.2935601868418792e-06
GC_7_44 b_7 NI_7 NS_44 0 5.9792832659446712e-08
GC_7_45 b_7 NI_7 NS_45 0 -3.0942233006109038e-10
GC_7_46 b_7 NI_7 NS_46 0 9.3377854094469354e-12
GC_7_47 b_7 NI_7 NS_47 0 -7.2720608954612445e-07
GC_7_48 b_7 NI_7 NS_48 0 -1.5722571216373884e-05
GC_7_49 b_7 NI_7 NS_49 0 -9.9778775287892488e-06
GC_7_50 b_7 NI_7 NS_50 0 -2.1078181903246291e-05
GC_7_51 b_7 NI_7 NS_51 0 -3.8198546514135727e-05
GC_7_52 b_7 NI_7 NS_52 0 -1.9856757526571437e-05
GC_7_53 b_7 NI_7 NS_53 0 -7.5906332078321399e-05
GC_7_54 b_7 NI_7 NS_54 0 -7.9824772490027647e-05
GC_7_55 b_7 NI_7 NS_55 0 -7.6276336396007878e-05
GC_7_56 b_7 NI_7 NS_56 0 2.2232889438398030e-04
GC_7_57 b_7 NI_7 NS_57 0 1.5515373960154716e-05
GC_7_58 b_7 NI_7 NS_58 0 -5.7943007494651015e-05
GC_7_59 b_7 NI_7 NS_59 0 -4.8366113771129896e-06
GC_7_60 b_7 NI_7 NS_60 0 1.3913723566528564e-05
GC_7_61 b_7 NI_7 NS_61 0 3.0534411449455201e-04
GC_7_62 b_7 NI_7 NS_62 0 -2.6784573495893725e-04
GC_7_63 b_7 NI_7 NS_63 0 4.2963844359766765e-05
GC_7_64 b_7 NI_7 NS_64 0 1.4101511282416920e-08
GC_7_65 b_7 NI_7 NS_65 0 -1.4707755419539942e-10
GC_7_66 b_7 NI_7 NS_66 0 1.3946692802478960e-11
GC_7_67 b_7 NI_7 NS_67 0 1.6536678491701663e-06
GC_7_68 b_7 NI_7 NS_68 0 7.0334548496977837e-06
GC_7_69 b_7 NI_7 NS_69 0 3.2641712444427585e-05
GC_7_70 b_7 NI_7 NS_70 0 2.1791256996051446e-05
GC_7_71 b_7 NI_7 NS_71 0 4.5840777204033669e-05
GC_7_72 b_7 NI_7 NS_72 0 -5.5994684995783240e-05
GC_7_73 b_7 NI_7 NS_73 0 7.2919507061638050e-05
GC_7_74 b_7 NI_7 NS_74 0 -1.2481997858989924e-04
GC_7_75 b_7 NI_7 NS_75 0 -1.8541625762494605e-04
GC_7_76 b_7 NI_7 NS_76 0 -7.4145717068885107e-05
GC_7_77 b_7 NI_7 NS_77 0 7.6332253356441662e-06
GC_7_78 b_7 NI_7 NS_78 0 3.5082934468758771e-06
GC_7_79 b_7 NI_7 NS_79 0 -5.3960457500944143e-05
GC_7_80 b_7 NI_7 NS_80 0 -3.1131045515411675e-05
GC_7_81 b_7 NI_7 NS_81 0 2.2333485082340444e-02
GC_7_82 b_7 NI_7 NS_82 0 8.9184338894236163e-03
GC_7_83 b_7 NI_7 NS_83 0 -1.1401600407329281e-02
GC_7_84 b_7 NI_7 NS_84 0 -5.3823441542970604e-06
GC_7_85 b_7 NI_7 NS_85 0 -9.5308344304798254e-08
GC_7_86 b_7 NI_7 NS_86 0 -1.2685910996488906e-09
GC_7_87 b_7 NI_7 NS_87 0 -3.3183157151447972e-03
GC_7_88 b_7 NI_7 NS_88 0 -2.3921302584309365e-03
GC_7_89 b_7 NI_7 NS_89 0 2.7239195437716969e-03
GC_7_90 b_7 NI_7 NS_90 0 1.1169875324060977e-02
GC_7_91 b_7 NI_7 NS_91 0 -3.6330705741111492e-04
GC_7_92 b_7 NI_7 NS_92 0 -1.7752735330577155e-02
GC_7_93 b_7 NI_7 NS_93 0 -2.2016949442888699e-02
GC_7_94 b_7 NI_7 NS_94 0 2.1338989335300419e-02
GC_7_95 b_7 NI_7 NS_95 0 2.8916848633880443e-02
GC_7_96 b_7 NI_7 NS_96 0 -1.8399470316659453e-02
GC_7_97 b_7 NI_7 NS_97 0 -2.4531764794582882e-03
GC_7_98 b_7 NI_7 NS_98 0 1.4162712486315101e-03
GC_7_99 b_7 NI_7 NS_99 0 -1.7821660735425411e-02
GC_7_100 b_7 NI_7 NS_100 0 -7.1344518936834840e-03
GC_7_101 b_7 NI_7 NS_101 0 -8.2237001685274022e-02
GC_7_102 b_7 NI_7 NS_102 0 6.5305852819415755e-02
GC_7_103 b_7 NI_7 NS_103 0 -1.0305226886049873e-02
GC_7_104 b_7 NI_7 NS_104 0 -2.4029859715820541e-06
GC_7_105 b_7 NI_7 NS_105 0 1.6307887535605273e-08
GC_7_106 b_7 NI_7 NS_106 0 1.6568107203015891e-09
GC_7_107 b_7 NI_7 NS_107 0 -3.9692405307444799e-04
GC_7_108 b_7 NI_7 NS_108 0 -1.4031043334391141e-03
GC_7_109 b_7 NI_7 NS_109 0 -6.9955150588786024e-03
GC_7_110 b_7 NI_7 NS_110 0 -3.7827359492864109e-03
GC_7_111 b_7 NI_7 NS_111 0 -9.0599083981290490e-03
GC_7_112 b_7 NI_7 NS_112 0 1.3124883430503342e-02
GC_7_113 b_7 NI_7 NS_113 0 -1.5228217957354139e-02
GC_7_114 b_7 NI_7 NS_114 0 2.8706591444978176e-02
GC_7_115 b_7 NI_7 NS_115 0 4.5065279293314185e-02
GC_7_116 b_7 NI_7 NS_116 0 1.6496171688892287e-02
GC_7_117 b_7 NI_7 NS_117 0 -2.1949566522532936e-03
GC_7_118 b_7 NI_7 NS_118 0 -1.3428667044198866e-03
GC_7_119 b_7 NI_7 NS_119 0 1.2861366874928644e-02
GC_7_120 b_7 NI_7 NS_120 0 6.9592344559018682e-03
GC_7_121 b_7 NI_7 NS_121 0 -9.3724215078567065e-04
GC_7_122 b_7 NI_7 NS_122 0 -1.7325126933718588e-02
GC_7_123 b_7 NI_7 NS_123 0 1.1756094412737820e-02
GC_7_124 b_7 NI_7 NS_124 0 2.9426120228631111e-06
GC_7_125 b_7 NI_7 NS_125 0 -5.0962309378903520e-07
GC_7_126 b_7 NI_7 NS_126 0 -2.9668137285065142e-08
GC_7_127 b_7 NI_7 NS_127 0 3.0719111104943685e-03
GC_7_128 b_7 NI_7 NS_128 0 1.2847115797605503e-03
GC_7_129 b_7 NI_7 NS_129 0 -2.9639193838224922e-03
GC_7_130 b_7 NI_7 NS_130 0 -9.9278284017269101e-03
GC_7_131 b_7 NI_7 NS_131 0 5.8579854535478976e-04
GC_7_132 b_7 NI_7 NS_132 0 1.3645082385554848e-02
GC_7_133 b_7 NI_7 NS_133 0 1.7411060835855217e-02
GC_7_134 b_7 NI_7 NS_134 0 -2.3905075600173912e-02
GC_7_135 b_7 NI_7 NS_135 0 -3.3221890743880371e-02
GC_7_136 b_7 NI_7 NS_136 0 2.1449496354453406e-02
GC_7_137 b_7 NI_7 NS_137 0 4.0698749363170259e-03
GC_7_138 b_7 NI_7 NS_138 0 -2.2340713099931399e-03
GC_7_139 b_7 NI_7 NS_139 0 1.5117889894520996e-02
GC_7_140 b_7 NI_7 NS_140 0 5.6202771396554633e-03
GC_7_141 b_7 NI_7 NS_141 0 -2.8556577271113448e-01
GC_7_142 b_7 NI_7 NS_142 0 1.2097570466705823e-01
GC_7_143 b_7 NI_7 NS_143 0 7.0770646840864317e-03
GC_7_144 b_7 NI_7 NS_144 0 5.7565181857973960e-05
GC_7_145 b_7 NI_7 NS_145 0 1.2985823924421718e-06
GC_7_146 b_7 NI_7 NS_146 0 1.4018775899321413e-08
GC_7_147 b_7 NI_7 NS_147 0 3.0464942524720588e-02
GC_7_148 b_7 NI_7 NS_148 0 4.1070361269665481e-03
GC_7_149 b_7 NI_7 NS_149 0 -7.3803962575599230e-03
GC_7_150 b_7 NI_7 NS_150 0 2.2172593675266340e-02
GC_7_151 b_7 NI_7 NS_151 0 -1.7062253783104074e-02
GC_7_152 b_7 NI_7 NS_152 0 -1.8682685512111830e-02
GC_7_153 b_7 NI_7 NS_153 0 4.4646589018879433e-02
GC_7_154 b_7 NI_7 NS_154 0 1.4294478899463782e-02
GC_7_155 b_7 NI_7 NS_155 0 8.1981818313159593e-02
GC_7_156 b_7 NI_7 NS_156 0 3.1414691112676703e-02
GC_7_157 b_7 NI_7 NS_157 0 -1.0082912228060001e-02
GC_7_158 b_7 NI_7 NS_158 0 -4.9140578261129206e-03
GC_7_159 b_7 NI_7 NS_159 0 -2.1489488726548763e-02
GC_7_160 b_7 NI_7 NS_160 0 -4.8797203984274062e-03
GC_7_161 b_7 NI_7 NS_161 0 1.1295688483407996e-04
GC_7_162 b_7 NI_7 NS_162 0 8.2945477082576122e-05
GC_7_163 b_7 NI_7 NS_163 0 -9.5451576287200189e-05
GC_7_164 b_7 NI_7 NS_164 0 -1.1416672263313228e-07
GC_7_165 b_7 NI_7 NS_165 0 -4.3387030287050156e-10
GC_7_166 b_7 NI_7 NS_166 0 -1.2075595162521273e-10
GC_7_167 b_7 NI_7 NS_167 0 -2.9066603421734840e-05
GC_7_168 b_7 NI_7 NS_168 0 -1.6184682557212674e-05
GC_7_169 b_7 NI_7 NS_169 0 2.8967662304576541e-05
GC_7_170 b_7 NI_7 NS_170 0 9.8864603401970365e-05
GC_7_171 b_7 NI_7 NS_171 0 2.9205669465846426e-07
GC_7_172 b_7 NI_7 NS_172 0 -1.4699327713335960e-04
GC_7_173 b_7 NI_7 NS_173 0 -1.6899333925139329e-04
GC_7_174 b_7 NI_7 NS_174 0 2.1090499791694210e-04
GC_7_175 b_7 NI_7 NS_175 0 2.7243837107477920e-04
GC_7_176 b_7 NI_7 NS_176 0 -2.1995137032994308e-04
GC_7_177 b_7 NI_7 NS_177 0 -2.5614900104793586e-05
GC_7_178 b_7 NI_7 NS_178 0 2.7761634542580783e-05
GC_7_179 b_7 NI_7 NS_179 0 -1.5191631439313684e-04
GC_7_180 b_7 NI_7 NS_180 0 -6.4140668310843765e-05
GC_7_181 b_7 NI_7 NS_181 0 -5.4693776099883236e-04
GC_7_182 b_7 NI_7 NS_182 0 4.9511188261016509e-04
GC_7_183 b_7 NI_7 NS_183 0 -7.8372628143930223e-05
GC_7_184 b_7 NI_7 NS_184 0 9.0352476105243056e-09
GC_7_185 b_7 NI_7 NS_185 0 3.0027638711902073e-10
GC_7_186 b_7 NI_7 NS_186 0 8.0533046243752736e-11
GC_7_187 b_7 NI_7 NS_187 0 -1.2560244064780396e-05
GC_7_188 b_7 NI_7 NS_188 0 -8.8756115475211013e-06
GC_7_189 b_7 NI_7 NS_189 0 -6.7306543272958476e-05
GC_7_190 b_7 NI_7 NS_190 0 -3.1843244938294189e-05
GC_7_191 b_7 NI_7 NS_191 0 -7.0775997861515056e-05
GC_7_192 b_7 NI_7 NS_192 0 1.1481870825892720e-04
GC_7_193 b_7 NI_7 NS_193 0 -1.3779794656960506e-04
GC_7_194 b_7 NI_7 NS_194 0 2.2324726954868476e-04
GC_7_195 b_7 NI_7 NS_195 0 3.5690612810441048e-04
GC_7_196 b_7 NI_7 NS_196 0 1.6256169708474339e-04
GC_7_197 b_7 NI_7 NS_197 0 -1.7294704905618621e-05
GC_7_198 b_7 NI_7 NS_198 0 -1.7940494303390717e-05
GC_7_199 b_7 NI_7 NS_199 0 1.0162292740936856e-04
GC_7_200 b_7 NI_7 NS_200 0 5.6167512421354907e-05
GC_7_201 b_7 NI_7 NS_201 0 2.7780708388510836e-04
GC_7_202 b_7 NI_7 NS_202 0 -1.2250103120979064e-05
GC_7_203 b_7 NI_7 NS_203 0 -9.4861499302946406e-06
GC_7_204 b_7 NI_7 NS_204 0 6.0731552451156132e-08
GC_7_205 b_7 NI_7 NS_205 0 -3.1317771972860439e-10
GC_7_206 b_7 NI_7 NS_206 0 8.9456590353495299e-12
GC_7_207 b_7 NI_7 NS_207 0 -7.0467252398542909e-07
GC_7_208 b_7 NI_7 NS_208 0 -1.5599737169766636e-05
GC_7_209 b_7 NI_7 NS_209 0 -9.9256357284097889e-06
GC_7_210 b_7 NI_7 NS_210 0 -2.0930532505578008e-05
GC_7_211 b_7 NI_7 NS_211 0 -3.7989342561761040e-05
GC_7_212 b_7 NI_7 NS_212 0 -1.9683745835306009e-05
GC_7_213 b_7 NI_7 NS_213 0 -7.5824501991868915e-05
GC_7_214 b_7 NI_7 NS_214 0 -7.9099395990473427e-05
GC_7_215 b_7 NI_7 NS_215 0 -7.4562448879335932e-05
GC_7_216 b_7 NI_7 NS_216 0 2.2166872018915479e-04
GC_7_217 b_7 NI_7 NS_217 0 1.5124434955054780e-05
GC_7_218 b_7 NI_7 NS_218 0 -5.7842961357215893e-05
GC_7_219 b_7 NI_7 NS_219 0 -4.6595009907653252e-06
GC_7_220 b_7 NI_7 NS_220 0 1.3855697755715459e-05
GC_7_221 b_7 NI_7 NS_221 0 3.0653426568902473e-04
GC_7_222 b_7 NI_7 NS_222 0 -2.6884033599544350e-04
GC_7_223 b_7 NI_7 NS_223 0 4.3094719103069400e-05
GC_7_224 b_7 NI_7 NS_224 0 1.3367636864314108e-08
GC_7_225 b_7 NI_7 NS_225 0 -1.4591751340557129e-10
GC_7_226 b_7 NI_7 NS_226 0 1.4531715036321401e-11
GC_7_227 b_7 NI_7 NS_227 0 1.8114016091243147e-06
GC_7_228 b_7 NI_7 NS_228 0 7.0832229582860302e-06
GC_7_229 b_7 NI_7 NS_229 0 3.2827978510239235e-05
GC_7_230 b_7 NI_7 NS_230 0 2.1661354227507276e-05
GC_7_231 b_7 NI_7 NS_231 0 4.5946585831196335e-05
GC_7_232 b_7 NI_7 NS_232 0 -5.6356955538016700e-05
GC_7_233 b_7 NI_7 NS_233 0 7.3626811598729523e-05
GC_7_234 b_7 NI_7 NS_234 0 -1.2529400709936130e-04
GC_7_235 b_7 NI_7 NS_235 0 -1.8750648006890335e-04
GC_7_236 b_7 NI_7 NS_236 0 -7.4918080160569510e-05
GC_7_237 b_7 NI_7 NS_237 0 8.1189043601180942e-06
GC_7_238 b_7 NI_7 NS_238 0 3.6709412360546730e-06
GC_7_239 b_7 NI_7 NS_239 0 -5.4185551642336151e-05
GC_7_240 b_7 NI_7 NS_240 0 -3.1100960358688675e-05
GD_7_1 b_7 NI_7 NA_1 0 1.9757259931334307e-05
GD_7_2 b_7 NI_7 NA_2 0 -3.9272282197895332e-06
GD_7_3 b_7 NI_7 NA_3 0 -6.9856716951854361e-05
GD_7_4 b_7 NI_7 NA_4 0 4.0802500649629713e-06
GD_7_5 b_7 NI_7 NA_5 0 6.1947474642984474e-03
GD_7_6 b_7 NI_7 NA_6 0 2.3344520397488963e-03
GD_7_7 b_7 NI_7 NA_7 0 -6.6185353254439314e-03
GD_7_8 b_7 NI_7 NA_8 0 5.6693579752425956e-02
GD_7_9 b_7 NI_7 NA_9 0 7.9448663504775118e-05
GD_7_10 b_7 NI_7 NA_10 0 -4.8736497492237166e-05
GD_7_11 b_7 NI_7 NA_11 0 -6.9107945941876872e-05
GD_7_12 b_7 NI_7 NA_12 0 4.7002113945810332e-06
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 5.0922304796729432e-05
GC_8_2 b_8 NI_8 NS_2 0 -3.8768879851388353e-05
GC_8_3 b_8 NI_8 NS_3 0 6.8058310931519460e-06
GC_8_4 b_8 NI_8 NS_4 0 -1.4678933388118026e-08
GC_8_5 b_8 NI_8 NS_5 0 -3.5984987794502828e-11
GC_8_6 b_8 NI_8 NS_6 0 8.7817190832386738e-13
GC_8_7 b_8 NI_8 NS_7 0 -3.9997170533247758e-07
GC_8_8 b_8 NI_8 NS_8 0 -1.0354840870727227e-06
GC_8_9 b_8 NI_8 NS_9 0 2.1268630337491299e-06
GC_8_10 b_8 NI_8 NS_10 0 2.5480814699178871e-06
GC_8_11 b_8 NI_8 NS_11 0 3.8281431402898081e-06
GC_8_12 b_8 NI_8 NS_12 0 -4.0076902610083228e-06
GC_8_13 b_8 NI_8 NS_13 0 9.5696479450842827e-06
GC_8_14 b_8 NI_8 NS_14 0 -1.5346626883144033e-05
GC_8_15 b_8 NI_8 NS_15 0 -2.5610122899577654e-05
GC_8_16 b_8 NI_8 NS_16 0 -8.5179429655716931e-06
GC_8_17 b_8 NI_8 NS_17 0 2.3607091123099380e-06
GC_8_18 b_8 NI_8 NS_18 0 2.6764566791704927e-07
GC_8_19 b_8 NI_8 NS_19 0 -6.9119891801749786e-06
GC_8_20 b_8 NI_8 NS_20 0 -3.8140224812499678e-06
GC_8_21 b_8 NI_8 NS_21 0 -8.6861196529398408e-05
GC_8_22 b_8 NI_8 NS_22 0 1.4645966944272327e-05
GC_8_23 b_8 NI_8 NS_23 0 -1.4880453250722978e-06
GC_8_24 b_8 NI_8 NS_24 0 -1.2743198584706806e-08
GC_8_25 b_8 NI_8 NS_25 0 2.5843959272213887e-10
GC_8_26 b_8 NI_8 NS_26 0 -1.6682804013659127e-11
GC_8_27 b_8 NI_8 NS_27 0 -1.1230021576452320e-06
GC_8_28 b_8 NI_8 NS_28 0 3.9730700117245459e-06
GC_8_29 b_8 NI_8 NS_29 0 2.2350121324021180e-06
GC_8_30 b_8 NI_8 NS_30 0 9.1477027438306674e-06
GC_8_31 b_8 NI_8 NS_31 0 1.0925656223202944e-05
GC_8_32 b_8 NI_8 NS_32 0 3.7171219761878228e-06
GC_8_33 b_8 NI_8 NS_33 0 1.4672172931112702e-05
GC_8_34 b_8 NI_8 NS_34 0 3.1019471994233983e-05
GC_8_35 b_8 NI_8 NS_35 0 3.7950164218659241e-05
GC_8_36 b_8 NI_8 NS_36 0 -6.4987152541086052e-05
GC_8_37 b_8 NI_8 NS_37 0 -7.1220145697854168e-06
GC_8_38 b_8 NI_8 NS_38 0 1.5944609030093089e-05
GC_8_39 b_8 NI_8 NS_39 0 -1.4986072843363618e-06
GC_8_40 b_8 NI_8 NS_40 0 -5.1723139022570671e-06
GC_8_41 b_8 NI_8 NS_41 0 3.0534162138949822e-04
GC_8_42 b_8 NI_8 NS_42 0 -2.6784547256392561e-04
GC_8_43 b_8 NI_8 NS_43 0 4.2963856641671385e-05
GC_8_44 b_8 NI_8 NS_44 0 1.4101248633886102e-08
GC_8_45 b_8 NI_8 NS_45 0 -1.4707387091607279e-10
GC_8_46 b_8 NI_8 NS_46 0 1.3946538889474264e-11
GC_8_47 b_8 NI_8 NS_47 0 1.6535510617389610e-06
GC_8_48 b_8 NI_8 NS_48 0 7.0335452705204600e-06
GC_8_49 b_8 NI_8 NS_49 0 3.2641608555240523e-05
GC_8_50 b_8 NI_8 NS_50 0 2.1791552353628925e-05
GC_8_51 b_8 NI_8 NS_51 0 4.5841507133548152e-05
GC_8_52 b_8 NI_8 NS_52 0 -5.5994157904633657e-05
GC_8_53 b_8 NI_8 NS_53 0 7.2920974293673679e-05
GC_8_54 b_8 NI_8 NS_54 0 -1.2481942338883546e-04
GC_8_55 b_8 NI_8 NS_55 0 -1.8541708907612647e-04
GC_8_56 b_8 NI_8 NS_56 0 -7.4147695752073650e-05
GC_8_57 b_8 NI_8 NS_57 0 7.6337243491298641e-06
GC_8_58 b_8 NI_8 NS_58 0 3.5085200629176176e-06
GC_8_59 b_8 NI_8 NS_59 0 -5.3960441175047136e-05
GC_8_60 b_8 NI_8 NS_60 0 -3.1131141088558436e-05
GC_8_61 b_8 NI_8 NS_61 0 2.8249440270747598e-04
GC_8_62 b_8 NI_8 NS_62 0 -1.3810042618752528e-05
GC_8_63 b_8 NI_8 NS_63 0 -9.2728558042537388e-06
GC_8_64 b_8 NI_8 NS_64 0 5.9696244784367656e-08
GC_8_65 b_8 NI_8 NS_65 0 -3.0906094163153654e-10
GC_8_66 b_8 NI_8 NS_66 0 9.3204269140457198e-12
GC_8_67 b_8 NI_8 NS_67 0 -7.6635919320991919e-07
GC_8_68 b_8 NI_8 NS_68 0 -1.5748718149639141e-05
GC_8_69 b_8 NI_8 NS_69 0 -1.0078797657654730e-05
GC_8_70 b_8 NI_8 NS_70 0 -2.1107423680928065e-05
GC_8_71 b_8 NI_8 NS_71 0 -3.8248667649133242e-05
GC_8_72 b_8 NI_8 NS_72 0 -1.9774688623254621e-05
GC_8_73 b_8 NI_8 NS_73 0 -7.5998900608222194e-05
GC_8_74 b_8 NI_8 NS_74 0 -7.9943369533168256e-05
GC_8_75 b_8 NI_8 NS_75 0 -7.6445579035574823e-05
GC_8_76 b_8 NI_8 NS_76 0 2.2266396074103716e-04
GC_8_77 b_8 NI_8 NS_77 0 1.5542652519110110e-05
GC_8_78 b_8 NI_8 NS_78 0 -5.8015181124038666e-05
GC_8_79 b_8 NI_8 NS_79 0 -4.8512122542565739e-06
GC_8_80 b_8 NI_8 NS_80 0 1.3939680235870520e-05
GC_8_81 b_8 NI_8 NS_81 0 -8.2237002117102137e-02
GC_8_82 b_8 NI_8 NS_82 0 6.5305853062585462e-02
GC_8_83 b_8 NI_8 NS_83 0 -1.0305226917226339e-02
GC_8_84 b_8 NI_8 NS_84 0 -2.4029859122670905e-06
GC_8_85 b_8 NI_8 NS_85 0 1.6307886457941093e-08
GC_8_86 b_8 NI_8 NS_86 0 1.6568107759413235e-09
GC_8_87 b_8 NI_8 NS_87 0 -3.9692419158303551e-04
GC_8_88 b_8 NI_8 NS_88 0 -1.4031044046410438e-03
GC_8_89 b_8 NI_8 NS_89 0 -6.9955152491419231e-03
GC_8_90 b_8 NI_8 NS_90 0 -3.7827359209492289e-03
GC_8_91 b_8 NI_8 NS_91 0 -9.0599084303843620e-03
GC_8_92 b_8 NI_8 NS_92 0 1.3124883863189675e-02
GC_8_93 b_8 NI_8 NS_93 0 -1.5228217851274994e-02
GC_8_94 b_8 NI_8 NS_94 0 2.8706592097895969e-02
GC_8_95 b_8 NI_8 NS_95 0 4.5065279952735335e-02
GC_8_96 b_8 NI_8 NS_96 0 1.6496170910624042e-02
GC_8_97 b_8 NI_8 NS_97 0 -2.1949567238097518e-03
GC_8_98 b_8 NI_8 NS_98 0 -1.3428664599567702e-03
GC_8_99 b_8 NI_8 NS_99 0 1.2861366894128383e-02
GC_8_100 b_8 NI_8 NS_100 0 6.9592344390310389e-03
GC_8_101 b_8 NI_8 NS_101 0 2.2333485084293284e-02
GC_8_102 b_8 NI_8 NS_102 0 8.9184338921983707e-03
GC_8_103 b_8 NI_8 NS_103 0 -1.1401600408274912e-02
GC_8_104 b_8 NI_8 NS_104 0 -5.3823441502440696e-06
GC_8_105 b_8 NI_8 NS_105 0 -9.5308344342151229e-08
GC_8_106 b_8 NI_8 NS_106 0 -1.2685911015145559e-09
GC_8_107 b_8 NI_8 NS_107 0 -3.3183157155340492e-03
GC_8_108 b_8 NI_8 NS_108 0 -2.3921302575102017e-03
GC_8_109 b_8 NI_8 NS_109 0 2.7239195453364101e-03
GC_8_110 b_8 NI_8 NS_110 0 1.1169875325987046e-02
GC_8_111 b_8 NI_8 NS_111 0 -3.6330705414728279e-04
GC_8_112 b_8 NI_8 NS_112 0 -1.7752735332879424e-02
GC_8_113 b_8 NI_8 NS_113 0 -2.2016949437053797e-02
GC_8_114 b_8 NI_8 NS_114 0 2.1338989327258542e-02
GC_8_115 b_8 NI_8 NS_115 0 2.8916848613793029e-02
GC_8_116 b_8 NI_8 NS_116 0 -1.8399470310471816e-02
GC_8_117 b_8 NI_8 NS_117 0 -2.4531764736285991e-03
GC_8_118 b_8 NI_8 NS_118 0 1.4162712460930320e-03
GC_8_119 b_8 NI_8 NS_119 0 -1.7821660735131032e-02
GC_8_120 b_8 NI_8 NS_120 0 -7.1344518915960791e-03
GC_8_121 b_8 NI_8 NS_121 0 -2.8556577260564170e-01
GC_8_122 b_8 NI_8 NS_122 0 1.2097570466138365e-01
GC_8_123 b_8 NI_8 NS_123 0 7.0770646832974777e-03
GC_8_124 b_8 NI_8 NS_124 0 5.7565181885888209e-05
GC_8_125 b_8 NI_8 NS_125 0 1.2985823916461685e-06
GC_8_126 b_8 NI_8 NS_126 0 1.4018775955621386e-08
GC_8_127 b_8 NI_8 NS_127 0 3.0464942510763079e-02
GC_8_128 b_8 NI_8 NS_128 0 4.1070361151387532e-03
GC_8_129 b_8 NI_8 NS_129 0 -7.3803962867941388e-03
GC_8_130 b_8 NI_8 NS_130 0 2.2172593674932080e-02
GC_8_131 b_8 NI_8 NS_131 0 -1.7062253800483457e-02
GC_8_132 b_8 NI_8 NS_132 0 -1.8682685482283010e-02
GC_8_133 b_8 NI_8 NS_133 0 4.4646588975949704e-02
GC_8_134 b_8 NI_8 NS_134 0 1.4294478945091137e-02
GC_8_135 b_8 NI_8 NS_135 0 8.1981818399922537e-02
GC_8_136 b_8 NI_8 NS_136 0 3.1414691106161768e-02
GC_8_137 b_8 NI_8 NS_137 0 -1.0082912249571925e-02
GC_8_138 b_8 NI_8 NS_138 0 -4.9140578126671006e-03
GC_8_139 b_8 NI_8 NS_139 0 -2.1489488728870142e-02
GC_8_140 b_8 NI_8 NS_140 0 -4.8797203983669043e-03
GC_8_141 b_8 NI_8 NS_141 0 -9.3724215078574318e-04
GC_8_142 b_8 NI_8 NS_142 0 -1.7325126933718585e-02
GC_8_143 b_8 NI_8 NS_143 0 1.1756094412737826e-02
GC_8_144 b_8 NI_8 NS_144 0 2.9426120228621324e-06
GC_8_145 b_8 NI_8 NS_145 0 -5.0962309378901127e-07
GC_8_146 b_8 NI_8 NS_146 0 -2.9668137285067015e-08
GC_8_147 b_8 NI_8 NS_147 0 3.0719111104943729e-03
GC_8_148 b_8 NI_8 NS_148 0 1.2847115797605493e-03
GC_8_149 b_8 NI_8 NS_149 0 -2.9639193838225017e-03
GC_8_150 b_8 NI_8 NS_150 0 -9.9278284017269066e-03
GC_8_151 b_8 NI_8 NS_151 0 5.8579854535479941e-04
GC_8_152 b_8 NI_8 NS_152 0 1.3645082385554853e-02
GC_8_153 b_8 NI_8 NS_153 0 1.7411060835855217e-02
GC_8_154 b_8 NI_8 NS_154 0 -2.3905075600173901e-02
GC_8_155 b_8 NI_8 NS_155 0 -3.3221890743880343e-02
GC_8_156 b_8 NI_8 NS_156 0 2.1449496354453396e-02
GC_8_157 b_8 NI_8 NS_157 0 4.0698749363170189e-03
GC_8_158 b_8 NI_8 NS_158 0 -2.2340713099931390e-03
GC_8_159 b_8 NI_8 NS_159 0 1.5117889894521005e-02
GC_8_160 b_8 NI_8 NS_160 0 5.6202771396554633e-03
GC_8_161 b_8 NI_8 NS_161 0 -5.4700630736864665e-04
GC_8_162 b_8 NI_8 NS_162 0 4.9510290645380826e-04
GC_8_163 b_8 NI_8 NS_163 0 -7.8370283245133047e-05
GC_8_164 b_8 NI_8 NS_164 0 9.0303558157988963e-09
GC_8_165 b_8 NI_8 NS_165 0 3.0029232059912873e-10
GC_8_166 b_8 NI_8 NS_166 0 8.0533182863992651e-11
GC_8_167 b_8 NI_8 NS_167 0 -1.2542339718070109e-05
GC_8_168 b_8 NI_8 NS_168 0 -8.8614480795574400e-06
GC_8_169 b_8 NI_8 NS_169 0 -6.7281719743211382e-05
GC_8_170 b_8 NI_8 NS_170 0 -3.1840155382627175e-05
GC_8_171 b_8 NI_8 NS_171 0 -7.0761526839265080e-05
GC_8_172 b_8 NI_8 NS_172 0 1.1477601938023793e-04
GC_8_173 b_8 NI_8 NS_173 0 -1.3778574473057975e-04
GC_8_174 b_8 NI_8 NS_174 0 2.2321532285458096e-04
GC_8_175 b_8 NI_8 NS_175 0 3.5686973575447736e-04
GC_8_176 b_8 NI_8 NS_176 0 1.6255711117117583e-04
GC_8_177 b_8 NI_8 NS_177 0 -1.7291809301621067e-05
GC_8_178 b_8 NI_8 NS_178 0 -1.7943729313510633e-05
GC_8_179 b_8 NI_8 NS_179 0 1.0162026241381898e-04
GC_8_180 b_8 NI_8 NS_180 0 5.6164392909121803e-05
GC_8_181 b_8 NI_8 NS_181 0 1.1295860957999061e-04
GC_8_182 b_8 NI_8 NS_182 0 8.2948154979246985e-05
GC_8_183 b_8 NI_8 NS_183 0 -9.5452145996015889e-05
GC_8_184 b_8 NI_8 NS_184 0 -1.1416549134760427e-07
GC_8_185 b_8 NI_8 NS_185 0 -4.3389909607732016e-10
GC_8_186 b_8 NI_8 NS_186 0 -1.2075666852436992e-10
GC_8_187 b_8 NI_8 NS_187 0 -2.9066900436932843e-05
GC_8_188 b_8 NI_8 NS_188 0 -1.6185056268689840e-05
GC_8_189 b_8 NI_8 NS_189 0 2.8967501300347830e-05
GC_8_190 b_8 NI_8 NS_190 0 9.8864437596006395e-05
GC_8_191 b_8 NI_8 NS_191 0 2.9105541260965561e-07
GC_8_192 b_8 NI_8 NS_192 0 -1.4699361475030347e-04
GC_8_193 b_8 NI_8 NS_193 0 -1.6899605726924643e-04
GC_8_194 b_8 NI_8 NS_194 0 2.1090410183706828e-04
GC_8_195 b_8 NI_8 NS_195 0 2.7243933392665187e-04
GC_8_196 b_8 NI_8 NS_196 0 -2.1994524868997983e-04
GC_8_197 b_8 NI_8 NS_197 0 -2.5615043947262666e-05
GC_8_198 b_8 NI_8 NS_198 0 2.7760261129273368e-05
GC_8_199 b_8 NI_8 NS_199 0 -1.5191569672424394e-04
GC_8_200 b_8 NI_8 NS_200 0 -6.4140001405985848e-05
GC_8_201 b_8 NI_8 NS_201 0 3.0653418678396179e-04
GC_8_202 b_8 NI_8 NS_202 0 -2.6883991117702971e-04
GC_8_203 b_8 NI_8 NS_203 0 4.3094616081745343e-05
GC_8_204 b_8 NI_8 NS_204 0 1.3368227447538744e-08
GC_8_205 b_8 NI_8 NS_205 0 -1.4592404995304150e-10
GC_8_206 b_8 NI_8 NS_206 0 1.4532028068205193e-11
GC_8_207 b_8 NI_8 NS_207 0 1.8116505436718663e-06
GC_8_208 b_8 NI_8 NS_208 0 7.0833099479955468e-06
GC_8_209 b_8 NI_8 NS_209 0 3.2828259682875197e-05
GC_8_210 b_8 NI_8 NS_210 0 2.1661244081668436e-05
GC_8_211 b_8 NI_8 NS_211 0 4.5946353490536149e-05
GC_8_212 b_8 NI_8 NS_212 0 -5.6357656261570595e-05
GC_8_213 b_8 NI_8 NS_213 0 7.3626025786069707e-05
GC_8_214 b_8 NI_8 NS_214 0 -1.2529469360062547e-04
GC_8_215 b_8 NI_8 NS_215 0 -1.8750628200790031e-04
GC_8_216 b_8 NI_8 NS_216 0 -7.4916452619383256e-05
GC_8_217 b_8 NI_8 NS_217 0 8.1186769826125205e-06
GC_8_218 b_8 NI_8 NS_218 0 3.6705872337105529e-06
GC_8_219 b_8 NI_8 NS_219 0 -5.4185473728654012e-05
GC_8_220 b_8 NI_8 NS_220 0 -3.1100851543840687e-05
GC_8_221 b_8 NI_8 NS_221 0 2.7679949274189366e-04
GC_8_222 b_8 NI_8 NS_222 0 -1.2052535148694732e-05
GC_8_223 b_8 NI_8 NS_223 0 -9.5072293465876136e-06
GC_8_224 b_8 NI_8 NS_224 0 6.0829925867838725e-08
GC_8_225 b_8 NI_8 NS_225 0 -3.1352473221155163e-10
GC_8_226 b_8 NI_8 NS_226 0 8.9636904157295970e-12
GC_8_227 b_8 NI_8 NS_227 0 -6.6497574178377544e-07
GC_8_228 b_8 NI_8 NS_228 0 -1.5571150330555896e-05
GC_8_229 b_8 NI_8 NS_229 0 -9.8226342205528997e-06
GC_8_230 b_8 NI_8 NS_230 0 -2.0899212882511418e-05
GC_8_231 b_8 NI_8 NS_231 0 -3.7936282424100298e-05
GC_8_232 b_8 NI_8 NS_232 0 -1.9764556219873195e-05
GC_8_233 b_8 NI_8 NS_233 0 -7.5725766778674312e-05
GC_8_234 b_8 NI_8 NS_234 0 -7.8970931115215893e-05
GC_8_235 b_8 NI_8 NS_235 0 -7.4379444878578177e-05
GC_8_236 b_8 NI_8 NS_236 0 2.2131546830836518e-04
GC_8_237 b_8 NI_8 NS_237 0 1.5094322300799678e-05
GC_8_238 b_8 NI_8 NS_238 0 -5.7767603465752146e-05
GC_8_239 b_8 NI_8 NS_239 0 -4.6444428821838573e-06
GC_8_240 b_8 NI_8 NS_240 0 1.3827759029105690e-05
GD_8_1 b_8 NI_8 NA_1 0 -3.9775991179505098e-06
GD_8_2 b_8 NI_8 NA_2 0 1.9756190420277364e-05
GD_8_3 b_8 NI_8 NA_3 0 4.0808617056373521e-06
GD_8_4 b_8 NI_8 NA_4 0 -7.0349371682824994e-05
GD_8_5 b_8 NI_8 NA_5 0 2.3344518686093029e-03
GD_8_6 b_8 NI_8 NA_6 0 6.1947474638148706e-03
GD_8_7 b_8 NI_8 NA_7 0 5.6693579678370000e-02
GD_8_8 b_8 NI_8 NA_8 0 -6.6185353254438854e-03
GD_8_9 b_8 NI_8 NA_9 0 -4.8688361207463915e-05
GD_8_10 b_8 NI_8 NA_10 0 7.9447560877128203e-05
GD_8_11 b_8 NI_8 NA_11 0 4.7004525765287765e-06
GD_8_12 b_8 NI_8 NA_12 0 -6.8612069487168189e-05
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 5.7390978472196079e-06
GC_9_2 b_9 NI_9 NS_2 0 1.3787316872853473e-06
GC_9_3 b_9 NI_9 NS_3 0 -8.6637357012641800e-07
GC_9_4 b_9 NI_9 NS_4 0 3.5224553343904405e-09
GC_9_5 b_9 NI_9 NS_5 0 5.0090022385165303e-11
GC_9_6 b_9 NI_9 NS_6 0 -5.2606201913128829e-13
GC_9_7 b_9 NI_9 NS_7 0 -4.1959944494275981e-07
GC_9_8 b_9 NI_9 NS_8 0 -3.4603311163766656e-07
GC_9_9 b_9 NI_9 NS_9 0 -2.5691669367213909e-07
GC_9_10 b_9 NI_9 NS_10 0 2.1863621766120423e-07
GC_9_11 b_9 NI_9 NS_11 0 -7.9604792207329838e-07
GC_9_12 b_9 NI_9 NS_12 0 -6.7621313136515386e-07
GC_9_13 b_9 NI_9 NS_13 0 -2.5375267671999934e-06
GC_9_14 b_9 NI_9 NS_14 0 -5.5017921379453530e-08
GC_9_15 b_9 NI_9 NS_15 0 3.8307271170020004e-07
GC_9_16 b_9 NI_9 NS_16 0 3.5238200844103892e-06
GC_9_17 b_9 NI_9 NS_17 0 1.6617774946858615e-07
GC_9_18 b_9 NI_9 NS_18 0 -8.5364105748222129e-07
GC_9_19 b_9 NI_9 NS_19 0 -5.6158082569454399e-07
GC_9_20 b_9 NI_9 NS_20 0 2.6962865853453207e-07
GC_9_21 b_9 NI_9 NS_21 0 2.0691345314184144e-05
GC_9_22 b_9 NI_9 NS_22 0 -5.0104182769148830e-06
GC_9_23 b_9 NI_9 NS_23 0 9.9579377396015020e-07
GC_9_24 b_9 NI_9 NS_24 0 -5.5012564767940408e-09
GC_9_25 b_9 NI_9 NS_25 0 -2.5924685435604894e-11
GC_9_26 b_9 NI_9 NS_26 0 -1.2333383506991129e-12
GC_9_27 b_9 NI_9 NS_27 0 -1.3186629654225303e-06
GC_9_28 b_9 NI_9 NS_28 0 -1.6811874878464046e-06
GC_9_29 b_9 NI_9 NS_29 0 -1.8034003428717991e-06
GC_9_30 b_9 NI_9 NS_30 0 1.3685277780664647e-07
GC_9_31 b_9 NI_9 NS_31 0 -2.4181787501519283e-06
GC_9_32 b_9 NI_9 NS_32 0 2.2165267222021415e-06
GC_9_33 b_9 NI_9 NS_33 0 -3.9553371628630241e-06
GC_9_34 b_9 NI_9 NS_34 0 -2.1598076618584207e-06
GC_9_35 b_9 NI_9 NS_35 0 1.2334142081022223e-06
GC_9_36 b_9 NI_9 NS_36 0 8.3243681164320260e-06
GC_9_37 b_9 NI_9 NS_37 0 -3.9465939055221754e-07
GC_9_38 b_9 NI_9 NS_38 0 -1.7930221500150909e-06
GC_9_39 b_9 NI_9 NS_39 0 -3.7110442774730541e-07
GC_9_40 b_9 NI_9 NS_40 0 1.7920434640260530e-07
GC_9_41 b_9 NI_9 NS_41 0 2.2540462022863969e-05
GC_9_42 b_9 NI_9 NS_42 0 -5.1376211092534144e-06
GC_9_43 b_9 NI_9 NS_43 0 3.6838722517184406e-07
GC_9_44 b_9 NI_9 NS_44 0 -8.1493942573161294e-09
GC_9_45 b_9 NI_9 NS_45 0 1.7606409927238712e-10
GC_9_46 b_9 NI_9 NS_46 0 -9.7890746400997934e-12
GC_9_47 b_9 NI_9 NS_47 0 -1.2143346670359238e-06
GC_9_48 b_9 NI_9 NS_48 0 -9.1148481915432079e-07
GC_9_49 b_9 NI_9 NS_49 0 -1.3990075973254999e-06
GC_9_50 b_9 NI_9 NS_50 0 -4.6289012470772894e-08
GC_9_51 b_9 NI_9 NS_51 0 -2.2031483324576186e-06
GC_9_52 b_9 NI_9 NS_52 0 2.3009464661419670e-08
GC_9_53 b_9 NI_9 NS_53 0 -4.7814127875165956e-06
GC_9_54 b_9 NI_9 NS_54 0 -4.5206613922041123e-07
GC_9_55 b_9 NI_9 NS_55 0 1.0105769195528552e-06
GC_9_56 b_9 NI_9 NS_56 0 7.1429856948233686e-06
GC_9_57 b_9 NI_9 NS_57 0 -3.5880409707351817e-07
GC_9_58 b_9 NI_9 NS_58 0 -1.8238538657411689e-06
GC_9_59 b_9 NI_9 NS_59 0 -1.0678623679011704e-06
GC_9_60 b_9 NI_9 NS_60 0 -3.9175124926740367e-07
GC_9_61 b_9 NI_9 NS_61 0 7.9173689463955098e-06
GC_9_62 b_9 NI_9 NS_62 0 -6.3418633442494048e-06
GC_9_63 b_9 NI_9 NS_63 0 4.7307430386273644e-07
GC_9_64 b_9 NI_9 NS_64 0 6.3738330768437887e-09
GC_9_65 b_9 NI_9 NS_65 0 -1.7569995758695236e-10
GC_9_66 b_9 NI_9 NS_66 0 8.2809626722172790e-12
GC_9_67 b_9 NI_9 NS_67 0 2.1359813233563007e-06
GC_9_68 b_9 NI_9 NS_68 0 -1.0057334842407916e-06
GC_9_69 b_9 NI_9 NS_69 0 2.8515665735692241e-06
GC_9_70 b_9 NI_9 NS_70 0 -1.3365743353395821e-06
GC_9_71 b_9 NI_9 NS_71 0 -2.5442370008941502e-07
GC_9_72 b_9 NI_9 NS_72 0 -3.4600117309024631e-06
GC_9_73 b_9 NI_9 NS_73 0 6.9380325851026979e-06
GC_9_74 b_9 NI_9 NS_74 0 -9.0883170900202075e-06
GC_9_75 b_9 NI_9 NS_75 0 -2.3892363422471707e-05
GC_9_76 b_9 NI_9 NS_76 0 -2.8584524701212824e-06
GC_9_77 b_9 NI_9 NS_77 0 5.9682591638931127e-06
GC_9_78 b_9 NI_9 NS_78 0 3.0695667226183084e-07
GC_9_79 b_9 NI_9 NS_79 0 -2.6280911429555245e-06
GC_9_80 b_9 NI_9 NS_80 0 1.4076505273487909e-06
GC_9_81 b_9 NI_9 NS_81 0 2.7806787162304171e-04
GC_9_82 b_9 NI_9 NS_82 0 -1.2586345914534690e-05
GC_9_83 b_9 NI_9 NS_83 0 -9.4421654407147865e-06
GC_9_84 b_9 NI_9 NS_84 0 6.0630184423795253e-08
GC_9_85 b_9 NI_9 NS_85 0 -3.1771024162602426e-10
GC_9_86 b_9 NI_9 NS_86 0 9.7760230307355103e-12
GC_9_87 b_9 NI_9 NS_87 0 -6.2007908928787734e-07
GC_9_88 b_9 NI_9 NS_88 0 -1.5605308694624964e-05
GC_9_89 b_9 NI_9 NS_89 0 -9.8498685703432411e-06
GC_9_90 b_9 NI_9 NS_90 0 -2.0984727374794569e-05
GC_9_91 b_9 NI_9 NS_91 0 -3.7922143369977857e-05
GC_9_92 b_9 NI_9 NS_92 0 -1.9808608657779218e-05
GC_9_93 b_9 NI_9 NS_93 0 -7.5514369191119674e-05
GC_9_94 b_9 NI_9 NS_94 0 -7.9383283150906119e-05
GC_9_95 b_9 NI_9 NS_95 0 -7.5463294631634552e-05
GC_9_96 b_9 NI_9 NS_96 0 2.2133252132671823e-04
GC_9_97 b_9 NI_9 NS_97 0 1.5336579952058152e-05
GC_9_98 b_9 NI_9 NS_98 0 -5.7741341368022671e-05
GC_9_99 b_9 NI_9 NS_99 0 -4.7436874531114934e-06
GC_9_100 b_9 NI_9 NS_100 0 1.3885238330345280e-05
GC_9_101 b_9 NI_9 NS_101 0 3.0487060545463673e-04
GC_9_102 b_9 NI_9 NS_102 0 -2.6795564239579905e-04
GC_9_103 b_9 NI_9 NS_103 0 4.3029677918844925e-05
GC_9_104 b_9 NI_9 NS_104 0 1.3275140730396054e-08
GC_9_105 b_9 NI_9 NS_105 0 -1.3642171731729853e-10
GC_9_106 b_9 NI_9 NS_106 0 1.3413647668954505e-11
GC_9_107 b_9 NI_9 NS_107 0 1.6673085993155116e-06
GC_9_108 b_9 NI_9 NS_108 0 7.0536130908585309e-06
GC_9_109 b_9 NI_9 NS_109 0 3.2663687313656756e-05
GC_9_110 b_9 NI_9 NS_110 0 2.1834068066124051e-05
GC_9_111 b_9 NI_9 NS_111 0 4.5895161296623844e-05
GC_9_112 b_9 NI_9 NS_112 0 -5.6019838141730546e-05
GC_9_113 b_9 NI_9 NS_113 0 7.3005719399870631e-05
GC_9_114 b_9 NI_9 NS_114 0 -1.2465455971853617e-04
GC_9_115 b_9 NI_9 NS_115 0 -1.8515939561345837e-04
GC_9_116 b_9 NI_9 NS_116 0 -7.4482521203583923e-05
GC_9_117 b_9 NI_9 NS_117 0 7.5437636130375665e-06
GC_9_118 b_9 NI_9 NS_118 0 3.5788425067525051e-06
GC_9_119 b_9 NI_9 NS_119 0 -5.3931892134989854e-05
GC_9_120 b_9 NI_9 NS_120 0 -3.1184820051210550e-05
GC_9_121 b_9 NI_9 NS_121 0 1.1295861105546993e-04
GC_9_122 b_9 NI_9 NS_122 0 8.2948154367615037e-05
GC_9_123 b_9 NI_9 NS_123 0 -9.5452145907623799e-05
GC_9_124 b_9 NI_9 NS_124 0 -1.1416549193369561e-07
GC_9_125 b_9 NI_9 NS_125 0 -4.3389909020998042e-10
GC_9_126 b_9 NI_9 NS_126 0 -1.2075667431791703e-10
GC_9_127 b_9 NI_9 NS_127 0 -2.9066900451074458e-05
GC_9_128 b_9 NI_9 NS_128 0 -1.6185056304081157e-05
GC_9_129 b_9 NI_9 NS_129 0 2.8967501275689410e-05
GC_9_130 b_9 NI_9 NS_130 0 9.8864437548317125e-05
GC_9_131 b_9 NI_9 NS_131 0 2.9105534634349433e-07
GC_9_132 b_9 NI_9 NS_132 0 -1.4699361478671152e-04
GC_9_133 b_9 NI_9 NS_133 0 -1.6899605723007659e-04
GC_9_134 b_9 NI_9 NS_134 0 2.1090410161937582e-04
GC_9_135 b_9 NI_9 NS_135 0 2.7243933329700650e-04
GC_9_136 b_9 NI_9 NS_136 0 -2.1994524863147189e-04
GC_9_137 b_9 NI_9 NS_137 0 -2.5615043815384776e-05
GC_9_138 b_9 NI_9 NS_138 0 2.7760261132743516e-05
GC_9_139 b_9 NI_9 NS_139 0 -1.5191569682340475e-04
GC_9_140 b_9 NI_9 NS_140 0 -6.4140001402287675e-05
GC_9_141 b_9 NI_9 NS_141 0 -5.4693776224337297e-04
GC_9_142 b_9 NI_9 NS_142 0 4.9511188287266236e-04
GC_9_143 b_9 NI_9 NS_143 0 -7.8372628189903824e-05
GC_9_144 b_9 NI_9 NS_144 0 9.0352485037519400e-09
GC_9_145 b_9 NI_9 NS_145 0 3.0027635543379612e-10
GC_9_146 b_9 NI_9 NS_146 0 8.0533051169209490e-11
GC_9_147 b_9 NI_9 NS_147 0 -1.2560244001534094e-05
GC_9_148 b_9 NI_9 NS_148 0 -8.8756115141360160e-06
GC_9_149 b_9 NI_9 NS_149 0 -6.7306543200356368e-05
GC_9_150 b_9 NI_9 NS_150 0 -3.1843244852164748e-05
GC_9_151 b_9 NI_9 NS_151 0 -7.0775997640748224e-05
GC_9_152 b_9 NI_9 NS_152 0 1.1481870820477744e-04
GC_9_153 b_9 NI_9 NS_153 0 -1.3779794618074166e-04
GC_9_154 b_9 NI_9 NS_154 0 2.2324726951687525e-04
GC_9_155 b_9 NI_9 NS_155 0 3.5690612782554766e-04
GC_9_156 b_9 NI_9 NS_156 0 1.6256169662721184e-04
GC_9_157 b_9 NI_9 NS_157 0 -1.7294704816653741e-05
GC_9_158 b_9 NI_9 NS_158 0 -1.7940494242141562e-05
GC_9_159 b_9 NI_9 NS_159 0 1.0162292741235845e-04
GC_9_160 b_9 NI_9 NS_160 0 5.6167512419856885e-05
GC_9_161 b_9 NI_9 NS_161 0 -1.4552043550153169e-03
GC_9_162 b_9 NI_9 NS_162 0 -1.7225745455679026e-02
GC_9_163 b_9 NI_9 NS_163 0 1.1743969835844900e-02
GC_9_164 b_9 NI_9 NS_164 0 2.9971100202435237e-06
GC_9_165 b_9 NI_9 NS_165 0 -5.0997794839438991e-07
GC_9_166 b_9 NI_9 NS_166 0 -2.9633812622701210e-08
GC_9_167 b_9 NI_9 NS_167 0 3.0965325744638024e-03
GC_9_168 b_9 NI_9 NS_168 0 1.3051952351373155e-03
GC_9_169 b_9 NI_9 NS_169 0 -2.9261117836365956e-03
GC_9_170 b_9 NI_9 NS_170 0 -9.9123400414394391e-03
GC_9_171 b_9 NI_9 NS_171 0 6.3753024716567343e-04
GC_9_172 b_9 NI_9 NS_172 0 1.3628526886658164e-02
GC_9_173 b_9 NI_9 NS_173 0 1.7509591131423193e-02
GC_9_174 b_9 NI_9 NS_174 0 -2.3852005511625213e-02
GC_9_175 b_9 NI_9 NS_175 0 -3.3177959769706430e-02
GC_9_176 b_9 NI_9 NS_176 0 2.1222688981119585e-02
GC_9_177 b_9 NI_9 NS_177 0 4.0624004815291064e-03
GC_9_178 b_9 NI_9 NS_178 0 -2.1854429728248317e-03
GC_9_179 b_9 NI_9 NS_179 0 1.5119317255816096e-02
GC_9_180 b_9 NI_9 NS_180 0 5.6106549878242934e-03
GC_9_181 b_9 NI_9 NS_181 0 -2.8564000535021833e-01
GC_9_182 b_9 NI_9 NS_182 0 1.2097605224131186e-01
GC_9_183 b_9 NI_9 NS_183 0 7.0824868764034149e-03
GC_9_184 b_9 NI_9 NS_184 0 5.7464553201005421e-05
GC_9_185 b_9 NI_9 NS_185 0 1.3019123280207871e-06
GC_9_186 b_9 NI_9 NS_186 0 1.3695319201275195e-08
GC_9_187 b_9 NI_9 NS_187 0 3.0465780908413641e-02
GC_9_188 b_9 NI_9 NS_188 0 4.1090451193687956e-03
GC_9_189 b_9 NI_9 NS_189 0 -7.3763971968879884e-03
GC_9_190 b_9 NI_9 NS_190 0 2.2180118949485742e-02
GC_9_191 b_9 NI_9 NS_191 0 -1.7056202386691761e-02
GC_9_192 b_9 NI_9 NS_192 0 -1.8685516755535279e-02
GC_9_193 b_9 NI_9 NS_193 0 4.4665646733334327e-02
GC_9_194 b_9 NI_9 NS_194 0 1.4315031528793093e-02
GC_9_195 b_9 NI_9 NS_195 0 8.2000100274753462e-02
GC_9_196 b_9 NI_9 NS_196 0 3.1380062919035015e-02
GC_9_197 b_9 NI_9 NS_197 0 -1.0089093262826811e-02
GC_9_198 b_9 NI_9 NS_198 0 -4.9101466682490462e-03
GC_9_199 b_9 NI_9 NS_199 0 -2.1483627566485634e-02
GC_9_200 b_9 NI_9 NS_200 0 -4.8833390641502767e-03
GC_9_201 b_9 NI_9 NS_201 0 2.2267872707234574e-02
GC_9_202 b_9 NI_9 NS_202 0 8.9573222676479283e-03
GC_9_203 b_9 NI_9 NS_203 0 -1.1409899591953671e-02
GC_9_204 b_9 NI_9 NS_204 0 -5.3357066209218500e-06
GC_9_205 b_9 NI_9 NS_205 0 -9.5823209710118688e-08
GC_9_206 b_9 NI_9 NS_206 0 -1.2410084341503947e-09
GC_9_207 b_9 NI_9 NS_207 0 -3.3142115015536498e-03
GC_9_208 b_9 NI_9 NS_208 0 -2.3908938231856640e-03
GC_9_209 b_9 NI_9 NS_209 0 2.7265908031992754e-03
GC_9_210 b_9 NI_9 NS_210 0 1.1171998927836282e-02
GC_9_211 b_9 NI_9 NS_211 0 -3.5268546161212048e-04
GC_9_212 b_9 NI_9 NS_212 0 -1.7759690683797038e-02
GC_9_213 b_9 NI_9 NS_213 0 -2.2020323746107354e-02
GC_9_214 b_9 NI_9 NS_214 0 2.1327619534720021e-02
GC_9_215 b_9 NI_9 NS_215 0 2.8910205978017089e-02
GC_9_216 b_9 NI_9 NS_216 0 -1.8399093090247787e-02
GC_9_217 b_9 NI_9 NS_217 0 -2.4511212692121453e-03
GC_9_218 b_9 NI_9 NS_218 0 1.4222330861585685e-03
GC_9_219 b_9 NI_9 NS_219 0 -1.7818694330355617e-02
GC_9_220 b_9 NI_9 NS_220 0 -7.1267653599122720e-03
GC_9_221 b_9 NI_9 NS_221 0 -8.2288462485228892e-02
GC_9_222 b_9 NI_9 NS_222 0 6.5322022208423369e-02
GC_9_223 b_9 NI_9 NS_223 0 -1.0307114067292350e-02
GC_9_224 b_9 NI_9 NS_224 0 -2.3858537991241015e-06
GC_9_225 b_9 NI_9 NS_225 0 1.6335227407096012e-08
GC_9_226 b_9 NI_9 NS_226 0 1.6410075214052320e-09
GC_9_227 b_9 NI_9 NS_227 0 -3.9597027682551818e-04
GC_9_228 b_9 NI_9 NS_228 0 -1.4000566629706723e-03
GC_9_229 b_9 NI_9 NS_229 0 -6.9917489107977192e-03
GC_9_230 b_9 NI_9 NS_230 0 -3.7822426750812022e-03
GC_9_231 b_9 NI_9 NS_231 0 -9.0594500218976869e-03
GC_9_232 b_9 NI_9 NS_232 0 1.3121191967177091e-02
GC_9_233 b_9 NI_9 NS_233 0 -1.5240953623193528e-02
GC_9_234 b_9 NI_9 NS_234 0 2.8718755465780857e-02
GC_9_235 b_9 NI_9 NS_235 0 4.5110989413125351e-02
GC_9_236 b_9 NI_9 NS_236 0 1.6488628398956279e-02
GC_9_237 b_9 NI_9 NS_237 0 -2.2090750093192433e-03
GC_9_238 b_9 NI_9 NS_238 0 -1.3391802446242637e-03
GC_9_239 b_9 NI_9 NS_239 0 1.2863710735179640e-02
GC_9_240 b_9 NI_9 NS_240 0 6.9572427906184732e-03
GD_9_1 b_9 NI_9 NA_1 0 -2.3046838042988428e-06
GD_9_2 b_9 NI_9 NA_2 0 -1.0364077490992301e-05
GD_9_3 b_9 NI_9 NA_3 0 -9.6649620208644518e-06
GD_9_4 b_9 NI_9 NA_4 0 1.1836312685296782e-05
GD_9_5 b_9 NI_9 NA_5 0 -6.8663486479112097e-05
GD_9_6 b_9 NI_9 NA_6 0 4.2508811434067072e-06
GD_9_7 b_9 NI_9 NA_7 0 7.9447560527822305e-05
GD_9_8 b_9 NI_9 NA_8 0 -4.8736496901073459e-05
GD_9_9 b_9 NI_9 NA_9 0 -6.3838861587847528e-03
GD_9_10 b_9 NI_9 NA_10 0 5.6719418020400640e-02
GD_9_11 b_9 NI_9 NA_11 0 6.2259707324474160e-03
GD_9_12 b_9 NI_9 NA_12 0 2.3474521306974614e-03
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 2.0691192645035641e-05
GC_10_2 b_10 NI_10 NS_2 0 -5.0103725317025265e-06
GC_10_3 b_10 NI_10 NS_3 0 9.9579002882639107e-07
GC_10_4 b_10 NI_10 NS_4 0 -5.5012620759976678e-09
GC_10_5 b_10 NI_10 NS_5 0 -2.5924610671857899e-11
GC_10_6 b_10 NI_10 NS_6 0 -1.2333465505248263e-12
GC_10_7 b_10 NI_10 NS_7 0 -1.3186728539131600e-06
GC_10_8 b_10 NI_10 NS_8 0 -1.6811812314031950e-06
GC_10_9 b_10 NI_10 NS_9 0 -1.8034084834098961e-06
GC_10_10 b_10 NI_10 NS_10 0 1.3687020187671202e-07
GC_10_11 b_10 NI_10 NS_11 0 -2.4181479820275404e-06
GC_10_12 b_10 NI_10 NS_12 0 2.2165537874112005e-06
GC_10_13 b_10 NI_10 NS_13 0 -3.9553009572672881e-06
GC_10_14 b_10 NI_10 NS_14 0 -2.1597698257946784e-06
GC_10_15 b_10 NI_10 NS_15 0 1.2334496055865885e-06
GC_10_16 b_10 NI_10 NS_16 0 8.3243088679273928e-06
GC_10_17 b_10 NI_10 NS_17 0 -3.9465728986527335e-07
GC_10_18 b_10 NI_10 NS_18 0 -1.7930156656051618e-06
GC_10_19 b_10 NI_10 NS_19 0 -3.7109478826758774e-07
GC_10_20 b_10 NI_10 NS_20 0 1.7920033006054919e-07
GC_10_21 b_10 NI_10 NS_21 0 5.6957081317909300e-06
GC_10_22 b_10 NI_10 NS_22 0 1.3939728452359954e-06
GC_10_23 b_10 NI_10 NS_23 0 -8.6838687784237528e-07
GC_10_24 b_10 NI_10 NS_24 0 3.5299819664848692e-09
GC_10_25 b_10 NI_10 NS_25 0 5.0050043093124610e-11
GC_10_26 b_10 NI_10 NS_26 0 -5.2578457448036197e-13
GC_10_27 b_10 NI_10 NS_27 0 -4.1796105125187352e-07
GC_10_28 b_10 NI_10 NS_28 0 -3.4615033616429947e-07
GC_10_29 b_10 NI_10 NS_29 0 -2.5593583049412240e-07
GC_10_30 b_10 NI_10 NS_30 0 2.1882227245907543e-07
GC_10_31 b_10 NI_10 NS_31 0 -7.9356267823765801e-07
GC_10_32 b_10 NI_10 NS_32 0 -6.7751045776571503e-07
GC_10_33 b_10 NI_10 NS_33 0 -2.5395447523424835e-06
GC_10_34 b_10 NI_10 NS_34 0 -5.4510433517351305e-08
GC_10_35 b_10 NI_10 NS_35 0 3.9405138171717458e-07
GC_10_36 b_10 NI_10 NS_36 0 3.5255764609214087e-06
GC_10_37 b_10 NI_10 NS_37 0 1.6398895174765606e-07
GC_10_38 b_10 NI_10 NS_38 0 -8.5380561359332002e-07
GC_10_39 b_10 NI_10 NS_39 0 -5.5850074828396323e-07
GC_10_40 b_10 NI_10 NS_40 0 2.6967844553775405e-07
GC_10_41 b_10 NI_10 NS_41 0 7.9171037199105126e-06
GC_10_42 b_10 NI_10 NS_42 0 -6.3407564546309457e-06
GC_10_43 b_10 NI_10 NS_43 0 4.7284624734746593e-07
GC_10_44 b_10 NI_10 NS_44 0 6.3751303999630724e-09
GC_10_45 b_10 NI_10 NS_45 0 -1.7572035765913081e-10
GC_10_46 b_10 NI_10 NS_46 0 8.2824505278467708e-12
GC_10_47 b_10 NI_10 NS_47 0 2.1357709326045701e-06
GC_10_48 b_10 NI_10 NS_48 0 -1.0057450487562881e-06
GC_10_49 b_10 NI_10 NS_49 0 2.8511711731659124e-06
GC_10_50 b_10 NI_10 NS_50 0 -1.3362567021655675e-06
GC_10_51 b_10 NI_10 NS_51 0 -2.5357602959870763e-07
GC_10_52 b_10 NI_10 NS_52 0 -3.4595027231948687e-06
GC_10_53 b_10 NI_10 NS_53 0 6.9393794367287138e-06
GC_10_54 b_10 NI_10 NS_54 0 -9.0892538037460291e-06
GC_10_55 b_10 NI_10 NS_55 0 -2.3895808695745000e-05
GC_10_56 b_10 NI_10 NS_56 0 -2.8566940611408663e-06
GC_10_57 b_10 NI_10 NS_57 0 5.9695861239536610e-06
GC_10_58 b_10 NI_10 NS_58 0 3.0591198151023560e-07
GC_10_59 b_10 NI_10 NS_59 0 -2.6278121901205887e-06
GC_10_60 b_10 NI_10 NS_60 0 1.4080032469442654e-06
GC_10_61 b_10 NI_10 NS_61 0 2.2539397004691460e-05
GC_10_62 b_10 NI_10 NS_62 0 -5.1374414550380930e-06
GC_10_63 b_10 NI_10 NS_63 0 3.6837557528412096e-07
GC_10_64 b_10 NI_10 NS_64 0 -8.1493388263504864e-09
GC_10_65 b_10 NI_10 NS_65 0 1.7606318337517197e-10
GC_10_66 b_10 NI_10 NS_66 0 -9.7889993222244253e-12
GC_10_67 b_10 NI_10 NS_67 0 -1.2142846311484010e-06
GC_10_68 b_10 NI_10 NS_68 0 -9.1145976239723391e-07
GC_10_69 b_10 NI_10 NS_69 0 -1.3989593425770613e-06
GC_10_70 b_10 NI_10 NS_70 0 -4.6250371912142176e-08
GC_10_71 b_10 NI_10 NS_71 0 -2.2030210113061749e-06
GC_10_72 b_10 NI_10 NS_72 0 2.2974992680673565e-08
GC_10_73 b_10 NI_10 NS_73 0 -4.7812860362606422e-06
GC_10_74 b_10 NI_10 NS_74 0 -4.5199504293283811e-07
GC_10_75 b_10 NI_10 NS_75 0 1.0107465530615555e-06
GC_10_76 b_10 NI_10 NS_76 0 7.1426260740383244e-06
GC_10_77 b_10 NI_10 NS_77 0 -3.5884008698306691e-07
GC_10_78 b_10 NI_10 NS_78 0 -1.8237682509264879e-06
GC_10_79 b_10 NI_10 NS_79 0 -1.0678367944055677e-06
GC_10_80 b_10 NI_10 NS_80 0 -3.9178573657480014e-07
GC_10_81 b_10 NI_10 NS_81 0 3.0487037429346065e-04
GC_10_82 b_10 NI_10 NS_82 0 -2.6795572098506549e-04
GC_10_83 b_10 NI_10 NS_83 0 4.3029734600109594e-05
GC_10_84 b_10 NI_10 NS_84 0 1.3274604688140648e-08
GC_10_85 b_10 NI_10 NS_85 0 -1.3641655192854776e-10
GC_10_86 b_10 NI_10 NS_86 0 1.3413385345429198e-11
GC_10_87 b_10 NI_10 NS_87 0 1.6671641423273872e-06
GC_10_88 b_10 NI_10 NS_88 0 7.0535561375674987e-06
GC_10_89 b_10 NI_10 NS_89 0 3.2663510671505017e-05
GC_10_90 b_10 NI_10 NS_90 0 2.1834098818946168e-05
GC_10_91 b_10 NI_10 NS_91 0 4.5895158745534811e-05
GC_10_92 b_10 NI_10 NS_92 0 -5.6019429034346753e-05
GC_10_93 b_10 NI_10 NS_93 0 7.3005783910184185e-05
GC_10_94 b_10 NI_10 NS_94 0 -1.2465399084920120e-04
GC_10_95 b_10 NI_10 NS_95 0 -1.8515862615629223e-04
GC_10_96 b_10 NI_10 NS_96 0 -7.4483189885910298e-05
GC_10_97 b_10 NI_10 NS_97 0 7.5436302491450120e-06
GC_10_98 b_10 NI_10 NS_98 0 3.5790286716566706e-06
GC_10_99 b_10 NI_10 NS_99 0 -5.3931860971922990e-05
GC_10_100 b_10 NI_10 NS_100 0 -3.1184917521333187e-05
GC_10_101 b_10 NI_10 NS_101 0 2.7705412605606467e-04
GC_10_102 b_10 NI_10 NS_102 0 -1.2387381110394262e-05
GC_10_103 b_10 NI_10 NS_103 0 -9.4633644510018811e-06
GC_10_104 b_10 NI_10 NS_104 0 6.0728928849303053e-08
GC_10_105 b_10 NI_10 NS_105 0 -3.1805478442232313e-10
GC_10_106 b_10 NI_10 NS_106 0 9.7939357125659492e-12
GC_10_107 b_10 NI_10 NS_107 0 -5.8027997103121449e-07
GC_10_108 b_10 NI_10 NS_108 0 -1.5576453625917426e-05
GC_10_109 b_10 NI_10 NS_109 0 -9.7465693696454706e-06
GC_10_110 b_10 NI_10 NS_110 0 -2.0953108988563895e-05
GC_10_111 b_10 NI_10 NS_111 0 -3.7868615365935905e-05
GC_10_112 b_10 NI_10 NS_112 0 -1.9889341190172082e-05
GC_10_113 b_10 NI_10 NS_113 0 -7.5415010438222032e-05
GC_10_114 b_10 NI_10 NS_114 0 -7.9253549038721613e-05
GC_10_115 b_10 NI_10 NS_115 0 -7.5278067049049913e-05
GC_10_116 b_10 NI_10 NS_116 0 2.2097702663396150e-04
GC_10_117 b_10 NI_10 NS_117 0 1.5306009280475845e-05
GC_10_118 b_10 NI_10 NS_118 0 -5.7665549226226596e-05
GC_10_119 b_10 NI_10 NS_119 0 -4.7284458127262936e-06
GC_10_120 b_10 NI_10 NS_120 0 1.3857052543977712e-05
GC_10_121 b_10 NI_10 NS_121 0 -5.4700630535832646e-04
GC_10_122 b_10 NI_10 NS_122 0 4.9510290645232323e-04
GC_10_123 b_10 NI_10 NS_123 0 -7.8370283293243732e-05
GC_10_124 b_10 NI_10 NS_124 0 9.0303565402375209e-09
GC_10_125 b_10 NI_10 NS_125 0 3.0029232396522675e-10
GC_10_126 b_10 NI_10 NS_126 0 8.0533178539707850e-11
GC_10_127 b_10 NI_10 NS_127 0 -1.2542339816083124e-05
GC_10_128 b_10 NI_10 NS_128 0 -8.8614482057009069e-06
GC_10_129 b_10 NI_10 NS_129 0 -6.7281719947213399e-05
GC_10_130 b_10 NI_10 NS_130 0 -3.1840155469184652e-05
GC_10_131 b_10 NI_10 NS_131 0 -7.0761527061274422e-05
GC_10_132 b_10 NI_10 NS_132 0 1.1477601947172771e-04
GC_10_133 b_10 NI_10 NS_133 0 -1.3778574511320684e-04
GC_10_134 b_10 NI_10 NS_134 0 2.2321532242238303e-04
GC_10_135 b_10 NI_10 NS_135 0 3.5686973517631441e-04
GC_10_136 b_10 NI_10 NS_136 0 1.6255711268310831e-04
GC_10_137 b_10 NI_10 NS_137 0 -1.7291809137883002e-05
GC_10_138 b_10 NI_10 NS_138 0 -1.7943729692750163e-05
GC_10_139 b_10 NI_10 NS_139 0 1.0162026247651601e-04
GC_10_140 b_10 NI_10 NS_140 0 5.6164393053275900e-05
GC_10_141 b_10 NI_10 NS_141 0 1.1295688141061621e-04
GC_10_142 b_10 NI_10 NS_142 0 8.2945478198952319e-05
GC_10_143 b_10 NI_10 NS_143 0 -9.5451576300802982e-05
GC_10_144 b_10 NI_10 NS_144 0 -1.1416672418962381e-07
GC_10_145 b_10 NI_10 NS_145 0 -4.3387028835237779e-10
GC_10_146 b_10 NI_10 NS_146 0 -1.2075594495359905e-10
GC_10_147 b_10 NI_10 NS_147 0 -2.9066603556922403e-05
GC_10_148 b_10 NI_10 NS_148 0 -1.6184682487769786e-05
GC_10_149 b_10 NI_10 NS_149 0 2.8967662116702258e-05
GC_10_150 b_10 NI_10 NS_150 0 9.8864603596073548e-05
GC_10_151 b_10 NI_10 NS_151 0 2.9205672354381258e-07
GC_10_152 b_10 NI_10 NS_152 0 -1.4699327668318588e-04
GC_10_153 b_10 NI_10 NS_153 0 -1.6899334006190416e-04
GC_10_154 b_10 NI_10 NS_154 0 2.1090499922032390e-04
GC_10_155 b_10 NI_10 NS_155 0 2.7243837506968387e-04
GC_10_156 b_10 NI_10 NS_156 0 -2.1995137041058165e-04
GC_10_157 b_10 NI_10 NS_157 0 -2.5614901102688424e-05
GC_10_158 b_10 NI_10 NS_158 0 2.7761634545572412e-05
GC_10_159 b_10 NI_10 NS_159 0 -1.5191631401453615e-04
GC_10_160 b_10 NI_10 NS_160 0 -6.4140668593203078e-05
GC_10_161 b_10 NI_10 NS_161 0 -2.8564002869835953e-01
GC_10_162 b_10 NI_10 NS_162 0 1.2097603305065899e-01
GC_10_163 b_10 NI_10 NS_163 0 7.0824901082775556e-03
GC_10_164 b_10 NI_10 NS_164 0 5.7464559620841052e-05
GC_10_165 b_10 NI_10 NS_165 0 1.3019119291359466e-06
GC_10_166 b_10 NI_10 NS_166 0 1.3695376744659098e-08
GC_10_167 b_10 NI_10 NS_167 0 3.0465752107894494e-02
GC_10_168 b_10 NI_10 NS_168 0 4.1090314984954775e-03
GC_10_169 b_10 NI_10 NS_169 0 -7.3764400359566393e-03
GC_10_170 b_10 NI_10 NS_170 0 2.2180134597622438e-02
GC_10_171 b_10 NI_10 NS_171 0 -1.7056159182509537e-02
GC_10_172 b_10 NI_10 NS_172 0 -1.8685423420253294e-02
GC_10_173 b_10 NI_10 NS_173 0 4.4665768057227523e-02
GC_10_174 b_10 NI_10 NS_174 0 1.4315101301281068e-02
GC_10_175 b_10 NI_10 NS_175 0 8.2000021972368164e-02
GC_10_176 b_10 NI_10 NS_176 0 3.1379880889758752e-02
GC_10_177 b_10 NI_10 NS_177 0 -1.0089045586302189e-02
GC_10_178 b_10 NI_10 NS_178 0 -4.9101180119019480e-03
GC_10_179 b_10 NI_10 NS_179 0 -2.1483638113516324e-02
GC_10_180 b_10 NI_10 NS_180 0 -4.8833464259343835e-03
GC_10_181 b_10 NI_10 NS_181 0 -1.4552043550153688e-03
GC_10_182 b_10 NI_10 NS_182 0 -1.7225745455679019e-02
GC_10_183 b_10 NI_10 NS_183 0 1.1743969835844897e-02
GC_10_184 b_10 NI_10 NS_184 0 2.9971100202442093e-06
GC_10_185 b_10 NI_10 NS_185 0 -5.0997794839438938e-07
GC_10_186 b_10 NI_10 NS_186 0 -2.9633812622700856e-08
GC_10_187 b_10 NI_10 NS_187 0 3.0965325744638015e-03
GC_10_188 b_10 NI_10 NS_188 0 1.3051952351373164e-03
GC_10_189 b_10 NI_10 NS_189 0 -2.9261117836365843e-03
GC_10_190 b_10 NI_10 NS_190 0 -9.9123400414394356e-03
GC_10_191 b_10 NI_10 NS_191 0 6.3753024716568221e-04
GC_10_192 b_10 NI_10 NS_192 0 1.3628526886658157e-02
GC_10_193 b_10 NI_10 NS_193 0 1.7509591131423207e-02
GC_10_194 b_10 NI_10 NS_194 0 -2.3852005511625217e-02
GC_10_195 b_10 NI_10 NS_195 0 -3.3177959769706437e-02
GC_10_196 b_10 NI_10 NS_196 0 2.1222688981119564e-02
GC_10_197 b_10 NI_10 NS_197 0 4.0624004815291107e-03
GC_10_198 b_10 NI_10 NS_198 0 -2.1854429728248282e-03
GC_10_199 b_10 NI_10 NS_199 0 1.5119317255816101e-02
GC_10_200 b_10 NI_10 NS_200 0 5.6106549878242934e-03
GC_10_201 b_10 NI_10 NS_201 0 -8.2288464694788621e-02
GC_10_202 b_10 NI_10 NS_202 0 6.5322022997245599e-02
GC_10_203 b_10 NI_10 NS_203 0 -1.0307114159569586e-02
GC_10_204 b_10 NI_10 NS_204 0 -2.3858535076404995e-06
GC_10_205 b_10 NI_10 NS_205 0 1.6335225056678213e-08
GC_10_206 b_10 NI_10 NS_206 0 1.6410076036530494e-09
GC_10_207 b_10 NI_10 NS_207 0 -3.9597042998080106e-04
GC_10_208 b_10 NI_10 NS_208 0 -1.4000566242028801e-03
GC_10_209 b_10 NI_10 NS_209 0 -6.9917490294911103e-03
GC_10_210 b_10 NI_10 NS_210 0 -3.7822424126441562e-03
GC_10_211 b_10 NI_10 NS_211 0 -9.0594497462318513e-03
GC_10_212 b_10 NI_10 NS_212 0 1.3121192334235773e-02
GC_10_213 b_10 NI_10 NS_213 0 -1.5240953398823445e-02
GC_10_214 b_10 NI_10 NS_214 0 2.8718756215261588e-02
GC_10_215 b_10 NI_10 NS_215 0 4.5110990633982911e-02
GC_10_216 b_10 NI_10 NS_216 0 1.6488627481823045e-02
GC_10_217 b_10 NI_10 NS_217 0 -2.2090752244941026e-03
GC_10_218 b_10 NI_10 NS_218 0 -1.3391800354162627e-03
GC_10_219 b_10 NI_10 NS_219 0 1.2863710852294810e-02
GC_10_220 b_10 NI_10 NS_220 0 6.9572427257932820e-03
GC_10_221 b_10 NI_10 NS_221 0 2.2274168818736589e-02
GC_10_222 b_10 NI_10 NS_222 0 8.9558653696552703e-03
GC_10_223 b_10 NI_10 NS_223 0 -1.1409760318263787e-02
GC_10_224 b_10 NI_10 NS_224 0 -5.3360829798493087e-06
GC_10_225 b_10 NI_10 NS_225 0 -9.5822584229290003e-08
GC_10_226 b_10 NI_10 NS_226 0 -1.2412247368594177e-09
GC_10_227 b_10 NI_10 NS_227 0 -3.3143876880205843e-03
GC_10_228 b_10 NI_10 NS_228 0 -2.3911424295166065e-03
GC_10_229 b_10 NI_10 NS_229 0 2.7261772326534050e-03
GC_10_230 b_10 NI_10 NS_230 0 1.1171778349198237e-02
GC_10_231 b_10 NI_10 NS_231 0 -3.5307692784337382e-04
GC_10_232 b_10 NI_10 NS_232 0 -1.7759589703801114e-02
GC_10_233 b_10 NI_10 NS_233 0 -2.2020926253592869e-02
GC_10_234 b_10 NI_10 NS_234 0 2.1326548385709781e-02
GC_10_235 b_10 NI_10 NS_235 0 2.8908354578924184e-02
GC_10_236 b_10 NI_10 NS_236 0 -1.8397055755763534e-02
GC_10_237 b_10 NI_10 NS_237 0 -2.4507582349978271e-03
GC_10_238 b_10 NI_10 NS_238 0 1.4218496269307454e-03
GC_10_239 b_10 NI_10 NS_239 0 -1.7818879423500012e-02
GC_10_240 b_10 NI_10 NS_240 0 -7.1265651977145709e-03
GD_10_1 b_10 NI_10 NA_1 0 -1.0364067804234872e-05
GD_10_2 b_10 NI_10 NA_2 0 -2.2799324788609173e-06
GD_10_3 b_10 NI_10 NA_3 0 1.1835727122594619e-05
GD_10_4 b_10 NI_10 NA_4 0 -9.6644135979843025e-06
GD_10_5 b_10 NI_10 NA_5 0 4.2506841281317482e-06
GD_10_6 b_10 NI_10 NA_6 0 -6.8166037152082881e-05
GD_10_7 b_10 NI_10 NA_7 0 -4.8688362054564848e-05
GD_10_8 b_10 NI_10 NA_8 0 7.9448663276090995e-05
GD_10_9 b_10 NI_10 NA_9 0 5.6719405138710724e-02
GD_10_10 b_10 NI_10 NA_10 0 -6.3838861587848048e-03
GD_10_11 b_10 NI_10 NA_11 0 2.3474522237801219e-03
GD_10_12 b_10 NI_10 NA_12 0 6.2239325459215612e-03
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 7.3320635119256587e-06
GC_11_2 b_11 NI_11 NS_2 0 -2.5195975340381514e-06
GC_11_3 b_11 NI_11 NS_3 0 1.5308897887445786e-07
GC_11_4 b_11 NI_11 NS_4 0 -4.0110863413750007e-09
GC_11_5 b_11 NI_11 NS_5 0 1.6388396100514402e-10
GC_11_6 b_11 NI_11 NS_6 0 -1.2217730138203231e-11
GC_11_7 b_11 NI_11 NS_7 0 -3.1665108632059984e-07
GC_11_8 b_11 NI_11 NS_8 0 -2.3698639691391637e-07
GC_11_9 b_11 NI_11 NS_9 0 -7.6390735673513434e-08
GC_11_10 b_11 NI_11 NS_10 0 9.2605558448058393e-08
GC_11_11 b_11 NI_11 NS_11 0 -7.8248627929574157e-07
GC_11_12 b_11 NI_11 NS_12 0 -4.1603027580655022e-07
GC_11_13 b_11 NI_11 NS_13 0 -9.7686390662721081e-07
GC_11_14 b_11 NI_11 NS_14 0 4.5613993082163198e-07
GC_11_15 b_11 NI_11 NS_15 0 2.6679549206624469e-07
GC_11_16 b_11 NI_11 NS_16 0 3.0984663476436894e-07
GC_11_17 b_11 NI_11 NS_17 0 -1.5150718620451382e-07
GC_11_18 b_11 NI_11 NS_18 0 -3.1207019848291174e-07
GC_11_19 b_11 NI_11 NS_19 0 -8.8431495986839893e-07
GC_11_20 b_11 NI_11 NS_20 0 -4.0325457058024189e-07
GC_11_21 b_11 NI_11 NS_21 0 -6.3363880136133440e-07
GC_11_22 b_11 NI_11 NS_22 0 -6.2720115017379480e-07
GC_11_23 b_11 NI_11 NS_23 0 -7.3992786262203136e-08
GC_11_24 b_11 NI_11 NS_24 0 4.6611086238831629e-09
GC_11_25 b_11 NI_11 NS_25 0 -1.7625101281892913e-10
GC_11_26 b_11 NI_11 NS_26 0 1.2487331173354975e-11
GC_11_27 b_11 NI_11 NS_27 0 9.0959400306971589e-07
GC_11_28 b_11 NI_11 NS_28 0 -8.4397985550099232e-07
GC_11_29 b_11 NI_11 NS_29 0 1.2588120029791293e-06
GC_11_30 b_11 NI_11 NS_30 0 -1.6665121740671311e-07
GC_11_31 b_11 NI_11 NS_31 0 -1.8644366632321290e-07
GC_11_32 b_11 NI_11 NS_32 0 -1.1990626431680742e-06
GC_11_33 b_11 NI_11 NS_33 0 2.8924862847882481e-06
GC_11_34 b_11 NI_11 NS_34 0 -4.1240289707414356e-06
GC_11_35 b_11 NI_11 NS_35 0 -8.7582609696884623e-06
GC_11_36 b_11 NI_11 NS_36 0 4.8511192175356670e-08
GC_11_37 b_11 NI_11 NS_37 0 2.1514258795915655e-06
GC_11_38 b_11 NI_11 NS_38 0 -3.9711471781788352e-07
GC_11_39 b_11 NI_11 NS_39 0 -8.8852819063033029e-07
GC_11_40 b_11 NI_11 NS_40 0 8.3679128487712826e-07
GC_11_41 b_11 NI_11 NS_41 0 5.6551598473692761e-06
GC_11_42 b_11 NI_11 NS_42 0 1.4060292192518661e-06
GC_11_43 b_11 NI_11 NS_43 0 -8.7122206510353899e-07
GC_11_44 b_11 NI_11 NS_44 0 3.5286918979685891e-09
GC_11_45 b_11 NI_11 NS_45 0 5.0023247508158485e-11
GC_11_46 b_11 NI_11 NS_46 0 -5.2267735037564020e-13
GC_11_47 b_11 NI_11 NS_47 0 -4.1810709630590889e-07
GC_11_48 b_11 NI_11 NS_48 0 -3.4338249522833054e-07
GC_11_49 b_11 NI_11 NS_49 0 -2.5300981267322165e-07
GC_11_50 b_11 NI_11 NS_50 0 2.2179396704874123e-07
GC_11_51 b_11 NI_11 NS_51 0 -7.9231987671029082e-07
GC_11_52 b_11 NI_11 NS_52 0 -6.7635771263564308e-07
GC_11_53 b_11 NI_11 NS_53 0 -2.5328283348336267e-06
GC_11_54 b_11 NI_11 NS_54 0 -3.6653809702571234e-08
GC_11_55 b_11 NI_11 NS_55 0 4.1620972890806052e-07
GC_11_56 b_11 NI_11 NS_56 0 3.4991362122943513e-06
GC_11_57 b_11 NI_11 NS_57 0 1.5924453386224219e-07
GC_11_58 b_11 NI_11 NS_58 0 -8.5029828952198551e-07
GC_11_59 b_11 NI_11 NS_59 0 -5.6118821927222438e-07
GC_11_60 b_11 NI_11 NS_60 0 2.6713390470856361e-07
GC_11_61 b_11 NI_11 NS_61 0 2.0604783570485272e-05
GC_11_62 b_11 NI_11 NS_62 0 -4.9935577892746953e-06
GC_11_63 b_11 NI_11 NS_63 0 9.9303255957749384e-07
GC_11_64 b_11 NI_11 NS_64 0 -5.4984994852284512e-09
GC_11_65 b_11 NI_11 NS_65 0 -2.5967349989590495e-11
GC_11_66 b_11 NI_11 NS_66 0 -1.2308357573067289e-12
GC_11_67 b_11 NI_11 NS_67 0 -1.3115854121946019e-06
GC_11_68 b_11 NI_11 NS_68 0 -1.6746877718185682e-06
GC_11_69 b_11 NI_11 NS_69 0 -1.7990787589851606e-06
GC_11_70 b_11 NI_11 NS_70 0 1.3848526790152708e-07
GC_11_71 b_11 NI_11 NS_71 0 -2.4070258456460363e-06
GC_11_72 b_11 NI_11 NS_72 0 2.2075749818517675e-06
GC_11_73 b_11 NI_11 NS_73 0 -3.9348572312664450e-06
GC_11_74 b_11 NI_11 NS_74 0 -2.1436724758979169e-06
GC_11_75 b_11 NI_11 NS_75 0 1.2291044267706858e-06
GC_11_76 b_11 NI_11 NS_76 0 8.2805547210346288e-06
GC_11_77 b_11 NI_11 NS_77 0 -3.9212386294308005e-07
GC_11_78 b_11 NI_11 NS_78 0 -1.7846281617456251e-06
GC_11_79 b_11 NI_11 NS_79 0 -3.6943300591297286e-07
GC_11_80 b_11 NI_11 NS_80 0 1.7726585106474835e-07
GC_11_81 b_11 NI_11 NS_81 0 -7.8387633795357336e-05
GC_11_82 b_11 NI_11 NS_82 0 1.3376513979630602e-05
GC_11_83 b_11 NI_11 NS_83 0 -1.3932390781742812e-06
GC_11_84 b_11 NI_11 NS_84 0 -1.3101589234341075e-08
GC_11_85 b_11 NI_11 NS_85 0 2.6342332131966400e-10
GC_11_86 b_11 NI_11 NS_86 0 -1.7097214224897069e-11
GC_11_87 b_11 NI_11 NS_87 0 -1.5337478877606512e-06
GC_11_88 b_11 NI_11 NS_88 0 3.6436028049769349e-06
GC_11_89 b_11 NI_11 NS_89 0 1.6182179152795021e-06
GC_11_90 b_11 NI_11 NS_90 0 8.9333690559039340e-06
GC_11_91 b_11 NI_11 NS_91 0 1.0127223119705450e-05
GC_11_92 b_11 NI_11 NS_92 0 3.9280734830836244e-06
GC_11_93 b_11 NI_11 NS_93 0 1.3025656661282496e-05
GC_11_94 b_11 NI_11 NS_94 0 2.9985128949224401e-05
GC_11_95 b_11 NI_11 NS_95 0 3.6900818534456587e-05
GC_11_96 b_11 NI_11 NS_96 0 -6.0920660378450721e-05
GC_11_97 b_11 NI_11 NS_97 0 -6.8802555083617864e-06
GC_11_98 b_11 NI_11 NS_98 0 1.5061063930782399e-05
GC_11_99 b_11 NI_11 NS_99 0 -1.5084569436846750e-06
GC_11_100 b_11 NI_11 NS_100 0 -4.9192660684890377e-06
GC_11_101 b_11 NI_11 NS_101 0 6.1496279513552165e-05
GC_11_102 b_11 NI_11 NS_102 0 -4.0968510987818591e-05
GC_11_103 b_11 NI_11 NS_103 0 7.0419746182253181e-06
GC_11_104 b_11 NI_11 NS_104 0 -1.5383549888936983e-08
GC_11_105 b_11 NI_11 NS_105 0 -2.8243307674114301e-11
GC_11_106 b_11 NI_11 NS_106 0 2.8286725162686319e-13
GC_11_107 b_11 NI_11 NS_107 0 -9.0513698786881370e-07
GC_11_108 b_11 NI_11 NS_108 0 -1.4038337236668178e-06
GC_11_109 b_11 NI_11 NS_109 0 1.3494589898731776e-06
GC_11_110 b_11 NI_11 NS_110 0 2.2662979080980320e-06
GC_11_111 b_11 NI_11 NS_111 0 2.9358433687896330e-06
GC_11_112 b_11 NI_11 NS_112 0 -3.4739240237580973e-06
GC_11_113 b_11 NI_11 NS_113 0 7.8879420402160429e-06
GC_11_114 b_11 NI_11 NS_114 0 -1.6508174204483424e-05
GC_11_115 b_11 NI_11 NS_115 0 -2.6704648623799613e-05
GC_11_116 b_11 NI_11 NS_116 0 -4.5356286417976216e-06
GC_11_117 b_11 NI_11 NS_117 0 2.5910947336487047e-06
GC_11_118 b_11 NI_11 NS_118 0 -5.5008396330162355e-07
GC_11_119 b_11 NI_11 NS_119 0 -7.0849924155030199e-06
GC_11_120 b_11 NI_11 NS_120 0 -3.6888955466615565e-06
GC_11_121 b_11 NI_11 NS_121 0 2.7679949342524380e-04
GC_11_122 b_11 NI_11 NS_122 0 -1.2052535487328645e-05
GC_11_123 b_11 NI_11 NS_123 0 -9.5072292852244710e-06
GC_11_124 b_11 NI_11 NS_124 0 6.0829925204118557e-08
GC_11_125 b_11 NI_11 NS_125 0 -3.1352473073178202e-10
GC_11_126 b_11 NI_11 NS_126 0 8.9636914427517287e-12
GC_11_127 b_11 NI_11 NS_127 0 -6.6497575405703954e-07
GC_11_128 b_11 NI_11 NS_128 0 -1.5571150353444075e-05
GC_11_129 b_11 NI_11 NS_129 0 -9.8226342515322370e-06
GC_11_130 b_11 NI_11 NS_130 0 -2.0899212907400959e-05
GC_11_131 b_11 NI_11 NS_131 0 -3.7936282468604853e-05
GC_11_132 b_11 NI_11 NS_132 0 -1.9764556206236927e-05
GC_11_133 b_11 NI_11 NS_133 0 -7.5725766781296536e-05
GC_11_134 b_11 NI_11 NS_134 0 -7.8970931124765396e-05
GC_11_135 b_11 NI_11 NS_135 0 -7.4379445021931714e-05
GC_11_136 b_11 NI_11 NS_136 0 2.2131546821256478e-04
GC_11_137 b_11 NI_11 NS_137 0 1.5094322324426538e-05
GC_11_138 b_11 NI_11 NS_138 0 -5.7767603422069247e-05
GC_11_139 b_11 NI_11 NS_139 0 -4.6444429310431241e-06
GC_11_140 b_11 NI_11 NS_140 0 1.3827759013040212e-05
GC_11_141 b_11 NI_11 NS_141 0 3.0653425718591586e-04
GC_11_142 b_11 NI_11 NS_142 0 -2.6884033384372134e-04
GC_11_143 b_11 NI_11 NS_143 0 4.3094718895175103e-05
GC_11_144 b_11 NI_11 NS_144 0 1.3367637485164449e-08
GC_11_145 b_11 NI_11 NS_145 0 -1.4591757609981580e-10
GC_11_146 b_11 NI_11 NS_146 0 1.4531717962074378e-11
GC_11_147 b_11 NI_11 NS_147 0 1.8114016000134280e-06
GC_11_148 b_11 NI_11 NS_148 0 7.0832232769391397e-06
GC_11_149 b_11 NI_11 NS_149 0 3.2827978653147476e-05
GC_11_150 b_11 NI_11 NS_150 0 2.1661354790301326e-05
GC_11_151 b_11 NI_11 NS_151 0 4.5946586622722143e-05
GC_11_152 b_11 NI_11 NS_152 0 -5.6356955123331968e-05
GC_11_153 b_11 NI_11 NS_153 0 7.3626812430193029e-05
GC_11_154 b_11 NI_11 NS_154 0 -1.2529400494813646e-04
GC_11_155 b_11 NI_11 NS_155 0 -1.8750647652978004e-04
GC_11_156 b_11 NI_11 NS_156 0 -7.4918083828874306e-05
GC_11_157 b_11 NI_11 NS_157 0 8.1189036546717761e-06
GC_11_158 b_11 NI_11 NS_158 0 3.6709421050132709e-06
GC_11_159 b_11 NI_11 NS_159 0 -5.4185551379471422e-05
GC_11_160 b_11 NI_11 NS_160 0 -3.1100960656261208e-05
GC_11_161 b_11 NI_11 NS_161 0 2.2274168818736589e-02
GC_11_162 b_11 NI_11 NS_162 0 8.9558653696552703e-03
GC_11_163 b_11 NI_11 NS_163 0 -1.1409760318263785e-02
GC_11_164 b_11 NI_11 NS_164 0 -5.3360829798495891e-06
GC_11_165 b_11 NI_11 NS_165 0 -9.5822584229266206e-08
GC_11_166 b_11 NI_11 NS_166 0 -1.2412247368604066e-09
GC_11_167 b_11 NI_11 NS_167 0 -3.3143876880205891e-03
GC_11_168 b_11 NI_11 NS_168 0 -2.3911424295166052e-03
GC_11_169 b_11 NI_11 NS_169 0 2.7261772326534119e-03
GC_11_170 b_11 NI_11 NS_170 0 1.1171778349198237e-02
GC_11_171 b_11 NI_11 NS_171 0 -3.5307692784337631e-04
GC_11_172 b_11 NI_11 NS_172 0 -1.7759589703801117e-02
GC_11_173 b_11 NI_11 NS_173 0 -2.2020926253592869e-02
GC_11_174 b_11 NI_11 NS_174 0 2.1326548385709757e-02
GC_11_175 b_11 NI_11 NS_175 0 2.8908354578924170e-02
GC_11_176 b_11 NI_11 NS_176 0 -1.8397055755763517e-02
GC_11_177 b_11 NI_11 NS_177 0 -2.4507582349978271e-03
GC_11_178 b_11 NI_11 NS_178 0 1.4218496269307417e-03
GC_11_179 b_11 NI_11 NS_179 0 -1.7818879423500012e-02
GC_11_180 b_11 NI_11 NS_180 0 -7.1265651977145674e-03
GC_11_181 b_11 NI_11 NS_181 0 -8.2288462498620471e-02
GC_11_182 b_11 NI_11 NS_182 0 6.5322022214093556e-02
GC_11_183 b_11 NI_11 NS_183 0 -1.0307114068140173e-02
GC_11_184 b_11 NI_11 NS_184 0 -2.3858537918053743e-06
GC_11_185 b_11 NI_11 NS_185 0 1.6335227246656692e-08
GC_11_186 b_11 NI_11 NS_186 0 1.6410075230771303e-09
GC_11_187 b_11 NI_11 NS_187 0 -3.9597027678169174e-04
GC_11_188 b_11 NI_11 NS_188 0 -1.4000566626429841e-03
GC_11_189 b_11 NI_11 NS_189 0 -6.9917489106644179e-03
GC_11_190 b_11 NI_11 NS_190 0 -3.7822426745787200e-03
GC_11_191 b_11 NI_11 NS_191 0 -9.0594500213065660e-03
GC_11_192 b_11 NI_11 NS_192 0 1.3121191967648098e-02
GC_11_193 b_11 NI_11 NS_193 0 -1.5240953623785794e-02
GC_11_194 b_11 NI_11 NS_194 0 2.8718755468089892e-02
GC_11_195 b_11 NI_11 NS_195 0 4.5110989419775836e-02
GC_11_196 b_11 NI_11 NS_196 0 1.6488628398225652e-02
GC_11_197 b_11 NI_11 NS_197 0 -2.2090750107975564e-03
GC_11_198 b_11 NI_11 NS_198 0 -1.3391802445669554e-03
GC_11_199 b_11 NI_11 NS_199 0 1.2863710736047005e-02
GC_11_200 b_11 NI_11 NS_200 0 6.9572427905245397e-03
GC_11_201 b_11 NI_11 NS_201 0 -1.0222218199022234e-03
GC_11_202 b_11 NI_11 NS_202 0 -1.7322667337562117e-02
GC_11_203 b_11 NI_11 NS_203 0 1.1757822321038440e-02
GC_11_204 b_11 NI_11 NS_204 0 2.8947521987479011e-06
GC_11_205 b_11 NI_11 NS_205 0 -5.0926480200552165e-07
GC_11_206 b_11 NI_11 NS_206 0 -2.9660693206967109e-08
GC_11_207 b_11 NI_11 NS_207 0 3.0704129206818977e-03
GC_11_208 b_11 NI_11 NS_208 0 1.2919122677458163e-03
GC_11_209 b_11 NI_11 NS_209 0 -2.9518617912495998e-03
GC_11_210 b_11 NI_11 NS_210 0 -9.9170147504578608e-03
GC_11_211 b_11 NI_11 NS_211 0 5.8893990155318553e-04
GC_11_212 b_11 NI_11 NS_212 0 1.3640194085604559e-02
GC_11_213 b_11 NI_11 NS_213 0 1.7423650847933028e-02
GC_11_214 b_11 NI_11 NS_214 0 -2.3868295329448192e-02
GC_11_215 b_11 NI_11 NS_215 0 -3.3167483068215389e-02
GC_11_216 b_11 NI_11 NS_216 0 2.1401806846109192e-02
GC_11_217 b_11 NI_11 NS_217 0 4.0587920128512681e-03
GC_11_218 b_11 NI_11 NS_218 0 -2.2320125572230726e-03
GC_11_219 b_11 NI_11 NS_219 0 1.5116274676881826e-02
GC_11_220 b_11 NI_11 NS_220 0 5.6072379775210174e-03
GC_11_221 b_11 NI_11 NS_221 0 -2.8699861301888163e-01
GC_11_222 b_11 NI_11 NS_222 0 1.2135733566209578e-01
GC_11_223 b_11 NI_11 NS_223 0 7.0298547325991752e-03
GC_11_224 b_11 NI_11 NS_224 0 5.7777308691342764e-05
GC_11_225 b_11 NI_11 NS_225 0 1.2954678207255965e-06
GC_11_226 b_11 NI_11 NS_226 0 1.4196126366674965e-08
GC_11_227 b_11 NI_11 NS_227 0 3.0514922368646502e-02
GC_11_228 b_11 NI_11 NS_228 0 4.1652927566380813e-03
GC_11_229 b_11 NI_11 NS_229 0 -7.3042423185197816e-03
GC_11_230 b_11 NI_11 NS_230 0 2.2210833277304599e-02
GC_11_231 b_11 NI_11 NS_231 0 -1.6943498694100917e-02
GC_11_232 b_11 NI_11 NS_232 0 -1.8718581784369616e-02
GC_11_233 b_11 NI_11 NS_233 0 4.4820937500064592e-02
GC_11_234 b_11 NI_11 NS_234 0 1.4501639766489303e-02
GC_11_235 b_11 NI_11 NS_235 0 8.2245805673077890e-02
GC_11_236 b_11 NI_11 NS_236 0 3.0932530814678252e-02
GC_11_237 b_11 NI_11 NS_237 0 -1.0134599971683741e-02
GC_11_238 b_11 NI_11 NS_238 0 -4.8138188428595227e-03
GC_11_239 b_11 NI_11 NS_239 0 -2.1451566498955427e-02
GC_11_240 b_11 NI_11 NS_240 0 -4.8857370374835538e-03
GD_11_1 b_11 NI_11 NA_1 0 -2.3872961867743070e-06
GD_11_2 b_11 NI_11 NA_2 0 6.5403357254194124e-06
GD_11_3 b_11 NI_11 NA_3 0 -2.2751425886264647e-06
GD_11_4 b_11 NI_11 NA_4 0 -1.0327428482952664e-05
GD_11_5 b_11 NI_11 NA_5 0 1.5822121425586232e-05
GD_11_6 b_11 NI_11 NA_6 0 -8.9720788191917314e-06
GD_11_7 b_11 NI_11 NA_7 0 -6.8612069661387471e-05
GD_11_8 b_11 NI_11 NA_8 0 4.7002133049589670e-06
GD_11_9 b_11 NI_11 NA_9 0 6.2239325459216514e-03
GD_11_10 b_11 NI_11 NA_10 0 2.3474521334049723e-03
GD_11_11 b_11 NI_11 NA_11 0 -6.6119414765316411e-03
GD_11_12 b_11 NI_11 NA_12 0 5.7256229496306169e-02
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -6.3290788378927718e-07
GC_12_2 b_12 NI_12 NS_2 0 -6.2866891910464745e-07
GC_12_3 b_12 NI_12 NS_3 0 -7.3718796085161488e-08
GC_12_4 b_12 NI_12 NS_4 0 4.6597127153938720e-09
GC_12_5 b_12 NI_12 NS_5 0 -1.7622882231889620e-10
GC_12_6 b_12 NI_12 NS_6 0 1.2485707011843411e-11
GC_12_7 b_12 NI_12 NS_7 0 9.0995538869945570e-07
GC_12_8 b_12 NI_12 NS_8 0 -8.4388375385126877e-07
GC_12_9 b_12 NI_12 NS_9 0 1.2594059199062994e-06
GC_12_10 b_12 NI_12 NS_10 0 -1.6700306022056056e-07
GC_12_11 b_12 NI_12 NS_11 0 -1.8724480129604691e-07
GC_12_12 b_12 NI_12 NS_12 0 -1.1999801867934967e-06
GC_12_13 b_12 NI_12 NS_13 0 2.8912206562769268e-06
GC_12_14 b_12 NI_12 NS_14 0 -4.1236267279435793e-06
GC_12_15 b_12 NI_12 NS_15 0 -8.7556921213651860e-06
GC_12_16 b_12 NI_12 NS_16 0 4.7054928053421935e-08
GC_12_17 b_12 NI_12 NS_17 0 2.1502533321987839e-06
GC_12_18 b_12 NI_12 NS_18 0 -3.9617857077803051e-07
GC_12_19 b_12 NI_12 NS_19 0 -8.8887426448317629e-07
GC_12_20 b_12 NI_12 NS_20 0 8.3645540967613525e-07
GC_12_21 b_12 NI_12 NS_21 0 7.3331183615713705e-06
GC_12_22 b_12 NI_12 NS_22 0 -2.5197815900965689e-06
GC_12_23 b_12 NI_12 NS_23 0 1.5310196321700546e-07
GC_12_24 b_12 NI_12 NS_24 0 -4.0111450393841471e-09
GC_12_25 b_12 NI_12 NS_25 0 1.6388492151532103e-10
GC_12_26 b_12 NI_12 NS_26 0 -1.2217805484311787e-11
GC_12_27 b_12 NI_12 NS_27 0 -3.1670347500463701e-07
GC_12_28 b_12 NI_12 NS_28 0 -2.3700965194203781e-07
GC_12_29 b_12 NI_12 NS_29 0 -7.6440590468033916e-08
GC_12_30 b_12 NI_12 NS_30 0 9.2571194281736848e-08
GC_12_31 b_12 NI_12 NS_31 0 -7.8260992580901296e-07
GC_12_32 b_12 NI_12 NS_32 0 -4.1598996545766936e-07
GC_12_33 b_12 NI_12 NS_33 0 -9.7698206334045851e-07
GC_12_34 b_12 NI_12 NS_34 0 4.5608518979317941e-07
GC_12_35 b_12 NI_12 NS_35 0 2.6664038813029764e-07
GC_12_36 b_12 NI_12 NS_36 0 3.1017418859141776e-07
GC_12_37 b_12 NI_12 NS_37 0 -1.5147396979805437e-07
GC_12_38 b_12 NI_12 NS_38 0 -3.1214805334718237e-07
GC_12_39 b_12 NI_12 NS_39 0 -8.8434226257387979e-07
GC_12_40 b_12 NI_12 NS_40 0 -4.0322299825756732e-07
GC_12_41 b_12 NI_12 NS_41 0 2.0605007071921828e-05
GC_12_42 b_12 NI_12 NS_42 0 -4.9936211052643231e-06
GC_12_43 b_12 NI_12 NS_43 0 9.9303793371084712e-07
GC_12_44 b_12 NI_12 NS_44 0 -5.4984967371157845e-09
GC_12_45 b_12 NI_12 NS_45 0 -2.5967407490769176e-11
GC_12_46 b_12 NI_12 NS_46 0 -1.2308300765102890e-12
GC_12_47 b_12 NI_12 NS_47 0 -1.3115724464306875e-06
GC_12_48 b_12 NI_12 NS_48 0 -1.6746979778810741e-06
GC_12_49 b_12 NI_12 NS_49 0 -1.7990700462192592e-06
GC_12_50 b_12 NI_12 NS_50 0 1.3846231364449422e-07
GC_12_51 b_12 NI_12 NS_51 0 -2.4070677722172857e-06
GC_12_52 b_12 NI_12 NS_52 0 2.2075384305251468e-06
GC_12_53 b_12 NI_12 NS_53 0 -3.9349091554389338e-06
GC_12_54 b_12 NI_12 NS_54 0 -2.1437294138403094e-06
GC_12_55 b_12 NI_12 NS_55 0 1.2290495648341703e-06
GC_12_56 b_12 NI_12 NS_56 0 8.2806510396724393e-06
GC_12_57 b_12 NI_12 NS_57 0 -3.9212471267388198e-07
GC_12_58 b_12 NI_12 NS_58 0 -1.7846417379064647e-06
GC_12_59 b_12 NI_12 NS_59 0 -3.6944482058148867e-07
GC_12_60 b_12 NI_12 NS_60 0 1.7727239498238500e-07
GC_12_61 b_12 NI_12 NS_61 0 5.6987573281481272e-06
GC_12_62 b_12 NI_12 NS_62 0 1.3907357992375358e-06
GC_12_63 b_12 NI_12 NS_63 0 -8.6920422367024303e-07
GC_12_64 b_12 NI_12 NS_64 0 3.5211619168848996e-09
GC_12_65 b_12 NI_12 NS_65 0 5.0063240303496537e-11
GC_12_66 b_12 NI_12 NS_66 0 -5.2297008142905652e-13
GC_12_67 b_12 NI_12 NS_67 0 -4.1974768109372614e-07
GC_12_68 b_12 NI_12 NS_68 0 -3.4327712256816691e-07
GC_12_69 b_12 NI_12 NS_69 0 -2.5399991669621554e-07
GC_12_70 b_12 NI_12 NS_70 0 2.2159700577989292e-07
GC_12_71 b_12 NI_12 NS_71 0 -7.9481937783193012e-07
GC_12_72 b_12 NI_12 NS_72 0 -6.7506845945513520e-07
GC_12_73 b_12 NI_12 NS_73 0 -2.5308339071263310e-06
GC_12_74 b_12 NI_12 NS_74 0 -3.7212592864869052e-08
GC_12_75 b_12 NI_12 NS_75 0 4.0514417156895624e-07
GC_12_76 b_12 NI_12 NS_76 0 3.4974523619603794e-06
GC_12_77 b_12 NI_12 NS_77 0 1.6145098651332762e-07
GC_12_78 b_12 NI_12 NS_78 0 -8.5014424438125345e-07
GC_12_79 b_12 NI_12 NS_79 0 -5.6427564799638657e-07
GC_12_80 b_12 NI_12 NS_80 0 2.6709321780139297e-07
GC_12_81 b_12 NI_12 NS_81 0 6.1561232496312854e-05
GC_12_82 b_12 NI_12 NS_82 0 -4.0958851303335263e-05
GC_12_83 b_12 NI_12 NS_83 0 7.0396238441792517e-06
GC_12_84 b_12 NI_12 NS_84 0 -1.5378936562559431e-08
GC_12_85 b_12 NI_12 NS_85 0 -2.8245671117932566e-11
GC_12_86 b_12 NI_12 NS_86 0 2.8279339416938707e-13
GC_12_87 b_12 NI_12 NS_87 0 -9.2347580134835979e-07
GC_12_88 b_12 NI_12 NS_88 0 -1.4177401810871660e-06
GC_12_89 b_12 NI_12 NS_89 0 1.3243137268732516e-06
GC_12_90 b_12 NI_12 NS_90 0 2.2639608902106843e-06
GC_12_91 b_12 NI_12 NS_91 0 2.9219975148668169e-06
GC_12_92 b_12 NI_12 NS_92 0 -3.4302899477628638e-06
GC_12_93 b_12 NI_12 NS_93 0 7.8764338850907101e-06
GC_12_94 b_12 NI_12 NS_94 0 -1.6473451780454270e-05
GC_12_95 b_12 NI_12 NS_95 0 -2.6664824402225746e-05
GC_12_96 b_12 NI_12 NS_96 0 -4.5354760750879556e-06
GC_12_97 b_12 NI_12 NS_97 0 2.5875753580031855e-06
GC_12_98 b_12 NI_12 NS_98 0 -5.4559824270517768e-07
GC_12_99 b_12 NI_12 NS_99 0 -7.0823181464555601e-06
GC_12_100 b_12 NI_12 NS_100 0 -3.6861006134273905e-06
GC_12_101 b_12 NI_12 NS_101 0 -7.8386261946403104e-05
GC_12_102 b_12 NI_12 NS_102 0 1.3378293153951663e-05
GC_12_103 b_12 NI_12 NS_103 0 -1.3935999271144057e-06
GC_12_104 b_12 NI_12 NS_104 0 -1.3100501299890116e-08
GC_12_105 b_12 NI_12 NS_105 0 2.6340784642751825e-10
GC_12_106 b_12 NI_12 NS_106 0 -1.7096271668709784e-11
GC_12_107 b_12 NI_12 NS_107 0 -1.5341826932945149e-06
GC_12_108 b_12 NI_12 NS_108 0 3.6435271177757809e-06
GC_12_109 b_12 NI_12 NS_109 0 1.6179622827286709e-06
GC_12_110 b_12 NI_12 NS_110 0 8.9335049960634538e-06
GC_12_111 b_12 NI_12 NS_111 0 1.0126601551899545e-05
GC_12_112 b_12 NI_12 NS_112 0 3.9283519349966383e-06
GC_12_113 b_12 NI_12 NS_113 0 1.3024106513905121e-05
GC_12_114 b_12 NI_12 NS_114 0 2.9985525527688097e-05
GC_12_115 b_12 NI_12 NS_115 0 3.6902719690009282e-05
GC_12_116 b_12 NI_12 NS_116 0 -6.0917486694685638e-05
GC_12_117 b_12 NI_12 NS_117 0 -6.8806255353126371e-06
GC_12_118 b_12 NI_12 NS_118 0 1.5060253555681945e-05
GC_12_119 b_12 NI_12 NS_119 0 -1.5080847490537638e-06
GC_12_120 b_12 NI_12 NS_120 0 -4.9189622965908964e-06
GC_12_121 b_12 NI_12 NS_121 0 3.0653417772478581e-04
GC_12_122 b_12 NI_12 NS_122 0 -2.6883990884266583e-04
GC_12_123 b_12 NI_12 NS_123 0 4.3094615836436782e-05
GC_12_124 b_12 NI_12 NS_124 0 1.3368228133868908e-08
GC_12_125 b_12 NI_12 NS_125 0 -1.4592405000296231e-10
GC_12_126 b_12 NI_12 NS_126 0 1.4532025229942466e-11
GC_12_127 b_12 NI_12 NS_127 0 1.8116506984137731e-06
GC_12_128 b_12 NI_12 NS_128 0 7.0833104131587975e-06
GC_12_129 b_12 NI_12 NS_129 0 3.2828260258652016e-05
GC_12_130 b_12 NI_12 NS_130 0 2.1661244590451996e-05
GC_12_131 b_12 NI_12 NS_131 0 4.5946354336465846e-05
GC_12_132 b_12 NI_12 NS_132 0 -5.6357656424812553e-05
GC_12_133 b_12 NI_12 NS_133 0 7.3626026507834545e-05
GC_12_134 b_12 NI_12 NS_134 0 -1.2529469236688772e-04
GC_12_135 b_12 NI_12 NS_135 0 -1.8750627923827927e-04
GC_12_136 b_12 NI_12 NS_136 0 -7.4916455071153611e-05
GC_12_137 b_12 NI_12 NS_137 0 8.1186763845942645e-06
GC_12_138 b_12 NI_12 NS_138 0 3.6705876998540959e-06
GC_12_139 b_12 NI_12 NS_139 0 -5.4185473401858401e-05
GC_12_140 b_12 NI_12 NS_140 0 -3.1100851790826563e-05
GC_12_141 b_12 NI_12 NS_141 0 2.7780708453021950e-04
GC_12_142 b_12 NI_12 NS_142 0 -1.2250103492826311e-05
GC_12_143 b_12 NI_12 NS_143 0 -9.4861498852765996e-06
GC_12_144 b_12 NI_12 NS_144 0 6.0731552473283756e-08
GC_12_145 b_12 NI_12 NS_145 0 -3.1317772365108767e-10
GC_12_146 b_12 NI_12 NS_146 0 8.9456590040487021e-12
GC_12_147 b_12 NI_12 NS_147 0 -7.0467245058718877e-07
GC_12_148 b_12 NI_12 NS_148 0 -1.5599737159566571e-05
GC_12_149 b_12 NI_12 NS_149 0 -9.9256356293910208e-06
GC_12_150 b_12 NI_12 NS_150 0 -2.0930532602158992e-05
GC_12_151 b_12 NI_12 NS_151 0 -3.7989342621725308e-05
GC_12_152 b_12 NI_12 NS_152 0 -1.9683745978959795e-05
GC_12_153 b_12 NI_12 NS_153 0 -7.5824501894951446e-05
GC_12_154 b_12 NI_12 NS_154 0 -7.9099396229594907e-05
GC_12_155 b_12 NI_12 NS_155 0 -7.4562449507106093e-05
GC_12_156 b_12 NI_12 NS_156 0 2.2166872013975204e-04
GC_12_157 b_12 NI_12 NS_157 0 1.5124435086401826e-05
GC_12_158 b_12 NI_12 NS_158 0 -5.7842961336570353e-05
GC_12_159 b_12 NI_12 NS_159 0 -4.6595010747284122e-06
GC_12_160 b_12 NI_12 NS_160 0 1.3855697769030026e-05
GC_12_161 b_12 NI_12 NS_161 0 -8.2288464694788621e-02
GC_12_162 b_12 NI_12 NS_162 0 6.5322022997245599e-02
GC_12_163 b_12 NI_12 NS_163 0 -1.0307114159569586e-02
GC_12_164 b_12 NI_12 NS_164 0 -2.3858535076404995e-06
GC_12_165 b_12 NI_12 NS_165 0 1.6335225056678213e-08
GC_12_166 b_12 NI_12 NS_166 0 1.6410076036530494e-09
GC_12_167 b_12 NI_12 NS_167 0 -3.9597042998080106e-04
GC_12_168 b_12 NI_12 NS_168 0 -1.4000566242028801e-03
GC_12_169 b_12 NI_12 NS_169 0 -6.9917490294911103e-03
GC_12_170 b_12 NI_12 NS_170 0 -3.7822424126441562e-03
GC_12_171 b_12 NI_12 NS_171 0 -9.0594497462318513e-03
GC_12_172 b_12 NI_12 NS_172 0 1.3121192334235773e-02
GC_12_173 b_12 NI_12 NS_173 0 -1.5240953398823445e-02
GC_12_174 b_12 NI_12 NS_174 0 2.8718756215261588e-02
GC_12_175 b_12 NI_12 NS_175 0 4.5110990633982911e-02
GC_12_176 b_12 NI_12 NS_176 0 1.6488627481823045e-02
GC_12_177 b_12 NI_12 NS_177 0 -2.2090752244941026e-03
GC_12_178 b_12 NI_12 NS_178 0 -1.3391800354162627e-03
GC_12_179 b_12 NI_12 NS_179 0 1.2863710852294810e-02
GC_12_180 b_12 NI_12 NS_180 0 6.9572427257932820e-03
GC_12_181 b_12 NI_12 NS_181 0 2.2267872707234619e-02
GC_12_182 b_12 NI_12 NS_182 0 8.9573222676478607e-03
GC_12_183 b_12 NI_12 NS_183 0 -1.1409899591953643e-02
GC_12_184 b_12 NI_12 NS_184 0 -5.3357066209233111e-06
GC_12_185 b_12 NI_12 NS_185 0 -9.5823209710086011e-08
GC_12_186 b_12 NI_12 NS_186 0 -1.2410084341522251e-09
GC_12_187 b_12 NI_12 NS_187 0 -3.3142115015536481e-03
GC_12_188 b_12 NI_12 NS_188 0 -2.3908938231856510e-03
GC_12_189 b_12 NI_12 NS_189 0 2.7265908031993036e-03
GC_12_190 b_12 NI_12 NS_190 0 1.1171998927836281e-02
GC_12_191 b_12 NI_12 NS_191 0 -3.5268546161212530e-04
GC_12_192 b_12 NI_12 NS_192 0 -1.7759690683797062e-02
GC_12_193 b_12 NI_12 NS_193 0 -2.2020323746107347e-02
GC_12_194 b_12 NI_12 NS_194 0 2.1327619534719986e-02
GC_12_195 b_12 NI_12 NS_195 0 2.8910205978017023e-02
GC_12_196 b_12 NI_12 NS_196 0 -1.8399093090247776e-02
GC_12_197 b_12 NI_12 NS_197 0 -2.4511212692121301e-03
GC_12_198 b_12 NI_12 NS_198 0 1.4222330861585661e-03
GC_12_199 b_12 NI_12 NS_199 0 -1.7818694330355617e-02
GC_12_200 b_12 NI_12 NS_200 0 -7.1267653599122668e-03
GC_12_201 b_12 NI_12 NS_201 0 -2.8699895172713702e-01
GC_12_202 b_12 NI_12 NS_202 0 1.2135745495950856e-01
GC_12_203 b_12 NI_12 NS_203 0 7.0298413472848547e-03
GC_12_204 b_12 NI_12 NS_204 0 5.7777328467957321e-05
GC_12_205 b_12 NI_12 NS_205 0 1.2954678402692023e-06
GC_12_206 b_12 NI_12 NS_206 0 1.4196095832331219e-08
GC_12_207 b_12 NI_12 NS_207 0 3.0514954728750588e-02
GC_12_208 b_12 NI_12 NS_208 0 4.1653131818644796e-03
GC_12_209 b_12 NI_12 NS_209 0 -7.3041991343619885e-03
GC_12_210 b_12 NI_12 NS_210 0 2.2210832243773123e-02
GC_12_211 b_12 NI_12 NS_211 0 -1.6943518811170524e-02
GC_12_212 b_12 NI_12 NS_212 0 -1.8718655752257899e-02
GC_12_213 b_12 NI_12 NS_213 0 4.4820829918844222e-02
GC_12_214 b_12 NI_12 NS_214 0 1.4501654652951437e-02
GC_12_215 b_12 NI_12 NS_215 0 8.2246059760329865e-02
GC_12_216 b_12 NI_12 NS_216 0 3.0932601360990644e-02
GC_12_217 b_12 NI_12 NS_217 0 -1.0134686762140580e-02
GC_12_218 b_12 NI_12 NS_218 0 -4.8138229160149884e-03
GC_12_219 b_12 NI_12 NS_219 0 -2.1451541440712946e-02
GC_12_220 b_12 NI_12 NS_220 0 -4.8857427933137578e-03
GC_12_221 b_12 NI_12 NS_221 0 -1.0222218199021406e-03
GC_12_222 b_12 NI_12 NS_222 0 -1.7322667337562141e-02
GC_12_223 b_12 NI_12 NS_223 0 1.1757822321038442e-02
GC_12_224 b_12 NI_12 NS_224 0 2.8947521987479596e-06
GC_12_225 b_12 NI_12 NS_225 0 -5.0926480200552260e-07
GC_12_226 b_12 NI_12 NS_226 0 -2.9660693206967926e-08
GC_12_227 b_12 NI_12 NS_227 0 3.0704129206818934e-03
GC_12_228 b_12 NI_12 NS_228 0 1.2919122677458135e-03
GC_12_229 b_12 NI_12 NS_229 0 -2.9518617912496089e-03
GC_12_230 b_12 NI_12 NS_230 0 -9.9170147504578556e-03
GC_12_231 b_12 NI_12 NS_231 0 5.8893990155318553e-04
GC_12_232 b_12 NI_12 NS_232 0 1.3640194085604570e-02
GC_12_233 b_12 NI_12 NS_233 0 1.7423650847933028e-02
GC_12_234 b_12 NI_12 NS_234 0 -2.3868295329448192e-02
GC_12_235 b_12 NI_12 NS_235 0 -3.3167483068215389e-02
GC_12_236 b_12 NI_12 NS_236 0 2.1401806846109192e-02
GC_12_237 b_12 NI_12 NS_237 0 4.0587920128512646e-03
GC_12_238 b_12 NI_12 NS_238 0 -2.2320125572230726e-03
GC_12_239 b_12 NI_12 NS_239 0 1.5116274676881819e-02
GC_12_240 b_12 NI_12 NS_240 0 5.6072379775210165e-03
GD_12_1 b_12 NI_12 NA_1 0 6.5411157714154100e-06
GD_12_2 b_12 NI_12 NA_2 0 -2.3878576207842484e-06
GD_12_3 b_12 NI_12 NA_3 0 -1.0327450587005908e-05
GD_12_4 b_12 NI_12 NA_4 0 -2.2999151906737156e-06
GD_12_5 b_12 NI_12 NA_5 0 -9.0215010429437939e-06
GD_12_6 b_12 NI_12 NA_6 0 1.5819161125309400e-05
GD_12_7 b_12 NI_12 NA_7 0 4.7004550697881715e-06
GD_12_8 b_12 NI_12 NA_8 0 -6.9107945848929060e-05
GD_12_9 b_12 NI_12 NA_9 0 2.3474522237801219e-03
GD_12_10 b_12 NI_12 NA_10 0 6.2259707324475279e-03
GD_12_11 b_12 NI_12 NA_11 0 5.7256341619874099e-02
GD_12_12 b_12 NI_12 NA_12 0 -6.6119414765317104e-03
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 4.5298699859481095e+00
GS_1_1 0 NS_1 NA_1 0 1.3906701219673681e+00
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 1.1221187714172293e+01
GS_2_1 0 NS_2 NA_1 0 1.3906701219673681e+00
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 1.8217191146854518e+01
GS_3_1 0 NS_3 NA_1 0 1.3906701219673681e+00
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 6.6287934454477863e+01
GS_4_1 0 NS_4 NA_1 0 1.3906701219673681e+00
*
* Real pole n. 5
CS_5 NS_5 0 9.9999999999999998e-13
RS_5 NS_5 0 5.4647183375290433e+02
GS_5_1 0 NS_5 NA_1 0 1.3906701219673681e+00
*
* Real pole n. 6
CS_6 NS_6 0 9.9999999999999998e-13
RS_6 NS_6 0 3.8169396682972065e+03
GS_6_1 0 NS_6 NA_1 0 1.3906701219673681e+00
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 2.1530817355819540e+01
RS_8 NS_8 0 2.1530817355819540e+01
GL_7 0 NS_7 NS_8 0 2.8893552838207953e-01
GL_8 0 NS_8 NS_7 0 -2.8893552838207953e-01
GS_7_1 0 NS_7 NA_1 0 1.3906701219673681e+00
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 1.7704391175337044e+01
RS_10 NS_10 0 1.7704391175337044e+01
GL_9 0 NS_9 NS_10 0 2.4113766587096394e-01
GL_10 0 NS_10 NS_9 0 -2.4113766587096394e-01
GS_9_1 0 NS_9 NA_1 0 1.3906701219673681e+00
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 1.5980319858751495e+01
RS_12 NS_12 0 1.5980319858751495e+01
GL_11 0 NS_11 NS_12 0 2.0836264676973826e-01
GL_12 0 NS_12 NS_11 0 -2.0836264676973826e-01
GS_11_1 0 NS_11 NA_1 0 1.3906701219673681e+00
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 1.5652313341768849e+01
RS_14 NS_14 0 1.5652313341768847e+01
GL_13 0 NS_13 NS_14 0 1.5274998946760082e-01
GL_14 0 NS_14 NS_13 0 -1.5274998946760082e-01
GS_13_1 0 NS_13 NA_1 0 1.3906701219673681e+00
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 1.5016887791939077e+01
RS_16 NS_16 0 1.5016887791939077e+01
GL_15 0 NS_15 NS_16 0 1.2573527610391108e-01
GL_16 0 NS_16 NS_15 0 -1.2573527610391108e-01
GS_15_1 0 NS_15 NA_1 0 1.3906701219673681e+00
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 1.9705893378385916e+01
RS_18 NS_18 0 1.9705893378385916e+01
GL_17 0 NS_17 NS_18 0 1.2264058452613225e-01
GL_18 0 NS_18 NS_17 0 -1.2264058452613225e-01
GS_17_1 0 NS_17 NA_1 0 1.3906701219673681e+00
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 1.7719166159098595e+01
RS_20 NS_20 0 1.7719166159098595e+01
GL_19 0 NS_19 NS_20 0 7.0127888352005202e-02
GL_20 0 NS_20 NS_19 0 -7.0127888352005202e-02
GS_19_1 0 NS_19 NA_1 0 1.3906701219673681e+00
*
* Real pole n. 21
CS_21 NS_21 0 9.9999999999999998e-13
RS_21 NS_21 0 4.5298699859481095e+00
GS_21_2 0 NS_21 NA_2 0 1.3906701219673681e+00
*
* Real pole n. 22
CS_22 NS_22 0 9.9999999999999998e-13
RS_22 NS_22 0 1.1221187714172293e+01
GS_22_2 0 NS_22 NA_2 0 1.3906701219673681e+00
*
* Real pole n. 23
CS_23 NS_23 0 9.9999999999999998e-13
RS_23 NS_23 0 1.8217191146854518e+01
GS_23_2 0 NS_23 NA_2 0 1.3906701219673681e+00
*
* Real pole n. 24
CS_24 NS_24 0 9.9999999999999998e-13
RS_24 NS_24 0 6.6287934454477863e+01
GS_24_2 0 NS_24 NA_2 0 1.3906701219673681e+00
*
* Real pole n. 25
CS_25 NS_25 0 9.9999999999999998e-13
RS_25 NS_25 0 5.4647183375290433e+02
GS_25_2 0 NS_25 NA_2 0 1.3906701219673681e+00
*
* Real pole n. 26
CS_26 NS_26 0 9.9999999999999998e-13
RS_26 NS_26 0 3.8169396682972065e+03
GS_26_2 0 NS_26 NA_2 0 1.3906701219673681e+00
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 2.1530817355819540e+01
RS_28 NS_28 0 2.1530817355819540e+01
GL_27 0 NS_27 NS_28 0 2.8893552838207953e-01
GL_28 0 NS_28 NS_27 0 -2.8893552838207953e-01
GS_27_2 0 NS_27 NA_2 0 1.3906701219673681e+00
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 1.7704391175337044e+01
RS_30 NS_30 0 1.7704391175337044e+01
GL_29 0 NS_29 NS_30 0 2.4113766587096394e-01
GL_30 0 NS_30 NS_29 0 -2.4113766587096394e-01
GS_29_2 0 NS_29 NA_2 0 1.3906701219673681e+00
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 1.5980319858751495e+01
RS_32 NS_32 0 1.5980319858751495e+01
GL_31 0 NS_31 NS_32 0 2.0836264676973826e-01
GL_32 0 NS_32 NS_31 0 -2.0836264676973826e-01
GS_31_2 0 NS_31 NA_2 0 1.3906701219673681e+00
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 1.5652313341768849e+01
RS_34 NS_34 0 1.5652313341768847e+01
GL_33 0 NS_33 NS_34 0 1.5274998946760082e-01
GL_34 0 NS_34 NS_33 0 -1.5274998946760082e-01
GS_33_2 0 NS_33 NA_2 0 1.3906701219673681e+00
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 1.5016887791939077e+01
RS_36 NS_36 0 1.5016887791939077e+01
GL_35 0 NS_35 NS_36 0 1.2573527610391108e-01
GL_36 0 NS_36 NS_35 0 -1.2573527610391108e-01
GS_35_2 0 NS_35 NA_2 0 1.3906701219673681e+00
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 1.9705893378385916e+01
RS_38 NS_38 0 1.9705893378385916e+01
GL_37 0 NS_37 NS_38 0 1.2264058452613225e-01
GL_38 0 NS_38 NS_37 0 -1.2264058452613225e-01
GS_37_2 0 NS_37 NA_2 0 1.3906701219673681e+00
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 1.7719166159098595e+01
RS_40 NS_40 0 1.7719166159098595e+01
GL_39 0 NS_39 NS_40 0 7.0127888352005202e-02
GL_40 0 NS_40 NS_39 0 -7.0127888352005202e-02
GS_39_2 0 NS_39 NA_2 0 1.3906701219673681e+00
*
* Real pole n. 41
CS_41 NS_41 0 9.9999999999999998e-13
RS_41 NS_41 0 4.5298699859481095e+00
GS_41_3 0 NS_41 NA_3 0 1.3906701219673681e+00
*
* Real pole n. 42
CS_42 NS_42 0 9.9999999999999998e-13
RS_42 NS_42 0 1.1221187714172293e+01
GS_42_3 0 NS_42 NA_3 0 1.3906701219673681e+00
*
* Real pole n. 43
CS_43 NS_43 0 9.9999999999999998e-13
RS_43 NS_43 0 1.8217191146854518e+01
GS_43_3 0 NS_43 NA_3 0 1.3906701219673681e+00
*
* Real pole n. 44
CS_44 NS_44 0 9.9999999999999998e-13
RS_44 NS_44 0 6.6287934454477863e+01
GS_44_3 0 NS_44 NA_3 0 1.3906701219673681e+00
*
* Real pole n. 45
CS_45 NS_45 0 9.9999999999999998e-13
RS_45 NS_45 0 5.4647183375290433e+02
GS_45_3 0 NS_45 NA_3 0 1.3906701219673681e+00
*
* Real pole n. 46
CS_46 NS_46 0 9.9999999999999998e-13
RS_46 NS_46 0 3.8169396682972065e+03
GS_46_3 0 NS_46 NA_3 0 1.3906701219673681e+00
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 2.1530817355819540e+01
RS_48 NS_48 0 2.1530817355819540e+01
GL_47 0 NS_47 NS_48 0 2.8893552838207953e-01
GL_48 0 NS_48 NS_47 0 -2.8893552838207953e-01
GS_47_3 0 NS_47 NA_3 0 1.3906701219673681e+00
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 1.7704391175337044e+01
RS_50 NS_50 0 1.7704391175337044e+01
GL_49 0 NS_49 NS_50 0 2.4113766587096394e-01
GL_50 0 NS_50 NS_49 0 -2.4113766587096394e-01
GS_49_3 0 NS_49 NA_3 0 1.3906701219673681e+00
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 1.5980319858751495e+01
RS_52 NS_52 0 1.5980319858751495e+01
GL_51 0 NS_51 NS_52 0 2.0836264676973826e-01
GL_52 0 NS_52 NS_51 0 -2.0836264676973826e-01
GS_51_3 0 NS_51 NA_3 0 1.3906701219673681e+00
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 1.5652313341768849e+01
RS_54 NS_54 0 1.5652313341768847e+01
GL_53 0 NS_53 NS_54 0 1.5274998946760082e-01
GL_54 0 NS_54 NS_53 0 -1.5274998946760082e-01
GS_53_3 0 NS_53 NA_3 0 1.3906701219673681e+00
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 1.5016887791939077e+01
RS_56 NS_56 0 1.5016887791939077e+01
GL_55 0 NS_55 NS_56 0 1.2573527610391108e-01
GL_56 0 NS_56 NS_55 0 -1.2573527610391108e-01
GS_55_3 0 NS_55 NA_3 0 1.3906701219673681e+00
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 1.9705893378385916e+01
RS_58 NS_58 0 1.9705893378385916e+01
GL_57 0 NS_57 NS_58 0 1.2264058452613225e-01
GL_58 0 NS_58 NS_57 0 -1.2264058452613225e-01
GS_57_3 0 NS_57 NA_3 0 1.3906701219673681e+00
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 1.7719166159098595e+01
RS_60 NS_60 0 1.7719166159098595e+01
GL_59 0 NS_59 NS_60 0 7.0127888352005202e-02
GL_60 0 NS_60 NS_59 0 -7.0127888352005202e-02
GS_59_3 0 NS_59 NA_3 0 1.3906701219673681e+00
*
* Real pole n. 61
CS_61 NS_61 0 9.9999999999999998e-13
RS_61 NS_61 0 4.5298699859481095e+00
GS_61_4 0 NS_61 NA_4 0 1.3906701219673681e+00
*
* Real pole n. 62
CS_62 NS_62 0 9.9999999999999998e-13
RS_62 NS_62 0 1.1221187714172293e+01
GS_62_4 0 NS_62 NA_4 0 1.3906701219673681e+00
*
* Real pole n. 63
CS_63 NS_63 0 9.9999999999999998e-13
RS_63 NS_63 0 1.8217191146854518e+01
GS_63_4 0 NS_63 NA_4 0 1.3906701219673681e+00
*
* Real pole n. 64
CS_64 NS_64 0 9.9999999999999998e-13
RS_64 NS_64 0 6.6287934454477863e+01
GS_64_4 0 NS_64 NA_4 0 1.3906701219673681e+00
*
* Real pole n. 65
CS_65 NS_65 0 9.9999999999999998e-13
RS_65 NS_65 0 5.4647183375290433e+02
GS_65_4 0 NS_65 NA_4 0 1.3906701219673681e+00
*
* Real pole n. 66
CS_66 NS_66 0 9.9999999999999998e-13
RS_66 NS_66 0 3.8169396682972065e+03
GS_66_4 0 NS_66 NA_4 0 1.3906701219673681e+00
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 2.1530817355819540e+01
RS_68 NS_68 0 2.1530817355819540e+01
GL_67 0 NS_67 NS_68 0 2.8893552838207953e-01
GL_68 0 NS_68 NS_67 0 -2.8893552838207953e-01
GS_67_4 0 NS_67 NA_4 0 1.3906701219673681e+00
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 1.7704391175337044e+01
RS_70 NS_70 0 1.7704391175337044e+01
GL_69 0 NS_69 NS_70 0 2.4113766587096394e-01
GL_70 0 NS_70 NS_69 0 -2.4113766587096394e-01
GS_69_4 0 NS_69 NA_4 0 1.3906701219673681e+00
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 1.5980319858751495e+01
RS_72 NS_72 0 1.5980319858751495e+01
GL_71 0 NS_71 NS_72 0 2.0836264676973826e-01
GL_72 0 NS_72 NS_71 0 -2.0836264676973826e-01
GS_71_4 0 NS_71 NA_4 0 1.3906701219673681e+00
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 1.5652313341768849e+01
RS_74 NS_74 0 1.5652313341768847e+01
GL_73 0 NS_73 NS_74 0 1.5274998946760082e-01
GL_74 0 NS_74 NS_73 0 -1.5274998946760082e-01
GS_73_4 0 NS_73 NA_4 0 1.3906701219673681e+00
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 1.5016887791939077e+01
RS_76 NS_76 0 1.5016887791939077e+01
GL_75 0 NS_75 NS_76 0 1.2573527610391108e-01
GL_76 0 NS_76 NS_75 0 -1.2573527610391108e-01
GS_75_4 0 NS_75 NA_4 0 1.3906701219673681e+00
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 1.9705893378385916e+01
RS_78 NS_78 0 1.9705893378385916e+01
GL_77 0 NS_77 NS_78 0 1.2264058452613225e-01
GL_78 0 NS_78 NS_77 0 -1.2264058452613225e-01
GS_77_4 0 NS_77 NA_4 0 1.3906701219673681e+00
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 1.7719166159098595e+01
RS_80 NS_80 0 1.7719166159098595e+01
GL_79 0 NS_79 NS_80 0 7.0127888352005202e-02
GL_80 0 NS_80 NS_79 0 -7.0127888352005202e-02
GS_79_4 0 NS_79 NA_4 0 1.3906701219673681e+00
*
* Real pole n. 81
CS_81 NS_81 0 9.9999999999999998e-13
RS_81 NS_81 0 4.5298699859481095e+00
GS_81_5 0 NS_81 NA_5 0 1.3906701219673681e+00
*
* Real pole n. 82
CS_82 NS_82 0 9.9999999999999998e-13
RS_82 NS_82 0 1.1221187714172293e+01
GS_82_5 0 NS_82 NA_5 0 1.3906701219673681e+00
*
* Real pole n. 83
CS_83 NS_83 0 9.9999999999999998e-13
RS_83 NS_83 0 1.8217191146854518e+01
GS_83_5 0 NS_83 NA_5 0 1.3906701219673681e+00
*
* Real pole n. 84
CS_84 NS_84 0 9.9999999999999998e-13
RS_84 NS_84 0 6.6287934454477863e+01
GS_84_5 0 NS_84 NA_5 0 1.3906701219673681e+00
*
* Real pole n. 85
CS_85 NS_85 0 9.9999999999999998e-13
RS_85 NS_85 0 5.4647183375290433e+02
GS_85_5 0 NS_85 NA_5 0 1.3906701219673681e+00
*
* Real pole n. 86
CS_86 NS_86 0 9.9999999999999998e-13
RS_86 NS_86 0 3.8169396682972065e+03
GS_86_5 0 NS_86 NA_5 0 1.3906701219673681e+00
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 2.1530817355819540e+01
RS_88 NS_88 0 2.1530817355819540e+01
GL_87 0 NS_87 NS_88 0 2.8893552838207953e-01
GL_88 0 NS_88 NS_87 0 -2.8893552838207953e-01
GS_87_5 0 NS_87 NA_5 0 1.3906701219673681e+00
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 1.7704391175337044e+01
RS_90 NS_90 0 1.7704391175337044e+01
GL_89 0 NS_89 NS_90 0 2.4113766587096394e-01
GL_90 0 NS_90 NS_89 0 -2.4113766587096394e-01
GS_89_5 0 NS_89 NA_5 0 1.3906701219673681e+00
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 1.5980319858751495e+01
RS_92 NS_92 0 1.5980319858751495e+01
GL_91 0 NS_91 NS_92 0 2.0836264676973826e-01
GL_92 0 NS_92 NS_91 0 -2.0836264676973826e-01
GS_91_5 0 NS_91 NA_5 0 1.3906701219673681e+00
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 1.5652313341768849e+01
RS_94 NS_94 0 1.5652313341768847e+01
GL_93 0 NS_93 NS_94 0 1.5274998946760082e-01
GL_94 0 NS_94 NS_93 0 -1.5274998946760082e-01
GS_93_5 0 NS_93 NA_5 0 1.3906701219673681e+00
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 1.5016887791939077e+01
RS_96 NS_96 0 1.5016887791939077e+01
GL_95 0 NS_95 NS_96 0 1.2573527610391108e-01
GL_96 0 NS_96 NS_95 0 -1.2573527610391108e-01
GS_95_5 0 NS_95 NA_5 0 1.3906701219673681e+00
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 1.9705893378385916e+01
RS_98 NS_98 0 1.9705893378385916e+01
GL_97 0 NS_97 NS_98 0 1.2264058452613225e-01
GL_98 0 NS_98 NS_97 0 -1.2264058452613225e-01
GS_97_5 0 NS_97 NA_5 0 1.3906701219673681e+00
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 1.7719166159098595e+01
RS_100 NS_100 0 1.7719166159098595e+01
GL_99 0 NS_99 NS_100 0 7.0127888352005202e-02
GL_100 0 NS_100 NS_99 0 -7.0127888352005202e-02
GS_99_5 0 NS_99 NA_5 0 1.3906701219673681e+00
*
* Real pole n. 101
CS_101 NS_101 0 9.9999999999999998e-13
RS_101 NS_101 0 4.5298699859481095e+00
GS_101_6 0 NS_101 NA_6 0 1.3906701219673681e+00
*
* Real pole n. 102
CS_102 NS_102 0 9.9999999999999998e-13
RS_102 NS_102 0 1.1221187714172293e+01
GS_102_6 0 NS_102 NA_6 0 1.3906701219673681e+00
*
* Real pole n. 103
CS_103 NS_103 0 9.9999999999999998e-13
RS_103 NS_103 0 1.8217191146854518e+01
GS_103_6 0 NS_103 NA_6 0 1.3906701219673681e+00
*
* Real pole n. 104
CS_104 NS_104 0 9.9999999999999998e-13
RS_104 NS_104 0 6.6287934454477863e+01
GS_104_6 0 NS_104 NA_6 0 1.3906701219673681e+00
*
* Real pole n. 105
CS_105 NS_105 0 9.9999999999999998e-13
RS_105 NS_105 0 5.4647183375290433e+02
GS_105_6 0 NS_105 NA_6 0 1.3906701219673681e+00
*
* Real pole n. 106
CS_106 NS_106 0 9.9999999999999998e-13
RS_106 NS_106 0 3.8169396682972065e+03
GS_106_6 0 NS_106 NA_6 0 1.3906701219673681e+00
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 2.1530817355819540e+01
RS_108 NS_108 0 2.1530817355819540e+01
GL_107 0 NS_107 NS_108 0 2.8893552838207953e-01
GL_108 0 NS_108 NS_107 0 -2.8893552838207953e-01
GS_107_6 0 NS_107 NA_6 0 1.3906701219673681e+00
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 1.7704391175337044e+01
RS_110 NS_110 0 1.7704391175337044e+01
GL_109 0 NS_109 NS_110 0 2.4113766587096394e-01
GL_110 0 NS_110 NS_109 0 -2.4113766587096394e-01
GS_109_6 0 NS_109 NA_6 0 1.3906701219673681e+00
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 1.5980319858751495e+01
RS_112 NS_112 0 1.5980319858751495e+01
GL_111 0 NS_111 NS_112 0 2.0836264676973826e-01
GL_112 0 NS_112 NS_111 0 -2.0836264676973826e-01
GS_111_6 0 NS_111 NA_6 0 1.3906701219673681e+00
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 1.5652313341768849e+01
RS_114 NS_114 0 1.5652313341768847e+01
GL_113 0 NS_113 NS_114 0 1.5274998946760082e-01
GL_114 0 NS_114 NS_113 0 -1.5274998946760082e-01
GS_113_6 0 NS_113 NA_6 0 1.3906701219673681e+00
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 1.5016887791939077e+01
RS_116 NS_116 0 1.5016887791939077e+01
GL_115 0 NS_115 NS_116 0 1.2573527610391108e-01
GL_116 0 NS_116 NS_115 0 -1.2573527610391108e-01
GS_115_6 0 NS_115 NA_6 0 1.3906701219673681e+00
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 1.9705893378385916e+01
RS_118 NS_118 0 1.9705893378385916e+01
GL_117 0 NS_117 NS_118 0 1.2264058452613225e-01
GL_118 0 NS_118 NS_117 0 -1.2264058452613225e-01
GS_117_6 0 NS_117 NA_6 0 1.3906701219673681e+00
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 1.7719166159098595e+01
RS_120 NS_120 0 1.7719166159098595e+01
GL_119 0 NS_119 NS_120 0 7.0127888352005202e-02
GL_120 0 NS_120 NS_119 0 -7.0127888352005202e-02
GS_119_6 0 NS_119 NA_6 0 1.3906701219673681e+00
*
* Real pole n. 121
CS_121 NS_121 0 9.9999999999999998e-13
RS_121 NS_121 0 4.5298699859481095e+00
GS_121_7 0 NS_121 NA_7 0 1.3906701219673681e+00
*
* Real pole n. 122
CS_122 NS_122 0 9.9999999999999998e-13
RS_122 NS_122 0 1.1221187714172293e+01
GS_122_7 0 NS_122 NA_7 0 1.3906701219673681e+00
*
* Real pole n. 123
CS_123 NS_123 0 9.9999999999999998e-13
RS_123 NS_123 0 1.8217191146854518e+01
GS_123_7 0 NS_123 NA_7 0 1.3906701219673681e+00
*
* Real pole n. 124
CS_124 NS_124 0 9.9999999999999998e-13
RS_124 NS_124 0 6.6287934454477863e+01
GS_124_7 0 NS_124 NA_7 0 1.3906701219673681e+00
*
* Real pole n. 125
CS_125 NS_125 0 9.9999999999999998e-13
RS_125 NS_125 0 5.4647183375290433e+02
GS_125_7 0 NS_125 NA_7 0 1.3906701219673681e+00
*
* Real pole n. 126
CS_126 NS_126 0 9.9999999999999998e-13
RS_126 NS_126 0 3.8169396682972065e+03
GS_126_7 0 NS_126 NA_7 0 1.3906701219673681e+00
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 2.1530817355819540e+01
RS_128 NS_128 0 2.1530817355819540e+01
GL_127 0 NS_127 NS_128 0 2.8893552838207953e-01
GL_128 0 NS_128 NS_127 0 -2.8893552838207953e-01
GS_127_7 0 NS_127 NA_7 0 1.3906701219673681e+00
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 1.7704391175337044e+01
RS_130 NS_130 0 1.7704391175337044e+01
GL_129 0 NS_129 NS_130 0 2.4113766587096394e-01
GL_130 0 NS_130 NS_129 0 -2.4113766587096394e-01
GS_129_7 0 NS_129 NA_7 0 1.3906701219673681e+00
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 1.5980319858751495e+01
RS_132 NS_132 0 1.5980319858751495e+01
GL_131 0 NS_131 NS_132 0 2.0836264676973826e-01
GL_132 0 NS_132 NS_131 0 -2.0836264676973826e-01
GS_131_7 0 NS_131 NA_7 0 1.3906701219673681e+00
*
* Complex pair n. 133/134
CS_133 NS_133 0 9.9999999999999998e-13
CS_134 NS_134 0 9.9999999999999998e-13
RS_133 NS_133 0 1.5652313341768849e+01
RS_134 NS_134 0 1.5652313341768847e+01
GL_133 0 NS_133 NS_134 0 1.5274998946760082e-01
GL_134 0 NS_134 NS_133 0 -1.5274998946760082e-01
GS_133_7 0 NS_133 NA_7 0 1.3906701219673681e+00
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 1.5016887791939077e+01
RS_136 NS_136 0 1.5016887791939077e+01
GL_135 0 NS_135 NS_136 0 1.2573527610391108e-01
GL_136 0 NS_136 NS_135 0 -1.2573527610391108e-01
GS_135_7 0 NS_135 NA_7 0 1.3906701219673681e+00
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 1.9705893378385916e+01
RS_138 NS_138 0 1.9705893378385916e+01
GL_137 0 NS_137 NS_138 0 1.2264058452613225e-01
GL_138 0 NS_138 NS_137 0 -1.2264058452613225e-01
GS_137_7 0 NS_137 NA_7 0 1.3906701219673681e+00
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 1.7719166159098595e+01
RS_140 NS_140 0 1.7719166159098595e+01
GL_139 0 NS_139 NS_140 0 7.0127888352005202e-02
GL_140 0 NS_140 NS_139 0 -7.0127888352005202e-02
GS_139_7 0 NS_139 NA_7 0 1.3906701219673681e+00
*
* Real pole n. 141
CS_141 NS_141 0 9.9999999999999998e-13
RS_141 NS_141 0 4.5298699859481095e+00
GS_141_8 0 NS_141 NA_8 0 1.3906701219673681e+00
*
* Real pole n. 142
CS_142 NS_142 0 9.9999999999999998e-13
RS_142 NS_142 0 1.1221187714172293e+01
GS_142_8 0 NS_142 NA_8 0 1.3906701219673681e+00
*
* Real pole n. 143
CS_143 NS_143 0 9.9999999999999998e-13
RS_143 NS_143 0 1.8217191146854518e+01
GS_143_8 0 NS_143 NA_8 0 1.3906701219673681e+00
*
* Real pole n. 144
CS_144 NS_144 0 9.9999999999999998e-13
RS_144 NS_144 0 6.6287934454477863e+01
GS_144_8 0 NS_144 NA_8 0 1.3906701219673681e+00
*
* Real pole n. 145
CS_145 NS_145 0 9.9999999999999998e-13
RS_145 NS_145 0 5.4647183375290433e+02
GS_145_8 0 NS_145 NA_8 0 1.3906701219673681e+00
*
* Real pole n. 146
CS_146 NS_146 0 9.9999999999999998e-13
RS_146 NS_146 0 3.8169396682972065e+03
GS_146_8 0 NS_146 NA_8 0 1.3906701219673681e+00
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 2.1530817355819540e+01
RS_148 NS_148 0 2.1530817355819540e+01
GL_147 0 NS_147 NS_148 0 2.8893552838207953e-01
GL_148 0 NS_148 NS_147 0 -2.8893552838207953e-01
GS_147_8 0 NS_147 NA_8 0 1.3906701219673681e+00
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 1.7704391175337044e+01
RS_150 NS_150 0 1.7704391175337044e+01
GL_149 0 NS_149 NS_150 0 2.4113766587096394e-01
GL_150 0 NS_150 NS_149 0 -2.4113766587096394e-01
GS_149_8 0 NS_149 NA_8 0 1.3906701219673681e+00
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 1.5980319858751495e+01
RS_152 NS_152 0 1.5980319858751495e+01
GL_151 0 NS_151 NS_152 0 2.0836264676973826e-01
GL_152 0 NS_152 NS_151 0 -2.0836264676973826e-01
GS_151_8 0 NS_151 NA_8 0 1.3906701219673681e+00
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 1.5652313341768849e+01
RS_154 NS_154 0 1.5652313341768847e+01
GL_153 0 NS_153 NS_154 0 1.5274998946760082e-01
GL_154 0 NS_154 NS_153 0 -1.5274998946760082e-01
GS_153_8 0 NS_153 NA_8 0 1.3906701219673681e+00
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 1.5016887791939077e+01
RS_156 NS_156 0 1.5016887791939077e+01
GL_155 0 NS_155 NS_156 0 1.2573527610391108e-01
GL_156 0 NS_156 NS_155 0 -1.2573527610391108e-01
GS_155_8 0 NS_155 NA_8 0 1.3906701219673681e+00
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 1.9705893378385916e+01
RS_158 NS_158 0 1.9705893378385916e+01
GL_157 0 NS_157 NS_158 0 1.2264058452613225e-01
GL_158 0 NS_158 NS_157 0 -1.2264058452613225e-01
GS_157_8 0 NS_157 NA_8 0 1.3906701219673681e+00
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 1.7719166159098595e+01
RS_160 NS_160 0 1.7719166159098595e+01
GL_159 0 NS_159 NS_160 0 7.0127888352005202e-02
GL_160 0 NS_160 NS_159 0 -7.0127888352005202e-02
GS_159_8 0 NS_159 NA_8 0 1.3906701219673681e+00
*
* Real pole n. 161
CS_161 NS_161 0 9.9999999999999998e-13
RS_161 NS_161 0 4.5298699859481095e+00
GS_161_9 0 NS_161 NA_9 0 1.3906701219673681e+00
*
* Real pole n. 162
CS_162 NS_162 0 9.9999999999999998e-13
RS_162 NS_162 0 1.1221187714172293e+01
GS_162_9 0 NS_162 NA_9 0 1.3906701219673681e+00
*
* Real pole n. 163
CS_163 NS_163 0 9.9999999999999998e-13
RS_163 NS_163 0 1.8217191146854518e+01
GS_163_9 0 NS_163 NA_9 0 1.3906701219673681e+00
*
* Real pole n. 164
CS_164 NS_164 0 9.9999999999999998e-13
RS_164 NS_164 0 6.6287934454477863e+01
GS_164_9 0 NS_164 NA_9 0 1.3906701219673681e+00
*
* Real pole n. 165
CS_165 NS_165 0 9.9999999999999998e-13
RS_165 NS_165 0 5.4647183375290433e+02
GS_165_9 0 NS_165 NA_9 0 1.3906701219673681e+00
*
* Real pole n. 166
CS_166 NS_166 0 9.9999999999999998e-13
RS_166 NS_166 0 3.8169396682972065e+03
GS_166_9 0 NS_166 NA_9 0 1.3906701219673681e+00
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 2.1530817355819540e+01
RS_168 NS_168 0 2.1530817355819540e+01
GL_167 0 NS_167 NS_168 0 2.8893552838207953e-01
GL_168 0 NS_168 NS_167 0 -2.8893552838207953e-01
GS_167_9 0 NS_167 NA_9 0 1.3906701219673681e+00
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 1.7704391175337044e+01
RS_170 NS_170 0 1.7704391175337044e+01
GL_169 0 NS_169 NS_170 0 2.4113766587096394e-01
GL_170 0 NS_170 NS_169 0 -2.4113766587096394e-01
GS_169_9 0 NS_169 NA_9 0 1.3906701219673681e+00
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 1.5980319858751495e+01
RS_172 NS_172 0 1.5980319858751495e+01
GL_171 0 NS_171 NS_172 0 2.0836264676973826e-01
GL_172 0 NS_172 NS_171 0 -2.0836264676973826e-01
GS_171_9 0 NS_171 NA_9 0 1.3906701219673681e+00
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 1.5652313341768849e+01
RS_174 NS_174 0 1.5652313341768847e+01
GL_173 0 NS_173 NS_174 0 1.5274998946760082e-01
GL_174 0 NS_174 NS_173 0 -1.5274998946760082e-01
GS_173_9 0 NS_173 NA_9 0 1.3906701219673681e+00
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 1.5016887791939077e+01
RS_176 NS_176 0 1.5016887791939077e+01
GL_175 0 NS_175 NS_176 0 1.2573527610391108e-01
GL_176 0 NS_176 NS_175 0 -1.2573527610391108e-01
GS_175_9 0 NS_175 NA_9 0 1.3906701219673681e+00
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 1.9705893378385916e+01
RS_178 NS_178 0 1.9705893378385916e+01
GL_177 0 NS_177 NS_178 0 1.2264058452613225e-01
GL_178 0 NS_178 NS_177 0 -1.2264058452613225e-01
GS_177_9 0 NS_177 NA_9 0 1.3906701219673681e+00
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 1.7719166159098595e+01
RS_180 NS_180 0 1.7719166159098595e+01
GL_179 0 NS_179 NS_180 0 7.0127888352005202e-02
GL_180 0 NS_180 NS_179 0 -7.0127888352005202e-02
GS_179_9 0 NS_179 NA_9 0 1.3906701219673681e+00
*
* Real pole n. 181
CS_181 NS_181 0 9.9999999999999998e-13
RS_181 NS_181 0 4.5298699859481095e+00
GS_181_10 0 NS_181 NA_10 0 1.3906701219673681e+00
*
* Real pole n. 182
CS_182 NS_182 0 9.9999999999999998e-13
RS_182 NS_182 0 1.1221187714172293e+01
GS_182_10 0 NS_182 NA_10 0 1.3906701219673681e+00
*
* Real pole n. 183
CS_183 NS_183 0 9.9999999999999998e-13
RS_183 NS_183 0 1.8217191146854518e+01
GS_183_10 0 NS_183 NA_10 0 1.3906701219673681e+00
*
* Real pole n. 184
CS_184 NS_184 0 9.9999999999999998e-13
RS_184 NS_184 0 6.6287934454477863e+01
GS_184_10 0 NS_184 NA_10 0 1.3906701219673681e+00
*
* Real pole n. 185
CS_185 NS_185 0 9.9999999999999998e-13
RS_185 NS_185 0 5.4647183375290433e+02
GS_185_10 0 NS_185 NA_10 0 1.3906701219673681e+00
*
* Real pole n. 186
CS_186 NS_186 0 9.9999999999999998e-13
RS_186 NS_186 0 3.8169396682972065e+03
GS_186_10 0 NS_186 NA_10 0 1.3906701219673681e+00
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 2.1530817355819540e+01
RS_188 NS_188 0 2.1530817355819540e+01
GL_187 0 NS_187 NS_188 0 2.8893552838207953e-01
GL_188 0 NS_188 NS_187 0 -2.8893552838207953e-01
GS_187_10 0 NS_187 NA_10 0 1.3906701219673681e+00
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 1.7704391175337044e+01
RS_190 NS_190 0 1.7704391175337044e+01
GL_189 0 NS_189 NS_190 0 2.4113766587096394e-01
GL_190 0 NS_190 NS_189 0 -2.4113766587096394e-01
GS_189_10 0 NS_189 NA_10 0 1.3906701219673681e+00
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 1.5980319858751495e+01
RS_192 NS_192 0 1.5980319858751495e+01
GL_191 0 NS_191 NS_192 0 2.0836264676973826e-01
GL_192 0 NS_192 NS_191 0 -2.0836264676973826e-01
GS_191_10 0 NS_191 NA_10 0 1.3906701219673681e+00
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 1.5652313341768849e+01
RS_194 NS_194 0 1.5652313341768847e+01
GL_193 0 NS_193 NS_194 0 1.5274998946760082e-01
GL_194 0 NS_194 NS_193 0 -1.5274998946760082e-01
GS_193_10 0 NS_193 NA_10 0 1.3906701219673681e+00
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 1.5016887791939077e+01
RS_196 NS_196 0 1.5016887791939077e+01
GL_195 0 NS_195 NS_196 0 1.2573527610391108e-01
GL_196 0 NS_196 NS_195 0 -1.2573527610391108e-01
GS_195_10 0 NS_195 NA_10 0 1.3906701219673681e+00
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 1.9705893378385916e+01
RS_198 NS_198 0 1.9705893378385916e+01
GL_197 0 NS_197 NS_198 0 1.2264058452613225e-01
GL_198 0 NS_198 NS_197 0 -1.2264058452613225e-01
GS_197_10 0 NS_197 NA_10 0 1.3906701219673681e+00
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 1.7719166159098595e+01
RS_200 NS_200 0 1.7719166159098595e+01
GL_199 0 NS_199 NS_200 0 7.0127888352005202e-02
GL_200 0 NS_200 NS_199 0 -7.0127888352005202e-02
GS_199_10 0 NS_199 NA_10 0 1.3906701219673681e+00
*
* Real pole n. 201
CS_201 NS_201 0 9.9999999999999998e-13
RS_201 NS_201 0 4.5298699859481095e+00
GS_201_11 0 NS_201 NA_11 0 1.3906701219673681e+00
*
* Real pole n. 202
CS_202 NS_202 0 9.9999999999999998e-13
RS_202 NS_202 0 1.1221187714172293e+01
GS_202_11 0 NS_202 NA_11 0 1.3906701219673681e+00
*
* Real pole n. 203
CS_203 NS_203 0 9.9999999999999998e-13
RS_203 NS_203 0 1.8217191146854518e+01
GS_203_11 0 NS_203 NA_11 0 1.3906701219673681e+00
*
* Real pole n. 204
CS_204 NS_204 0 9.9999999999999998e-13
RS_204 NS_204 0 6.6287934454477863e+01
GS_204_11 0 NS_204 NA_11 0 1.3906701219673681e+00
*
* Real pole n. 205
CS_205 NS_205 0 9.9999999999999998e-13
RS_205 NS_205 0 5.4647183375290433e+02
GS_205_11 0 NS_205 NA_11 0 1.3906701219673681e+00
*
* Real pole n. 206
CS_206 NS_206 0 9.9999999999999998e-13
RS_206 NS_206 0 3.8169396682972065e+03
GS_206_11 0 NS_206 NA_11 0 1.3906701219673681e+00
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 2.1530817355819540e+01
RS_208 NS_208 0 2.1530817355819540e+01
GL_207 0 NS_207 NS_208 0 2.8893552838207953e-01
GL_208 0 NS_208 NS_207 0 -2.8893552838207953e-01
GS_207_11 0 NS_207 NA_11 0 1.3906701219673681e+00
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 1.7704391175337044e+01
RS_210 NS_210 0 1.7704391175337044e+01
GL_209 0 NS_209 NS_210 0 2.4113766587096394e-01
GL_210 0 NS_210 NS_209 0 -2.4113766587096394e-01
GS_209_11 0 NS_209 NA_11 0 1.3906701219673681e+00
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 1.5980319858751495e+01
RS_212 NS_212 0 1.5980319858751495e+01
GL_211 0 NS_211 NS_212 0 2.0836264676973826e-01
GL_212 0 NS_212 NS_211 0 -2.0836264676973826e-01
GS_211_11 0 NS_211 NA_11 0 1.3906701219673681e+00
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 1.5652313341768849e+01
RS_214 NS_214 0 1.5652313341768847e+01
GL_213 0 NS_213 NS_214 0 1.5274998946760082e-01
GL_214 0 NS_214 NS_213 0 -1.5274998946760082e-01
GS_213_11 0 NS_213 NA_11 0 1.3906701219673681e+00
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 1.5016887791939077e+01
RS_216 NS_216 0 1.5016887791939077e+01
GL_215 0 NS_215 NS_216 0 1.2573527610391108e-01
GL_216 0 NS_216 NS_215 0 -1.2573527610391108e-01
GS_215_11 0 NS_215 NA_11 0 1.3906701219673681e+00
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 1.9705893378385916e+01
RS_218 NS_218 0 1.9705893378385916e+01
GL_217 0 NS_217 NS_218 0 1.2264058452613225e-01
GL_218 0 NS_218 NS_217 0 -1.2264058452613225e-01
GS_217_11 0 NS_217 NA_11 0 1.3906701219673681e+00
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 1.7719166159098595e+01
RS_220 NS_220 0 1.7719166159098595e+01
GL_219 0 NS_219 NS_220 0 7.0127888352005202e-02
GL_220 0 NS_220 NS_219 0 -7.0127888352005202e-02
GS_219_11 0 NS_219 NA_11 0 1.3906701219673681e+00
*
* Real pole n. 221
CS_221 NS_221 0 9.9999999999999998e-13
RS_221 NS_221 0 4.5298699859481095e+00
GS_221_12 0 NS_221 NA_12 0 1.3906701219673681e+00
*
* Real pole n. 222
CS_222 NS_222 0 9.9999999999999998e-13
RS_222 NS_222 0 1.1221187714172293e+01
GS_222_12 0 NS_222 NA_12 0 1.3906701219673681e+00
*
* Real pole n. 223
CS_223 NS_223 0 9.9999999999999998e-13
RS_223 NS_223 0 1.8217191146854518e+01
GS_223_12 0 NS_223 NA_12 0 1.3906701219673681e+00
*
* Real pole n. 224
CS_224 NS_224 0 9.9999999999999998e-13
RS_224 NS_224 0 6.6287934454477863e+01
GS_224_12 0 NS_224 NA_12 0 1.3906701219673681e+00
*
* Real pole n. 225
CS_225 NS_225 0 9.9999999999999998e-13
RS_225 NS_225 0 5.4647183375290433e+02
GS_225_12 0 NS_225 NA_12 0 1.3906701219673681e+00
*
* Real pole n. 226
CS_226 NS_226 0 9.9999999999999998e-13
RS_226 NS_226 0 3.8169396682972065e+03
GS_226_12 0 NS_226 NA_12 0 1.3906701219673681e+00
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 2.1530817355819540e+01
RS_228 NS_228 0 2.1530817355819540e+01
GL_227 0 NS_227 NS_228 0 2.8893552838207953e-01
GL_228 0 NS_228 NS_227 0 -2.8893552838207953e-01
GS_227_12 0 NS_227 NA_12 0 1.3906701219673681e+00
*
* Complex pair n. 229/230
CS_229 NS_229 0 9.9999999999999998e-13
CS_230 NS_230 0 9.9999999999999998e-13
RS_229 NS_229 0 1.7704391175337044e+01
RS_230 NS_230 0 1.7704391175337044e+01
GL_229 0 NS_229 NS_230 0 2.4113766587096394e-01
GL_230 0 NS_230 NS_229 0 -2.4113766587096394e-01
GS_229_12 0 NS_229 NA_12 0 1.3906701219673681e+00
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 1.5980319858751495e+01
RS_232 NS_232 0 1.5980319858751495e+01
GL_231 0 NS_231 NS_232 0 2.0836264676973826e-01
GL_232 0 NS_232 NS_231 0 -2.0836264676973826e-01
GS_231_12 0 NS_231 NA_12 0 1.3906701219673681e+00
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 1.5652313341768849e+01
RS_234 NS_234 0 1.5652313341768847e+01
GL_233 0 NS_233 NS_234 0 1.5274998946760082e-01
GL_234 0 NS_234 NS_233 0 -1.5274998946760082e-01
GS_233_12 0 NS_233 NA_12 0 1.3906701219673681e+00
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 1.5016887791939077e+01
RS_236 NS_236 0 1.5016887791939077e+01
GL_235 0 NS_235 NS_236 0 1.2573527610391108e-01
GL_236 0 NS_236 NS_235 0 -1.2573527610391108e-01
GS_235_12 0 NS_235 NA_12 0 1.3906701219673681e+00
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 1.9705893378385916e+01
RS_238 NS_238 0 1.9705893378385916e+01
GL_237 0 NS_237 NS_238 0 1.2264058452613225e-01
GL_238 0 NS_238 NS_237 0 -1.2264058452613225e-01
GS_237_12 0 NS_237 NA_12 0 1.3906701219673681e+00
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 1.7719166159098595e+01
RS_240 NS_240 0 1.7719166159098595e+01
GL_239 0 NS_239 NS_240 0 7.0127888352005202e-02
GL_240 0 NS_240 NS_239 0 -7.0127888352005202e-02
GS_239_12 0 NS_239 NA_12 0 1.3906701219673681e+00
*
******************************


.ends
*******************
* End of subcircuit
*******************
