**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [12 6 56] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_3_BoardVia_withStub
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 -6.3310249348106792e-02
GC_1_2 b_1 NI_1 NS_2 0 1.5489071479615136e-02
GC_1_3 b_1 NI_1 NS_3 0 3.7815962075700093e-03
GC_1_4 b_1 NI_1 NS_4 0 2.3857091210699190e-03
GC_1_5 b_1 NI_1 NS_5 0 1.2285349351785909e-02
GC_1_6 b_1 NI_1 NS_6 0 -1.1042949136476257e-03
GC_1_7 b_1 NI_1 NS_7 0 7.0928419201913076e-04
GC_1_8 b_1 NI_1 NS_8 0 1.7664716366658372e-03
GC_1_9 b_1 NI_1 NS_9 0 1.1726170902720113e-02
GC_1_10 b_1 NI_1 NS_10 0 8.1088721873762513e-03
GC_1_11 b_1 NI_1 NS_11 0 4.3589557693481286e-04
GC_1_12 b_1 NI_1 NS_12 0 9.1058784458553890e-04
GC_1_13 b_1 NI_1 NS_13 0 5.5740303151044389e-03
GC_1_14 b_1 NI_1 NS_14 0 -9.4376752971391518e-04
GC_1_15 b_1 NI_1 NS_15 0 1.0411245133568699e-04
GC_1_16 b_1 NI_1 NS_16 0 1.5028948048868996e-03
GC_1_17 b_1 NI_1 NS_17 0 8.1095499515330249e-03
GC_1_18 b_1 NI_1 NS_18 0 -4.9462221923222754e-04
GC_1_19 b_1 NI_1 NS_19 0 4.0456181613621961e-03
GC_1_20 b_1 NI_1 NS_20 0 3.4129156498171991e-03
GC_1_21 b_1 NI_1 NS_21 0 1.2551091452211885e-04
GC_1_22 b_1 NI_1 NS_22 0 5.7540042747057855e-05
GC_1_23 b_1 NI_1 NS_23 0 2.8879262839855966e-03
GC_1_24 b_1 NI_1 NS_24 0 6.6305753940859640e-03
GC_1_25 b_1 NI_1 NS_25 0 6.0995952426757866e-04
GC_1_26 b_1 NI_1 NS_26 0 8.8109255891160508e-05
GC_1_27 b_1 NI_1 NS_27 0 -1.3121095151922990e-04
GC_1_28 b_1 NI_1 NS_28 0 1.4439945021934582e-04
GC_1_29 b_1 NI_1 NS_29 0 6.3593264160131323e-05
GC_1_30 b_1 NI_1 NS_30 0 1.2894602167955172e-04
GC_1_31 b_1 NI_1 NS_31 0 3.2635760814943166e-05
GC_1_32 b_1 NI_1 NS_32 0 1.8295988437350249e-05
GC_1_33 b_1 NI_1 NS_33 0 -4.5547032556436234e-04
GC_1_34 b_1 NI_1 NS_34 0 4.5993484435320380e-03
GC_1_35 b_1 NI_1 NS_35 0 -6.8590665240567845e-07
GC_1_36 b_1 NI_1 NS_36 0 -4.2179232692269116e-05
GC_1_37 b_1 NI_1 NS_37 0 8.2402630911276463e-04
GC_1_38 b_1 NI_1 NS_38 0 8.7513436907590391e-04
GC_1_39 b_1 NI_1 NS_39 0 -2.1024110883265945e-03
GC_1_40 b_1 NI_1 NS_40 0 1.4125821056477747e-03
GC_1_41 b_1 NI_1 NS_41 0 1.2559340909011878e-04
GC_1_42 b_1 NI_1 NS_42 0 1.6557673878857474e-04
GC_1_43 b_1 NI_1 NS_43 0 4.5742598168811985e-08
GC_1_44 b_1 NI_1 NS_44 0 -1.3727376573707185e-06
GC_1_45 b_1 NI_1 NS_45 0 7.2120788122911843e-06
GC_1_46 b_1 NI_1 NS_46 0 1.8004024483835741e-05
GC_1_47 b_1 NI_1 NS_47 0 2.5815460776128663e-04
GC_1_48 b_1 NI_1 NS_48 0 -8.5169801914699396e-05
GC_1_49 b_1 NI_1 NS_49 0 3.2492230381986094e-06
GC_1_50 b_1 NI_1 NS_50 0 3.1900127830695705e-05
GC_1_51 b_1 NI_1 NS_51 0 9.5893189209557935e-06
GC_1_52 b_1 NI_1 NS_52 0 2.5417050618643812e-06
GC_1_53 b_1 NI_1 NS_53 0 -1.6055914192190649e-05
GC_1_54 b_1 NI_1 NS_54 0 1.7587350959668492e-05
GC_1_55 b_1 NI_1 NS_55 0 3.1002571521558607e-05
GC_1_56 b_1 NI_1 NS_56 0 -1.7395933000908362e-05
GC_1_57 b_1 NI_1 NS_57 0 -1.5506986626855889e-02
GC_1_58 b_1 NI_1 NS_58 0 1.2182092646436240e-02
GC_1_59 b_1 NI_1 NS_59 0 -2.2350826156665648e-03
GC_1_60 b_1 NI_1 NS_60 0 1.2891383970963137e-03
GC_1_61 b_1 NI_1 NS_61 0 -2.0941791550019928e-03
GC_1_62 b_1 NI_1 NS_62 0 4.4904251475437647e-03
GC_1_63 b_1 NI_1 NS_63 0 -1.0314936662724013e-03
GC_1_64 b_1 NI_1 NS_64 0 -2.9828055445532083e-03
GC_1_65 b_1 NI_1 NS_65 0 -1.2456170311631390e-02
GC_1_66 b_1 NI_1 NS_66 0 -3.1962467646465429e-03
GC_1_67 b_1 NI_1 NS_67 0 3.4147725722953609e-04
GC_1_68 b_1 NI_1 NS_68 0 -1.9124658127477439e-04
GC_1_69 b_1 NI_1 NS_69 0 3.4168713016576448e-03
GC_1_70 b_1 NI_1 NS_70 0 -2.1288944255163920e-04
GC_1_71 b_1 NI_1 NS_71 0 7.7650908752570098e-04
GC_1_72 b_1 NI_1 NS_72 0 7.4827476423032437e-04
GC_1_73 b_1 NI_1 NS_73 0 4.5561429187660468e-03
GC_1_74 b_1 NI_1 NS_74 0 -1.8590671235830386e-03
GC_1_75 b_1 NI_1 NS_75 0 -8.8966181897233280e-04
GC_1_76 b_1 NI_1 NS_76 0 -2.9542410422275149e-04
GC_1_77 b_1 NI_1 NS_77 0 -1.3763886874762265e-04
GC_1_78 b_1 NI_1 NS_78 0 2.4470474728122513e-07
GC_1_79 b_1 NI_1 NS_79 0 6.1739101357005787e-03
GC_1_80 b_1 NI_1 NS_80 0 -2.1833436137421035e-04
GC_1_81 b_1 NI_1 NS_81 0 -8.0641780117096499e-04
GC_1_82 b_1 NI_1 NS_82 0 -1.6305320855992316e-04
GC_1_83 b_1 NI_1 NS_83 0 -9.2428603678946719e-05
GC_1_84 b_1 NI_1 NS_84 0 5.0339566512763872e-05
GC_1_85 b_1 NI_1 NS_85 0 -2.1532831514699892e-04
GC_1_86 b_1 NI_1 NS_86 0 2.0220368589888598e-04
GC_1_87 b_1 NI_1 NS_87 0 -1.5103864256728333e-04
GC_1_88 b_1 NI_1 NS_88 0 -6.2868059979265500e-05
GC_1_89 b_1 NI_1 NS_89 0 -1.0615296539246589e-03
GC_1_90 b_1 NI_1 NS_90 0 9.8325178790836820e-04
GC_1_91 b_1 NI_1 NS_91 0 -4.1832230681170165e-05
GC_1_92 b_1 NI_1 NS_92 0 7.8578848690040803e-05
GC_1_93 b_1 NI_1 NS_93 0 -9.0811809111353270e-05
GC_1_94 b_1 NI_1 NS_94 0 -2.4836285925629092e-04
GC_1_95 b_1 NI_1 NS_95 0 3.0488610919346646e-05
GC_1_96 b_1 NI_1 NS_96 0 -6.5365301005044368e-04
GC_1_97 b_1 NI_1 NS_97 0 1.6334965855561976e-04
GC_1_98 b_1 NI_1 NS_98 0 1.3708115485054238e-04
GC_1_99 b_1 NI_1 NS_99 0 9.6295166841799058e-07
GC_1_100 b_1 NI_1 NS_100 0 7.1860456718614654e-07
GC_1_101 b_1 NI_1 NS_101 0 1.4807160975745252e-06
GC_1_102 b_1 NI_1 NS_102 0 -6.0732255439116969e-06
GC_1_103 b_1 NI_1 NS_103 0 -1.0954991206418223e-04
GC_1_104 b_1 NI_1 NS_104 0 2.4349477768981441e-05
GC_1_105 b_1 NI_1 NS_105 0 4.0184396146067342e-06
GC_1_106 b_1 NI_1 NS_106 0 -1.3923577451945675e-05
GC_1_107 b_1 NI_1 NS_107 0 1.0945361948776527e-05
GC_1_108 b_1 NI_1 NS_108 0 -3.7775688070779525e-06
GC_1_109 b_1 NI_1 NS_109 0 1.3782754853249001e-05
GC_1_110 b_1 NI_1 NS_110 0 2.6818741354552976e-05
GC_1_111 b_1 NI_1 NS_111 0 -7.6320503897100191e-06
GC_1_112 b_1 NI_1 NS_112 0 -4.5971950534550427e-05
GC_1_113 b_1 NI_1 NS_113 0 -3.0061678552903925e-02
GC_1_114 b_1 NI_1 NS_114 0 1.7198922485858555e-03
GC_1_115 b_1 NI_1 NS_115 0 3.6993481782388389e-03
GC_1_116 b_1 NI_1 NS_116 0 2.5857513434126194e-03
GC_1_117 b_1 NI_1 NS_117 0 -5.7084431512846798e-03
GC_1_118 b_1 NI_1 NS_118 0 -6.5718121671517055e-03
GC_1_119 b_1 NI_1 NS_119 0 3.6822857173963129e-03
GC_1_120 b_1 NI_1 NS_120 0 1.5264879083309931e-03
GC_1_121 b_1 NI_1 NS_121 0 1.0503292478052081e-02
GC_1_122 b_1 NI_1 NS_122 0 -1.1738965848328817e-02
GC_1_123 b_1 NI_1 NS_123 0 -3.1359001327151934e-04
GC_1_124 b_1 NI_1 NS_124 0 3.7815499838037296e-04
GC_1_125 b_1 NI_1 NS_125 0 8.9978538010014771e-03
GC_1_126 b_1 NI_1 NS_126 0 3.2733639668066812e-03
GC_1_127 b_1 NI_1 NS_127 0 3.0707357152287047e-04
GC_1_128 b_1 NI_1 NS_128 0 2.1644017065025711e-03
GC_1_129 b_1 NI_1 NS_129 0 6.9122911817218911e-03
GC_1_130 b_1 NI_1 NS_130 0 -9.4757062618381943e-05
GC_1_131 b_1 NI_1 NS_131 0 2.1100430980769665e-03
GC_1_132 b_1 NI_1 NS_132 0 3.5101180094774002e-03
GC_1_133 b_1 NI_1 NS_133 0 2.4907149336465129e-04
GC_1_134 b_1 NI_1 NS_134 0 7.6313269789032544e-05
GC_1_135 b_1 NI_1 NS_135 0 -2.9575680320302546e-03
GC_1_136 b_1 NI_1 NS_136 0 1.0405969697251089e-02
GC_1_137 b_1 NI_1 NS_137 0 1.1307156915983676e-03
GC_1_138 b_1 NI_1 NS_138 0 2.1733352820325037e-04
GC_1_139 b_1 NI_1 NS_139 0 -3.3581849914669283e-04
GC_1_140 b_1 NI_1 NS_140 0 1.3357878838939858e-04
GC_1_141 b_1 NI_1 NS_141 0 -1.0068490823996658e-04
GC_1_142 b_1 NI_1 NS_142 0 2.6008483043971759e-04
GC_1_143 b_1 NI_1 NS_143 0 -5.6162723457417680e-05
GC_1_144 b_1 NI_1 NS_144 0 1.6912398887399511e-05
GC_1_145 b_1 NI_1 NS_145 0 -1.5928408893947934e-03
GC_1_146 b_1 NI_1 NS_146 0 -4.3090501890842552e-03
GC_1_147 b_1 NI_1 NS_147 0 1.0073688950404938e-04
GC_1_148 b_1 NI_1 NS_148 0 -2.1165660277760593e-05
GC_1_149 b_1 NI_1 NS_149 0 -4.4324151069342671e-04
GC_1_150 b_1 NI_1 NS_150 0 1.5110486192685148e-03
GC_1_151 b_1 NI_1 NS_151 0 -2.4284296528715804e-04
GC_1_152 b_1 NI_1 NS_152 0 2.2524629335645922e-03
GC_1_153 b_1 NI_1 NS_153 0 3.5591338445224562e-05
GC_1_154 b_1 NI_1 NS_154 0 9.5883026259153967e-05
GC_1_155 b_1 NI_1 NS_155 0 -1.1070332931803911e-07
GC_1_156 b_1 NI_1 NS_156 0 -2.0307617894100640e-07
GC_1_157 b_1 NI_1 NS_157 0 4.0069034497285557e-06
GC_1_158 b_1 NI_1 NS_158 0 2.9542911482612969e-06
GC_1_159 b_1 NI_1 NS_159 0 3.1009779820251092e-05
GC_1_160 b_1 NI_1 NS_160 0 -4.7582579358292751e-05
GC_1_161 b_1 NI_1 NS_161 0 3.9521651290588850e-06
GC_1_162 b_1 NI_1 NS_162 0 7.8537545182054178e-06
GC_1_163 b_1 NI_1 NS_163 0 5.7934194423664700e-06
GC_1_164 b_1 NI_1 NS_164 0 -8.5733407083817506e-07
GC_1_165 b_1 NI_1 NS_165 0 -2.0764588293281909e-06
GC_1_166 b_1 NI_1 NS_166 0 1.2093767465677475e-05
GC_1_167 b_1 NI_1 NS_167 0 8.5478539842394908e-06
GC_1_168 b_1 NI_1 NS_168 0 -1.6952655547687951e-05
GC_1_169 b_1 NI_1 NS_169 0 6.0535066632412191e-02
GC_1_170 b_1 NI_1 NS_170 0 -8.1708332951175157e-04
GC_1_171 b_1 NI_1 NS_171 0 -1.9120438285759487e-03
GC_1_172 b_1 NI_1 NS_172 0 2.2999153625500486e-03
GC_1_173 b_1 NI_1 NS_173 0 2.9401047194300362e-03
GC_1_174 b_1 NI_1 NS_174 0 1.1664003224791924e-04
GC_1_175 b_1 NI_1 NS_175 0 -4.9470419708674811e-03
GC_1_176 b_1 NI_1 NS_176 0 5.4589942198300168e-04
GC_1_177 b_1 NI_1 NS_177 0 -5.8274075655746840e-03
GC_1_178 b_1 NI_1 NS_178 0 1.1489937746495092e-02
GC_1_179 b_1 NI_1 NS_179 0 -5.6786859385071331e-04
GC_1_180 b_1 NI_1 NS_180 0 -1.0385963228401762e-04
GC_1_181 b_1 NI_1 NS_181 0 1.3568965921493940e-03
GC_1_182 b_1 NI_1 NS_182 0 -3.5525847751272017e-03
GC_1_183 b_1 NI_1 NS_183 0 7.0463864870200059e-04
GC_1_184 b_1 NI_1 NS_184 0 1.4367273921531067e-03
GC_1_185 b_1 NI_1 NS_185 0 -9.5147356303626148e-04
GC_1_186 b_1 NI_1 NS_186 0 1.0489586295444029e-03
GC_1_187 b_1 NI_1 NS_187 0 -5.9662103493487873e-03
GC_1_188 b_1 NI_1 NS_188 0 4.7372473498887626e-04
GC_1_189 b_1 NI_1 NS_189 0 -4.9267151388732972e-05
GC_1_190 b_1 NI_1 NS_190 0 -7.2311259961202324e-05
GC_1_191 b_1 NI_1 NS_191 0 3.0653951500635873e-04
GC_1_192 b_1 NI_1 NS_192 0 4.4832666209713998e-03
GC_1_193 b_1 NI_1 NS_193 0 -3.7029353569310831e-04
GC_1_194 b_1 NI_1 NS_194 0 -2.3078703100623188e-04
GC_1_195 b_1 NI_1 NS_195 0 -2.6502668606234649e-04
GC_1_196 b_1 NI_1 NS_196 0 -2.0110847216929799e-05
GC_1_197 b_1 NI_1 NS_197 0 -3.1761625275762489e-04
GC_1_198 b_1 NI_1 NS_198 0 3.4796407774774165e-04
GC_1_199 b_1 NI_1 NS_199 0 -1.9068453977067436e-04
GC_1_200 b_1 NI_1 NS_200 0 -3.0658727717185580e-05
GC_1_201 b_1 NI_1 NS_201 0 -6.4936291446574456e-03
GC_1_202 b_1 NI_1 NS_202 0 -1.2733897529665888e-03
GC_1_203 b_1 NI_1 NS_203 0 -1.1274157778041306e-05
GC_1_204 b_1 NI_1 NS_204 0 2.5829096361098794e-05
GC_1_205 b_1 NI_1 NS_205 0 -1.0252021384560210e-04
GC_1_206 b_1 NI_1 NS_206 0 7.0577862335119402e-04
GC_1_207 b_1 NI_1 NS_207 0 -6.8789583060754271e-04
GC_1_208 b_1 NI_1 NS_208 0 -2.1624420222072418e-03
GC_1_209 b_1 NI_1 NS_209 0 1.8350642472146714e-04
GC_1_210 b_1 NI_1 NS_210 0 8.9580574777626041e-05
GC_1_211 b_1 NI_1 NS_211 0 3.4689152015799329e-06
GC_1_212 b_1 NI_1 NS_212 0 2.7662353647993308e-06
GC_1_213 b_1 NI_1 NS_213 0 -6.0387414023949989e-06
GC_1_214 b_1 NI_1 NS_214 0 -1.1214784910992943e-05
GC_1_215 b_1 NI_1 NS_215 0 -5.9285862572646555e-05
GC_1_216 b_1 NI_1 NS_216 0 2.0581797754294084e-04
GC_1_217 b_1 NI_1 NS_217 0 -1.3231783038377544e-05
GC_1_218 b_1 NI_1 NS_218 0 -2.6512655682270976e-05
GC_1_219 b_1 NI_1 NS_219 0 -6.9061028904578899e-06
GC_1_220 b_1 NI_1 NS_220 0 9.9048500586287887e-06
GC_1_221 b_1 NI_1 NS_221 0 -9.5811569449001355e-06
GC_1_222 b_1 NI_1 NS_222 0 -4.8954932939036001e-05
GC_1_223 b_1 NI_1 NS_223 0 -1.0044599841741471e-05
GC_1_224 b_1 NI_1 NS_224 0 7.9771044770541569e-05
GC_1_225 b_1 NI_1 NS_225 0 3.9255922856516287e-02
GC_1_226 b_1 NI_1 NS_226 0 8.4906406420230860e-05
GC_1_227 b_1 NI_1 NS_227 0 5.3213037231660395e-03
GC_1_228 b_1 NI_1 NS_228 0 7.7864468082188825e-05
GC_1_229 b_1 NI_1 NS_229 0 -3.9292101639273758e-03
GC_1_230 b_1 NI_1 NS_230 0 3.0866355596600348e-03
GC_1_231 b_1 NI_1 NS_231 0 -1.7463966475125313e-03
GC_1_232 b_1 NI_1 NS_232 0 7.6522113254450528e-03
GC_1_233 b_1 NI_1 NS_233 0 -9.4884937240900247e-03
GC_1_234 b_1 NI_1 NS_234 0 -5.9785944858842168e-03
GC_1_235 b_1 NI_1 NS_235 0 -2.6382611877958777e-04
GC_1_236 b_1 NI_1 NS_236 0 -1.1882059360638273e-04
GC_1_237 b_1 NI_1 NS_237 0 7.6099315043868469e-03
GC_1_238 b_1 NI_1 NS_238 0 2.6309735783637111e-04
GC_1_239 b_1 NI_1 NS_239 0 7.0235856596889592e-05
GC_1_240 b_1 NI_1 NS_240 0 2.2030319256351959e-03
GC_1_241 b_1 NI_1 NS_241 0 -1.1519151613035392e-03
GC_1_242 b_1 NI_1 NS_242 0 1.6540954058413577e-03
GC_1_243 b_1 NI_1 NS_243 0 1.1223345824186053e-03
GC_1_244 b_1 NI_1 NS_244 0 5.4039141022992456e-03
GC_1_245 b_1 NI_1 NS_245 0 2.9250243053735900e-04
GC_1_246 b_1 NI_1 NS_246 0 9.8879282896959615e-05
GC_1_247 b_1 NI_1 NS_247 0 -9.7263860482745407e-03
GC_1_248 b_1 NI_1 NS_248 0 4.0457099531822482e-03
GC_1_249 b_1 NI_1 NS_249 0 1.1626125657069914e-03
GC_1_250 b_1 NI_1 NS_250 0 3.4034004408314042e-04
GC_1_251 b_1 NI_1 NS_251 0 -3.7366477906806495e-04
GC_1_252 b_1 NI_1 NS_252 0 6.2673808995336691e-05
GC_1_253 b_1 NI_1 NS_253 0 -1.9765313112296226e-04
GC_1_254 b_1 NI_1 NS_254 0 2.5834166597390784e-04
GC_1_255 b_1 NI_1 NS_255 0 -8.3960394057373065e-05
GC_1_256 b_1 NI_1 NS_256 0 7.4307383211529304e-06
GC_1_257 b_1 NI_1 NS_257 0 -8.7301582356035402e-03
GC_1_258 b_1 NI_1 NS_258 0 -9.8459004977780578e-03
GC_1_259 b_1 NI_1 NS_259 0 1.0100869528502163e-04
GC_1_260 b_1 NI_1 NS_260 0 -5.6669580292447506e-05
GC_1_261 b_1 NI_1 NS_261 0 -4.8209041000271078e-04
GC_1_262 b_1 NI_1 NS_262 0 2.3272483731544579e-03
GC_1_263 b_1 NI_1 NS_263 0 5.9199581256005095e-03
GC_1_264 b_1 NI_1 NS_264 0 -1.5671446125292715e-04
GC_1_265 b_1 NI_1 NS_265 0 4.4812749839564879e-04
GC_1_266 b_1 NI_1 NS_266 0 4.0248478939157337e-04
GC_1_267 b_1 NI_1 NS_267 0 2.5527359346412804e-06
GC_1_268 b_1 NI_1 NS_268 0 3.5557784946817286e-06
GC_1_269 b_1 NI_1 NS_269 0 5.6281754698261320e-06
GC_1_270 b_1 NI_1 NS_270 0 -1.6198824868779577e-05
GC_1_271 b_1 NI_1 NS_271 0 -3.1726559552725046e-04
GC_1_272 b_1 NI_1 NS_272 0 -1.2513953714946598e-05
GC_1_273 b_1 NI_1 NS_273 0 1.9844323073033128e-05
GC_1_274 b_1 NI_1 NS_274 0 -2.8636864359067070e-05
GC_1_275 b_1 NI_1 NS_275 0 -1.7002672156315179e-05
GC_1_276 b_1 NI_1 NS_276 0 1.0656877357609322e-07
GC_1_277 b_1 NI_1 NS_277 0 5.0687603539298289e-05
GC_1_278 b_1 NI_1 NS_278 0 -3.5673429346591790e-05
GC_1_279 b_1 NI_1 NS_279 0 -8.7190713155247350e-05
GC_1_280 b_1 NI_1 NS_280 0 2.8753954698110163e-05
GC_1_281 b_1 NI_1 NS_281 0 -6.3897974355345598e-03
GC_1_282 b_1 NI_1 NS_282 0 -2.5326893473840860e-04
GC_1_283 b_1 NI_1 NS_283 0 -1.3426740229843860e-03
GC_1_284 b_1 NI_1 NS_284 0 3.0615288795078103e-03
GC_1_285 b_1 NI_1 NS_285 0 -9.8183977847618909e-04
GC_1_286 b_1 NI_1 NS_286 0 -2.2450650996151855e-03
GC_1_287 b_1 NI_1 NS_287 0 -5.0728768600041109e-03
GC_1_288 b_1 NI_1 NS_288 0 -5.7632622973394091e-03
GC_1_289 b_1 NI_1 NS_289 0 7.2881496558373244e-03
GC_1_290 b_1 NI_1 NS_290 0 -1.4230082272091206e-03
GC_1_291 b_1 NI_1 NS_291 0 -3.1156989322422764e-04
GC_1_292 b_1 NI_1 NS_292 0 4.3384388254961986e-04
GC_1_293 b_1 NI_1 NS_293 0 4.2215432821092243e-03
GC_1_294 b_1 NI_1 NS_294 0 -2.5833428306949349e-03
GC_1_295 b_1 NI_1 NS_295 0 8.0837411603041796e-04
GC_1_296 b_1 NI_1 NS_296 0 1.1386264035180395e-03
GC_1_297 b_1 NI_1 NS_297 0 4.4334332003021545e-04
GC_1_298 b_1 NI_1 NS_298 0 2.1270323315511286e-03
GC_1_299 b_1 NI_1 NS_299 0 -3.1835499923509639e-03
GC_1_300 b_1 NI_1 NS_300 0 1.1322991748356709e-03
GC_1_301 b_1 NI_1 NS_301 0 -2.3049875329692973e-04
GC_1_302 b_1 NI_1 NS_302 0 3.3301933494902477e-05
GC_1_303 b_1 NI_1 NS_303 0 3.3068057230815121e-03
GC_1_304 b_1 NI_1 NS_304 0 -8.6570998081859874e-04
GC_1_305 b_1 NI_1 NS_305 0 -1.1627426536231730e-03
GC_1_306 b_1 NI_1 NS_306 0 -8.8280599746789858e-05
GC_1_307 b_1 NI_1 NS_307 0 -1.5568734989219082e-04
GC_1_308 b_1 NI_1 NS_308 0 8.3490840879539137e-05
GC_1_309 b_1 NI_1 NS_309 0 -3.1787777221401538e-04
GC_1_310 b_1 NI_1 NS_310 0 2.4792683837209574e-04
GC_1_311 b_1 NI_1 NS_311 0 -2.0513994572314751e-04
GC_1_312 b_1 NI_1 NS_312 0 -1.0639250177408491e-04
GC_1_313 b_1 NI_1 NS_313 0 2.5969343421787749e-03
GC_1_314 b_1 NI_1 NS_314 0 1.2344002523850316e-03
GC_1_315 b_1 NI_1 NS_315 0 -6.1292942481213213e-05
GC_1_316 b_1 NI_1 NS_316 0 1.4455674590555979e-04
GC_1_317 b_1 NI_1 NS_317 0 -3.7073854381347750e-04
GC_1_318 b_1 NI_1 NS_318 0 -1.0402169006624505e-03
GC_1_319 b_1 NI_1 NS_319 0 -7.5674654860369154e-04
GC_1_320 b_1 NI_1 NS_320 0 1.0343240174498982e-03
GC_1_321 b_1 NI_1 NS_321 0 -7.8345589657751394e-07
GC_1_322 b_1 NI_1 NS_322 0 -2.2586606462684895e-04
GC_1_323 b_1 NI_1 NS_323 0 2.1316300591053416e-06
GC_1_324 b_1 NI_1 NS_324 0 1.1252689307369839e-06
GC_1_325 b_1 NI_1 NS_325 0 2.5045368743114579e-06
GC_1_326 b_1 NI_1 NS_326 0 1.6565171746220648e-06
GC_1_327 b_1 NI_1 NS_327 0 1.1025839531434864e-04
GC_1_328 b_1 NI_1 NS_328 0 -2.9691556780927628e-05
GC_1_329 b_1 NI_1 NS_329 0 -4.9179546928213117e-06
GC_1_330 b_1 NI_1 NS_330 0 1.9215066764747525e-06
GC_1_331 b_1 NI_1 NS_331 0 1.1896375179735491e-05
GC_1_332 b_1 NI_1 NS_332 0 -1.0032959266326280e-06
GC_1_333 b_1 NI_1 NS_333 0 -2.2105309166184037e-05
GC_1_334 b_1 NI_1 NS_334 0 1.6304046014983336e-05
GC_1_335 b_1 NI_1 NS_335 0 3.8049426923099907e-05
GC_1_336 b_1 NI_1 NS_336 0 -6.5227122792403257e-06
GC_1_337 b_1 NI_1 NS_337 0 8.7304398110492842e-02
GC_1_338 b_1 NI_1 NS_338 0 -6.0122120130227865e-04
GC_1_339 b_1 NI_1 NS_339 0 4.0530896420456920e-03
GC_1_340 b_1 NI_1 NS_340 0 -1.5490071474400134e-03
GC_1_341 b_1 NI_1 NS_341 0 7.8453436217614469e-05
GC_1_342 b_1 NI_1 NS_342 0 5.5038400272815263e-03
GC_1_343 b_1 NI_1 NS_343 0 -1.2061496917228133e-03
GC_1_344 b_1 NI_1 NS_344 0 1.1589545008597293e-02
GC_1_345 b_1 NI_1 NS_345 0 -1.5625989539401065e-02
GC_1_346 b_1 NI_1 NS_346 0 5.5669629573620524e-03
GC_1_347 b_1 NI_1 NS_347 0 1.0316180314248067e-04
GC_1_348 b_1 NI_1 NS_348 0 6.3074953734998596e-05
GC_1_349 b_1 NI_1 NS_349 0 2.9428163021857820e-03
GC_1_350 b_1 NI_1 NS_350 0 6.1115288388415262e-04
GC_1_351 b_1 NI_1 NS_351 0 2.5123131252883661e-04
GC_1_352 b_1 NI_1 NS_352 0 2.0083417416859963e-03
GC_1_353 b_1 NI_1 NS_353 0 -6.7042076153042999e-03
GC_1_354 b_1 NI_1 NS_354 0 6.5997323108380737e-03
GC_1_355 b_1 NI_1 NS_355 0 -1.7608760307409390e-04
GC_1_356 b_1 NI_1 NS_356 0 6.1387843672537426e-03
GC_1_357 b_1 NI_1 NS_357 0 3.5322564792497450e-04
GC_1_358 b_1 NI_1 NS_358 0 8.5689308268302878e-05
GC_1_359 b_1 NI_1 NS_359 0 -1.9433940848696703e-02
GC_1_360 b_1 NI_1 NS_360 0 9.2620152803144645e-04
GC_1_361 b_1 NI_1 NS_361 0 1.2635821915315934e-03
GC_1_362 b_1 NI_1 NS_362 0 5.8042423561586109e-04
GC_1_363 b_1 NI_1 NS_363 0 -5.2180237914985325e-04
GC_1_364 b_1 NI_1 NS_364 0 -2.3816938882803467e-04
GC_1_365 b_1 NI_1 NS_365 0 -4.6673986766808124e-04
GC_1_366 b_1 NI_1 NS_366 0 2.2032709024474189e-04
GC_1_367 b_1 NI_1 NS_367 0 -1.9651045295069811e-04
GC_1_368 b_1 NI_1 NS_368 0 -7.9602561658700307e-06
GC_1_369 b_1 NI_1 NS_369 0 -7.8911477551059338e-03
GC_1_370 b_1 NI_1 NS_370 0 -1.4291063158346601e-02
GC_1_371 b_1 NI_1 NS_371 0 2.0902396211504187e-04
GC_1_372 b_1 NI_1 NS_372 0 -3.7711964779354848e-05
GC_1_373 b_1 NI_1 NS_373 0 -2.1997658538194919e-03
GC_1_374 b_1 NI_1 NS_374 0 2.7833234031235023e-03
GC_1_375 b_1 NI_1 NS_375 0 8.0639162651205184e-03
GC_1_376 b_1 NI_1 NS_376 0 -2.7509416758558403e-03
GC_1_377 b_1 NI_1 NS_377 0 -2.3262065734145818e-04
GC_1_378 b_1 NI_1 NS_378 0 4.2506571793018207e-04
GC_1_379 b_1 NI_1 NS_379 0 1.2389195699655526e-06
GC_1_380 b_1 NI_1 NS_380 0 5.6803064886259305e-06
GC_1_381 b_1 NI_1 NS_381 0 2.0723810303456439e-06
GC_1_382 b_1 NI_1 NS_382 0 -2.5087260721122597e-05
GC_1_383 b_1 NI_1 NS_383 0 -5.1687721697917140e-04
GC_1_384 b_1 NI_1 NS_384 0 1.0480751537484485e-04
GC_1_385 b_1 NI_1 NS_385 0 2.2190710886306289e-05
GC_1_386 b_1 NI_1 NS_386 0 -4.9175704823591366e-05
GC_1_387 b_1 NI_1 NS_387 0 -3.0195695432570882e-05
GC_1_388 b_1 NI_1 NS_388 0 -1.3421877435301727e-05
GC_1_389 b_1 NI_1 NS_389 0 1.1106904931523290e-04
GC_1_390 b_1 NI_1 NS_390 0 -5.2454594377982342e-05
GC_1_391 b_1 NI_1 NS_391 0 -1.8572327369162139e-04
GC_1_392 b_1 NI_1 NS_392 0 2.4900950676945171e-05
GC_1_393 b_1 NI_1 NS_393 0 -3.7701362339135576e-02
GC_1_394 b_1 NI_1 NS_394 0 -9.0949517691750158e-05
GC_1_395 b_1 NI_1 NS_395 0 -3.4758651154029091e-04
GC_1_396 b_1 NI_1 NS_396 0 2.3768057867345556e-03
GC_1_397 b_1 NI_1 NS_397 0 -2.4923580644026617e-03
GC_1_398 b_1 NI_1 NS_398 0 -1.4025237067787841e-03
GC_1_399 b_1 NI_1 NS_399 0 -5.5894393074071326e-03
GC_1_400 b_1 NI_1 NS_400 0 -6.1963786255559749e-03
GC_1_401 b_1 NI_1 NS_401 0 7.9811227553670001e-03
GC_1_402 b_1 NI_1 NS_402 0 -9.6907931229293122e-03
GC_1_403 b_1 NI_1 NS_403 0 3.0169147990353549e-05
GC_1_404 b_1 NI_1 NS_404 0 5.5634538323816101e-04
GC_1_405 b_1 NI_1 NS_405 0 5.1817747285674374e-03
GC_1_406 b_1 NI_1 NS_406 0 -2.0646373902267917e-03
GC_1_407 b_1 NI_1 NS_407 0 4.0474550878669542e-04
GC_1_408 b_1 NI_1 NS_408 0 4.6321923703218426e-04
GC_1_409 b_1 NI_1 NS_409 0 8.7973404643494992e-04
GC_1_410 b_1 NI_1 NS_410 0 2.1873013167585170e-03
GC_1_411 b_1 NI_1 NS_411 0 -1.4206434910884479e-06
GC_1_412 b_1 NI_1 NS_412 0 7.6879833359357494e-05
GC_1_413 b_1 NI_1 NS_413 0 -1.5187627701659066e-04
GC_1_414 b_1 NI_1 NS_414 0 1.0322612231403160e-04
GC_1_415 b_1 NI_1 NS_415 0 6.5162768212804188e-04
GC_1_416 b_1 NI_1 NS_416 0 -4.1065977893970061e-03
GC_1_417 b_1 NI_1 NS_417 0 -8.1744060234876061e-04
GC_1_418 b_1 NI_1 NS_418 0 2.7486033360018522e-04
GC_1_419 b_1 NI_1 NS_419 0 -2.9096148470410479e-06
GC_1_420 b_1 NI_1 NS_420 0 -3.0287635173618993e-05
GC_1_421 b_1 NI_1 NS_421 0 -2.2523373499288614e-04
GC_1_422 b_1 NI_1 NS_422 0 -8.7724037907094919e-05
GC_1_423 b_1 NI_1 NS_423 0 -7.0284200181686704e-05
GC_1_424 b_1 NI_1 NS_424 0 -1.4317018525551164e-04
GC_1_425 b_1 NI_1 NS_425 0 9.2805573396012742e-03
GC_1_426 b_1 NI_1 NS_426 0 8.0023686719510876e-04
GC_1_427 b_1 NI_1 NS_427 0 -5.9514575065446854e-05
GC_1_428 b_1 NI_1 NS_428 0 1.3298812055328061e-04
GC_1_429 b_1 NI_1 NS_429 0 -5.7895331746160735e-04
GC_1_430 b_1 NI_1 NS_430 0 -1.7065018604399294e-03
GC_1_431 b_1 NI_1 NS_431 0 -5.2353237639927823e-04
GC_1_432 b_1 NI_1 NS_432 0 2.3359122362130945e-03
GC_1_433 b_1 NI_1 NS_433 0 -4.6952452662668391e-04
GC_1_434 b_1 NI_1 NS_434 0 -2.9728910195318353e-04
GC_1_435 b_1 NI_1 NS_435 0 -1.2103062000064702e-07
GC_1_436 b_1 NI_1 NS_436 0 -1.3562405209712993e-06
GC_1_437 b_1 NI_1 NS_437 0 5.3033514290186201e-06
GC_1_438 b_1 NI_1 NS_438 0 1.3704186934937423e-05
GC_1_439 b_1 NI_1 NS_439 0 1.6474620008059029e-04
GC_1_440 b_1 NI_1 NS_440 0 -1.4824621166139305e-04
GC_1_441 b_1 NI_1 NS_441 0 -4.9275000607265716e-08
GC_1_442 b_1 NI_1 NS_442 0 2.5780093194336360e-05
GC_1_443 b_1 NI_1 NS_443 0 1.3619426543817380e-05
GC_1_444 b_1 NI_1 NS_444 0 -7.5222429833219099e-07
GC_1_445 b_1 NI_1 NS_445 0 -3.5922423279688798e-05
GC_1_446 b_1 NI_1 NS_446 0 3.8364746744661563e-05
GC_1_447 b_1 NI_1 NS_447 0 6.8212066014166224e-05
GC_1_448 b_1 NI_1 NS_448 0 -3.3336323581733796e-05
GC_1_449 b_1 NI_1 NS_449 0 4.6820193732603418e-03
GC_1_450 b_1 NI_1 NS_450 0 1.3455451164585714e-04
GC_1_451 b_1 NI_1 NS_451 0 -1.7937763128380327e-04
GC_1_452 b_1 NI_1 NS_452 0 -1.8179982547129929e-04
GC_1_453 b_1 NI_1 NS_453 0 1.1938773449165252e-04
GC_1_454 b_1 NI_1 NS_454 0 -2.8494641304722485e-04
GC_1_455 b_1 NI_1 NS_455 0 1.1086842889311116e-03
GC_1_456 b_1 NI_1 NS_456 0 -7.6331996237435939e-04
GC_1_457 b_1 NI_1 NS_457 0 1.6985078722210026e-03
GC_1_458 b_1 NI_1 NS_458 0 5.0716159345712427e-04
GC_1_459 b_1 NI_1 NS_459 0 -3.8893313591423283e-04
GC_1_460 b_1 NI_1 NS_460 0 2.1793810144347183e-04
GC_1_461 b_1 NI_1 NS_461 0 1.3070139610563624e-03
GC_1_462 b_1 NI_1 NS_462 0 -6.5820893135344020e-04
GC_1_463 b_1 NI_1 NS_463 0 1.2840784158055494e-03
GC_1_464 b_1 NI_1 NS_464 0 -5.6987637296701734e-05
GC_1_465 b_1 NI_1 NS_465 0 1.1039119511435033e-03
GC_1_466 b_1 NI_1 NS_466 0 2.3356345754324704e-03
GC_1_467 b_1 NI_1 NS_467 0 1.4822839493100256e-03
GC_1_468 b_1 NI_1 NS_468 0 8.8246726381578254e-05
GC_1_469 b_1 NI_1 NS_469 0 4.2063044098903274e-04
GC_1_470 b_1 NI_1 NS_470 0 1.9173293128911900e-04
GC_1_471 b_1 NI_1 NS_471 0 -1.2679167005962027e-04
GC_1_472 b_1 NI_1 NS_472 0 9.1803020593375587e-03
GC_1_473 b_1 NI_1 NS_473 0 -7.3660576921313903e-04
GC_1_474 b_1 NI_1 NS_474 0 -7.3117782619602485e-04
GC_1_475 b_1 NI_1 NS_475 0 -9.6407865161853414e-04
GC_1_476 b_1 NI_1 NS_476 0 -9.3676360296166046e-05
GC_1_477 b_1 NI_1 NS_477 0 -4.0627976559117683e-04
GC_1_478 b_1 NI_1 NS_478 0 -4.1332466723800943e-04
GC_1_479 b_1 NI_1 NS_479 0 -8.3705885274521074e-05
GC_1_480 b_1 NI_1 NS_480 0 -3.0450248692062368e-06
GC_1_481 b_1 NI_1 NS_481 0 -5.0694599385178920e-03
GC_1_482 b_1 NI_1 NS_482 0 -1.3984832079484862e-03
GC_1_483 b_1 NI_1 NS_483 0 1.2594835053276655e-05
GC_1_484 b_1 NI_1 NS_484 0 -2.2330847103727287e-05
GC_1_485 b_1 NI_1 NS_485 0 2.6398337700645897e-05
GC_1_486 b_1 NI_1 NS_486 0 2.9797190786171604e-04
GC_1_487 b_1 NI_1 NS_487 0 1.3575794346346558e-03
GC_1_488 b_1 NI_1 NS_488 0 -2.1416889199484504e-03
GC_1_489 b_1 NI_1 NS_489 0 6.4852876906359343e-05
GC_1_490 b_1 NI_1 NS_490 0 1.4315027374490149e-04
GC_1_491 b_1 NI_1 NS_491 0 -1.9190585949319157e-06
GC_1_492 b_1 NI_1 NS_492 0 1.8204297699116964e-06
GC_1_493 b_1 NI_1 NS_493 0 -1.3029505583220473e-06
GC_1_494 b_1 NI_1 NS_494 0 -7.5787941747992455e-06
GC_1_495 b_1 NI_1 NS_495 0 -1.1522831343387060e-04
GC_1_496 b_1 NI_1 NS_496 0 8.3892111363134876e-05
GC_1_497 b_1 NI_1 NS_497 0 2.6508552590208090e-06
GC_1_498 b_1 NI_1 NS_498 0 -1.7725512114219494e-05
GC_1_499 b_1 NI_1 NS_499 0 -1.1609215501703752e-05
GC_1_500 b_1 NI_1 NS_500 0 -1.4127494152241257e-05
GC_1_501 b_1 NI_1 NS_501 0 5.3961300645233244e-05
GC_1_502 b_1 NI_1 NS_502 0 -2.0720651495049425e-05
GC_1_503 b_1 NI_1 NS_503 0 -9.3365193213947972e-05
GC_1_504 b_1 NI_1 NS_504 0 5.0058813617999195e-06
GC_1_505 b_1 NI_1 NS_505 0 5.5660533841558543e-03
GC_1_506 b_1 NI_1 NS_506 0 -1.0145321138746868e-04
GC_1_507 b_1 NI_1 NS_507 0 1.9992950229116697e-04
GC_1_508 b_1 NI_1 NS_508 0 1.6140516246580022e-05
GC_1_509 b_1 NI_1 NS_509 0 1.0372911734717554e-04
GC_1_510 b_1 NI_1 NS_510 0 2.4325577023126175e-04
GC_1_511 b_1 NI_1 NS_511 0 -3.1611090393726524e-04
GC_1_512 b_1 NI_1 NS_512 0 1.2476672671577979e-03
GC_1_513 b_1 NI_1 NS_513 0 -1.7128848404918901e-03
GC_1_514 b_1 NI_1 NS_514 0 5.6251575511968150e-04
GC_1_515 b_1 NI_1 NS_515 0 3.8290556158616592e-04
GC_1_516 b_1 NI_1 NS_516 0 -9.3814592350528682e-04
GC_1_517 b_1 NI_1 NS_517 0 -5.3111055563097352e-04
GC_1_518 b_1 NI_1 NS_518 0 -1.0183091500536913e-03
GC_1_519 b_1 NI_1 NS_519 0 5.9511083819859651e-04
GC_1_520 b_1 NI_1 NS_520 0 -3.8076081417931339e-04
GC_1_521 b_1 NI_1 NS_521 0 1.3702353233698930e-03
GC_1_522 b_1 NI_1 NS_522 0 1.0770191555477609e-03
GC_1_523 b_1 NI_1 NS_523 0 -7.6306369664594191e-04
GC_1_524 b_1 NI_1 NS_524 0 2.2130015074534946e-03
GC_1_525 b_1 NI_1 NS_525 0 -2.1002614300633763e-04
GC_1_526 b_1 NI_1 NS_526 0 -2.7445049667742039e-06
GC_1_527 b_1 NI_1 NS_527 0 -2.8947164745072042e-03
GC_1_528 b_1 NI_1 NS_528 0 1.8290981455397367e-03
GC_1_529 b_1 NI_1 NS_529 0 3.4458234987817864e-04
GC_1_530 b_1 NI_1 NS_530 0 3.5811355743281222e-04
GC_1_531 b_1 NI_1 NS_531 0 -8.0098250863461142e-04
GC_1_532 b_1 NI_1 NS_532 0 8.1147455517494588e-05
GC_1_533 b_1 NI_1 NS_533 0 -5.4047661649014888e-04
GC_1_534 b_1 NI_1 NS_534 0 -1.0269537315843089e-04
GC_1_535 b_1 NI_1 NS_535 0 -8.9800300916849761e-05
GC_1_536 b_1 NI_1 NS_536 0 -5.5939958532596070e-05
GC_1_537 b_1 NI_1 NS_537 0 -1.2217264408033964e-03
GC_1_538 b_1 NI_1 NS_538 0 -5.7137305867577459e-03
GC_1_539 b_1 NI_1 NS_539 0 5.1376449979148510e-05
GC_1_540 b_1 NI_1 NS_540 0 -2.2848655436121097e-05
GC_1_541 b_1 NI_1 NS_541 0 -1.1269313238573633e-03
GC_1_542 b_1 NI_1 NS_542 0 4.1506642030035237e-04
GC_1_543 b_1 NI_1 NS_543 0 2.1247866607420379e-03
GC_1_544 b_1 NI_1 NS_544 0 4.3545860347383411e-04
GC_1_545 b_1 NI_1 NS_545 0 -8.8815121691124865e-05
GC_1_546 b_1 NI_1 NS_546 0 1.6625290195650504e-04
GC_1_547 b_1 NI_1 NS_547 0 -1.0222119359328299e-06
GC_1_548 b_1 NI_1 NS_548 0 1.2395205605004254e-06
GC_1_549 b_1 NI_1 NS_549 0 5.6207858849345201e-06
GC_1_550 b_1 NI_1 NS_550 0 -1.9364294416793295e-06
GC_1_551 b_1 NI_1 NS_551 0 -1.3162829318790983e-04
GC_1_552 b_1 NI_1 NS_552 0 -7.4360257118673005e-05
GC_1_553 b_1 NI_1 NS_553 0 1.7462363966848644e-05
GC_1_554 b_1 NI_1 NS_554 0 -2.1723022339221642e-06
GC_1_555 b_1 NI_1 NS_555 0 -6.0489143191667170e-06
GC_1_556 b_1 NI_1 NS_556 0 -1.1046712097852097e-05
GC_1_557 b_1 NI_1 NS_557 0 4.1274347070368523e-05
GC_1_558 b_1 NI_1 NS_558 0 4.4225436589773846e-05
GC_1_559 b_1 NI_1 NS_559 0 -4.3629130832430513e-05
GC_1_560 b_1 NI_1 NS_560 0 -7.7747881122318269e-05
GC_1_561 b_1 NI_1 NS_561 0 3.2345193180308866e-02
GC_1_562 b_1 NI_1 NS_562 0 -2.1059964198199675e-05
GC_1_563 b_1 NI_1 NS_563 0 2.3040074279731865e-04
GC_1_564 b_1 NI_1 NS_564 0 -5.6559446719547522e-04
GC_1_565 b_1 NI_1 NS_565 0 7.6516420633372868e-04
GC_1_566 b_1 NI_1 NS_566 0 3.5584541722963304e-04
GC_1_567 b_1 NI_1 NS_567 0 1.8691430500484981e-03
GC_1_568 b_1 NI_1 NS_568 0 1.9497909510207770e-03
GC_1_569 b_1 NI_1 NS_569 0 -3.8033075040036312e-04
GC_1_570 b_1 NI_1 NS_570 0 4.2106693176441725e-03
GC_1_571 b_1 NI_1 NS_571 0 -2.3257555751737388e-04
GC_1_572 b_1 NI_1 NS_572 0 5.7504164784109727e-04
GC_1_573 b_1 NI_1 NS_573 0 1.0508309566411684e-03
GC_1_574 b_1 NI_1 NS_574 0 5.8664605060386541e-04
GC_1_575 b_1 NI_1 NS_575 0 1.0300021625476348e-03
GC_1_576 b_1 NI_1 NS_576 0 2.8732096166688093e-04
GC_1_577 b_1 NI_1 NS_577 0 3.6921704063288710e-05
GC_1_578 b_1 NI_1 NS_578 0 5.3304317228772399e-03
GC_1_579 b_1 NI_1 NS_579 0 1.0929009073900302e-03
GC_1_580 b_1 NI_1 NS_580 0 1.9270998397397155e-03
GC_1_581 b_1 NI_1 NS_581 0 3.3144581941211464e-04
GC_1_582 b_1 NI_1 NS_582 0 1.5942086079007609e-04
GC_1_583 b_1 NI_1 NS_583 0 -6.7849043611652405e-03
GC_1_584 b_1 NI_1 NS_584 0 8.9135615988947276e-03
GC_1_585 b_1 NI_1 NS_585 0 -1.5271809998202091e-04
GC_1_586 b_1 NI_1 NS_586 0 -2.6374402912206479e-04
GC_1_587 b_1 NI_1 NS_587 0 -7.3644263703290420e-04
GC_1_588 b_1 NI_1 NS_588 0 -9.9349715198550150e-05
GC_1_589 b_1 NI_1 NS_589 0 -3.7092847757952153e-04
GC_1_590 b_1 NI_1 NS_590 0 -1.4108233965267212e-04
GC_1_591 b_1 NI_1 NS_591 0 -1.1156669776775876e-04
GC_1_592 b_1 NI_1 NS_592 0 2.2538329030908995e-05
GC_1_593 b_1 NI_1 NS_593 0 -8.3646600483860273e-03
GC_1_594 b_1 NI_1 NS_594 0 -4.3034895441377901e-03
GC_1_595 b_1 NI_1 NS_595 0 5.9660640416596389e-05
GC_1_596 b_1 NI_1 NS_596 0 -6.2654333391271797e-05
GC_1_597 b_1 NI_1 NS_597 0 -2.5759488961755192e-04
GC_1_598 b_1 NI_1 NS_598 0 1.5037226128031709e-03
GC_1_599 b_1 NI_1 NS_599 0 3.0373757556187804e-03
GC_1_600 b_1 NI_1 NS_600 0 -4.5808894921764093e-03
GC_1_601 b_1 NI_1 NS_601 0 7.2403686094357452e-05
GC_1_602 b_1 NI_1 NS_602 0 3.4665172275284993e-04
GC_1_603 b_1 NI_1 NS_603 0 1.4136709581725163e-06
GC_1_604 b_1 NI_1 NS_604 0 3.8101517481046541e-06
GC_1_605 b_1 NI_1 NS_605 0 -5.1045094275053428e-06
GC_1_606 b_1 NI_1 NS_606 0 -1.9812760349810145e-05
GC_1_607 b_1 NI_1 NS_607 0 -3.0450303987782497e-04
GC_1_608 b_1 NI_1 NS_608 0 2.7827138924364027e-04
GC_1_609 b_1 NI_1 NS_609 0 1.3734273722926002e-06
GC_1_610 b_1 NI_1 NS_610 0 -4.7309306613019768e-05
GC_1_611 b_1 NI_1 NS_611 0 -3.4617224131402949e-05
GC_1_612 b_1 NI_1 NS_612 0 -7.0181506825475590e-06
GC_1_613 b_1 NI_1 NS_613 0 9.6426075407993395e-05
GC_1_614 b_1 NI_1 NS_614 0 -9.7333428518469852e-05
GC_1_615 b_1 NI_1 NS_615 0 -1.8916155324037959e-04
GC_1_616 b_1 NI_1 NS_616 0 9.9144720726442311e-05
GC_1_617 b_1 NI_1 NS_617 0 -7.7620210888951482e-03
GC_1_618 b_1 NI_1 NS_618 0 -9.4331735254380155e-05
GC_1_619 b_1 NI_1 NS_619 0 2.4035115825599392e-04
GC_1_620 b_1 NI_1 NS_620 0 2.9997188130974188e-04
GC_1_621 b_1 NI_1 NS_621 0 -3.6393067352241828e-04
GC_1_622 b_1 NI_1 NS_622 0 2.9345792259034603e-04
GC_1_623 b_1 NI_1 NS_623 0 -1.7710689390551702e-03
GC_1_624 b_1 NI_1 NS_624 0 2.2436576938405755e-04
GC_1_625 b_1 NI_1 NS_625 0 -1.2042529903520790e-03
GC_1_626 b_1 NI_1 NS_626 0 -2.5335848451696810e-03
GC_1_627 b_1 NI_1 NS_627 0 6.1732082219518561e-04
GC_1_628 b_1 NI_1 NS_628 0 -4.9215614304204652e-04
GC_1_629 b_1 NI_1 NS_629 0 7.0860718599525586e-04
GC_1_630 b_1 NI_1 NS_630 0 -1.6586984946251378e-03
GC_1_631 b_1 NI_1 NS_631 0 3.1036444299956388e-04
GC_1_632 b_1 NI_1 NS_632 0 -1.4334112915044531e-04
GC_1_633 b_1 NI_1 NS_633 0 1.2872285744243933e-03
GC_1_634 b_1 NI_1 NS_634 0 9.4271671193600485e-04
GC_1_635 b_1 NI_1 NS_635 0 -4.8374934929036324e-04
GC_1_636 b_1 NI_1 NS_636 0 7.3696491810889533e-04
GC_1_637 b_1 NI_1 NS_637 0 -8.7836481995061665e-05
GC_1_638 b_1 NI_1 NS_638 0 7.6888173462283179e-05
GC_1_639 b_1 NI_1 NS_639 0 -2.7511100083400719e-03
GC_1_640 b_1 NI_1 NS_640 0 -6.7960325354598659e-04
GC_1_641 b_1 NI_1 NS_641 0 -1.7801832522632991e-06
GC_1_642 b_1 NI_1 NS_642 0 5.7095899183584001e-04
GC_1_643 b_1 NI_1 NS_643 0 -3.9126304968047348e-04
GC_1_644 b_1 NI_1 NS_644 0 -7.5098841359436404e-05
GC_1_645 b_1 NI_1 NS_645 0 -3.6757492688339655e-04
GC_1_646 b_1 NI_1 NS_646 0 -1.4754985017814110e-04
GC_1_647 b_1 NI_1 NS_647 0 -6.3669568592445537e-05
GC_1_648 b_1 NI_1 NS_648 0 -9.7178864548417757e-05
GC_1_649 b_1 NI_1 NS_649 0 3.2029717163245749e-03
GC_1_650 b_1 NI_1 NS_650 0 -4.5270884572621885e-03
GC_1_651 b_1 NI_1 NS_651 0 2.0866877919822675e-05
GC_1_652 b_1 NI_1 NS_652 0 4.9503424064673713e-05
GC_1_653 b_1 NI_1 NS_653 0 -9.9415350544265432e-04
GC_1_654 b_1 NI_1 NS_654 0 -4.6610164850786304e-04
GC_1_655 b_1 NI_1 NS_655 0 1.0041225959387917e-03
GC_1_656 b_1 NI_1 NS_656 0 1.6132437760498187e-03
GC_1_657 b_1 NI_1 NS_657 0 -2.5067919362715388e-04
GC_1_658 b_1 NI_1 NS_658 0 1.2755644886112914e-05
GC_1_659 b_1 NI_1 NS_659 0 -1.5638223732629776e-06
GC_1_660 b_1 NI_1 NS_660 0 -1.1825436905847892e-06
GC_1_661 b_1 NI_1 NS_661 0 7.4144411416747233e-06
GC_1_662 b_1 NI_1 NS_662 0 7.1981130207087539e-06
GC_1_663 b_1 NI_1 NS_663 0 -7.1480713803349815e-05
GC_1_664 b_1 NI_1 NS_664 0 -1.6319146682746777e-04
GC_1_665 b_1 NI_1 NS_665 0 1.5574851173472834e-05
GC_1_666 b_1 NI_1 NS_666 0 1.7159357074963415e-05
GC_1_667 b_1 NI_1 NS_667 0 8.4181572052298210e-06
GC_1_668 b_1 NI_1 NS_668 0 -6.4349542198406466e-06
GC_1_669 b_1 NI_1 NS_669 0 5.2095429431655241e-06
GC_1_670 b_1 NI_1 NS_670 0 6.1062621703107065e-05
GC_1_671 b_1 NI_1 NS_671 0 2.0450563760568257e-05
GC_1_672 b_1 NI_1 NS_672 0 -8.8654192363125776e-05
GD_1_1 b_1 NI_1 NA_1 0 -1.1467324481976099e-01
GD_1_2 b_1 NI_1 NA_2 0 1.4108445671211355e-02
GD_1_3 b_1 NI_1 NA_3 0 -1.7791070396064364e-04
GD_1_4 b_1 NI_1 NA_4 0 -6.0404051628888143e-02
GD_1_5 b_1 NI_1 NA_5 0 -4.3599531985803915e-02
GD_1_6 b_1 NI_1 NA_6 0 2.3305025613108098e-03
GD_1_7 b_1 NI_1 NA_7 0 -8.1417525917378455e-02
GD_1_8 b_1 NI_1 NA_8 0 4.0846446920761524e-02
GD_1_9 b_1 NI_1 NA_9 0 -1.1601535750839389e-02
GD_1_10 b_1 NI_1 NA_10 0 1.7248625842619383e-03
GD_1_11 b_1 NI_1 NA_11 0 -4.0811928009420316e-02
GD_1_12 b_1 NI_1 NA_12 0 1.7846885875167594e-02
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 -1.5506986626876924e-02
GC_2_2 b_2 NI_2 NS_2 0 1.2182092646436993e-02
GC_2_3 b_2 NI_2 NS_3 0 -2.2350826156666993e-03
GC_2_4 b_2 NI_2 NS_4 0 1.2891383970957742e-03
GC_2_5 b_2 NI_2 NS_5 0 -2.0941791550015895e-03
GC_2_6 b_2 NI_2 NS_6 0 4.4904251475433232e-03
GC_2_7 b_2 NI_2 NS_7 0 -1.0314936662711568e-03
GC_2_8 b_2 NI_2 NS_8 0 -2.9828055445542483e-03
GC_2_9 b_2 NI_2 NS_9 0 -1.2456170311629797e-02
GC_2_10 b_2 NI_2 NS_10 0 -3.1962467646477386e-03
GC_2_11 b_2 NI_2 NS_11 0 3.4147725723090115e-04
GC_2_12 b_2 NI_2 NS_12 0 -1.9124658127345979e-04
GC_2_13 b_2 NI_2 NS_13 0 3.4168713016583807e-03
GC_2_14 b_2 NI_2 NS_14 0 -2.1288944255216881e-04
GC_2_15 b_2 NI_2 NS_15 0 7.7650908752560459e-04
GC_2_16 b_2 NI_2 NS_16 0 7.4827476423017431e-04
GC_2_17 b_2 NI_2 NS_17 0 4.5561429187667849e-03
GC_2_18 b_2 NI_2 NS_18 0 -1.8590671235842718e-03
GC_2_19 b_2 NI_2 NS_19 0 -8.8966181897166786e-04
GC_2_20 b_2 NI_2 NS_20 0 -2.9542410422332102e-04
GC_2_21 b_2 NI_2 NS_21 0 -1.3763886874765027e-04
GC_2_22 b_2 NI_2 NS_22 0 2.4470474732531521e-07
GC_2_23 b_2 NI_2 NS_23 0 6.1739101357029163e-03
GC_2_24 b_2 NI_2 NS_24 0 -2.1833436137610299e-04
GC_2_25 b_2 NI_2 NS_25 0 -8.0641780117117663e-04
GC_2_26 b_2 NI_2 NS_26 0 -1.6305320855984051e-04
GC_2_27 b_2 NI_2 NS_27 0 -9.2428603678830655e-05
GC_2_28 b_2 NI_2 NS_28 0 5.0339566512784207e-05
GC_2_29 b_2 NI_2 NS_29 0 -2.1532831514692278e-04
GC_2_30 b_2 NI_2 NS_30 0 2.0220368589879284e-04
GC_2_31 b_2 NI_2 NS_31 0 -1.5103864256724734e-04
GC_2_32 b_2 NI_2 NS_32 0 -6.2868059979280977e-05
GC_2_33 b_2 NI_2 NS_33 0 -1.0615296539215643e-03
GC_2_34 b_2 NI_2 NS_34 0 9.8325178790927632e-04
GC_2_35 b_2 NI_2 NS_35 0 -4.1832230681196145e-05
GC_2_36 b_2 NI_2 NS_36 0 7.8578848690061322e-05
GC_2_37 b_2 NI_2 NS_37 0 -9.0811809111266805e-05
GC_2_38 b_2 NI_2 NS_38 0 -2.4836285925684576e-04
GC_2_39 b_2 NI_2 NS_39 0 3.0488610919434608e-05
GC_2_40 b_2 NI_2 NS_40 0 -6.5365301004863122e-04
GC_2_41 b_2 NI_2 NS_41 0 1.6334965855556278e-04
GC_2_42 b_2 NI_2 NS_42 0 1.3708115485048356e-04
GC_2_43 b_2 NI_2 NS_43 0 9.6295166841737373e-07
GC_2_44 b_2 NI_2 NS_44 0 7.1860456718627772e-07
GC_2_45 b_2 NI_2 NS_45 0 1.4807160975786346e-06
GC_2_46 b_2 NI_2 NS_46 0 -6.0732255439109303e-06
GC_2_47 b_2 NI_2 NS_47 0 -1.0954991206421212e-04
GC_2_48 b_2 NI_2 NS_48 0 2.4349477768896020e-05
GC_2_49 b_2 NI_2 NS_49 0 4.0184396146151308e-06
GC_2_50 b_2 NI_2 NS_50 0 -1.3923577451941402e-05
GC_2_51 b_2 NI_2 NS_51 0 1.0945361948780334e-05
GC_2_52 b_2 NI_2 NS_52 0 -3.7775688070847639e-06
GC_2_53 b_2 NI_2 NS_53 0 1.3782754853263920e-05
GC_2_54 b_2 NI_2 NS_54 0 2.6818741354575585e-05
GC_2_55 b_2 NI_2 NS_55 0 -7.6320503897203902e-06
GC_2_56 b_2 NI_2 NS_56 0 -4.5971950534591146e-05
GC_2_57 b_2 NI_2 NS_57 0 -9.0977813245553624e-02
GC_2_58 b_2 NI_2 NS_58 0 8.1314517547627068e-03
GC_2_59 b_2 NI_2 NS_59 0 -1.5994169007266609e-04
GC_2_60 b_2 NI_2 NS_60 0 -1.1851109395686408e-03
GC_2_61 b_2 NI_2 NS_61 0 -1.3692608254135190e-03
GC_2_62 b_2 NI_2 NS_62 0 -1.3642040029422319e-03
GC_2_63 b_2 NI_2 NS_63 0 1.6058821495374086e-03
GC_2_64 b_2 NI_2 NS_64 0 2.4456583238871487e-03
GC_2_65 b_2 NI_2 NS_65 0 9.4553862145875210e-03
GC_2_66 b_2 NI_2 NS_66 0 -1.1367126023233917e-03
GC_2_67 b_2 NI_2 NS_67 0 6.5712916163003867e-04
GC_2_68 b_2 NI_2 NS_68 0 -5.4801842966670765e-04
GC_2_69 b_2 NI_2 NS_69 0 -6.8251419766470292e-04
GC_2_70 b_2 NI_2 NS_70 0 -2.2904482973653234e-03
GC_2_71 b_2 NI_2 NS_71 0 5.9704649637978054e-04
GC_2_72 b_2 NI_2 NS_72 0 2.7777466547850732e-04
GC_2_73 b_2 NI_2 NS_73 0 7.0977046804564204e-04
GC_2_74 b_2 NI_2 NS_74 0 -1.8893794997087245e-03
GC_2_75 b_2 NI_2 NS_75 0 1.5737233114593674e-03
GC_2_76 b_2 NI_2 NS_76 0 -1.6965529662778616e-03
GC_2_77 b_2 NI_2 NS_77 0 3.5511683716995895e-05
GC_2_78 b_2 NI_2 NS_78 0 -2.6394392994469139e-05
GC_2_79 b_2 NI_2 NS_79 0 4.0032651227775396e-03
GC_2_80 b_2 NI_2 NS_80 0 2.8618216001398463e-03
GC_2_81 b_2 NI_2 NS_81 0 1.3775868230604655e-04
GC_2_82 b_2 NI_2 NS_82 0 -3.6127767362863121e-05
GC_2_83 b_2 NI_2 NS_83 0 -8.8731015525357328e-05
GC_2_84 b_2 NI_2 NS_84 0 4.8754810031469012e-05
GC_2_85 b_2 NI_2 NS_85 0 2.0339937959234513e-04
GC_2_86 b_2 NI_2 NS_86 0 -1.6628215497694747e-04
GC_2_87 b_2 NI_2 NS_87 0 2.6901981226018073e-04
GC_2_88 b_2 NI_2 NS_88 0 -7.1228751471121037e-05
GC_2_89 b_2 NI_2 NS_89 0 -9.3289871053525084e-03
GC_2_90 b_2 NI_2 NS_90 0 2.3240041343204790e-03
GC_2_91 b_2 NI_2 NS_91 0 -1.7650775922122282e-04
GC_2_92 b_2 NI_2 NS_92 0 -2.1747545996984348e-04
GC_2_93 b_2 NI_2 NS_93 0 3.5331723932515045e-03
GC_2_94 b_2 NI_2 NS_94 0 9.3320660300466303e-04
GC_2_95 b_2 NI_2 NS_95 0 3.1730754228623662e-03
GC_2_96 b_2 NI_2 NS_96 0 -1.8928136572296311e-03
GC_2_97 b_2 NI_2 NS_97 0 1.0316556481403615e-03
GC_2_98 b_2 NI_2 NS_98 0 1.9373227006860559e-04
GC_2_99 b_2 NI_2 NS_99 0 -6.1201691732619915e-07
GC_2_100 b_2 NI_2 NS_100 0 -1.9794208940313557e-06
GC_2_101 b_2 NI_2 NS_101 0 -2.0861050559599726e-05
GC_2_102 b_2 NI_2 NS_102 0 -1.5907044021443898e-05
GC_2_103 b_2 NI_2 NS_103 0 -5.8024408835097597e-05
GC_2_104 b_2 NI_2 NS_104 0 -2.4340685859651988e-05
GC_2_105 b_2 NI_2 NS_105 0 -3.6170478464430640e-05
GC_2_106 b_2 NI_2 NS_106 0 -7.8784779394288881e-06
GC_2_107 b_2 NI_2 NS_107 0 -2.5448188140666252e-05
GC_2_108 b_2 NI_2 NS_108 0 -2.9247743852263230e-06
GC_2_109 b_2 NI_2 NS_109 0 1.6420100958241404e-04
GC_2_110 b_2 NI_2 NS_110 0 -1.3817454853235720e-04
GC_2_111 b_2 NI_2 NS_111 0 -2.8887190126695902e-04
GC_2_112 b_2 NI_2 NS_112 0 1.3634141561118428e-04
GC_2_113 b_2 NI_2 NS_113 0 5.8904813671195821e-02
GC_2_114 b_2 NI_2 NS_114 0 -7.7058472661237958e-04
GC_2_115 b_2 NI_2 NS_115 0 -1.8477663733946677e-03
GC_2_116 b_2 NI_2 NS_116 0 2.3852737836362933e-03
GC_2_117 b_2 NI_2 NS_117 0 2.9557673877871706e-03
GC_2_118 b_2 NI_2 NS_118 0 1.3870493842873898e-04
GC_2_119 b_2 NI_2 NS_119 0 -5.2073017576513680e-03
GC_2_120 b_2 NI_2 NS_120 0 3.6875906355964238e-04
GC_2_121 b_2 NI_2 NS_121 0 -5.9150297396432733e-03
GC_2_122 b_2 NI_2 NS_122 0 1.1177472469110553e-02
GC_2_123 b_2 NI_2 NS_123 0 -6.2312734181520116e-04
GC_2_124 b_2 NI_2 NS_124 0 -1.0715164626851945e-05
GC_2_125 b_2 NI_2 NS_125 0 1.5956146972998749e-03
GC_2_126 b_2 NI_2 NS_126 0 -3.9321062194472671e-03
GC_2_127 b_2 NI_2 NS_127 0 8.7691057710740305e-04
GC_2_128 b_2 NI_2 NS_128 0 1.5833254259818674e-03
GC_2_129 b_2 NI_2 NS_129 0 -8.9525702965536161e-04
GC_2_130 b_2 NI_2 NS_130 0 1.0681648792983714e-03
GC_2_131 b_2 NI_2 NS_131 0 -6.1601864062879423e-03
GC_2_132 b_2 NI_2 NS_132 0 4.4880520179613637e-04
GC_2_133 b_2 NI_2 NS_133 0 -7.6801113580174981e-05
GC_2_134 b_2 NI_2 NS_134 0 -9.6447244105362612e-05
GC_2_135 b_2 NI_2 NS_135 0 1.1955370131195252e-03
GC_2_136 b_2 NI_2 NS_136 0 4.8946183370804320e-03
GC_2_137 b_2 NI_2 NS_137 0 -5.2880103799279573e-04
GC_2_138 b_2 NI_2 NS_138 0 -3.1099948303371622e-04
GC_2_139 b_2 NI_2 NS_139 0 -3.3143186335694689e-04
GC_2_140 b_2 NI_2 NS_140 0 3.7071894161047354e-05
GC_2_141 b_2 NI_2 NS_141 0 -4.0297072770120192e-04
GC_2_142 b_2 NI_2 NS_142 0 4.5626748235621779e-04
GC_2_143 b_2 NI_2 NS_143 0 -2.7267673881582174e-04
GC_2_144 b_2 NI_2 NS_144 0 -5.2040472670711656e-05
GC_2_145 b_2 NI_2 NS_145 0 -6.7125275555275825e-03
GC_2_146 b_2 NI_2 NS_146 0 -1.2772742053174799e-03
GC_2_147 b_2 NI_2 NS_147 0 -8.9489728982564908e-06
GC_2_148 b_2 NI_2 NS_148 0 6.1599928232405318e-05
GC_2_149 b_2 NI_2 NS_149 0 -2.9817067265101974e-04
GC_2_150 b_2 NI_2 NS_150 0 5.7412853251855272e-04
GC_2_151 b_2 NI_2 NS_151 0 -2.5290935943304621e-04
GC_2_152 b_2 NI_2 NS_152 0 -2.6220952131041481e-03
GC_2_153 b_2 NI_2 NS_153 0 1.7046023056426879e-04
GC_2_154 b_2 NI_2 NS_154 0 1.1461022660858142e-04
GC_2_155 b_2 NI_2 NS_155 0 2.7258146709332989e-06
GC_2_156 b_2 NI_2 NS_156 0 1.6411699713431926e-06
GC_2_157 b_2 NI_2 NS_157 0 -8.9952760822309473e-06
GC_2_158 b_2 NI_2 NS_158 0 -7.6723026928190184e-06
GC_2_159 b_2 NI_2 NS_159 0 -5.3983039488681891e-05
GC_2_160 b_2 NI_2 NS_160 0 1.8907607765443596e-04
GC_2_161 b_2 NI_2 NS_161 0 -1.1985776192311854e-05
GC_2_162 b_2 NI_2 NS_162 0 -1.8676540732271451e-05
GC_2_163 b_2 NI_2 NS_163 0 -9.3935389493916321e-06
GC_2_164 b_2 NI_2 NS_164 0 7.5934348583198117e-06
GC_2_165 b_2 NI_2 NS_165 0 -7.7891775382643339e-06
GC_2_166 b_2 NI_2 NS_166 0 -5.3546497357605064e-05
GC_2_167 b_2 NI_2 NS_167 0 -1.5897269635651836e-05
GC_2_168 b_2 NI_2 NS_168 0 7.9137096494024886e-05
GC_2_169 b_2 NI_2 NS_169 0 -1.2798903194295684e-02
GC_2_170 b_2 NI_2 NS_170 0 -1.3735151895688182e-03
GC_2_171 b_2 NI_2 NS_171 0 -7.7962845981666942e-04
GC_2_172 b_2 NI_2 NS_172 0 -1.0572048332984690e-03
GC_2_173 b_2 NI_2 NS_173 0 -1.1036283190315804e-03
GC_2_174 b_2 NI_2 NS_174 0 1.5093200932891971e-03
GC_2_175 b_2 NI_2 NS_175 0 7.0972612306937548e-04
GC_2_176 b_2 NI_2 NS_176 0 -2.1293394780239487e-04
GC_2_177 b_2 NI_2 NS_177 0 -3.8917604739495976e-03
GC_2_178 b_2 NI_2 NS_178 0 -8.6536570789337817e-03
GC_2_179 b_2 NI_2 NS_179 0 8.6157430509371176e-05
GC_2_180 b_2 NI_2 NS_180 0 2.5385781240002979e-05
GC_2_181 b_2 NI_2 NS_181 0 2.1257436803678660e-03
GC_2_182 b_2 NI_2 NS_182 0 -2.2730706406083735e-03
GC_2_183 b_2 NI_2 NS_183 0 6.7197057485494937e-04
GC_2_184 b_2 NI_2 NS_184 0 3.0585337893493478e-04
GC_2_185 b_2 NI_2 NS_185 0 7.3461482351454136e-04
GC_2_186 b_2 NI_2 NS_186 0 -2.0411679363500162e-03
GC_2_187 b_2 NI_2 NS_187 0 1.4968514691158970e-03
GC_2_188 b_2 NI_2 NS_188 0 -2.0038818705841359e-03
GC_2_189 b_2 NI_2 NS_189 0 7.7292631871118696e-06
GC_2_190 b_2 NI_2 NS_190 0 2.0772088152379693e-06
GC_2_191 b_2 NI_2 NS_191 0 6.7007287899464689e-03
GC_2_192 b_2 NI_2 NS_192 0 1.4714120732038408e-03
GC_2_193 b_2 NI_2 NS_193 0 -6.0566693759519012e-05
GC_2_194 b_2 NI_2 NS_194 0 2.0744099576978610e-07
GC_2_195 b_2 NI_2 NS_195 0 -3.0959080065083821e-05
GC_2_196 b_2 NI_2 NS_196 0 4.5355675120075711e-05
GC_2_197 b_2 NI_2 NS_197 0 2.4627682350200484e-04
GC_2_198 b_2 NI_2 NS_198 0 -2.2727999067520104e-04
GC_2_199 b_2 NI_2 NS_199 0 2.9855239985703658e-04
GC_2_200 b_2 NI_2 NS_200 0 -7.5248850481225886e-05
GC_2_201 b_2 NI_2 NS_201 0 -8.5166146043966565e-03
GC_2_202 b_2 NI_2 NS_202 0 2.5929244226599265e-03
GC_2_203 b_2 NI_2 NS_203 0 -1.8240805603958311e-04
GC_2_204 b_2 NI_2 NS_204 0 -2.0481532344429135e-04
GC_2_205 b_2 NI_2 NS_205 0 3.4833247209246584e-03
GC_2_206 b_2 NI_2 NS_206 0 7.8743780957204752e-04
GC_2_207 b_2 NI_2 NS_207 0 2.8067326936712842e-03
GC_2_208 b_2 NI_2 NS_208 0 -1.3090522347963818e-03
GC_2_209 b_2 NI_2 NS_209 0 8.0134483786085248e-04
GC_2_210 b_2 NI_2 NS_210 0 1.4275697876460773e-04
GC_2_211 b_2 NI_2 NS_211 0 -1.8181429149265241e-06
GC_2_212 b_2 NI_2 NS_212 0 -2.7381198883077553e-06
GC_2_213 b_2 NI_2 NS_213 0 -1.8801006871482599e-05
GC_2_214 b_2 NI_2 NS_214 0 -1.8315029431094277e-05
GC_2_215 b_2 NI_2 NS_215 0 -8.3260898781688396e-05
GC_2_216 b_2 NI_2 NS_216 0 -4.4662709256309957e-06
GC_2_217 b_2 NI_2 NS_217 0 -3.3079741706845261e-05
GC_2_218 b_2 NI_2 NS_218 0 -1.3760385736903524e-05
GC_2_219 b_2 NI_2 NS_219 0 -1.5576296403275328e-05
GC_2_220 b_2 NI_2 NS_220 0 -1.0832312980412678e-05
GC_2_221 b_2 NI_2 NS_221 0 1.8926518007384858e-04
GC_2_222 b_2 NI_2 NS_222 0 -9.7087313836390388e-05
GC_2_223 b_2 NI_2 NS_223 0 -3.0963968265402294e-04
GC_2_224 b_2 NI_2 NS_224 0 5.9902708952897910e-05
GC_2_225 b_2 NI_2 NS_225 0 -5.8437431343390349e-03
GC_2_226 b_2 NI_2 NS_226 0 -2.5992688754311420e-04
GC_2_227 b_2 NI_2 NS_227 0 -1.3292982173812654e-03
GC_2_228 b_2 NI_2 NS_228 0 3.0355052147258707e-03
GC_2_229 b_2 NI_2 NS_229 0 -9.5126401772886217e-04
GC_2_230 b_2 NI_2 NS_230 0 -2.2008466563582531e-03
GC_2_231 b_2 NI_2 NS_231 0 -5.0103479130262901e-03
GC_2_232 b_2 NI_2 NS_232 0 -5.7005805576151531e-03
GC_2_233 b_2 NI_2 NS_233 0 7.2765678784787770e-03
GC_2_234 b_2 NI_2 NS_234 0 -1.0999239210184204e-03
GC_2_235 b_2 NI_2 NS_235 0 -9.0613370144799042e-05
GC_2_236 b_2 NI_2 NS_236 0 -3.3558464459356500e-05
GC_2_237 b_2 NI_2 NS_237 0 4.0156481686962940e-03
GC_2_238 b_2 NI_2 NS_238 0 -2.3759595544820635e-03
GC_2_239 b_2 NI_2 NS_239 0 7.9215622525377095e-04
GC_2_240 b_2 NI_2 NS_240 0 1.1360894362744736e-03
GC_2_241 b_2 NI_2 NS_241 0 3.0544221532282165e-04
GC_2_242 b_2 NI_2 NS_242 0 2.2186151797784766e-03
GC_2_243 b_2 NI_2 NS_243 0 -3.3756750504005143e-03
GC_2_244 b_2 NI_2 NS_244 0 1.0898686606649439e-03
GC_2_245 b_2 NI_2 NS_245 0 -2.1849272191892775e-04
GC_2_246 b_2 NI_2 NS_246 0 5.6866315100945298e-06
GC_2_247 b_2 NI_2 NS_247 0 2.9342657956879107e-03
GC_2_248 b_2 NI_2 NS_248 0 -4.5477697113913596e-04
GC_2_249 b_2 NI_2 NS_249 0 -1.0827613662088675e-03
GC_2_250 b_2 NI_2 NS_250 0 -1.8172426413043505e-04
GC_2_251 b_2 NI_2 NS_251 0 -1.5170823785683378e-04
GC_2_252 b_2 NI_2 NS_252 0 8.3132763297186107e-05
GC_2_253 b_2 NI_2 NS_253 0 -3.1767124285327129e-04
GC_2_254 b_2 NI_2 NS_254 0 2.8571134671271248e-04
GC_2_255 b_2 NI_2 NS_255 0 -2.0423523715244309e-04
GC_2_256 b_2 NI_2 NS_256 0 -8.7120834806874703e-05
GC_2_257 b_2 NI_2 NS_257 0 2.1318505270863301e-03
GC_2_258 b_2 NI_2 NS_258 0 4.0851511497377355e-07
GC_2_259 b_2 NI_2 NS_259 0 -2.6501039890291786e-05
GC_2_260 b_2 NI_2 NS_260 0 1.2289428691585565e-04
GC_2_261 b_2 NI_2 NS_261 0 -4.6833155305236904e-04
GC_2_262 b_2 NI_2 NS_262 0 -7.2111847405659658e-04
GC_2_263 b_2 NI_2 NS_263 0 -7.0385127645733589e-04
GC_2_264 b_2 NI_2 NS_264 0 1.0700920481879689e-03
GC_2_265 b_2 NI_2 NS_265 0 8.2099507453667724e-05
GC_2_266 b_2 NI_2 NS_266 0 -6.0920722711557747e-05
GC_2_267 b_2 NI_2 NS_267 0 1.0117574893062332e-06
GC_2_268 b_2 NI_2 NS_268 0 -4.8294358437036080e-07
GC_2_269 b_2 NI_2 NS_269 0 -1.0041469975110893e-06
GC_2_270 b_2 NI_2 NS_270 0 2.5545879802866204e-06
GC_2_271 b_2 NI_2 NS_271 0 1.0881026975625784e-04
GC_2_272 b_2 NI_2 NS_272 0 -3.9564429648707290e-06
GC_2_273 b_2 NI_2 NS_273 0 -5.4194295292896328e-06
GC_2_274 b_2 NI_2 NS_274 0 7.8767466564094813e-06
GC_2_275 b_2 NI_2 NS_275 0 -6.9514270065032798e-06
GC_2_276 b_2 NI_2 NS_276 0 -1.6376175821333215e-06
GC_2_277 b_2 NI_2 NS_277 0 -7.1184987483110955e-06
GC_2_278 b_2 NI_2 NS_278 0 7.1693213654211799e-07
GC_2_279 b_2 NI_2 NS_279 0 9.7273291412771540e-06
GC_2_280 b_2 NI_2 NS_280 0 4.0972988851983995e-06
GC_2_281 b_2 NI_2 NS_281 0 1.2032637891326652e-02
GC_2_282 b_2 NI_2 NS_282 0 -7.2270226862523727e-04
GC_2_283 b_2 NI_2 NS_283 0 -1.1910284465163061e-03
GC_2_284 b_2 NI_2 NS_284 0 -1.1286308443557984e-03
GC_2_285 b_2 NI_2 NS_285 0 9.9826007770359437e-04
GC_2_286 b_2 NI_2 NS_286 0 3.4854179319811278e-04
GC_2_287 b_2 NI_2 NS_287 0 4.5306469299292631e-03
GC_2_288 b_2 NI_2 NS_288 0 1.2211091454261331e-03
GC_2_289 b_2 NI_2 NS_289 0 -6.6820236634093748e-03
GC_2_290 b_2 NI_2 NS_290 0 3.5747103329934827e-03
GC_2_291 b_2 NI_2 NS_291 0 -1.6137197653311473e-04
GC_2_292 b_2 NI_2 NS_292 0 6.3875543864493284e-04
GC_2_293 b_2 NI_2 NS_293 0 3.8026641848807757e-05
GC_2_294 b_2 NI_2 NS_294 0 -3.6917289180761590e-03
GC_2_295 b_2 NI_2 NS_295 0 8.0985043945372946e-04
GC_2_296 b_2 NI_2 NS_296 0 4.8595397565357541e-04
GC_2_297 b_2 NI_2 NS_297 0 1.5118653123269419e-04
GC_2_298 b_2 NI_2 NS_298 0 1.5726199271812067e-03
GC_2_299 b_2 NI_2 NS_299 0 1.2904708773208043e-03
GC_2_300 b_2 NI_2 NS_300 0 -1.5030878472658594e-03
GC_2_301 b_2 NI_2 NS_301 0 9.3449949980499450e-05
GC_2_302 b_2 NI_2 NS_302 0 -1.9605129453983336e-05
GC_2_303 b_2 NI_2 NS_303 0 5.6161683856529481e-04
GC_2_304 b_2 NI_2 NS_304 0 2.5506483565814636e-03
GC_2_305 b_2 NI_2 NS_305 0 3.2641404145827997e-04
GC_2_306 b_2 NI_2 NS_306 0 1.0814512994666462e-04
GC_2_307 b_2 NI_2 NS_307 0 -1.7961350877249935e-04
GC_2_308 b_2 NI_2 NS_308 0 -4.0826359738045761e-05
GC_2_309 b_2 NI_2 NS_309 0 1.2862152786601898e-04
GC_2_310 b_2 NI_2 NS_310 0 -2.6556661984788289e-04
GC_2_311 b_2 NI_2 NS_311 0 3.4747760964609018e-04
GC_2_312 b_2 NI_2 NS_312 0 -1.4933843406638329e-04
GC_2_313 b_2 NI_2 NS_313 0 -1.5144877905474152e-02
GC_2_314 b_2 NI_2 NS_314 0 2.3793619515232517e-03
GC_2_315 b_2 NI_2 NS_315 0 -2.1725120545999863e-04
GC_2_316 b_2 NI_2 NS_316 0 -2.8037863194055259e-04
GC_2_317 b_2 NI_2 NS_317 0 4.4112449348026189e-03
GC_2_318 b_2 NI_2 NS_318 0 1.4099792854977400e-03
GC_2_319 b_2 NI_2 NS_319 0 6.8708671874440535e-03
GC_2_320 b_2 NI_2 NS_320 0 -5.2392284240824162e-03
GC_2_321 b_2 NI_2 NS_321 0 1.1178129382874537e-03
GC_2_322 b_2 NI_2 NS_322 0 1.3642544628383389e-04
GC_2_323 b_2 NI_2 NS_323 0 -1.8415218408715050e-07
GC_2_324 b_2 NI_2 NS_324 0 -4.9394087234034317e-06
GC_2_325 b_2 NI_2 NS_325 0 -4.1493492266966181e-05
GC_2_326 b_2 NI_2 NS_326 0 -3.9763491122337783e-05
GC_2_327 b_2 NI_2 NS_327 0 -3.7080463241726284e-04
GC_2_328 b_2 NI_2 NS_328 0 3.3286600653227035e-04
GC_2_329 b_2 NI_2 NS_329 0 -5.4693408707161545e-05
GC_2_330 b_2 NI_2 NS_330 0 -5.5405343873079692e-05
GC_2_331 b_2 NI_2 NS_331 0 -4.9200192694147581e-05
GC_2_332 b_2 NI_2 NS_332 0 -1.0547459974038942e-05
GC_2_333 b_2 NI_2 NS_333 0 3.0569263639511698e-04
GC_2_334 b_2 NI_2 NS_334 0 -2.8722204617325858e-04
GC_2_335 b_2 NI_2 NS_335 0 -5.6334344393852407e-04
GC_2_336 b_2 NI_2 NS_336 0 2.8088331574910866e-04
GC_2_337 b_2 NI_2 NS_337 0 -3.7744081428320628e-02
GC_2_338 b_2 NI_2 NS_338 0 -9.0932264974363363e-05
GC_2_339 b_2 NI_2 NS_339 0 -3.0858689607588381e-04
GC_2_340 b_2 NI_2 NS_340 0 2.4212140736379673e-03
GC_2_341 b_2 NI_2 NS_341 0 -2.5417475313668026e-03
GC_2_342 b_2 NI_2 NS_342 0 -1.4090481662053524e-03
GC_2_343 b_2 NI_2 NS_343 0 -5.7681344956312820e-03
GC_2_344 b_2 NI_2 NS_344 0 -6.2456448783011227e-03
GC_2_345 b_2 NI_2 NS_345 0 8.1080997461525760e-03
GC_2_346 b_2 NI_2 NS_346 0 -9.8242341333045456e-03
GC_2_347 b_2 NI_2 NS_347 0 3.5721824755487587e-04
GC_2_348 b_2 NI_2 NS_348 0 4.3932322268290243e-04
GC_2_349 b_2 NI_2 NS_349 0 5.3359142992848692e-03
GC_2_350 b_2 NI_2 NS_350 0 -2.2773339839649077e-03
GC_2_351 b_2 NI_2 NS_351 0 5.2666382728458353e-04
GC_2_352 b_2 NI_2 NS_352 0 5.6600073516314595e-04
GC_2_353 b_2 NI_2 NS_353 0 1.0159074818498609e-03
GC_2_354 b_2 NI_2 NS_354 0 2.3597400573428630e-03
GC_2_355 b_2 NI_2 NS_355 0 -1.6045620962957811e-04
GC_2_356 b_2 NI_2 NS_356 0 6.9411562632446522e-05
GC_2_357 b_2 NI_2 NS_357 0 -1.7845474784793821e-04
GC_2_358 b_2 NI_2 NS_358 0 7.8033621587528143e-05
GC_2_359 b_2 NI_2 NS_359 0 1.0261232391520620e-03
GC_2_360 b_2 NI_2 NS_360 0 -3.4202526036767682e-03
GC_2_361 b_2 NI_2 NS_361 0 -8.9230910426334154e-04
GC_2_362 b_2 NI_2 NS_362 0 1.7320729742708270e-04
GC_2_363 b_2 NI_2 NS_363 0 -3.2388660653932076e-05
GC_2_364 b_2 NI_2 NS_364 0 3.6437987106815913e-05
GC_2_365 b_2 NI_2 NS_365 0 -2.3531942786654962e-04
GC_2_366 b_2 NI_2 NS_366 0 -2.8014087548916443e-05
GC_2_367 b_2 NI_2 NS_367 0 -9.9213685850764691e-05
GC_2_368 b_2 NI_2 NS_368 0 -1.3351814043004309e-04
GC_2_369 b_2 NI_2 NS_369 0 8.0871988385383346e-03
GC_2_370 b_2 NI_2 NS_370 0 -3.6638662879715661e-05
GC_2_371 b_2 NI_2 NS_371 0 -5.7313388012246619e-05
GC_2_372 b_2 NI_2 NS_372 0 1.2753681639952495e-04
GC_2_373 b_2 NI_2 NS_373 0 -4.6378670170156984e-04
GC_2_374 b_2 NI_2 NS_374 0 -1.4512536239931031e-03
GC_2_375 b_2 NI_2 NS_375 0 -2.0239529926207605e-04
GC_2_376 b_2 NI_2 NS_376 0 2.0288549986203380e-03
GC_2_377 b_2 NI_2 NS_377 0 -3.9067901948651619e-04
GC_2_378 b_2 NI_2 NS_378 0 -6.7787755302829849e-05
GC_2_379 b_2 NI_2 NS_379 0 -2.1470203941047615e-06
GC_2_380 b_2 NI_2 NS_380 0 -2.3909737711553593e-06
GC_2_381 b_2 NI_2 NS_381 0 5.7483737556602762e-06
GC_2_382 b_2 NI_2 NS_382 0 1.4820634674124796e-05
GC_2_383 b_2 NI_2 NS_383 0 1.7966600367815691e-04
GC_2_384 b_2 NI_2 NS_384 0 -1.6573033964209369e-04
GC_2_385 b_2 NI_2 NS_385 0 -8.1028247294888182e-07
GC_2_386 b_2 NI_2 NS_386 0 2.7997753219469377e-05
GC_2_387 b_2 NI_2 NS_387 0 5.2009873171537571e-06
GC_2_388 b_2 NI_2 NS_388 0 4.7376995611873553e-07
GC_2_389 b_2 NI_2 NS_389 0 -1.9362264172633481e-05
GC_2_390 b_2 NI_2 NS_390 0 1.8911107066380537e-05
GC_2_391 b_2 NI_2 NS_391 0 4.0892770381791909e-05
GC_2_392 b_2 NI_2 NS_392 0 -1.0329265962740696e-05
GC_2_393 b_2 NI_2 NS_393 0 3.5910367315370006e-02
GC_2_394 b_2 NI_2 NS_394 0 -3.1429226743116351e-04
GC_2_395 b_2 NI_2 NS_395 0 -9.8606758519924841e-04
GC_2_396 b_2 NI_2 NS_396 0 -7.4407239656688179e-04
GC_2_397 b_2 NI_2 NS_397 0 1.3776247464895245e-03
GC_2_398 b_2 NI_2 NS_398 0 -5.8709030361679031e-04
GC_2_399 b_2 NI_2 NS_399 0 5.8524960557296366e-03
GC_2_400 b_2 NI_2 NS_400 0 1.0117589782778539e-03
GC_2_401 b_2 NI_2 NS_401 0 -2.3683178004464860e-03
GC_2_402 b_2 NI_2 NS_402 0 1.0272689602108422e-02
GC_2_403 b_2 NI_2 NS_403 0 -6.2157140848124581e-04
GC_2_404 b_2 NI_2 NS_404 0 5.6000171216505834e-04
GC_2_405 b_2 NI_2 NS_405 0 -1.2606988330544264e-03
GC_2_406 b_2 NI_2 NS_406 0 -1.0364921425745149e-03
GC_2_407 b_2 NI_2 NS_407 0 7.4875507557964815e-04
GC_2_408 b_2 NI_2 NS_408 0 4.8267935796432064e-04
GC_2_409 b_2 NI_2 NS_409 0 4.9234937065087316e-04
GC_2_410 b_2 NI_2 NS_410 0 5.3901312214264755e-03
GC_2_411 b_2 NI_2 NS_411 0 3.5274397044072326e-04
GC_2_412 b_2 NI_2 NS_412 0 1.7455762014508528e-04
GC_2_413 b_2 NI_2 NS_413 0 1.2493285449655209e-04
GC_2_414 b_2 NI_2 NS_414 0 -9.6936990730175519e-05
GC_2_415 b_2 NI_2 NS_415 0 -5.3911521061942962e-03
GC_2_416 b_2 NI_2 NS_416 0 6.9711323626780661e-03
GC_2_417 b_2 NI_2 NS_417 0 6.0619714866474940e-04
GC_2_418 b_2 NI_2 NS_418 0 -9.4366346682414083e-05
GC_2_419 b_2 NI_2 NS_419 0 -3.9814487410865391e-04
GC_2_420 b_2 NI_2 NS_420 0 8.4054051878745059e-06
GC_2_421 b_2 NI_2 NS_421 0 -2.3339141158860369e-05
GC_2_422 b_2 NI_2 NS_422 0 9.1540846724558558e-05
GC_2_423 b_2 NI_2 NS_423 0 1.1974575860353532e-04
GC_2_424 b_2 NI_2 NS_424 0 2.7722550734262570e-05
GC_2_425 b_2 NI_2 NS_425 0 -1.4763940327448932e-02
GC_2_426 b_2 NI_2 NS_426 0 -2.3762289663708806e-03
GC_2_427 b_2 NI_2 NS_427 0 -4.2613218751495339e-05
GC_2_428 b_2 NI_2 NS_428 0 -2.3098353251976034e-04
GC_2_429 b_2 NI_2 NS_429 0 2.2834434537556884e-03
GC_2_430 b_2 NI_2 NS_430 0 2.8685343114613704e-03
GC_2_431 b_2 NI_2 NS_431 0 5.0342847802196129e-03
GC_2_432 b_2 NI_2 NS_432 0 -5.9581456547060513e-03
GC_2_433 b_2 NI_2 NS_433 0 5.1150303657497293e-04
GC_2_434 b_2 NI_2 NS_434 0 5.9032712986196469e-04
GC_2_435 b_2 NI_2 NS_435 0 1.4572920346555583e-06
GC_2_436 b_2 NI_2 NS_436 0 1.6908306902629452e-06
GC_2_437 b_2 NI_2 NS_437 0 -2.7054273301182909e-05
GC_2_438 b_2 NI_2 NS_438 0 -2.9496064331014186e-05
GC_2_439 b_2 NI_2 NS_439 0 -2.5735080158091194e-04
GC_2_440 b_2 NI_2 NS_440 0 4.3914125023757463e-04
GC_2_441 b_2 NI_2 NS_441 0 -3.6131219803848330e-05
GC_2_442 b_2 NI_2 NS_442 0 -5.5776953002303133e-05
GC_2_443 b_2 NI_2 NS_443 0 -4.1377972421378297e-05
GC_2_444 b_2 NI_2 NS_444 0 -8.0878654923995936e-06
GC_2_445 b_2 NI_2 NS_445 0 2.2984231418617104e-04
GC_2_446 b_2 NI_2 NS_446 0 -1.7204653426358075e-04
GC_2_447 b_2 NI_2 NS_447 0 -4.1222525109965876e-04
GC_2_448 b_2 NI_2 NS_448 0 1.5602551283213739e-04
GC_2_449 b_2 NI_2 NS_449 0 6.8933819317503727e-03
GC_2_450 b_2 NI_2 NS_450 0 -1.0644520660846400e-04
GC_2_451 b_2 NI_2 NS_451 0 2.0352845610884781e-04
GC_2_452 b_2 NI_2 NS_452 0 1.3318975982334664e-05
GC_2_453 b_2 NI_2 NS_453 0 1.1210497364431358e-04
GC_2_454 b_2 NI_2 NS_454 0 2.4840970216949122e-04
GC_2_455 b_2 NI_2 NS_455 0 -2.9209880167927859e-04
GC_2_456 b_2 NI_2 NS_456 0 1.2655702757038954e-03
GC_2_457 b_2 NI_2 NS_457 0 -1.6527243209257488e-03
GC_2_458 b_2 NI_2 NS_458 0 6.1720321042298923e-04
GC_2_459 b_2 NI_2 NS_459 0 2.2969805698199675e-05
GC_2_460 b_2 NI_2 NS_460 0 -6.7241150208234969e-04
GC_2_461 b_2 NI_2 NS_461 0 -5.0508664300412474e-04
GC_2_462 b_2 NI_2 NS_462 0 -9.5467609399853661e-04
GC_2_463 b_2 NI_2 NS_463 0 5.8454731615165231e-04
GC_2_464 b_2 NI_2 NS_464 0 -3.7083277568575773e-04
GC_2_465 b_2 NI_2 NS_465 0 1.4122577837842661e-03
GC_2_466 b_2 NI_2 NS_466 0 1.0497249932325463e-03
GC_2_467 b_2 NI_2 NS_467 0 -7.0611981297312009e-04
GC_2_468 b_2 NI_2 NS_468 0 2.2659496004005944e-03
GC_2_469 b_2 NI_2 NS_469 0 -1.9643866248952670e-04
GC_2_470 b_2 NI_2 NS_470 0 -3.9496959101416074e-05
GC_2_471 b_2 NI_2 NS_471 0 -2.8171317767972390e-03
GC_2_472 b_2 NI_2 NS_472 0 1.8507465934647161e-03
GC_2_473 b_2 NI_2 NS_473 0 3.4238746154189085e-04
GC_2_474 b_2 NI_2 NS_474 0 3.9183739306485326e-04
GC_2_475 b_2 NI_2 NS_475 0 -7.2355628482098221e-04
GC_2_476 b_2 NI_2 NS_476 0 6.4083023710125039e-05
GC_2_477 b_2 NI_2 NS_477 0 -4.8192077080339046e-04
GC_2_478 b_2 NI_2 NS_478 0 -8.8720984604284827e-06
GC_2_479 b_2 NI_2 NS_479 0 -1.0675296667504022e-04
GC_2_480 b_2 NI_2 NS_480 0 -3.9732297252156082e-05
GC_2_481 b_2 NI_2 NS_481 0 -1.2492284418026678e-03
GC_2_482 b_2 NI_2 NS_482 0 -5.7938783285331292e-03
GC_2_483 b_2 NI_2 NS_483 0 5.3639413469965472e-05
GC_2_484 b_2 NI_2 NS_484 0 -2.3815449607207535e-05
GC_2_485 b_2 NI_2 NS_485 0 -1.1841675076423774e-03
GC_2_486 b_2 NI_2 NS_486 0 4.7077786491225653e-04
GC_2_487 b_2 NI_2 NS_487 0 2.2133158999129033e-03
GC_2_488 b_2 NI_2 NS_488 0 9.0375708429624136e-04
GC_2_489 b_2 NI_2 NS_489 0 -5.5571860225568295e-05
GC_2_490 b_2 NI_2 NS_490 0 8.5588308608980121e-05
GC_2_491 b_2 NI_2 NS_491 0 -1.8478033189025696e-06
GC_2_492 b_2 NI_2 NS_492 0 6.1298819363354745e-07
GC_2_493 b_2 NI_2 NS_493 0 4.5507247070893123e-06
GC_2_494 b_2 NI_2 NS_494 0 -3.6783055166436088e-06
GC_2_495 b_2 NI_2 NS_495 0 -1.4969050344462400e-04
GC_2_496 b_2 NI_2 NS_496 0 -7.6982179370024587e-05
GC_2_497 b_2 NI_2 NS_497 0 1.1121307654470358e-05
GC_2_498 b_2 NI_2 NS_498 0 -2.1018406954451733e-06
GC_2_499 b_2 NI_2 NS_499 0 6.6808464656059868e-06
GC_2_500 b_2 NI_2 NS_500 0 -1.1074127821071045e-05
GC_2_501 b_2 NI_2 NS_501 0 3.3025178294525827e-05
GC_2_502 b_2 NI_2 NS_502 0 4.5271129853185612e-05
GC_2_503 b_2 NI_2 NS_503 0 -2.7214012701539643e-05
GC_2_504 b_2 NI_2 NS_504 0 -8.3981291250880585e-05
GC_2_505 b_2 NI_2 NS_505 0 -4.8613628801469164e-03
GC_2_506 b_2 NI_2 NS_506 0 1.2504095849436104e-05
GC_2_507 b_2 NI_2 NS_507 0 -8.5592895262749435e-05
GC_2_508 b_2 NI_2 NS_508 0 8.1985214466445805e-05
GC_2_509 b_2 NI_2 NS_509 0 -1.5105019694404019e-04
GC_2_510 b_2 NI_2 NS_510 0 -5.6342206206584492e-05
GC_2_511 b_2 NI_2 NS_511 0 -3.4950084920867120e-04
GC_2_512 b_2 NI_2 NS_512 0 -8.4344312354503979e-04
GC_2_513 b_2 NI_2 NS_513 0 8.4168984435091044e-04
GC_2_514 b_2 NI_2 NS_514 0 -8.5660294286593684e-04
GC_2_515 b_2 NI_2 NS_515 0 -8.3025956917493932e-05
GC_2_516 b_2 NI_2 NS_516 0 -3.0335263408558141e-04
GC_2_517 b_2 NI_2 NS_517 0 -5.2232730692755370e-05
GC_2_518 b_2 NI_2 NS_518 0 -3.6360763275085296e-04
GC_2_519 b_2 NI_2 NS_519 0 2.5710647125127965e-04
GC_2_520 b_2 NI_2 NS_520 0 -4.3842628548464765e-04
GC_2_521 b_2 NI_2 NS_521 0 7.1113824972634989e-04
GC_2_522 b_2 NI_2 NS_522 0 2.6094297775467080e-04
GC_2_523 b_2 NI_2 NS_523 0 -9.1662656257158288e-04
GC_2_524 b_2 NI_2 NS_524 0 -6.4155290721427905e-04
GC_2_525 b_2 NI_2 NS_525 0 1.1410892663369088e-04
GC_2_526 b_2 NI_2 NS_526 0 5.8382742747894538e-05
GC_2_527 b_2 NI_2 NS_527 0 3.8663637365475589e-03
GC_2_528 b_2 NI_2 NS_528 0 -1.7525553831201095e-03
GC_2_529 b_2 NI_2 NS_529 0 -4.3608719419699365e-04
GC_2_530 b_2 NI_2 NS_530 0 3.2550078920472501e-04
GC_2_531 b_2 NI_2 NS_531 0 -3.1011544371371125e-04
GC_2_532 b_2 NI_2 NS_532 0 4.5865175709288027e-04
GC_2_533 b_2 NI_2 NS_533 0 -4.7654157987813751e-05
GC_2_534 b_2 NI_2 NS_534 0 -4.6737828820807764e-04
GC_2_535 b_2 NI_2 NS_535 0 1.8169937734192193e-04
GC_2_536 b_2 NI_2 NS_536 0 -1.7472912262262396e-05
GC_2_537 b_2 NI_2 NS_537 0 7.9546172492166493e-04
GC_2_538 b_2 NI_2 NS_538 0 4.7628415835891252e-03
GC_2_539 b_2 NI_2 NS_539 0 -1.0855606152513290e-04
GC_2_540 b_2 NI_2 NS_540 0 1.8723149207928162e-04
GC_2_541 b_2 NI_2 NS_541 0 1.6604547346938626e-03
GC_2_542 b_2 NI_2 NS_542 0 -8.3590331480120803e-04
GC_2_543 b_2 NI_2 NS_543 0 -3.1566913070166101e-03
GC_2_544 b_2 NI_2 NS_544 0 -1.3331616079304890e-03
GC_2_545 b_2 NI_2 NS_545 0 -5.1394661386951819e-04
GC_2_546 b_2 NI_2 NS_546 0 4.8358058258116110e-04
GC_2_547 b_2 NI_2 NS_547 0 5.2981377580914924e-06
GC_2_548 b_2 NI_2 NS_548 0 -5.9206901969566402e-06
GC_2_549 b_2 NI_2 NS_549 0 1.0611129974088318e-06
GC_2_550 b_2 NI_2 NS_550 0 6.1285182886373804e-05
GC_2_551 b_2 NI_2 NS_551 0 3.0114607947007545e-04
GC_2_552 b_2 NI_2 NS_552 0 -1.6904585293554415e-04
GC_2_553 b_2 NI_2 NS_553 0 4.7392356731492710e-05
GC_2_554 b_2 NI_2 NS_554 0 7.3875693362933088e-05
GC_2_555 b_2 NI_2 NS_555 0 1.1853743967797268e-05
GC_2_556 b_2 NI_2 NS_556 0 4.5739162550090911e-05
GC_2_557 b_2 NI_2 NS_557 0 1.7738831963380643e-04
GC_2_558 b_2 NI_2 NS_558 0 -1.9777833066230035e-04
GC_2_559 b_2 NI_2 NS_559 0 -3.1917549713475626e-04
GC_2_560 b_2 NI_2 NS_560 0 2.1291102533670426e-04
GC_2_561 b_2 NI_2 NS_561 0 -6.3518825150371584e-03
GC_2_562 b_2 NI_2 NS_562 0 -1.0081876760133912e-04
GC_2_563 b_2 NI_2 NS_563 0 2.5384877415705756e-04
GC_2_564 b_2 NI_2 NS_564 0 2.9809391808544895e-04
GC_2_565 b_2 NI_2 NS_565 0 -3.5932983007142455e-04
GC_2_566 b_2 NI_2 NS_566 0 3.0721814472934672e-04
GC_2_567 b_2 NI_2 NS_567 0 -1.7649585074817652e-03
GC_2_568 b_2 NI_2 NS_568 0 2.7455024735818247e-04
GC_2_569 b_2 NI_2 NS_569 0 -1.2020526483094219e-03
GC_2_570 b_2 NI_2 NS_570 0 -2.4964273512982208e-03
GC_2_571 b_2 NI_2 NS_571 0 5.9946031205910578e-04
GC_2_572 b_2 NI_2 NS_572 0 -4.4721532436221053e-04
GC_2_573 b_2 NI_2 NS_573 0 7.3554217786908074e-04
GC_2_574 b_2 NI_2 NS_574 0 -1.7145084796334603e-03
GC_2_575 b_2 NI_2 NS_575 0 3.8518369841138275e-04
GC_2_576 b_2 NI_2 NS_576 0 -1.9544643462083493e-04
GC_2_577 b_2 NI_2 NS_577 0 1.4905749938434827e-03
GC_2_578 b_2 NI_2 NS_578 0 1.1008207424833586e-03
GC_2_579 b_2 NI_2 NS_579 0 -5.3474494476073208e-04
GC_2_580 b_2 NI_2 NS_580 0 9.0367037034468837e-04
GC_2_581 b_2 NI_2 NS_581 0 -1.1872172573019986e-04
GC_2_582 b_2 NI_2 NS_582 0 4.4347108448606650e-05
GC_2_583 b_2 NI_2 NS_583 0 -2.5664879608193413e-03
GC_2_584 b_2 NI_2 NS_584 0 -5.0936308984211366e-04
GC_2_585 b_2 NI_2 NS_585 0 3.1108016566690817e-05
GC_2_586 b_2 NI_2 NS_586 0 6.2462264487415237e-04
GC_2_587 b_2 NI_2 NS_587 0 -3.8495822163254291e-04
GC_2_588 b_2 NI_2 NS_588 0 1.3247920809456584e-05
GC_2_589 b_2 NI_2 NS_589 0 -4.1481098937186178e-04
GC_2_590 b_2 NI_2 NS_590 0 -9.6518399696319567e-05
GC_2_591 b_2 NI_2 NS_591 0 -8.4349460368413762e-05
GC_2_592 b_2 NI_2 NS_592 0 -9.2948657357268328e-05
GC_2_593 b_2 NI_2 NS_593 0 2.9607833226215890e-03
GC_2_594 b_2 NI_2 NS_594 0 -4.5932897099369178e-03
GC_2_595 b_2 NI_2 NS_595 0 1.6884833381500761e-05
GC_2_596 b_2 NI_2 NS_596 0 4.3792659461857264e-05
GC_2_597 b_2 NI_2 NS_597 0 -1.0129361422474090e-03
GC_2_598 b_2 NI_2 NS_598 0 -4.1718160094560212e-04
GC_2_599 b_2 NI_2 NS_599 0 7.6169041996018412e-04
GC_2_600 b_2 NI_2 NS_600 0 1.6985234613869475e-03
GC_2_601 b_2 NI_2 NS_601 0 -1.9284682913115242e-04
GC_2_602 b_2 NI_2 NS_602 0 6.9016590704690882e-05
GC_2_603 b_2 NI_2 NS_603 0 -3.5285770419473263e-06
GC_2_604 b_2 NI_2 NS_604 0 -9.4886666779542527e-07
GC_2_605 b_2 NI_2 NS_605 0 1.0819846895330371e-05
GC_2_606 b_2 NI_2 NS_606 0 7.0055322870835496e-06
GC_2_607 b_2 NI_2 NS_607 0 -5.8573627167801826e-05
GC_2_608 b_2 NI_2 NS_608 0 -2.2009852464768839e-04
GC_2_609 b_2 NI_2 NS_609 0 2.3120321964674558e-05
GC_2_610 b_2 NI_2 NS_610 0 1.6594776746843874e-05
GC_2_611 b_2 NI_2 NS_611 0 1.7087941099968626e-05
GC_2_612 b_2 NI_2 NS_612 0 -9.4796204582707297e-06
GC_2_613 b_2 NI_2 NS_613 0 1.6240348733158148e-05
GC_2_614 b_2 NI_2 NS_614 0 4.8356424693522560e-05
GC_2_615 b_2 NI_2 NS_615 0 6.5092655283588074e-06
GC_2_616 b_2 NI_2 NS_616 0 -7.6064802322646535e-05
GC_2_617 b_2 NI_2 NS_617 0 6.5332306778082020e-03
GC_2_618 b_2 NI_2 NS_618 0 -4.6004791693508609e-06
GC_2_619 b_2 NI_2 NS_619 0 -2.2451200675513387e-04
GC_2_620 b_2 NI_2 NS_620 0 1.0290603925402305e-05
GC_2_621 b_2 NI_2 NS_621 0 -5.1957644364984904e-06
GC_2_622 b_2 NI_2 NS_622 0 -2.8521714318300884e-04
GC_2_623 b_2 NI_2 NS_623 0 9.2569461080844150e-04
GC_2_624 b_2 NI_2 NS_624 0 -9.7941643978760313e-04
GC_2_625 b_2 NI_2 NS_625 0 1.8408054698002944e-03
GC_2_626 b_2 NI_2 NS_626 0 1.3644773320635769e-03
GC_2_627 b_2 NI_2 NS_627 0 -6.0706432119539226e-04
GC_2_628 b_2 NI_2 NS_628 0 3.6954344488114376e-04
GC_2_629 b_2 NI_2 NS_629 0 -1.6228634437263468e-05
GC_2_630 b_2 NI_2 NS_630 0 1.6181464691945936e-04
GC_2_631 b_2 NI_2 NS_631 0 3.6050867524336919e-04
GC_2_632 b_2 NI_2 NS_632 0 -1.7203513699822252e-04
GC_2_633 b_2 NI_2 NS_633 0 1.5310678048170959e-03
GC_2_634 b_2 NI_2 NS_634 0 1.6236685147743299e-03
GC_2_635 b_2 NI_2 NS_635 0 -4.2217538500447150e-04
GC_2_636 b_2 NI_2 NS_636 0 6.3770821157185837e-06
GC_2_637 b_2 NI_2 NS_637 0 7.1412911020107294e-05
GC_2_638 b_2 NI_2 NS_638 0 8.0109964101663356e-06
GC_2_639 b_2 NI_2 NS_639 0 1.3339226480310886e-03
GC_2_640 b_2 NI_2 NS_640 0 2.3726207126616968e-03
GC_2_641 b_2 NI_2 NS_641 0 -8.7320947498269376e-05
GC_2_642 b_2 NI_2 NS_642 0 1.0173817586041512e-04
GC_2_643 b_2 NI_2 NS_643 0 -2.9829627394234573e-04
GC_2_644 b_2 NI_2 NS_644 0 2.7549361649724683e-04
GC_2_645 b_2 NI_2 NS_645 0 2.6288256347032482e-05
GC_2_646 b_2 NI_2 NS_646 0 -1.7328847209552829e-04
GC_2_647 b_2 NI_2 NS_647 0 1.1221792263806579e-04
GC_2_648 b_2 NI_2 NS_648 0 4.2270672723523392e-05
GC_2_649 b_2 NI_2 NS_649 0 -3.9389346470361389e-03
GC_2_650 b_2 NI_2 NS_650 0 2.5330233660196448e-03
GC_2_651 b_2 NI_2 NS_651 0 -8.1070847226315276e-05
GC_2_652 b_2 NI_2 NS_652 0 2.3559984152372804e-06
GC_2_653 b_2 NI_2 NS_653 0 1.6437105092909825e-03
GC_2_654 b_2 NI_2 NS_654 0 6.6062319480681678e-04
GC_2_655 b_2 NI_2 NS_655 0 -1.3701144339382403e-03
GC_2_656 b_2 NI_2 NS_656 0 -2.7717461229871485e-03
GC_2_657 b_2 NI_2 NS_657 0 -9.2689362393121635e-05
GC_2_658 b_2 NI_2 NS_658 0 3.8985275793156668e-04
GC_2_659 b_2 NI_2 NS_659 0 4.9482637786735591e-06
GC_2_660 b_2 NI_2 NS_660 0 -1.1087045889509808e-06
GC_2_661 b_2 NI_2 NS_661 0 -1.4236523276791935e-05
GC_2_662 b_2 NI_2 NS_662 0 2.4194250673175203e-05
GC_2_663 b_2 NI_2 NS_663 0 2.2701005965866758e-04
GC_2_664 b_2 NI_2 NS_664 0 6.8932487833522896e-05
GC_2_665 b_2 NI_2 NS_665 0 1.8021726190300823e-06
GC_2_666 b_2 NI_2 NS_666 0 3.3011302570030702e-05
GC_2_667 b_2 NI_2 NS_667 0 -1.4465508678393518e-05
GC_2_668 b_2 NI_2 NS_668 0 2.8840373491436287e-05
GC_2_669 b_2 NI_2 NS_669 0 1.3309326230905643e-04
GC_2_670 b_2 NI_2 NS_670 0 -1.2730198132296619e-04
GC_2_671 b_2 NI_2 NS_671 0 -2.3862282960066222e-04
GC_2_672 b_2 NI_2 NS_672 0 1.3943998138661452e-04
GD_2_1 b_2 NI_2 NA_1 0 1.4108445671219128e-02
GD_2_2 b_2 NI_2 NA_2 0 1.2534658725686457e-01
GD_2_3 b_2 NI_2 NA_3 0 -5.8445864033969050e-02
GD_2_4 b_2 NI_2 NA_4 0 1.1471403074311859e-02
GD_2_5 b_2 NI_2 NA_5 0 2.9162948474695007e-03
GD_2_6 b_2 NI_2 NA_6 0 -2.0018996693913955e-02
GD_2_7 b_2 NI_2 NA_7 0 4.0311334785694625e-02
GD_2_8 b_2 NI_2 NA_8 0 -4.7215764370695842e-02
GD_2_9 b_2 NI_2 NA_9 0 -5.2820242334684876e-04
GD_2_10 b_2 NI_2 NA_10 0 3.9415667803263908e-03
GD_2_11 b_2 NI_2 NA_11 0 1.5285228591889808e-02
GD_2_12 b_2 NI_2 NA_12 0 -1.2519126254088653e-02
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 -3.0061678552868780e-02
GC_3_2 b_3 NI_3 NS_2 0 1.7198922485852435e-03
GC_3_3 b_3 NI_3 NS_3 0 3.6993481782394925e-03
GC_3_4 b_3 NI_3 NS_4 0 2.5857513434127143e-03
GC_3_5 b_3 NI_3 NS_5 0 -5.7084431512842366e-03
GC_3_6 b_3 NI_3 NS_6 0 -6.5718121671506534e-03
GC_3_7 b_3 NI_3 NS_7 0 3.6822857173954789e-03
GC_3_8 b_3 NI_3 NS_8 0 1.5264879083350198e-03
GC_3_9 b_3 NI_3 NS_9 0 1.0503292478048057e-02
GC_3_10 b_3 NI_3 NS_10 0 -1.1738965848324085e-02
GC_3_11 b_3 NI_3 NS_11 0 -3.1359001327008787e-04
GC_3_12 b_3 NI_3 NS_12 0 3.7815499837699345e-04
GC_3_13 b_3 NI_3 NS_13 0 8.9978538009992289e-03
GC_3_14 b_3 NI_3 NS_14 0 3.2733639668079476e-03
GC_3_15 b_3 NI_3 NS_15 0 3.0707357152310352e-04
GC_3_16 b_3 NI_3 NS_16 0 2.1644017065029415e-03
GC_3_17 b_3 NI_3 NS_17 0 6.9122911817196871e-03
GC_3_18 b_3 NI_3 NS_18 0 -9.4757062615213159e-05
GC_3_19 b_3 NI_3 NS_19 0 2.1100430980749070e-03
GC_3_20 b_3 NI_3 NS_20 0 3.5101180094787346e-03
GC_3_21 b_3 NI_3 NS_21 0 2.4907149336475255e-04
GC_3_22 b_3 NI_3 NS_22 0 7.6313269788912713e-05
GC_3_23 b_3 NI_3 NS_23 0 -2.9575680320381090e-03
GC_3_24 b_3 NI_3 NS_24 0 1.0405969697255154e-02
GC_3_25 b_3 NI_3 NS_25 0 1.1307156915990580e-03
GC_3_26 b_3 NI_3 NS_26 0 2.1733352820311235e-04
GC_3_27 b_3 NI_3 NS_27 0 -3.3581849914702297e-04
GC_3_28 b_3 NI_3 NS_28 0 1.3357878838928886e-04
GC_3_29 b_3 NI_3 NS_29 0 -1.0068490824022127e-04
GC_3_30 b_3 NI_3 NS_30 0 2.6008483044003835e-04
GC_3_31 b_3 NI_3 NS_31 0 -5.6162723457585467e-05
GC_3_32 b_3 NI_3 NS_32 0 1.6912398887465918e-05
GC_3_33 b_3 NI_3 NS_33 0 -1.5928408894039477e-03
GC_3_34 b_3 NI_3 NS_34 0 -4.3090501890928343e-03
GC_3_35 b_3 NI_3 NS_35 0 1.0073688950415506e-04
GC_3_36 b_3 NI_3 NS_36 0 -2.1165660277797066e-05
GC_3_37 b_3 NI_3 NS_37 0 -4.4324151069423693e-04
GC_3_38 b_3 NI_3 NS_38 0 1.5110486192706286e-03
GC_3_39 b_3 NI_3 NS_39 0 -2.4284296528299387e-04
GC_3_40 b_3 NI_3 NS_40 0 2.2524629335597584e-03
GC_3_41 b_3 NI_3 NS_41 0 3.5591338445405516e-05
GC_3_42 b_3 NI_3 NS_42 0 9.5883026259629308e-05
GC_3_43 b_3 NI_3 NS_43 0 -1.1070332931778496e-07
GC_3_44 b_3 NI_3 NS_44 0 -2.0307617893383492e-07
GC_3_45 b_3 NI_3 NS_45 0 4.0069034497164482e-06
GC_3_46 b_3 NI_3 NS_46 0 2.9542911482460244e-06
GC_3_47 b_3 NI_3 NS_47 0 3.1009779820116461e-05
GC_3_48 b_3 NI_3 NS_48 0 -4.7582579357984296e-05
GC_3_49 b_3 NI_3 NS_49 0 3.9521651290419672e-06
GC_3_50 b_3 NI_3 NS_50 0 7.8537545181724395e-06
GC_3_51 b_3 NI_3 NS_51 0 5.7934194423373685e-06
GC_3_52 b_3 NI_3 NS_52 0 -8.5733407084049360e-07
GC_3_53 b_3 NI_3 NS_53 0 -2.0764588292910486e-06
GC_3_54 b_3 NI_3 NS_54 0 1.2093767465601042e-05
GC_3_55 b_3 NI_3 NS_55 0 8.5478539841460428e-06
GC_3_56 b_3 NI_3 NS_56 0 -1.6952655547589756e-05
GC_3_57 b_3 NI_3 NS_57 0 5.8904813671215479e-02
GC_3_58 b_3 NI_3 NS_58 0 -7.7058472661268662e-04
GC_3_59 b_3 NI_3 NS_59 0 -1.8477663733942962e-03
GC_3_60 b_3 NI_3 NS_60 0 2.3852737836363648e-03
GC_3_61 b_3 NI_3 NS_61 0 2.9557673877873931e-03
GC_3_62 b_3 NI_3 NS_62 0 1.3870493842929238e-04
GC_3_63 b_3 NI_3 NS_63 0 -5.2073017576517453e-03
GC_3_64 b_3 NI_3 NS_64 0 3.6875906356174281e-04
GC_3_65 b_3 NI_3 NS_65 0 -5.9150297396448216e-03
GC_3_66 b_3 NI_3 NS_66 0 1.1177472469113088e-02
GC_3_67 b_3 NI_3 NS_67 0 -6.2312734181708376e-04
GC_3_68 b_3 NI_3 NS_68 0 -1.0715164632992204e-05
GC_3_69 b_3 NI_3 NS_69 0 1.5956146972993656e-03
GC_3_70 b_3 NI_3 NS_70 0 -3.9321062194462245e-03
GC_3_71 b_3 NI_3 NS_71 0 8.7691057710770999e-04
GC_3_72 b_3 NI_3 NS_72 0 1.5833254259819429e-03
GC_3_73 b_3 NI_3 NS_73 0 -8.9525702965525731e-04
GC_3_74 b_3 NI_3 NS_74 0 1.0681648793013543e-03
GC_3_75 b_3 NI_3 NS_75 0 -6.1601864062889771e-03
GC_3_76 b_3 NI_3 NS_76 0 4.4880520179807769e-04
GC_3_77 b_3 NI_3 NS_77 0 -7.6801113580115242e-05
GC_3_78 b_3 NI_3 NS_78 0 -9.6447244105482566e-05
GC_3_79 b_3 NI_3 NS_79 0 1.1955370131150726e-03
GC_3_80 b_3 NI_3 NS_80 0 4.8946183370859953e-03
GC_3_81 b_3 NI_3 NS_81 0 -5.2880103799230599e-04
GC_3_82 b_3 NI_3 NS_82 0 -3.1099948303397735e-04
GC_3_83 b_3 NI_3 NS_83 0 -3.3143186335715609e-04
GC_3_84 b_3 NI_3 NS_84 0 3.7071894161078104e-05
GC_3_85 b_3 NI_3 NS_85 0 -4.0297072770120366e-04
GC_3_86 b_3 NI_3 NS_86 0 4.5626748235648071e-04
GC_3_87 b_3 NI_3 NS_87 0 -2.7267673881586240e-04
GC_3_88 b_3 NI_3 NS_88 0 -5.2040472670612092e-05
GC_3_89 b_3 NI_3 NS_89 0 -6.7125275555387489e-03
GC_3_90 b_3 NI_3 NS_90 0 -1.2772742053178264e-03
GC_3_91 b_3 NI_3 NS_91 0 -8.9489728982356979e-06
GC_3_92 b_3 NI_3 NS_92 0 6.1599928232296424e-05
GC_3_93 b_3 NI_3 NS_93 0 -2.9817067265028752e-04
GC_3_94 b_3 NI_3 NS_94 0 5.7412853252032116e-04
GC_3_95 b_3 NI_3 NS_95 0 -2.5290935943350547e-04
GC_3_96 b_3 NI_3 NS_96 0 -2.6220952131110983e-03
GC_3_97 b_3 NI_3 NS_97 0 1.7046023056462240e-04
GC_3_98 b_3 NI_3 NS_98 0 1.1461022660873432e-04
GC_3_99 b_3 NI_3 NS_99 0 2.7258146709366811e-06
GC_3_100 b_3 NI_3 NS_100 0 1.6411699713442885e-06
GC_3_101 b_3 NI_3 NS_101 0 -8.9952760822540476e-06
GC_3_102 b_3 NI_3 NS_102 0 -7.6723026928206972e-06
GC_3_103 b_3 NI_3 NS_103 0 -5.3983039488507924e-05
GC_3_104 b_3 NI_3 NS_104 0 1.8907607765480258e-04
GC_3_105 b_3 NI_3 NS_105 0 -1.1985776192355350e-05
GC_3_106 b_3 NI_3 NS_106 0 -1.8676540732283726e-05
GC_3_107 b_3 NI_3 NS_107 0 -9.3935389494078291e-06
GC_3_108 b_3 NI_3 NS_108 0 7.5934348583482847e-06
GC_3_109 b_3 NI_3 NS_109 0 -7.7891775383150560e-06
GC_3_110 b_3 NI_3 NS_110 0 -5.3546497357698563e-05
GC_3_111 b_3 NI_3 NS_111 0 -1.5897269635619354e-05
GC_3_112 b_3 NI_3 NS_112 0 7.9137096494190877e-05
GC_3_113 b_3 NI_3 NS_113 0 -1.9831653589567472e-02
GC_3_114 b_3 NI_3 NS_114 0 1.4980049510268326e-02
GC_3_115 b_3 NI_3 NS_115 0 8.3191373700100477e-03
GC_3_116 b_3 NI_3 NS_116 0 1.3388313318701752e-03
GC_3_117 b_3 NI_3 NS_117 0 9.9266241581687543e-03
GC_3_118 b_3 NI_3 NS_118 0 5.2662762738067822e-03
GC_3_119 b_3 NI_3 NS_119 0 -3.1032396492007399e-03
GC_3_120 b_3 NI_3 NS_120 0 8.5536253966760015e-03
GC_3_121 b_3 NI_3 NS_121 0 -3.0116495696150256e-03
GC_3_122 b_3 NI_3 NS_122 0 4.4654007125132129e-03
GC_3_123 b_3 NI_3 NS_123 0 1.0372541279033059e-04
GC_3_124 b_3 NI_3 NS_124 0 1.0275997741687052e-03
GC_3_125 b_3 NI_3 NS_125 0 1.1666252115683283e-02
GC_3_126 b_3 NI_3 NS_126 0 -2.2579156220219648e-03
GC_3_127 b_3 NI_3 NS_127 0 1.6560996142643613e-05
GC_3_128 b_3 NI_3 NS_128 0 3.3819925704405927e-03
GC_3_129 b_3 NI_3 NS_129 0 3.3878896842682140e-03
GC_3_130 b_3 NI_3 NS_130 0 1.5595227640346403e-03
GC_3_131 b_3 NI_3 NS_131 0 3.1820062013416142e-03
GC_3_132 b_3 NI_3 NS_132 0 7.6032781054045338e-03
GC_3_133 b_3 NI_3 NS_133 0 3.2716546138672790e-04
GC_3_134 b_3 NI_3 NS_134 0 2.5218686457107765e-04
GC_3_135 b_3 NI_3 NS_135 0 -6.6790616836194952e-03
GC_3_136 b_3 NI_3 NS_136 0 9.5092304009987590e-04
GC_3_137 b_3 NI_3 NS_137 0 1.1896631559105326e-03
GC_3_138 b_3 NI_3 NS_138 0 9.6700962174392079e-04
GC_3_139 b_3 NI_3 NS_139 0 -2.5700474892163968e-04
GC_3_140 b_3 NI_3 NS_140 0 2.3605962752840370e-05
GC_3_141 b_3 NI_3 NS_141 0 -1.6929447931299029e-04
GC_3_142 b_3 NI_3 NS_142 0 1.2508690338039515e-04
GC_3_143 b_3 NI_3 NS_143 0 -5.5063507162005878e-05
GC_3_144 b_3 NI_3 NS_144 0 -4.3388828817828780e-05
GC_3_145 b_3 NI_3 NS_145 0 3.2016517659980473e-05
GC_3_146 b_3 NI_3 NS_146 0 -3.2129527676983973e-03
GC_3_147 b_3 NI_3 NS_147 0 1.1104783844985688e-04
GC_3_148 b_3 NI_3 NS_148 0 3.9589903912866557e-05
GC_3_149 b_3 NI_3 NS_149 0 -9.1858734302535661e-04
GC_3_150 b_3 NI_3 NS_150 0 1.1188656055821167e-03
GC_3_151 b_3 NI_3 NS_151 0 2.9932977831156602e-03
GC_3_152 b_3 NI_3 NS_152 0 4.3537729960042232e-03
GC_3_153 b_3 NI_3 NS_153 0 -2.7154620384415129e-05
GC_3_154 b_3 NI_3 NS_154 0 -3.7496132673397694e-05
GC_3_155 b_3 NI_3 NS_155 0 -1.5271141186308355e-06
GC_3_156 b_3 NI_3 NS_156 0 -1.1178565905019278e-06
GC_3_157 b_3 NI_3 NS_157 0 1.1247242640059570e-05
GC_3_158 b_3 NI_3 NS_158 0 8.6817243860901188e-06
GC_3_159 b_3 NI_3 NS_159 0 2.0961163886001723e-06
GC_3_160 b_3 NI_3 NS_160 0 -2.2467508971357760e-04
GC_3_161 b_3 NI_3 NS_161 0 1.8580945442475934e-05
GC_3_162 b_3 NI_3 NS_162 0 2.0323355415632612e-05
GC_3_163 b_3 NI_3 NS_163 0 1.6216031122509201e-05
GC_3_164 b_3 NI_3 NS_164 0 -1.1698880865250408e-05
GC_3_165 b_3 NI_3 NS_165 0 1.3474650644604439e-05
GC_3_166 b_3 NI_3 NS_166 0 6.6280509166160483e-05
GC_3_167 b_3 NI_3 NS_167 0 1.0749158398608779e-05
GC_3_168 b_3 NI_3 NS_168 0 -1.0486893042091272e-04
GC_3_169 b_3 NI_3 NS_169 0 -3.9239711967129047e-02
GC_3_170 b_3 NI_3 NS_170 0 1.1912590977744983e-02
GC_3_171 b_3 NI_3 NS_171 0 -2.9631647745846481e-03
GC_3_172 b_3 NI_3 NS_172 0 3.8370699507883446e-03
GC_3_173 b_3 NI_3 NS_173 0 -4.5209998938928447e-03
GC_3_174 b_3 NI_3 NS_174 0 2.0762529289841953e-03
GC_3_175 b_3 NI_3 NS_175 0 -4.6100700842438731e-03
GC_3_176 b_3 NI_3 NS_176 0 -9.0087771136975660e-03
GC_3_177 b_3 NI_3 NS_177 0 -2.2016986909280745e-03
GC_3_178 b_3 NI_3 NS_178 0 -8.6781035757114815e-03
GC_3_179 b_3 NI_3 NS_179 0 7.2684118588135988e-04
GC_3_180 b_3 NI_3 NS_180 0 -1.4323299987929045e-04
GC_3_181 b_3 NI_3 NS_181 0 6.8572941190360309e-03
GC_3_182 b_3 NI_3 NS_182 0 -5.0622900790423539e-04
GC_3_183 b_3 NI_3 NS_183 0 1.2644404686549490e-03
GC_3_184 b_3 NI_3 NS_184 0 1.4479564218832332e-03
GC_3_185 b_3 NI_3 NS_185 0 4.3732778280134573e-03
GC_3_186 b_3 NI_3 NS_186 0 1.6167447990985443e-03
GC_3_187 b_3 NI_3 NS_187 0 -2.2047009088209122e-03
GC_3_188 b_3 NI_3 NS_188 0 9.4748631449837525e-04
GC_3_189 b_3 NI_3 NS_189 0 -2.4089088171210156e-04
GC_3_190 b_3 NI_3 NS_190 0 2.9282183121520413e-06
GC_3_191 b_3 NI_3 NS_191 0 5.3978745791555599e-03
GC_3_192 b_3 NI_3 NS_192 0 -2.1314084227527052e-03
GC_3_193 b_3 NI_3 NS_193 0 -1.2310588939635266e-03
GC_3_194 b_3 NI_3 NS_194 0 -2.2056253294854981e-04
GC_3_195 b_3 NI_3 NS_195 0 -1.7998280294237901e-04
GC_3_196 b_3 NI_3 NS_196 0 2.3497368635757447e-05
GC_3_197 b_3 NI_3 NS_197 0 -4.1235200157247696e-04
GC_3_198 b_3 NI_3 NS_198 0 2.8860449762701477e-04
GC_3_199 b_3 NI_3 NS_199 0 -2.2729731722031447e-04
GC_3_200 b_3 NI_3 NS_200 0 -1.2617695839982449e-04
GC_3_201 b_3 NI_3 NS_201 0 1.0266668770112870e-03
GC_3_202 b_3 NI_3 NS_202 0 -1.6449325450807728e-04
GC_3_203 b_3 NI_3 NS_203 0 -4.2568704220306658e-05
GC_3_204 b_3 NI_3 NS_204 0 1.2650722765239920e-04
GC_3_205 b_3 NI_3 NS_205 0 -5.3924316988106940e-04
GC_3_206 b_3 NI_3 NS_206 0 -7.0337230304038127e-04
GC_3_207 b_3 NI_3 NS_207 0 2.7149552122342690e-03
GC_3_208 b_3 NI_3 NS_208 0 -1.2023563682534940e-03
GC_3_209 b_3 NI_3 NS_209 0 5.3558155907298439e-06
GC_3_210 b_3 NI_3 NS_210 0 -6.7699487457956260e-05
GC_3_211 b_3 NI_3 NS_211 0 1.0049583684831394e-06
GC_3_212 b_3 NI_3 NS_212 0 1.7508605250485764e-07
GC_3_213 b_3 NI_3 NS_213 0 -8.6957305514603539e-06
GC_3_214 b_3 NI_3 NS_214 0 -2.5581890871166456e-06
GC_3_215 b_3 NI_3 NS_215 0 -1.7822793407318773e-05
GC_3_216 b_3 NI_3 NS_216 0 1.3447638870789946e-04
GC_3_217 b_3 NI_3 NS_217 0 -1.1934955497169143e-05
GC_3_218 b_3 NI_3 NS_218 0 -8.8811559122570617e-06
GC_3_219 b_3 NI_3 NS_219 0 -2.5113739551193155e-06
GC_3_220 b_3 NI_3 NS_220 0 2.8261283412666609e-06
GC_3_221 b_3 NI_3 NS_221 0 -1.0100739494328153e-05
GC_3_222 b_3 NI_3 NS_222 0 -3.2439834344379941e-05
GC_3_223 b_3 NI_3 NS_223 0 -3.6959740104510360e-06
GC_3_224 b_3 NI_3 NS_224 0 4.9034476039718582e-05
GC_3_225 b_3 NI_3 NS_225 0 3.4757877230650082e-02
GC_3_226 b_3 NI_3 NS_226 0 1.4285908315952319e-03
GC_3_227 b_3 NI_3 NS_227 0 5.8246829355908655e-03
GC_3_228 b_3 NI_3 NS_228 0 1.1407472833037606e-03
GC_3_229 b_3 NI_3 NS_229 0 -4.4989329353635867e-03
GC_3_230 b_3 NI_3 NS_230 0 -3.3622288087814772e-03
GC_3_231 b_3 NI_3 NS_231 0 4.1888735887330858e-03
GC_3_232 b_3 NI_3 NS_232 0 9.8493817124333319e-03
GC_3_233 b_3 NI_3 NS_233 0 4.6730983945938184e-04
GC_3_234 b_3 NI_3 NS_234 0 -4.9714329890041646e-03
GC_3_235 b_3 NI_3 NS_235 0 -3.4611869274358290e-04
GC_3_236 b_3 NI_3 NS_236 0 3.9560643956182033e-04
GC_3_237 b_3 NI_3 NS_237 0 9.6488309528016559e-03
GC_3_238 b_3 NI_3 NS_238 0 3.5231083082222416e-03
GC_3_239 b_3 NI_3 NS_239 0 5.3910614606901422e-04
GC_3_240 b_3 NI_3 NS_240 0 3.3158879071447981e-03
GC_3_241 b_3 NI_3 NS_241 0 2.4550411785967856e-03
GC_3_242 b_3 NI_3 NS_242 0 4.4743865182051996e-03
GC_3_243 b_3 NI_3 NS_243 0 3.0647654859360480e-03
GC_3_244 b_3 NI_3 NS_244 0 7.6251244386716412e-03
GC_3_245 b_3 NI_3 NS_245 0 4.3958183871922095e-04
GC_3_246 b_3 NI_3 NS_246 0 1.1146693101658695e-04
GC_3_247 b_3 NI_3 NS_247 0 -1.5839669244084531e-02
GC_3_248 b_3 NI_3 NS_248 0 1.3005523545575871e-02
GC_3_249 b_3 NI_3 NS_249 0 1.9133503178615026e-03
GC_3_250 b_3 NI_3 NS_250 0 3.9897100395983346e-04
GC_3_251 b_3 NI_3 NS_251 0 -7.3988404221788328e-04
GC_3_252 b_3 NI_3 NS_252 0 -4.3012283592819766e-07
GC_3_253 b_3 NI_3 NS_253 0 -4.0116847401071927e-04
GC_3_254 b_3 NI_3 NS_254 0 4.6161814261200072e-04
GC_3_255 b_3 NI_3 NS_255 0 -1.8700759973486810e-04
GC_3_256 b_3 NI_3 NS_256 0 4.4962329795653251e-05
GC_3_257 b_3 NI_3 NS_257 0 -8.4930949933743564e-03
GC_3_258 b_3 NI_3 NS_258 0 -1.1959306376013879e-02
GC_3_259 b_3 NI_3 NS_259 0 2.3586608241740509e-04
GC_3_260 b_3 NI_3 NS_260 0 -7.3130540341046835e-05
GC_3_261 b_3 NI_3 NS_261 0 -1.6032663930487250e-03
GC_3_262 b_3 NI_3 NS_262 0 3.5605087776995276e-03
GC_3_263 b_3 NI_3 NS_263 0 3.8194174490022068e-03
GC_3_264 b_3 NI_3 NS_264 0 -1.1618800347937897e-03
GC_3_265 b_3 NI_3 NS_265 0 9.7128552002293873e-05
GC_3_266 b_3 NI_3 NS_266 0 4.4580671647250739e-04
GC_3_267 b_3 NI_3 NS_267 0 -1.4552407116620744e-06
GC_3_268 b_3 NI_3 NS_268 0 3.2419541331391929e-06
GC_3_269 b_3 NI_3 NS_269 0 5.0113612610637621e-06
GC_3_270 b_3 NI_3 NS_270 0 -1.0945075609609469e-05
GC_3_271 b_3 NI_3 NS_271 0 -2.2221420917017915e-04
GC_3_272 b_3 NI_3 NS_272 0 -1.4552022294567150e-05
GC_3_273 b_3 NI_3 NS_273 0 1.6328445474129360e-05
GC_3_274 b_3 NI_3 NS_274 0 -1.8600795521781785e-05
GC_3_275 b_3 NI_3 NS_275 0 -8.0767790051587809e-06
GC_3_276 b_3 NI_3 NS_276 0 -9.2024029862440512e-06
GC_3_277 b_3 NI_3 NS_277 0 4.9664954267494876e-05
GC_3_278 b_3 NI_3 NS_278 0 -1.0182248542215168e-05
GC_3_279 b_3 NI_3 NS_279 0 -7.6913548773706179e-05
GC_3_280 b_3 NI_3 NS_280 0 -9.5243839755829584e-06
GC_3_281 b_3 NI_3 NS_281 0 2.6597972873215942e-02
GC_3_282 b_3 NI_3 NS_282 0 -8.3746175878945484e-04
GC_3_283 b_3 NI_3 NS_283 0 -1.8272418774958029e-03
GC_3_284 b_3 NI_3 NS_284 0 3.8984134861737249e-03
GC_3_285 b_3 NI_3 NS_285 0 1.0402788885113211e-03
GC_3_286 b_3 NI_3 NS_286 0 -3.2871410829277999e-04
GC_3_287 b_3 NI_3 NS_287 0 -9.8877834306809222e-03
GC_3_288 b_3 NI_3 NS_288 0 -3.7811999428766546e-03
GC_3_289 b_3 NI_3 NS_289 0 -1.5496381115098217e-03
GC_3_290 b_3 NI_3 NS_290 0 2.3303385167901280e-03
GC_3_291 b_3 NI_3 NS_291 0 -4.1464690174440317e-04
GC_3_292 b_3 NI_3 NS_292 0 -2.4631858878832199e-05
GC_3_293 b_3 NI_3 NS_293 0 5.6562834173204532e-03
GC_3_294 b_3 NI_3 NS_294 0 -6.1506372459033693e-03
GC_3_295 b_3 NI_3 NS_295 0 1.1720249732534778e-03
GC_3_296 b_3 NI_3 NS_296 0 1.7308458933911999e-03
GC_3_297 b_3 NI_3 NS_297 0 4.7278939376054597e-04
GC_3_298 b_3 NI_3 NS_298 0 1.8533894887272802e-03
GC_3_299 b_3 NI_3 NS_299 0 -5.0851002786971248e-03
GC_3_300 b_3 NI_3 NS_300 0 1.5509155084458820e-04
GC_3_301 b_3 NI_3 NS_301 0 -2.3040988039775857e-04
GC_3_302 b_3 NI_3 NS_302 0 -2.7503614060036473e-05
GC_3_303 b_3 NI_3 NS_303 0 2.4868171775528753e-03
GC_3_304 b_3 NI_3 NS_304 0 2.8878410974242166e-03
GC_3_305 b_3 NI_3 NS_305 0 -1.1638277521306849e-03
GC_3_306 b_3 NI_3 NS_306 0 -1.4323730973361825e-04
GC_3_307 b_3 NI_3 NS_307 0 -3.9402696983495487e-04
GC_3_308 b_3 NI_3 NS_308 0 6.4033254267303706e-05
GC_3_309 b_3 NI_3 NS_309 0 -5.7285674020434157e-04
GC_3_310 b_3 NI_3 NS_310 0 5.0309144512043552e-04
GC_3_311 b_3 NI_3 NS_311 0 -3.5340939021322420e-04
GC_3_312 b_3 NI_3 NS_312 0 -1.2701656279969981e-04
GC_3_313 b_3 NI_3 NS_313 0 -6.1998991962183164e-04
GC_3_314 b_3 NI_3 NS_314 0 -8.3127016708574764e-04
GC_3_315 b_3 NI_3 NS_315 0 -3.7576784601940825e-05
GC_3_316 b_3 NI_3 NS_316 0 1.6148703380101646e-04
GC_3_317 b_3 NI_3 NS_317 0 -7.1504344039869392e-04
GC_3_318 b_3 NI_3 NS_318 0 -5.5142715209372363e-04
GC_3_319 b_3 NI_3 NS_319 0 -1.0252926936737637e-03
GC_3_320 b_3 NI_3 NS_320 0 -9.6717133990087488e-04
GC_3_321 b_3 NI_3 NS_321 0 5.6909722820807386e-05
GC_3_322 b_3 NI_3 NS_322 0 -7.7398421222819964e-05
GC_3_323 b_3 NI_3 NS_323 0 1.4545001979756636e-06
GC_3_324 b_3 NI_3 NS_324 0 1.8107271753375866e-07
GC_3_325 b_3 NI_3 NS_325 0 -3.1829227494769057e-06
GC_3_326 b_3 NI_3 NS_326 0 4.6012058864385526e-06
GC_3_327 b_3 NI_3 NS_327 0 6.1819659496186583e-05
GC_3_328 b_3 NI_3 NS_328 0 1.3721932440267267e-05
GC_3_329 b_3 NI_3 NS_329 0 -5.1515587828730154e-06
GC_3_330 b_3 NI_3 NS_330 0 5.3360972907858041e-06
GC_3_331 b_3 NI_3 NS_331 0 1.0608991543826854e-06
GC_3_332 b_3 NI_3 NS_332 0 2.1639646630789377e-06
GC_3_333 b_3 NI_3 NS_333 0 -2.5173884000859833e-05
GC_3_334 b_3 NI_3 NS_334 0 -1.9972854348936507e-05
GC_3_335 b_3 NI_3 NS_335 0 2.2885449489045223e-05
GC_3_336 b_3 NI_3 NS_336 0 3.8354284660585508e-05
GC_3_337 b_3 NI_3 NS_337 0 3.8795067795002788e-02
GC_3_338 b_3 NI_3 NS_338 0 1.9750542861049323e-04
GC_3_339 b_3 NI_3 NS_339 0 5.2441381790848196e-03
GC_3_340 b_3 NI_3 NS_340 0 -5.0639849259763439e-05
GC_3_341 b_3 NI_3 NS_341 0 -3.8439901486909730e-03
GC_3_342 b_3 NI_3 NS_342 0 2.9963247926827505e-03
GC_3_343 b_3 NI_3 NS_343 0 -1.1812884697321769e-03
GC_3_344 b_3 NI_3 NS_344 0 7.1585111778294588e-03
GC_3_345 b_3 NI_3 NS_345 0 -8.4626749362280984e-03
GC_3_346 b_3 NI_3 NS_346 0 -5.6478453618081393e-03
GC_3_347 b_3 NI_3 NS_347 0 -1.6913173611875719e-04
GC_3_348 b_3 NI_3 NS_348 0 -1.8144928396313860e-04
GC_3_349 b_3 NI_3 NS_349 0 8.2792212334503075e-03
GC_3_350 b_3 NI_3 NS_350 0 5.1720878020746419e-04
GC_3_351 b_3 NI_3 NS_351 0 2.7691025390372850e-04
GC_3_352 b_3 NI_3 NS_352 0 2.3814244004106357e-03
GC_3_353 b_3 NI_3 NS_353 0 -7.2951634884542329e-04
GC_3_354 b_3 NI_3 NS_354 0 3.1567003907452275e-03
GC_3_355 b_3 NI_3 NS_355 0 6.1194599778338231e-04
GC_3_356 b_3 NI_3 NS_356 0 5.3578776252227543e-03
GC_3_357 b_3 NI_3 NS_357 0 3.3841060791704405e-04
GC_3_358 b_3 NI_3 NS_358 0 1.7577813560610734e-04
GC_3_359 b_3 NI_3 NS_359 0 -1.0819859358057420e-02
GC_3_360 b_3 NI_3 NS_360 0 5.3913820168369486e-03
GC_3_361 b_3 NI_3 NS_361 0 9.9973975282424557e-04
GC_3_362 b_3 NI_3 NS_362 0 4.5517616987643514e-04
GC_3_363 b_3 NI_3 NS_363 0 -5.4244451223299452e-04
GC_3_364 b_3 NI_3 NS_364 0 1.8787830252016255e-06
GC_3_365 b_3 NI_3 NS_365 0 -2.7958400500446352e-04
GC_3_366 b_3 NI_3 NS_366 0 2.1243215299784139e-04
GC_3_367 b_3 NI_3 NS_367 0 -1.3207582852796956e-04
GC_3_368 b_3 NI_3 NS_368 0 1.2753242153168290e-05
GC_3_369 b_3 NI_3 NS_369 0 -8.0524317465706079e-03
GC_3_370 b_3 NI_3 NS_370 0 -1.1297655016082316e-02
GC_3_371 b_3 NI_3 NS_371 0 1.4347883842292662e-04
GC_3_372 b_3 NI_3 NS_372 0 -4.5514726057740350e-05
GC_3_373 b_3 NI_3 NS_373 0 -1.1618775368565002e-03
GC_3_374 b_3 NI_3 NS_374 0 2.3711141662525921e-03
GC_3_375 b_3 NI_3 NS_375 0 6.1320464700326737e-03
GC_3_376 b_3 NI_3 NS_376 0 -2.1279855864912193e-04
GC_3_377 b_3 NI_3 NS_377 0 1.3792545076888270e-04
GC_3_378 b_3 NI_3 NS_378 0 3.3187763860133491e-04
GC_3_379 b_3 NI_3 NS_379 0 -2.2625934404591355e-08
GC_3_380 b_3 NI_3 NS_380 0 4.3694038747223382e-06
GC_3_381 b_3 NI_3 NS_381 0 4.1984813915330730e-06
GC_3_382 b_3 NI_3 NS_382 0 -1.9601858204853222e-05
GC_3_383 b_3 NI_3 NS_383 0 -3.6146939135683784e-04
GC_3_384 b_3 NI_3 NS_384 0 7.4582472429852981e-05
GC_3_385 b_3 NI_3 NS_385 0 1.8606664139765353e-05
GC_3_386 b_3 NI_3 NS_386 0 -3.6500753531034451e-05
GC_3_387 b_3 NI_3 NS_387 0 -2.0254702025635266e-05
GC_3_388 b_3 NI_3 NS_388 0 -1.2254882260356872e-05
GC_3_389 b_3 NI_3 NS_389 0 8.2425155540495791e-05
GC_3_390 b_3 NI_3 NS_390 0 -3.4698500511904721e-05
GC_3_391 b_3 NI_3 NS_391 0 -1.3711722737264393e-04
GC_3_392 b_3 NI_3 NS_392 0 1.1500336898388507e-05
GC_3_393 b_3 NI_3 NS_393 0 -4.7108844398448145e-03
GC_3_394 b_3 NI_3 NS_394 0 -2.7057613611155900e-04
GC_3_395 b_3 NI_3 NS_395 0 -1.2981495452321619e-03
GC_3_396 b_3 NI_3 NS_396 0 2.9646937939682683e-03
GC_3_397 b_3 NI_3 NS_397 0 -9.0101273618555032e-04
GC_3_398 b_3 NI_3 NS_398 0 -2.1585934591383687e-03
GC_3_399 b_3 NI_3 NS_399 0 -4.8241010355929287e-03
GC_3_400 b_3 NI_3 NS_400 0 -5.2327791563048136e-03
GC_3_401 b_3 NI_3 NS_401 0 6.6113530061491441e-03
GC_3_402 b_3 NI_3 NS_402 0 -1.2399264939440809e-03
GC_3_403 b_3 NI_3 NS_403 0 -2.7231652955136753e-04
GC_3_404 b_3 NI_3 NS_404 0 -5.8239358582231165e-05
GC_3_405 b_3 NI_3 NS_405 0 3.9896801950786457e-03
GC_3_406 b_3 NI_3 NS_406 0 -2.5678389338220373e-03
GC_3_407 b_3 NI_3 NS_407 0 7.3641777279544521e-04
GC_3_408 b_3 NI_3 NS_408 0 1.0236524976487396e-03
GC_3_409 b_3 NI_3 NS_409 0 7.3404456570473197e-04
GC_3_410 b_3 NI_3 NS_410 0 2.3515104468575612e-03
GC_3_411 b_3 NI_3 NS_411 0 -3.0485347367975070e-03
GC_3_412 b_3 NI_3 NS_412 0 1.0842577934819988e-03
GC_3_413 b_3 NI_3 NS_413 0 -1.9783189680260403e-04
GC_3_414 b_3 NI_3 NS_414 0 -8.6295389436529197e-06
GC_3_415 b_3 NI_3 NS_415 0 2.3282267874746403e-03
GC_3_416 b_3 NI_3 NS_416 0 5.7151092053750224e-04
GC_3_417 b_3 NI_3 NS_417 0 -7.9255932660393733e-04
GC_3_418 b_3 NI_3 NS_418 0 -1.0153501657718157e-04
GC_3_419 b_3 NI_3 NS_419 0 -2.7113352381981880e-04
GC_3_420 b_3 NI_3 NS_420 0 6.1973332087673886e-05
GC_3_421 b_3 NI_3 NS_421 0 -3.4873616518603070e-04
GC_3_422 b_3 NI_3 NS_422 0 1.9196022250090548e-04
GC_3_423 b_3 NI_3 NS_423 0 -1.6152454343237152e-04
GC_3_424 b_3 NI_3 NS_424 0 -1.0442915857269730e-04
GC_3_425 b_3 NI_3 NS_425 0 7.8243403052909979e-04
GC_3_426 b_3 NI_3 NS_426 0 -4.3737885597626414e-04
GC_3_427 b_3 NI_3 NS_427 0 -4.1987216208890414e-05
GC_3_428 b_3 NI_3 NS_428 0 8.3393285725222337e-05
GC_3_429 b_3 NI_3 NS_429 0 -2.9876630299329300e-04
GC_3_430 b_3 NI_3 NS_430 0 -6.1646384840924686e-04
GC_3_431 b_3 NI_3 NS_431 0 2.0354368494803518e-04
GC_3_432 b_3 NI_3 NS_432 0 9.6545422648546041e-04
GC_3_433 b_3 NI_3 NS_433 0 -3.6004383183062449e-06
GC_3_434 b_3 NI_3 NS_434 0 -1.0300740019429488e-04
GC_3_435 b_3 NI_3 NS_435 0 2.2385732610515298e-07
GC_3_436 b_3 NI_3 NS_436 0 -1.3347125162164964e-08
GC_3_437 b_3 NI_3 NS_437 0 7.6529026010712048e-07
GC_3_438 b_3 NI_3 NS_438 0 4.8152492440170139e-06
GC_3_439 b_3 NI_3 NS_439 0 3.3833487260309777e-05
GC_3_440 b_3 NI_3 NS_440 0 -6.0533840475386246e-05
GC_3_441 b_3 NI_3 NS_441 0 -2.4540247750453978e-07
GC_3_442 b_3 NI_3 NS_442 0 9.1689172100903894e-06
GC_3_443 b_3 NI_3 NS_443 0 1.7848319040101912e-06
GC_3_444 b_3 NI_3 NS_444 0 4.1267889077220437e-07
GC_3_445 b_3 NI_3 NS_445 0 -1.7052453410867674e-05
GC_3_446 b_3 NI_3 NS_446 0 -3.6587089270963734e-06
GC_3_447 b_3 NI_3 NS_447 0 2.0952939396638547e-05
GC_3_448 b_3 NI_3 NS_448 0 1.2817498122742270e-05
GC_3_449 b_3 NI_3 NS_449 0 1.1882631102780858e-02
GC_3_450 b_3 NI_3 NS_450 0 1.4764342989849902e-04
GC_3_451 b_3 NI_3 NS_451 0 -5.3398686662567910e-05
GC_3_452 b_3 NI_3 NS_452 0 -4.2102087572411988e-04
GC_3_453 b_3 NI_3 NS_453 0 3.8317487005423066e-04
GC_3_454 b_3 NI_3 NS_454 0 -3.7460189626749819e-05
GC_3_455 b_3 NI_3 NS_455 0 1.4796056176757100e-03
GC_3_456 b_3 NI_3 NS_456 0 -6.7680496528912035e-06
GC_3_457 b_3 NI_3 NS_457 0 7.6812323413465427e-04
GC_3_458 b_3 NI_3 NS_458 0 1.4996449982135540e-03
GC_3_459 b_3 NI_3 NS_459 0 -6.6989975854354000e-04
GC_3_460 b_3 NI_3 NS_460 0 2.0341095115855912e-04
GC_3_461 b_3 NI_3 NS_461 0 1.5028186362201917e-03
GC_3_462 b_3 NI_3 NS_462 0 -1.1499122455190084e-03
GC_3_463 b_3 NI_3 NS_463 0 1.8186828969274204e-03
GC_3_464 b_3 NI_3 NS_464 0 5.9667258851829440e-05
GC_3_465 b_3 NI_3 NS_465 0 8.4398209843193265e-05
GC_3_466 b_3 NI_3 NS_466 0 2.7198332830241402e-03
GC_3_467 b_3 NI_3 NS_467 0 2.9815000925612705e-03
GC_3_468 b_3 NI_3 NS_468 0 2.1941592177839638e-04
GC_3_469 b_3 NI_3 NS_469 0 6.0527599184169781e-04
GC_3_470 b_3 NI_3 NS_470 0 2.8814940486928390e-04
GC_3_471 b_3 NI_3 NS_471 0 -7.2197180976825632e-04
GC_3_472 b_3 NI_3 NS_472 0 1.1775135480006738e-02
GC_3_473 b_3 NI_3 NS_473 0 -8.4249396361382018e-04
GC_3_474 b_3 NI_3 NS_474 0 -1.0914240584630475e-03
GC_3_475 b_3 NI_3 NS_475 0 -1.3554585215737177e-03
GC_3_476 b_3 NI_3 NS_476 0 -1.1284117149359157e-05
GC_3_477 b_3 NI_3 NS_477 0 -5.1981516851475854e-04
GC_3_478 b_3 NI_3 NS_478 0 -4.4011104029983880e-04
GC_3_479 b_3 NI_3 NS_479 0 -1.3884847390338966e-04
GC_3_480 b_3 NI_3 NS_480 0 3.8054941467917635e-05
GC_3_481 b_3 NI_3 NS_481 0 -6.2717937525885942e-03
GC_3_482 b_3 NI_3 NS_482 0 -1.5195153023956527e-03
GC_3_483 b_3 NI_3 NS_483 0 3.3755317059853481e-05
GC_3_484 b_3 NI_3 NS_484 0 -4.5268963098559990e-05
GC_3_485 b_3 NI_3 NS_485 0 1.0857337631758424e-04
GC_3_486 b_3 NI_3 NS_486 0 7.5451808165084226e-04
GC_3_487 b_3 NI_3 NS_487 0 9.3791498969820054e-04
GC_3_488 b_3 NI_3 NS_488 0 -3.1098494944362593e-03
GC_3_489 b_3 NI_3 NS_489 0 1.9400010600651156e-05
GC_3_490 b_3 NI_3 NS_490 0 8.1218386609909838e-05
GC_3_491 b_3 NI_3 NS_491 0 -2.1435995809600158e-07
GC_3_492 b_3 NI_3 NS_492 0 1.4075854965984279e-06
GC_3_493 b_3 NI_3 NS_493 0 -1.6694584153746925e-06
GC_3_494 b_3 NI_3 NS_494 0 -9.7022253062420737e-06
GC_3_495 b_3 NI_3 NS_495 0 -1.2083548515373456e-04
GC_3_496 b_3 NI_3 NS_496 0 1.1974123843470761e-04
GC_3_497 b_3 NI_3 NS_497 0 1.1021616179792643e-06
GC_3_498 b_3 NI_3 NS_498 0 -2.0671068150217233e-05
GC_3_499 b_3 NI_3 NS_499 0 -1.5485134567425916e-05
GC_3_500 b_3 NI_3 NS_500 0 -4.9914990418652355e-06
GC_3_501 b_3 NI_3 NS_501 0 4.0908954193349478e-05
GC_3_502 b_3 NI_3 NS_502 0 -4.3805200845016154e-05
GC_3_503 b_3 NI_3 NS_503 0 -8.1823357208589306e-05
GC_3_504 b_3 NI_3 NS_504 0 4.5837541200951684e-05
GC_3_505 b_3 NI_3 NS_505 0 8.0622616758193755e-03
GC_3_506 b_3 NI_3 NS_506 0 -1.5147958968031347e-04
GC_3_507 b_3 NI_3 NS_507 0 3.0541915684610541e-04
GC_3_508 b_3 NI_3 NS_508 0 1.6335775894025058e-04
GC_3_509 b_3 NI_3 NS_509 0 -7.9987552418869212e-05
GC_3_510 b_3 NI_3 NS_510 0 3.3356406188108392e-04
GC_3_511 b_3 NI_3 NS_511 0 -9.2575855701806085e-04
GC_3_512 b_3 NI_3 NS_512 0 1.2090068577257826e-03
GC_3_513 b_3 NI_3 NS_513 0 -1.5895623139253023e-03
GC_3_514 b_3 NI_3 NS_514 0 -3.8700471426876337e-04
GC_3_515 b_3 NI_3 NS_515 0 1.1951301586369402e-04
GC_3_516 b_3 NI_3 NS_516 0 -3.3159016631971553e-04
GC_3_517 b_3 NI_3 NS_517 0 6.1336311602017984e-06
GC_3_518 b_3 NI_3 NS_518 0 -1.5464995924781321e-03
GC_3_519 b_3 NI_3 NS_519 0 9.7343882697028270e-04
GC_3_520 b_3 NI_3 NS_520 0 -6.1912788012133174e-04
GC_3_521 b_3 NI_3 NS_521 0 1.9281476701842007e-03
GC_3_522 b_3 NI_3 NS_522 0 1.8630683813450784e-03
GC_3_523 b_3 NI_3 NS_523 0 -4.4927500655998754e-04
GC_3_524 b_3 NI_3 NS_524 0 2.7060367652649926e-03
GC_3_525 b_3 NI_3 NS_525 0 -3.2995533555222055e-04
GC_3_526 b_3 NI_3 NS_526 0 -2.9811296601143056e-05
GC_3_527 b_3 NI_3 NS_527 0 -2.4211673695573991e-03
GC_3_528 b_3 NI_3 NS_528 0 2.7066650125625318e-03
GC_3_529 b_3 NI_3 NS_529 0 3.2268182754218024e-04
GC_3_530 b_3 NI_3 NS_530 0 3.1889536375258928e-04
GC_3_531 b_3 NI_3 NS_531 0 -1.0964657468361604e-03
GC_3_532 b_3 NI_3 NS_532 0 2.9468117661322500e-04
GC_3_533 b_3 NI_3 NS_533 0 -7.2148819670719128e-04
GC_3_534 b_3 NI_3 NS_534 0 -1.8717931940762171e-05
GC_3_535 b_3 NI_3 NS_535 0 -1.2988785710845664e-04
GC_3_536 b_3 NI_3 NS_536 0 -6.6050004640614817e-05
GC_3_537 b_3 NI_3 NS_537 0 -7.5857983995373211e-04
GC_3_538 b_3 NI_3 NS_538 0 -5.5940445553690089e-03
GC_3_539 b_3 NI_3 NS_539 0 5.8518715740415440e-05
GC_3_540 b_3 NI_3 NS_540 0 -3.8795707393095432e-05
GC_3_541 b_3 NI_3 NS_541 0 -1.2958630157918916e-03
GC_3_542 b_3 NI_3 NS_542 0 5.4380859927678998e-04
GC_3_543 b_3 NI_3 NS_543 0 1.5320740886254744e-03
GC_3_544 b_3 NI_3 NS_544 0 -6.5140497972946844e-05
GC_3_545 b_3 NI_3 NS_545 0 -1.4958657324575569e-04
GC_3_546 b_3 NI_3 NS_546 0 1.8029244868943386e-04
GC_3_547 b_3 NI_3 NS_547 0 -9.0707459757118283e-07
GC_3_548 b_3 NI_3 NS_548 0 4.2021229901586795e-07
GC_3_549 b_3 NI_3 NS_549 0 6.0058677843031992e-06
GC_3_550 b_3 NI_3 NS_550 0 -2.4411451994465545e-06
GC_3_551 b_3 NI_3 NS_551 0 -8.8381023001193486e-05
GC_3_552 b_3 NI_3 NS_552 0 -1.9622247307829556e-05
GC_3_553 b_3 NI_3 NS_553 0 1.3051385205854760e-05
GC_3_554 b_3 NI_3 NS_554 0 -6.5008808585741517e-06
GC_3_555 b_3 NI_3 NS_555 0 -4.8254306562479425e-06
GC_3_556 b_3 NI_3 NS_556 0 -5.1549035295303231e-06
GC_3_557 b_3 NI_3 NS_557 0 2.1021661776705647e-05
GC_3_558 b_3 NI_3 NS_558 0 -9.2628863186051368e-06
GC_3_559 b_3 NI_3 NS_559 0 -4.0870480982460701e-05
GC_3_560 b_3 NI_3 NS_560 0 1.2329322907518139e-06
GC_3_561 b_3 NI_3 NS_561 0 2.6865503605721174e-02
GC_3_562 b_3 NI_3 NS_562 0 -9.1147608017663412e-06
GC_3_563 b_3 NI_3 NS_563 0 7.2304462123803221e-04
GC_3_564 b_3 NI_3 NS_564 0 -6.2661469541228575e-04
GC_3_565 b_3 NI_3 NS_565 0 3.6818239143610108e-04
GC_3_566 b_3 NI_3 NS_566 0 1.0225473640243558e-03
GC_3_567 b_3 NI_3 NS_567 0 8.8921276972481591e-04
GC_3_568 b_3 NI_3 NS_568 0 2.2914004338157961e-03
GC_3_569 b_3 NI_3 NS_569 0 -2.2939181483884667e-03
GC_3_570 b_3 NI_3 NS_570 0 2.2457940546062915e-03
GC_3_571 b_3 NI_3 NS_571 0 -2.2456681869007783e-04
GC_3_572 b_3 NI_3 NS_572 0 1.5650219517208993e-04
GC_3_573 b_3 NI_3 NS_573 0 1.9356349081290874e-03
GC_3_574 b_3 NI_3 NS_574 0 -6.1778877852016422e-04
GC_3_575 b_3 NI_3 NS_575 0 1.3680151610096500e-03
GC_3_576 b_3 NI_3 NS_576 0 4.3539802342574044e-04
GC_3_577 b_3 NI_3 NS_577 0 -5.6560418246883479e-04
GC_3_578 b_3 NI_3 NS_578 0 3.9670545029505374e-03
GC_3_579 b_3 NI_3 NS_579 0 1.5711343398204230e-03
GC_3_580 b_3 NI_3 NS_580 0 1.9963452962697354e-03
GC_3_581 b_3 NI_3 NS_581 0 4.2452545424467527e-04
GC_3_582 b_3 NI_3 NS_582 0 2.6692915130683610e-04
GC_3_583 b_3 NI_3 NS_583 0 -4.6616642530292410e-03
GC_3_584 b_3 NI_3 NS_584 0 8.8629447378391468e-03
GC_3_585 b_3 NI_3 NS_585 0 -3.5175343472628574e-04
GC_3_586 b_3 NI_3 NS_586 0 -5.7005744886923671e-04
GC_3_587 b_3 NI_3 NS_587 0 -9.6580447283145846e-04
GC_3_588 b_3 NI_3 NS_588 0 4.9223777711217521e-05
GC_3_589 b_3 NI_3 NS_589 0 -4.5987323190145281e-04
GC_3_590 b_3 NI_3 NS_590 0 -1.3566619392528636e-04
GC_3_591 b_3 NI_3 NS_591 0 -1.5010314340278900e-04
GC_3_592 b_3 NI_3 NS_592 0 1.6853737736492646e-05
GC_3_593 b_3 NI_3 NS_593 0 -9.1781170042699763e-03
GC_3_594 b_3 NI_3 NS_594 0 -4.4385164887259044e-03
GC_3_595 b_3 NI_3 NS_595 0 4.8783912430632938e-05
GC_3_596 b_3 NI_3 NS_596 0 -6.2366839353456821e-05
GC_3_597 b_3 NI_3 NS_597 0 -1.2650838807188561e-04
GC_3_598 b_3 NI_3 NS_598 0 1.4402378597647243e-03
GC_3_599 b_3 NI_3 NS_599 0 3.7609136743046666e-03
GC_3_600 b_3 NI_3 NS_600 0 -4.1553736394126439e-03
GC_3_601 b_3 NI_3 NS_601 0 8.2575235934030791e-05
GC_3_602 b_3 NI_3 NS_602 0 3.0350562369069526e-04
GC_3_603 b_3 NI_3 NS_603 0 1.0518228281473313e-06
GC_3_604 b_3 NI_3 NS_604 0 3.7403128709402183e-06
GC_3_605 b_3 NI_3 NS_605 0 -2.3233031573927304e-06
GC_3_606 b_3 NI_3 NS_606 0 -1.6481915753630129e-05
GC_3_607 b_3 NI_3 NS_607 0 -2.4524358388571026e-04
GC_3_608 b_3 NI_3 NS_608 0 1.8847931204362046e-04
GC_3_609 b_3 NI_3 NS_609 0 4.3947344507322293e-06
GC_3_610 b_3 NI_3 NS_610 0 -3.5957957946230073e-05
GC_3_611 b_3 NI_3 NS_611 0 -2.5741989974368039e-05
GC_3_612 b_3 NI_3 NS_612 0 -6.6870901752615989e-06
GC_3_613 b_3 NI_3 NS_613 0 6.8713426889766731e-05
GC_3_614 b_3 NI_3 NS_614 0 -6.7102354468995073e-05
GC_3_615 b_3 NI_3 NS_615 0 -1.3336769739707931e-04
GC_3_616 b_3 NI_3 NS_616 0 6.7183059052034445e-05
GC_3_617 b_3 NI_3 NS_617 0 1.8343209445956577e-03
GC_3_618 b_3 NI_3 NS_618 0 -1.4045422862653644e-04
GC_3_619 b_3 NI_3 NS_619 0 1.7043545740904326e-04
GC_3_620 b_3 NI_3 NS_620 0 5.6335193925874296e-04
GC_3_621 b_3 NI_3 NS_621 0 -5.2540736870451319e-04
GC_3_622 b_3 NI_3 NS_622 0 -8.3983885507483046e-06
GC_3_623 b_3 NI_3 NS_623 0 -1.6439500113466048e-03
GC_3_624 b_3 NI_3 NS_624 0 -2.9679517304510329e-04
GC_3_625 b_3 NI_3 NS_625 0 6.6223652284030032e-04
GC_3_626 b_3 NI_3 NS_626 0 -1.9688513874594094e-03
GC_3_627 b_3 NI_3 NS_627 0 -1.9852777234227338e-04
GC_3_628 b_3 NI_3 NS_628 0 -2.6793605110241541e-04
GC_3_629 b_3 NI_3 NS_629 0 1.2415093807381272e-03
GC_3_630 b_3 NI_3 NS_630 0 -1.2282972748894707e-03
GC_3_631 b_3 NI_3 NS_631 0 7.4733383889136152e-04
GC_3_632 b_3 NI_3 NS_632 0 -2.2160304251822474e-04
GC_3_633 b_3 NI_3 NS_633 0 1.8707857116173673e-03
GC_3_634 b_3 NI_3 NS_634 0 2.0314576518510839e-03
GC_3_635 b_3 NI_3 NS_635 0 -4.3013844366037379e-04
GC_3_636 b_3 NI_3 NS_636 0 2.2303045855759955e-03
GC_3_637 b_3 NI_3 NS_637 0 -1.8781921884157340e-04
GC_3_638 b_3 NI_3 NS_638 0 -1.1098050345265320e-05
GC_3_639 b_3 NI_3 NS_639 0 -1.7978773910401560e-03
GC_3_640 b_3 NI_3 NS_640 0 1.9533684365708502e-03
GC_3_641 b_3 NI_3 NS_641 0 6.4382667788426295e-06
GC_3_642 b_3 NI_3 NS_642 0 2.4502003338131592e-04
GC_3_643 b_3 NI_3 NS_643 0 -6.4434296997726767e-04
GC_3_644 b_3 NI_3 NS_644 0 1.1840981343235214e-04
GC_3_645 b_3 NI_3 NS_645 0 -4.2460554636692543e-04
GC_3_646 b_3 NI_3 NS_646 0 2.4659134874611803e-05
GC_3_647 b_3 NI_3 NS_647 0 -9.2256356567707603e-05
GC_3_648 b_3 NI_3 NS_648 0 -5.5463596042368376e-05
GC_3_649 b_3 NI_3 NS_649 0 -7.9526760555186115e-04
GC_3_650 b_3 NI_3 NS_650 0 -3.2736039530614695e-03
GC_3_651 b_3 NI_3 NS_651 0 2.8720098436949133e-05
GC_3_652 b_3 NI_3 NS_652 0 -7.4296749632365476e-06
GC_3_653 b_3 NI_3 NS_653 0 -7.0063770688854449e-04
GC_3_654 b_3 NI_3 NS_654 0 2.4396799489524433e-04
GC_3_655 b_3 NI_3 NS_655 0 1.2436848992139202e-03
GC_3_656 b_3 NI_3 NS_656 0 -2.9690449212347475e-04
GC_3_657 b_3 NI_3 NS_657 0 -9.2697154098483021e-05
GC_3_658 b_3 NI_3 NS_658 0 1.2856424565508342e-04
GC_3_659 b_3 NI_3 NS_659 0 -1.9757713894089986e-07
GC_3_660 b_3 NI_3 NS_660 0 2.0347467125289411e-07
GC_3_661 b_3 NI_3 NS_661 0 2.7512744182652251e-06
GC_3_662 b_3 NI_3 NS_662 0 3.3178900145481107e-07
GC_3_663 b_3 NI_3 NS_663 0 -6.5912927937626059e-05
GC_3_664 b_3 NI_3 NS_664 0 -2.4386784367678006e-05
GC_3_665 b_3 NI_3 NS_665 0 6.1590259149054160e-06
GC_3_666 b_3 NI_3 NS_666 0 -7.4028698065730108e-07
GC_3_667 b_3 NI_3 NS_667 0 -3.7118713092084124e-06
GC_3_668 b_3 NI_3 NS_668 0 -9.2754915850706763e-07
GC_3_669 b_3 NI_3 NS_669 0 4.8541134545791483e-06
GC_3_670 b_3 NI_3 NS_670 0 -1.0376135443648932e-05
GC_3_671 b_3 NI_3 NS_671 0 -1.4136928671128219e-05
GC_3_672 b_3 NI_3 NS_672 0 1.1979204006423040e-05
GD_3_1 b_3 NI_3 NA_1 0 -1.7791070397795390e-04
GD_3_2 b_3 NI_3 NA_2 0 -5.8445864033957462e-02
GD_3_3 b_3 NI_3 NA_3 0 -1.4960139313291909e-01
GD_3_4 b_3 NI_3 NA_4 0 3.7780276852587447e-02
GD_3_5 b_3 NI_3 NA_5 0 -6.6182539289818057e-02
GD_3_6 b_3 NI_3 NA_6 0 -1.8764971022874888e-02
GD_3_7 b_3 NI_3 NA_7 0 -4.4479508840138758e-02
GD_3_8 b_3 NI_3 NA_8 0 3.0795733089736496e-03
GD_3_9 b_3 NI_3 NA_9 0 -2.0309520865165086e-02
GD_3_10 b_3 NI_3 NA_10 0 -3.4648378884948082e-03
GD_3_11 b_3 NI_3 NA_11 0 -3.1130932126012111e-02
GD_3_12 b_3 NI_3 NA_12 0 1.3438244043632161e-03
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 6.0535066632422030e-02
GC_4_2 b_4 NI_4 NS_2 0 -8.1708332951199887e-04
GC_4_3 b_4 NI_4 NS_3 0 -1.9120438285757468e-03
GC_4_4 b_4 NI_4 NS_4 0 2.2999153625501896e-03
GC_4_5 b_4 NI_4 NS_5 0 2.9401047194299330e-03
GC_4_6 b_4 NI_4 NS_6 0 1.1664003224815722e-04
GC_4_7 b_4 NI_4 NS_7 0 -4.9470419708676095e-03
GC_4_8 b_4 NI_4 NS_8 0 5.4589942198381050e-04
GC_4_9 b_4 NI_4 NS_9 0 -5.8274075655755479e-03
GC_4_10 b_4 NI_4 NS_10 0 1.1489937746496558e-02
GC_4_11 b_4 NI_4 NS_11 0 -5.6786859384979824e-04
GC_4_12 b_4 NI_4 NS_12 0 -1.0385963228499942e-04
GC_4_13 b_4 NI_4 NS_13 0 1.3568965921485132e-03
GC_4_14 b_4 NI_4 NS_14 0 -3.5525847751266566e-03
GC_4_15 b_4 NI_4 NS_15 0 7.0463864870206347e-04
GC_4_16 b_4 NI_4 NS_16 0 1.4367273921532847e-03
GC_4_17 b_4 NI_4 NS_17 0 -9.5147356303743882e-04
GC_4_18 b_4 NI_4 NS_18 0 1.0489586295451519e-03
GC_4_19 b_4 NI_4 NS_19 0 -5.9662103493495124e-03
GC_4_20 b_4 NI_4 NS_20 0 4.7372473498894543e-04
GC_4_21 b_4 NI_4 NS_21 0 -4.9267151388715360e-05
GC_4_22 b_4 NI_4 NS_22 0 -7.2311259961209588e-05
GC_4_23 b_4 NI_4 NS_23 0 3.0653951500463143e-04
GC_4_24 b_4 NI_4 NS_24 0 4.4832666209717051e-03
GC_4_25 b_4 NI_4 NS_25 0 -3.7029353569301349e-04
GC_4_26 b_4 NI_4 NS_26 0 -2.3078703100620589e-04
GC_4_27 b_4 NI_4 NS_27 0 -2.6502668606240450e-04
GC_4_28 b_4 NI_4 NS_28 0 -2.0110847216954681e-05
GC_4_29 b_4 NI_4 NS_29 0 -3.1761625275766062e-04
GC_4_30 b_4 NI_4 NS_30 0 3.4796407774779342e-04
GC_4_31 b_4 NI_4 NS_31 0 -1.9068453977069352e-04
GC_4_32 b_4 NI_4 NS_32 0 -3.0658727717170239e-05
GC_4_33 b_4 NI_4 NS_33 0 -6.4936291446599211e-03
GC_4_34 b_4 NI_4 NS_34 0 -1.2733897529683719e-03
GC_4_35 b_4 NI_4 NS_35 0 -1.1274157778021927e-05
GC_4_36 b_4 NI_4 NS_36 0 2.5829096361076741e-05
GC_4_37 b_4 NI_4 NS_37 0 -1.0252021384567813e-04
GC_4_38 b_4 NI_4 NS_38 0 7.0577862335170273e-04
GC_4_39 b_4 NI_4 NS_39 0 -6.8789583060646598e-04
GC_4_40 b_4 NI_4 NS_40 0 -2.1624420222088308e-03
GC_4_41 b_4 NI_4 NS_41 0 1.8350642472152873e-04
GC_4_42 b_4 NI_4 NS_42 0 8.9580574777718916e-05
GC_4_43 b_4 NI_4 NS_43 0 3.4689152015806927e-06
GC_4_44 b_4 NI_4 NS_44 0 2.7662353648002071e-06
GC_4_45 b_4 NI_4 NS_45 0 -6.0387414024006249e-06
GC_4_46 b_4 NI_4 NS_46 0 -1.1214784910998217e-05
GC_4_47 b_4 NI_4 NS_47 0 -5.9285862572674643e-05
GC_4_48 b_4 NI_4 NS_48 0 2.0581797754306357e-04
GC_4_49 b_4 NI_4 NS_49 0 -1.3231783038386167e-05
GC_4_50 b_4 NI_4 NS_50 0 -2.6512655682282608e-05
GC_4_51 b_4 NI_4 NS_51 0 -6.9061028904662450e-06
GC_4_52 b_4 NI_4 NS_52 0 9.9048500586323090e-06
GC_4_53 b_4 NI_4 NS_53 0 -9.5811569449009182e-06
GC_4_54 b_4 NI_4 NS_54 0 -4.8954932939067253e-05
GC_4_55 b_4 NI_4 NS_55 0 -1.0044599841755782e-05
GC_4_56 b_4 NI_4 NS_56 0 7.9771044770588189e-05
GC_4_57 b_4 NI_4 NS_57 0 -1.2798903194289640e-02
GC_4_58 b_4 NI_4 NS_58 0 -1.3735151895689769e-03
GC_4_59 b_4 NI_4 NS_59 0 -7.7962845981644998e-04
GC_4_60 b_4 NI_4 NS_60 0 -1.0572048332984385e-03
GC_4_61 b_4 NI_4 NS_61 0 -1.1036283190314316e-03
GC_4_62 b_4 NI_4 NS_62 0 1.5093200932895336e-03
GC_4_63 b_4 NI_4 NS_63 0 7.0972612306895654e-04
GC_4_64 b_4 NI_4 NS_64 0 -2.1293394780094906e-04
GC_4_65 b_4 NI_4 NS_65 0 -3.8917604739517656e-03
GC_4_66 b_4 NI_4 NS_66 0 -8.6536570789324738e-03
GC_4_67 b_4 NI_4 NS_67 0 8.6157430512906515e-05
GC_4_68 b_4 NI_4 NS_68 0 2.5385781239928525e-05
GC_4_69 b_4 NI_4 NS_69 0 2.1257436803667346e-03
GC_4_70 b_4 NI_4 NS_70 0 -2.2730706406085704e-03
GC_4_71 b_4 NI_4 NS_71 0 6.7197057485488692e-04
GC_4_72 b_4 NI_4 NS_72 0 3.0585337893505009e-04
GC_4_73 b_4 NI_4 NS_73 0 7.3461482351343049e-04
GC_4_74 b_4 NI_4 NS_74 0 -2.0411679363497529e-03
GC_4_75 b_4 NI_4 NS_75 0 1.4968514691151462e-03
GC_4_76 b_4 NI_4 NS_76 0 -2.0038818705840891e-03
GC_4_77 b_4 NI_4 NS_77 0 7.7292631871702437e-06
GC_4_78 b_4 NI_4 NS_78 0 2.0772088151994810e-06
GC_4_79 b_4 NI_4 NS_79 0 6.7007287899427401e-03
GC_4_80 b_4 NI_4 NS_80 0 1.4714120732037699e-03
GC_4_81 b_4 NI_4 NS_81 0 -6.0566693759215009e-05
GC_4_82 b_4 NI_4 NS_82 0 2.0744099581541182e-07
GC_4_83 b_4 NI_4 NS_83 0 -3.0959080065209738e-05
GC_4_84 b_4 NI_4 NS_84 0 4.5355675119951732e-05
GC_4_85 b_4 NI_4 NS_85 0 2.4627682350181407e-04
GC_4_86 b_4 NI_4 NS_86 0 -2.2727999067512024e-04
GC_4_87 b_4 NI_4 NS_87 0 2.9855239985695202e-04
GC_4_88 b_4 NI_4 NS_88 0 -7.5248850481228610e-05
GC_4_89 b_4 NI_4 NS_89 0 -8.5166146043975169e-03
GC_4_90 b_4 NI_4 NS_90 0 2.5929244226529031e-03
GC_4_91 b_4 NI_4 NS_91 0 -1.8240805603949168e-04
GC_4_92 b_4 NI_4 NS_92 0 -2.0481532344429509e-04
GC_4_93 b_4 NI_4 NS_93 0 3.4833247209234801e-03
GC_4_94 b_4 NI_4 NS_94 0 7.8743780957288387e-04
GC_4_95 b_4 NI_4 NS_95 0 2.8067326936751708e-03
GC_4_96 b_4 NI_4 NS_96 0 -1.3090522347969148e-03
GC_4_97 b_4 NI_4 NS_97 0 8.0134483786074178e-04
GC_4_98 b_4 NI_4 NS_98 0 1.4275697876488572e-04
GC_4_99 b_4 NI_4 NS_99 0 -1.8181429149290391e-06
GC_4_100 b_4 NI_4 NS_100 0 -2.7381198883037547e-06
GC_4_101 b_4 NI_4 NS_101 0 -1.8801006871483680e-05
GC_4_102 b_4 NI_4 NS_102 0 -1.8315029431109391e-05
GC_4_103 b_4 NI_4 NS_103 0 -8.3260898781884976e-05
GC_4_104 b_4 NI_4 NS_104 0 -4.4662709254962294e-06
GC_4_105 b_4 NI_4 NS_105 0 -3.3079741706843695e-05
GC_4_106 b_4 NI_4 NS_106 0 -1.3760385736931465e-05
GC_4_107 b_4 NI_4 NS_107 0 -1.5576296403285581e-05
GC_4_108 b_4 NI_4 NS_108 0 -1.0832312980421589e-05
GC_4_109 b_4 NI_4 NS_109 0 1.8926518007387826e-04
GC_4_110 b_4 NI_4 NS_110 0 -9.7087313836421803e-05
GC_4_111 b_4 NI_4 NS_111 0 -3.0963968265408496e-04
GC_4_112 b_4 NI_4 NS_112 0 5.9902708952928864e-05
GC_4_113 b_4 NI_4 NS_113 0 -3.9239711967164234e-02
GC_4_114 b_4 NI_4 NS_114 0 1.1912590977745536e-02
GC_4_115 b_4 NI_4 NS_115 0 -2.9631647745848345e-03
GC_4_116 b_4 NI_4 NS_116 0 3.8370699507880492e-03
GC_4_117 b_4 NI_4 NS_117 0 -4.5209998938927276e-03
GC_4_118 b_4 NI_4 NS_118 0 2.0762529289838688e-03
GC_4_119 b_4 NI_4 NS_119 0 -4.6100700842439373e-03
GC_4_120 b_4 NI_4 NS_120 0 -9.0087771136988081e-03
GC_4_121 b_4 NI_4 NS_121 0 -2.2016986909285199e-03
GC_4_122 b_4 NI_4 NS_122 0 -8.6781035757144947e-03
GC_4_123 b_4 NI_4 NS_123 0 7.2684118588306804e-04
GC_4_124 b_4 NI_4 NS_124 0 -1.4323299987784014e-04
GC_4_125 b_4 NI_4 NS_125 0 6.8572941190363796e-03
GC_4_126 b_4 NI_4 NS_126 0 -5.0622900790650409e-04
GC_4_127 b_4 NI_4 NS_127 0 1.2644404686545639e-03
GC_4_128 b_4 NI_4 NS_128 0 1.4479564218829843e-03
GC_4_129 b_4 NI_4 NS_129 0 4.3732778280137878e-03
GC_4_130 b_4 NI_4 NS_130 0 1.6167447990951408e-03
GC_4_131 b_4 NI_4 NS_131 0 -2.2047009088198657e-03
GC_4_132 b_4 NI_4 NS_132 0 9.4748631449664681e-04
GC_4_133 b_4 NI_4 NS_133 0 -2.4089088171214276e-04
GC_4_134 b_4 NI_4 NS_134 0 2.9282183122564554e-06
GC_4_135 b_4 NI_4 NS_135 0 5.3978745791590857e-03
GC_4_136 b_4 NI_4 NS_136 0 -2.1314084227576900e-03
GC_4_137 b_4 NI_4 NS_137 0 -1.2310588939639206e-03
GC_4_138 b_4 NI_4 NS_138 0 -2.2056253294829278e-04
GC_4_139 b_4 NI_4 NS_139 0 -1.7998280294215973e-04
GC_4_140 b_4 NI_4 NS_140 0 2.3497368635751690e-05
GC_4_141 b_4 NI_4 NS_141 0 -4.1235200157240019e-04
GC_4_142 b_4 NI_4 NS_142 0 2.8860449762683929e-04
GC_4_143 b_4 NI_4 NS_143 0 -2.2729731722027062e-04
GC_4_144 b_4 NI_4 NS_144 0 -1.2617695839986352e-04
GC_4_145 b_4 NI_4 NS_145 0 1.0266668770185471e-03
GC_4_146 b_4 NI_4 NS_146 0 -1.6449325450880329e-04
GC_4_147 b_4 NI_4 NS_147 0 -4.2568704220304923e-05
GC_4_148 b_4 NI_4 NS_148 0 1.2650722765244601e-04
GC_4_149 b_4 NI_4 NS_149 0 -5.3924316988157128e-04
GC_4_150 b_4 NI_4 NS_150 0 -7.0337230304131672e-04
GC_4_151 b_4 NI_4 NS_151 0 2.7149552122351294e-03
GC_4_152 b_4 NI_4 NS_152 0 -1.2023563682492307e-03
GC_4_153 b_4 NI_4 NS_153 0 5.3558155904755019e-06
GC_4_154 b_4 NI_4 NS_154 0 -6.7699487458003802e-05
GC_4_155 b_4 NI_4 NS_155 0 1.0049583684796537e-06
GC_4_156 b_4 NI_4 NS_156 0 1.7508605250424508e-07
GC_4_157 b_4 NI_4 NS_157 0 -8.6957305514440790e-06
GC_4_158 b_4 NI_4 NS_158 0 -2.5581890871147630e-06
GC_4_159 b_4 NI_4 NS_159 0 -1.7822793407443345e-05
GC_4_160 b_4 NI_4 NS_160 0 1.3447638870765777e-04
GC_4_161 b_4 NI_4 NS_161 0 -1.1934955497138982e-05
GC_4_162 b_4 NI_4 NS_162 0 -8.8811559122492046e-06
GC_4_163 b_4 NI_4 NS_163 0 -2.5113739551108981e-06
GC_4_164 b_4 NI_4 NS_164 0 2.8261283412485171e-06
GC_4_165 b_4 NI_4 NS_165 0 -1.0100739494280852e-05
GC_4_166 b_4 NI_4 NS_166 0 -3.2439834344324457e-05
GC_4_167 b_4 NI_4 NS_167 0 -3.6959740104947704e-06
GC_4_168 b_4 NI_4 NS_168 0 4.9034476039613590e-05
GC_4_169 b_4 NI_4 NS_169 0 -6.0818432819240043e-02
GC_4_170 b_4 NI_4 NS_170 0 7.5807118575123428e-03
GC_4_171 b_4 NI_4 NS_171 0 -9.8091228911859063e-04
GC_4_172 b_4 NI_4 NS_172 0 -2.0294191659633852e-03
GC_4_173 b_4 NI_4 NS_173 0 2.4005451058554895e-04
GC_4_174 b_4 NI_4 NS_174 0 -1.4488913961279112e-03
GC_4_175 b_4 NI_4 NS_175 0 5.8552229702910049e-03
GC_4_176 b_4 NI_4 NS_176 0 4.6818704388598992e-03
GC_4_177 b_4 NI_4 NS_177 0 3.2519505645615125e-03
GC_4_178 b_4 NI_4 NS_178 0 7.6747495563929593e-03
GC_4_179 b_4 NI_4 NS_179 0 4.1950978996390965e-04
GC_4_180 b_4 NI_4 NS_180 0 -5.5380253428973685e-04
GC_4_181 b_4 NI_4 NS_181 0 -1.5857941757957824e-03
GC_4_182 b_4 NI_4 NS_182 0 -4.7820897565462881e-03
GC_4_183 b_4 NI_4 NS_183 0 8.7936987609945033e-04
GC_4_184 b_4 NI_4 NS_184 0 7.3538508584163010e-04
GC_4_185 b_4 NI_4 NS_185 0 -3.7702003859717063e-05
GC_4_186 b_4 NI_4 NS_186 0 1.2505451594484944e-03
GC_4_187 b_4 NI_4 NS_187 0 2.1544852266436633e-03
GC_4_188 b_4 NI_4 NS_188 0 -1.7211664957633083e-03
GC_4_189 b_4 NI_4 NS_189 0 7.5761862631838474e-05
GC_4_190 b_4 NI_4 NS_190 0 -7.2013779600476938e-05
GC_4_191 b_4 NI_4 NS_191 0 -3.6572228129933058e-04
GC_4_192 b_4 NI_4 NS_192 0 5.8773739282680032e-03
GC_4_193 b_4 NI_4 NS_193 0 3.7425992133361421e-04
GC_4_194 b_4 NI_4 NS_194 0 -8.8468399123390581e-05
GC_4_195 b_4 NI_4 NS_195 0 -2.9595758259527065e-04
GC_4_196 b_4 NI_4 NS_196 0 8.4649971156855606e-06
GC_4_197 b_4 NI_4 NS_197 0 1.6864720608622189e-04
GC_4_198 b_4 NI_4 NS_198 0 5.1596647535398090e-05
GC_4_199 b_4 NI_4 NS_199 0 2.3074272175940889e-04
GC_4_200 b_4 NI_4 NS_200 0 2.1179152119868600e-05
GC_4_201 b_4 NI_4 NS_201 0 -1.5670645308070181e-02
GC_4_202 b_4 NI_4 NS_202 0 5.5070763462703538e-05
GC_4_203 b_4 NI_4 NS_203 0 -1.2232371087629335e-04
GC_4_204 b_4 NI_4 NS_204 0 -2.9338052622987477e-04
GC_4_205 b_4 NI_4 NS_205 0 3.6041695465826302e-03
GC_4_206 b_4 NI_4 NS_206 0 2.6869019027340115e-03
GC_4_207 b_4 NI_4 NS_207 0 5.2228650763106350e-03
GC_4_208 b_4 NI_4 NS_208 0 -4.7087506325030502e-03
GC_4_209 b_4 NI_4 NS_209 0 1.0073459075107840e-03
GC_4_210 b_4 NI_4 NS_210 0 4.6760000054408348e-04
GC_4_211 b_4 NI_4 NS_211 0 -5.2107294566976143e-07
GC_4_212 b_4 NI_4 NS_212 0 2.8267133927803731e-07
GC_4_213 b_4 NI_4 NS_213 0 -2.3463638791729242e-05
GC_4_214 b_4 NI_4 NS_214 0 -2.9841307406882994e-05
GC_4_215 b_4 NI_4 NS_215 0 -1.9304958890799937e-04
GC_4_216 b_4 NI_4 NS_216 0 1.9972681376553879e-04
GC_4_217 b_4 NI_4 NS_217 0 -3.8427502397604370e-05
GC_4_218 b_4 NI_4 NS_218 0 -4.0874776374536988e-05
GC_4_219 b_4 NI_4 NS_219 0 -3.4843707435899823e-05
GC_4_220 b_4 NI_4 NS_220 0 -8.6530495471663253e-06
GC_4_221 b_4 NI_4 NS_221 0 2.2545845373708341e-04
GC_4_222 b_4 NI_4 NS_222 0 -1.4606603983484301e-04
GC_4_223 b_4 NI_4 NS_223 0 -3.8771615367328203e-04
GC_4_224 b_4 NI_4 NS_224 0 1.1466486548714784e-04
GC_4_225 b_4 NI_4 NS_225 0 2.6989211300671719e-02
GC_4_226 b_4 NI_4 NS_226 0 -8.4386319150217331e-04
GC_4_227 b_4 NI_4 NS_227 0 -1.9460633039185076e-03
GC_4_228 b_4 NI_4 NS_228 0 3.7443949577555757e-03
GC_4_229 b_4 NI_4 NS_229 0 1.0569242403267122e-03
GC_4_230 b_4 NI_4 NS_230 0 -3.7916553289240511e-04
GC_4_231 b_4 NI_4 NS_231 0 -9.3446228957584816e-03
GC_4_232 b_4 NI_4 NS_232 0 -3.7940206932798896e-03
GC_4_233 b_4 NI_4 NS_233 0 -1.3066320561323161e-03
GC_4_234 b_4 NI_4 NS_234 0 2.7861828183319108e-03
GC_4_235 b_4 NI_4 NS_235 0 -2.9107677086610232e-04
GC_4_236 b_4 NI_4 NS_236 0 2.3487895642100836e-04
GC_4_237 b_4 NI_4 NS_237 0 5.2061840433455832e-03
GC_4_238 b_4 NI_4 NS_238 0 -5.5271193144066037e-03
GC_4_239 b_4 NI_4 NS_239 0 8.5166089350641747e-04
GC_4_240 b_4 NI_4 NS_240 0 1.5028430640703493e-03
GC_4_241 b_4 NI_4 NS_241 0 2.8189484599622320e-04
GC_4_242 b_4 NI_4 NS_242 0 1.3819754804295507e-03
GC_4_243 b_4 NI_4 NS_243 0 -4.8241587449047206e-03
GC_4_244 b_4 NI_4 NS_244 0 -1.6647652561091448e-04
GC_4_245 b_4 NI_4 NS_245 0 -1.8588142242706166e-04
GC_4_246 b_4 NI_4 NS_246 0 -4.5725509494538588e-06
GC_4_247 b_4 NI_4 NS_247 0 2.1097177417264855e-03
GC_4_248 b_4 NI_4 NS_248 0 1.9641640314517223e-03
GC_4_249 b_4 NI_4 NS_249 0 -9.6364450439150214e-04
GC_4_250 b_4 NI_4 NS_250 0 -1.4031939445820899e-04
GC_4_251 b_4 NI_4 NS_251 0 -2.4112531614903606e-04
GC_4_252 b_4 NI_4 NS_252 0 -8.4638617697790332e-06
GC_4_253 b_4 NI_4 NS_253 0 -4.1669281871319964e-04
GC_4_254 b_4 NI_4 NS_254 0 3.2033563921056983e-04
GC_4_255 b_4 NI_4 NS_255 0 -2.1999514476167892e-04
GC_4_256 b_4 NI_4 NS_256 0 -9.5169664529578225e-05
GC_4_257 b_4 NI_4 NS_257 0 8.3068316000220704e-04
GC_4_258 b_4 NI_4 NS_258 0 -4.0393455624720070e-04
GC_4_259 b_4 NI_4 NS_259 0 -1.7883384735859075e-05
GC_4_260 b_4 NI_4 NS_260 0 1.0993220563713222e-04
GC_4_261 b_4 NI_4 NS_261 0 -5.5298481693346040e-04
GC_4_262 b_4 NI_4 NS_262 0 -4.2752852314276852e-04
GC_4_263 b_4 NI_4 NS_263 0 -2.0470058215678330e-03
GC_4_264 b_4 NI_4 NS_264 0 1.3332881979306708e-04
GC_4_265 b_4 NI_4 NS_265 0 -2.9643042164940427e-05
GC_4_266 b_4 NI_4 NS_266 0 -3.3649383177491123e-05
GC_4_267 b_4 NI_4 NS_267 0 1.3157909568518273e-06
GC_4_268 b_4 NI_4 NS_268 0 -9.2372066177586760e-07
GC_4_269 b_4 NI_4 NS_269 0 1.1669231170803827e-06
GC_4_270 b_4 NI_4 NS_270 0 1.8590746820232203e-06
GC_4_271 b_4 NI_4 NS_271 0 6.5307997702787902e-05
GC_4_272 b_4 NI_4 NS_272 0 -3.7685260909283676e-05
GC_4_273 b_4 NI_4 NS_273 0 -4.5025443450322969e-08
GC_4_274 b_4 NI_4 NS_274 0 7.2192038472186848e-06
GC_4_275 b_4 NI_4 NS_275 0 -8.0829895935449439e-07
GC_4_276 b_4 NI_4 NS_276 0 -6.0596552944332953e-07
GC_4_277 b_4 NI_4 NS_277 0 -7.8439897250440056e-06
GC_4_278 b_4 NI_4 NS_278 0 1.8834634144447677e-05
GC_4_279 b_4 NI_4 NS_279 0 2.1496455210599123e-05
GC_4_280 b_4 NI_4 NS_280 0 -2.4033905025388407e-05
GC_4_281 b_4 NI_4 NS_281 0 5.2611173122921002e-03
GC_4_282 b_4 NI_4 NS_282 0 -1.4446755189497684e-03
GC_4_283 b_4 NI_4 NS_283 0 -1.5058079172478396e-03
GC_4_284 b_4 NI_4 NS_284 0 -1.4352623017341456e-03
GC_4_285 b_4 NI_4 NS_285 0 -3.9263870268734413e-04
GC_4_286 b_4 NI_4 NS_286 0 8.0826351442799145e-04
GC_4_287 b_4 NI_4 NS_287 0 4.7945383371956109e-03
GC_4_288 b_4 NI_4 NS_288 0 -4.7617583962850313e-04
GC_4_289 b_4 NI_4 NS_289 0 -3.9753895549588282e-03
GC_4_290 b_4 NI_4 NS_290 0 -1.7587520754782048e-03
GC_4_291 b_4 NI_4 NS_291 0 -1.3886792395549136e-04
GC_4_292 b_4 NI_4 NS_292 0 7.2685637820118392e-04
GC_4_293 b_4 NI_4 NS_293 0 9.1338579209485331e-04
GC_4_294 b_4 NI_4 NS_294 0 -2.7491081364170744e-03
GC_4_295 b_4 NI_4 NS_295 0 1.0979251236178530e-03
GC_4_296 b_4 NI_4 NS_296 0 6.0131867554932394e-04
GC_4_297 b_4 NI_4 NS_297 0 9.0939266746785830e-04
GC_4_298 b_4 NI_4 NS_298 0 1.1361251319690485e-03
GC_4_299 b_4 NI_4 NS_299 0 1.7045646241894263e-03
GC_4_300 b_4 NI_4 NS_300 0 -2.4860657744305366e-03
GC_4_301 b_4 NI_4 NS_301 0 9.7859251360283132e-05
GC_4_302 b_4 NI_4 NS_302 0 -5.8372778425798439e-05
GC_4_303 b_4 NI_4 NS_303 0 3.5051835049586329e-03
GC_4_304 b_4 NI_4 NS_304 0 5.0803000828476249e-03
GC_4_305 b_4 NI_4 NS_305 0 3.3688937898242118e-04
GC_4_306 b_4 NI_4 NS_306 0 -1.5566461414926015e-05
GC_4_307 b_4 NI_4 NS_307 0 -2.3857886335985602e-04
GC_4_308 b_4 NI_4 NS_308 0 -1.6350139988313338e-07
GC_4_309 b_4 NI_4 NS_309 0 1.9882301834672457e-04
GC_4_310 b_4 NI_4 NS_310 0 -1.9992883678419224e-04
GC_4_311 b_4 NI_4 NS_311 0 3.6454801651638686e-04
GC_4_312 b_4 NI_4 NS_312 0 -9.7169942370181568e-05
GC_4_313 b_4 NI_4 NS_313 0 -1.5278548446068328e-02
GC_4_314 b_4 NI_4 NS_314 0 1.8372239903463388e-03
GC_4_315 b_4 NI_4 NS_315 0 -2.2191141534569104e-04
GC_4_316 b_4 NI_4 NS_316 0 -3.1094019685639734e-04
GC_4_317 b_4 NI_4 NS_317 0 4.7744086698169484e-03
GC_4_318 b_4 NI_4 NS_318 0 1.9067385497154917e-03
GC_4_319 b_4 NI_4 NS_319 0 5.4014192378234634e-03
GC_4_320 b_4 NI_4 NS_320 0 -4.1644053390029198e-03
GC_4_321 b_4 NI_4 NS_321 0 1.1613846415988798e-03
GC_4_322 b_4 NI_4 NS_322 0 3.7782698335559850e-04
GC_4_323 b_4 NI_4 NS_323 0 -3.3728978004524926e-06
GC_4_324 b_4 NI_4 NS_324 0 -2.8875224737229977e-06
GC_4_325 b_4 NI_4 NS_325 0 -3.7912087523905887e-05
GC_4_326 b_4 NI_4 NS_326 0 -3.3743935094596988e-05
GC_4_327 b_4 NI_4 NS_327 0 -2.3296012894842165e-04
GC_4_328 b_4 NI_4 NS_328 0 2.1070988092929390e-04
GC_4_329 b_4 NI_4 NS_329 0 -5.5623602755961638e-05
GC_4_330 b_4 NI_4 NS_330 0 -4.1523025595019690e-05
GC_4_331 b_4 NI_4 NS_331 0 -3.6381468076481535e-05
GC_4_332 b_4 NI_4 NS_332 0 -1.2374187497504261e-05
GC_4_333 b_4 NI_4 NS_333 0 2.9572101839388969e-04
GC_4_334 b_4 NI_4 NS_334 0 -2.2809499656839476e-04
GC_4_335 b_4 NI_4 NS_335 0 -5.2276230576959624e-04
GC_4_336 b_4 NI_4 NS_336 0 1.9857930666267846e-04
GC_4_337 b_4 NI_4 NS_337 0 -8.2280834145474074e-03
GC_4_338 b_4 NI_4 NS_338 0 -2.3837370115162415e-04
GC_4_339 b_4 NI_4 NS_339 0 -1.3510034806756791e-03
GC_4_340 b_4 NI_4 NS_340 0 2.9662468753485246e-03
GC_4_341 b_4 NI_4 NS_341 0 -9.2138232963093235e-04
GC_4_342 b_4 NI_4 NS_342 0 -2.2289397577293199e-03
GC_4_343 b_4 NI_4 NS_343 0 -4.8028512757119736e-03
GC_4_344 b_4 NI_4 NS_344 0 -5.4465581545350434e-03
GC_4_345 b_4 NI_4 NS_345 0 6.6780373885698225e-03
GC_4_346 b_4 NI_4 NS_346 0 -1.5237086673317920e-03
GC_4_347 b_4 NI_4 NS_347 0 1.6747671394367507e-04
GC_4_348 b_4 NI_4 NS_348 0 -3.0856848388568779e-05
GC_4_349 b_4 NI_4 NS_349 0 4.0263033397165242e-03
GC_4_350 b_4 NI_4 NS_350 0 -2.6519574755887450e-03
GC_4_351 b_4 NI_4 NS_351 0 6.9140887688245458e-04
GC_4_352 b_4 NI_4 NS_352 0 1.0151562673964862e-03
GC_4_353 b_4 NI_4 NS_353 0 7.1352989709989076e-04
GC_4_354 b_4 NI_4 NS_354 0 2.1040188619612823e-03
GC_4_355 b_4 NI_4 NS_355 0 -3.0951634400905367e-03
GC_4_356 b_4 NI_4 NS_356 0 8.4633238507211155e-04
GC_4_357 b_4 NI_4 NS_357 0 -1.9656287550763439e-04
GC_4_358 b_4 NI_4 NS_358 0 -3.6504364565889678e-06
GC_4_359 b_4 NI_4 NS_359 0 2.5992903858759629e-03
GC_4_360 b_4 NI_4 NS_360 0 5.4805897875661029e-05
GC_4_361 b_4 NI_4 NS_361 0 -7.9285856059737550e-04
GC_4_362 b_4 NI_4 NS_362 0 -1.2485858719580637e-04
GC_4_363 b_4 NI_4 NS_363 0 -2.1064989308783221e-04
GC_4_364 b_4 NI_4 NS_364 0 5.0355621137772227e-05
GC_4_365 b_4 NI_4 NS_365 0 -2.6612980420952378e-04
GC_4_366 b_4 NI_4 NS_366 0 1.3769874454962552e-04
GC_4_367 b_4 NI_4 NS_367 0 -1.2376747751925138e-04
GC_4_368 b_4 NI_4 NS_368 0 -8.5167744465394895e-05
GC_4_369 b_4 NI_4 NS_369 0 7.8164186086159318e-04
GC_4_370 b_4 NI_4 NS_370 0 -7.9134408292500327e-04
GC_4_371 b_4 NI_4 NS_371 0 -3.9438199385855825e-05
GC_4_372 b_4 NI_4 NS_372 0 6.8819462196139630e-05
GC_4_373 b_4 NI_4 NS_373 0 -1.9211240642430234e-04
GC_4_374 b_4 NI_4 NS_374 0 -4.7540070049969694e-04
GC_4_375 b_4 NI_4 NS_375 0 4.9724636543216664e-04
GC_4_376 b_4 NI_4 NS_376 0 1.2130326488493327e-03
GC_4_377 b_4 NI_4 NS_377 0 8.9668980479304893e-06
GC_4_378 b_4 NI_4 NS_378 0 2.0842974941574848e-07
GC_4_379 b_4 NI_4 NS_379 0 -1.6851757960209650e-06
GC_4_380 b_4 NI_4 NS_380 0 -3.7129175061898085e-07
GC_4_381 b_4 NI_4 NS_381 0 4.4123157210418153e-06
GC_4_382 b_4 NI_4 NS_382 0 4.5135015225276798e-06
GC_4_383 b_4 NI_4 NS_383 0 1.6767756935924137e-05
GC_4_384 b_4 NI_4 NS_384 0 -8.8235344594712002e-05
GC_4_385 b_4 NI_4 NS_385 0 3.9265157875443603e-06
GC_4_386 b_4 NI_4 NS_386 0 8.3148982085252731e-06
GC_4_387 b_4 NI_4 NS_387 0 -4.7725574122671133e-08
GC_4_388 b_4 NI_4 NS_388 0 -2.8866313194585851e-06
GC_4_389 b_4 NI_4 NS_389 0 1.1959584208702612e-05
GC_4_390 b_4 NI_4 NS_390 0 1.1578073844377463e-05
GC_4_391 b_4 NI_4 NS_391 0 -8.7168575127969246e-06
GC_4_392 b_4 NI_4 NS_392 0 -1.6252124349344176e-05
GC_4_393 b_4 NI_4 NS_393 0 1.1842650810295671e-02
GC_4_394 b_4 NI_4 NS_394 0 -7.2521038553273139e-04
GC_4_395 b_4 NI_4 NS_395 0 -1.1313545394729674e-03
GC_4_396 b_4 NI_4 NS_396 0 -1.1311517575342846e-03
GC_4_397 b_4 NI_4 NS_397 0 9.5330693731841799e-04
GC_4_398 b_4 NI_4 NS_398 0 3.3415515629537702e-04
GC_4_399 b_4 NI_4 NS_399 0 4.1690772209937443e-03
GC_4_400 b_4 NI_4 NS_400 0 1.0302037479534261e-03
GC_4_401 b_4 NI_4 NS_401 0 -5.8912814116804596e-03
GC_4_402 b_4 NI_4 NS_402 0 3.3053768409972649e-03
GC_4_403 b_4 NI_4 NS_403 0 -4.9250640759408715e-04
GC_4_404 b_4 NI_4 NS_404 0 3.5152937801975162e-04
GC_4_405 b_4 NI_4 NS_405 0 2.6535154767793083e-04
GC_4_406 b_4 NI_4 NS_406 0 -3.2422231045397387e-03
GC_4_407 b_4 NI_4 NS_407 0 6.2509022745123896e-04
GC_4_408 b_4 NI_4 NS_408 0 4.1636414722859196e-04
GC_4_409 b_4 NI_4 NS_409 0 2.4331667145754493e-04
GC_4_410 b_4 NI_4 NS_410 0 1.5777783061693500e-03
GC_4_411 b_4 NI_4 NS_411 0 9.3434572320541314e-04
GC_4_412 b_4 NI_4 NS_412 0 -1.1539185529056075e-03
GC_4_413 b_4 NI_4 NS_413 0 5.9006497812741167e-05
GC_4_414 b_4 NI_4 NS_414 0 -9.8351545604671147e-06
GC_4_415 b_4 NI_4 NS_415 0 8.5116331058274263e-04
GC_4_416 b_4 NI_4 NS_416 0 2.4042279701405713e-03
GC_4_417 b_4 NI_4 NS_417 0 1.2560314525202331e-04
GC_4_418 b_4 NI_4 NS_418 0 5.7032581258317247e-05
GC_4_419 b_4 NI_4 NS_419 0 -2.0477979791696561e-04
GC_4_420 b_4 NI_4 NS_420 0 1.7448236318028497e-05
GC_4_421 b_4 NI_4 NS_421 0 1.0462875316985487e-04
GC_4_422 b_4 NI_4 NS_422 0 -1.3838927664821019e-04
GC_4_423 b_4 NI_4 NS_423 0 2.0754026954036039e-04
GC_4_424 b_4 NI_4 NS_424 0 -2.2819396009707637e-05
GC_4_425 b_4 NI_4 NS_425 0 -9.4772238826392099e-03
GC_4_426 b_4 NI_4 NS_426 0 5.7440921416814774e-04
GC_4_427 b_4 NI_4 NS_427 0 -1.1239263406409256e-04
GC_4_428 b_4 NI_4 NS_428 0 -1.6637232888435128e-04
GC_4_429 b_4 NI_4 NS_429 0 2.5983750767696813e-03
GC_4_430 b_4 NI_4 NS_430 0 1.4392307009514834e-03
GC_4_431 b_4 NI_4 NS_431 0 2.8563323868147309e-03
GC_4_432 b_4 NI_4 NS_432 0 -2.4036037360852273e-03
GC_4_433 b_4 NI_4 NS_433 0 5.7602435479319652e-04
GC_4_434 b_4 NI_4 NS_434 0 3.3119793354136241e-04
GC_4_435 b_4 NI_4 NS_435 0 -9.6470845240151036e-07
GC_4_436 b_4 NI_4 NS_436 0 -9.6680916382199984e-07
GC_4_437 b_4 NI_4 NS_437 0 -1.5589765477560651e-05
GC_4_438 b_4 NI_4 NS_438 0 -1.2977505443487446e-05
GC_4_439 b_4 NI_4 NS_439 0 -7.9312499640558692e-05
GC_4_440 b_4 NI_4 NS_440 0 1.0143600172930184e-04
GC_4_441 b_4 NI_4 NS_441 0 -2.4181462017810817e-05
GC_4_442 b_4 NI_4 NS_442 0 -1.9458132785039453e-05
GC_4_443 b_4 NI_4 NS_443 0 -1.7406629508542091e-05
GC_4_444 b_4 NI_4 NS_444 0 -7.7274045355825316e-06
GC_4_445 b_4 NI_4 NS_445 0 1.8336965072920510e-04
GC_4_446 b_4 NI_4 NS_446 0 -8.5640317900231652e-05
GC_4_447 b_4 NI_4 NS_447 0 -3.0286086554602711e-04
GC_4_448 b_4 NI_4 NS_448 0 4.9418538355000207e-05
GC_4_449 b_4 NI_4 NS_449 0 8.3541258382879863e-03
GC_4_450 b_4 NI_4 NS_450 0 -1.5596779753311102e-04
GC_4_451 b_4 NI_4 NS_451 0 2.9992008258201486e-04
GC_4_452 b_4 NI_4 NS_452 0 1.6281321917316073e-04
GC_4_453 b_4 NI_4 NS_453 0 -7.2501531760149534e-05
GC_4_454 b_4 NI_4 NS_454 0 3.3259414805535245e-04
GC_4_455 b_4 NI_4 NS_455 0 -8.9291454119784432e-04
GC_4_456 b_4 NI_4 NS_456 0 1.2037554243241237e-03
GC_4_457 b_4 NI_4 NS_457 0 -1.5304361208724837e-03
GC_4_458 b_4 NI_4 NS_458 0 -2.8040310377887273e-04
GC_4_459 b_4 NI_4 NS_459 0 -7.1976696991134990e-05
GC_4_460 b_4 NI_4 NS_460 0 -4.3687741543183928e-04
GC_4_461 b_4 NI_4 NS_461 0 -1.3282069440219160e-05
GC_4_462 b_4 NI_4 NS_462 0 -1.3372988690781810e-03
GC_4_463 b_4 NI_4 NS_463 0 8.4212323447788293e-04
GC_4_464 b_4 NI_4 NS_464 0 -4.9874178830056765e-04
GC_4_465 b_4 NI_4 NS_465 0 1.7715174851959225e-03
GC_4_466 b_4 NI_4 NS_466 0 1.6514170984603066e-03
GC_4_467 b_4 NI_4 NS_467 0 -4.2767996000230680e-04
GC_4_468 b_4 NI_4 NS_468 0 2.6322706769465625e-03
GC_4_469 b_4 NI_4 NS_469 0 -2.2164509615889169e-04
GC_4_470 b_4 NI_4 NS_470 0 -3.6807200594322628e-05
GC_4_471 b_4 NI_4 NS_471 0 -2.7962257153377758e-03
GC_4_472 b_4 NI_4 NS_472 0 2.2968638823877524e-03
GC_4_473 b_4 NI_4 NS_473 0 2.5995171705707503e-04
GC_4_474 b_4 NI_4 NS_474 0 3.1486733049427179e-04
GC_4_475 b_4 NI_4 NS_475 0 -8.7293648607054237e-04
GC_4_476 b_4 NI_4 NS_476 0 5.9799869603380964e-05
GC_4_477 b_4 NI_4 NS_477 0 -4.4767132611177085e-04
GC_4_478 b_4 NI_4 NS_478 0 -4.9558419342544723e-06
GC_4_479 b_4 NI_4 NS_479 0 -1.0010037658399066e-04
GC_4_480 b_4 NI_4 NS_480 0 -2.7372519025534829e-05
GC_4_481 b_4 NI_4 NS_481 0 -9.3885194285084057e-04
GC_4_482 b_4 NI_4 NS_482 0 -4.9262550703068715e-03
GC_4_483 b_4 NI_4 NS_483 0 4.9795896337567164e-05
GC_4_484 b_4 NI_4 NS_484 0 -3.2849116563761617e-05
GC_4_485 b_4 NI_4 NS_485 0 -1.0385789816076522e-03
GC_4_486 b_4 NI_4 NS_486 0 6.1131235076380334e-04
GC_4_487 b_4 NI_4 NS_487 0 1.3134074791262571e-03
GC_4_488 b_4 NI_4 NS_488 0 -3.7140542409262077e-05
GC_4_489 b_4 NI_4 NS_489 0 -1.1646922975184790e-04
GC_4_490 b_4 NI_4 NS_490 0 1.1464536013124625e-04
GC_4_491 b_4 NI_4 NS_491 0 -8.6928792501576774e-07
GC_4_492 b_4 NI_4 NS_492 0 7.0669456043097715e-07
GC_4_493 b_4 NI_4 NS_493 0 -6.8625981140483941e-07
GC_4_494 b_4 NI_4 NS_494 0 -3.6740313875714558e-06
GC_4_495 b_4 NI_4 NS_495 0 -5.5523096424230983e-05
GC_4_496 b_4 NI_4 NS_496 0 9.0751851989159499e-06
GC_4_497 b_4 NI_4 NS_497 0 -4.6765968020468784e-07
GC_4_498 b_4 NI_4 NS_498 0 -4.3128747410743420e-06
GC_4_499 b_4 NI_4 NS_499 0 -8.7701489183852265e-07
GC_4_500 b_4 NI_4 NS_500 0 -4.6204918300566405e-06
GC_4_501 b_4 NI_4 NS_501 0 1.9695804147559234e-05
GC_4_502 b_4 NI_4 NS_502 0 1.2629825504408031e-05
GC_4_503 b_4 NI_4 NS_503 0 -2.3089587112974992e-05
GC_4_504 b_4 NI_4 NS_504 0 -2.7862051852029891e-05
GC_4_505 b_4 NI_4 NS_505 0 -4.8220290292238874e-03
GC_4_506 b_4 NI_4 NS_506 0 8.1014462567417299e-06
GC_4_507 b_4 NI_4 NS_507 0 -1.8579110550171675e-04
GC_4_508 b_4 NI_4 NS_508 0 7.5669461402395928e-05
GC_4_509 b_4 NI_4 NS_509 0 -1.1905336900613564e-04
GC_4_510 b_4 NI_4 NS_510 0 -1.7175623636041137e-04
GC_4_511 b_4 NI_4 NS_511 0 4.4306678526383631e-05
GC_4_512 b_4 NI_4 NS_512 0 -1.0739952950733543e-03
GC_4_513 b_4 NI_4 NS_513 0 1.0894129461494560e-03
GC_4_514 b_4 NI_4 NS_514 0 -5.0462019153918583e-05
GC_4_515 b_4 NI_4 NS_515 0 -1.4218737152429860e-04
GC_4_516 b_4 NI_4 NS_516 0 7.4389031958401307e-05
GC_4_517 b_4 NI_4 NS_517 0 -4.1158124747220679e-04
GC_4_518 b_4 NI_4 NS_518 0 -3.2487793676991722e-04
GC_4_519 b_4 NI_4 NS_519 0 3.8850714071465099e-04
GC_4_520 b_4 NI_4 NS_520 0 -4.6949377487971836e-04
GC_4_521 b_4 NI_4 NS_521 0 2.0966579713653819e-04
GC_4_522 b_4 NI_4 NS_522 0 1.0461961465598284e-03
GC_4_523 b_4 NI_4 NS_523 0 -1.4394810726183131e-03
GC_4_524 b_4 NI_4 NS_524 0 -1.3501915266895552e-03
GC_4_525 b_4 NI_4 NS_525 0 1.2089471799869636e-04
GC_4_526 b_4 NI_4 NS_526 0 5.9695122355743779e-05
GC_4_527 b_4 NI_4 NS_527 0 3.7622566574762768e-03
GC_4_528 b_4 NI_4 NS_528 0 -2.2908599282003379e-03
GC_4_529 b_4 NI_4 NS_529 0 -4.7923894773774743e-04
GC_4_530 b_4 NI_4 NS_530 0 3.2762336628876411e-04
GC_4_531 b_4 NI_4 NS_531 0 -4.3239448104811080e-04
GC_4_532 b_4 NI_4 NS_532 0 4.7632357880427129e-04
GC_4_533 b_4 NI_4 NS_533 0 -4.9976557412764536e-05
GC_4_534 b_4 NI_4 NS_534 0 -5.0453787232199469e-04
GC_4_535 b_4 NI_4 NS_535 0 1.6528289762708949e-04
GC_4_536 b_4 NI_4 NS_536 0 -1.5927763877036886e-05
GC_4_537 b_4 NI_4 NS_537 0 1.7151528197458781e-03
GC_4_538 b_4 NI_4 NS_538 0 3.6008122969227014e-03
GC_4_539 b_4 NI_4 NS_539 0 -1.1146193223280208e-04
GC_4_540 b_4 NI_4 NS_540 0 1.7564959984267298e-04
GC_4_541 b_4 NI_4 NS_541 0 1.5058143802241376e-03
GC_4_542 b_4 NI_4 NS_542 0 -7.2804425506133551e-04
GC_4_543 b_4 NI_4 NS_543 0 -2.3375350693180543e-03
GC_4_544 b_4 NI_4 NS_544 0 -5.8274616820692450e-04
GC_4_545 b_4 NI_4 NS_545 0 -7.2179203897080962e-04
GC_4_546 b_4 NI_4 NS_546 0 5.0053665904014276e-04
GC_4_547 b_4 NI_4 NS_547 0 4.8217365205937500e-06
GC_4_548 b_4 NI_4 NS_548 0 -4.3372150851124209e-06
GC_4_549 b_4 NI_4 NS_549 0 -1.1612599990686002e-06
GC_4_550 b_4 NI_4 NS_550 0 5.5955075002358601e-05
GC_4_551 b_4 NI_4 NS_551 0 2.2287175037177833e-04
GC_4_552 b_4 NI_4 NS_552 0 -1.5966784911228404e-04
GC_4_553 b_4 NI_4 NS_553 0 4.8453017270866098e-05
GC_4_554 b_4 NI_4 NS_554 0 7.3424305143475761e-05
GC_4_555 b_4 NI_4 NS_555 0 7.1263624059530908e-06
GC_4_556 b_4 NI_4 NS_556 0 3.8255164872408591e-05
GC_4_557 b_4 NI_4 NS_557 0 2.1947760902529443e-04
GC_4_558 b_4 NI_4 NS_558 0 -1.6130824447481814e-04
GC_4_559 b_4 NI_4 NS_559 0 -3.6770304792301911e-04
GC_4_560 b_4 NI_4 NS_560 0 1.3817210153537152e-04
GC_4_561 b_4 NI_4 NS_561 0 1.5858636601444537e-03
GC_4_562 b_4 NI_4 NS_562 0 -1.3930469552208511e-04
GC_4_563 b_4 NI_4 NS_563 0 1.6660069711449312e-04
GC_4_564 b_4 NI_4 NS_564 0 5.6245497460988595e-04
GC_4_565 b_4 NI_4 NS_565 0 -5.2813873839790927e-04
GC_4_566 b_4 NI_4 NS_566 0 -1.1100270235502406e-05
GC_4_567 b_4 NI_4 NS_567 0 -1.6224592255486558e-03
GC_4_568 b_4 NI_4 NS_568 0 -2.9776274694617979e-04
GC_4_569 b_4 NI_4 NS_569 0 5.9819465835813268e-04
GC_4_570 b_4 NI_4 NS_570 0 -1.9505061449112584e-03
GC_4_571 b_4 NI_4 NS_571 0 -1.5459692254231479e-05
GC_4_572 b_4 NI_4 NS_572 0 -1.9708618841355241e-04
GC_4_573 b_4 NI_4 NS_573 0 1.1849199735914830e-03
GC_4_574 b_4 NI_4 NS_574 0 -1.2359309433804316e-03
GC_4_575 b_4 NI_4 NS_575 0 7.3022842895235863e-04
GC_4_576 b_4 NI_4 NS_576 0 -2.3178773431841156e-04
GC_4_577 b_4 NI_4 NS_577 0 1.8185155508737905e-03
GC_4_578 b_4 NI_4 NS_578 0 1.9867095240929614e-03
GC_4_579 b_4 NI_4 NS_579 0 -5.4998114947572808e-04
GC_4_580 b_4 NI_4 NS_580 0 2.1768067422879172e-03
GC_4_581 b_4 NI_4 NS_581 0 -1.7623390754204879e-04
GC_4_582 b_4 NI_4 NS_582 0 -1.3365964921591280e-05
GC_4_583 b_4 NI_4 NS_583 0 -1.7125346298857199e-03
GC_4_584 b_4 NI_4 NS_584 0 1.3173825088645789e-03
GC_4_585 b_4 NI_4 NS_585 0 -1.3141239330172483e-05
GC_4_586 b_4 NI_4 NS_586 0 2.9410002192192699e-04
GC_4_587 b_4 NI_4 NS_587 0 -5.4947397875090983e-04
GC_4_588 b_4 NI_4 NS_588 0 9.6961764525919036e-05
GC_4_589 b_4 NI_4 NS_589 0 -3.4944923352631167e-04
GC_4_590 b_4 NI_4 NS_590 0 1.8528832096961622e-06
GC_4_591 b_4 NI_4 NS_591 0 -7.7701770086029443e-05
GC_4_592 b_4 NI_4 NS_592 0 -4.2295818295627514e-05
GC_4_593 b_4 NI_4 NS_593 0 -4.8350120676219922e-04
GC_4_594 b_4 NI_4 NS_594 0 -2.6842009504624178e-03
GC_4_595 b_4 NI_4 NS_595 0 1.8486442492201550e-05
GC_4_596 b_4 NI_4 NS_596 0 -6.2174111641037304e-06
GC_4_597 b_4 NI_4 NS_597 0 -6.3530729613604233e-04
GC_4_598 b_4 NI_4 NS_598 0 1.9393675084698847e-04
GC_4_599 b_4 NI_4 NS_599 0 9.7894910789429420e-04
GC_4_600 b_4 NI_4 NS_600 0 -3.1189658230046293e-04
GC_4_601 b_4 NI_4 NS_601 0 -1.0361976580204264e-04
GC_4_602 b_4 NI_4 NS_602 0 5.9585767990028749e-05
GC_4_603 b_4 NI_4 NS_603 0 -1.2427407089017877e-06
GC_4_604 b_4 NI_4 NS_604 0 7.7525633150601748e-07
GC_4_605 b_4 NI_4 NS_605 0 3.9412766755316030e-06
GC_4_606 b_4 NI_4 NS_606 0 -3.1970582338253176e-07
GC_4_607 b_4 NI_4 NS_607 0 -5.0436767265441377e-05
GC_4_608 b_4 NI_4 NS_608 0 -5.8783799963088863e-05
GC_4_609 b_4 NI_4 NS_609 0 1.1300242728689475e-05
GC_4_610 b_4 NI_4 NS_610 0 2.8132194829211404e-07
GC_4_611 b_4 NI_4 NS_611 0 3.1110831360953645e-06
GC_4_612 b_4 NI_4 NS_612 0 -3.6760171352308174e-06
GC_4_613 b_4 NI_4 NS_613 0 1.9556764542855390e-05
GC_4_614 b_4 NI_4 NS_614 0 -1.9747561453474472e-06
GC_4_615 b_4 NI_4 NS_615 0 -2.3715436457460311e-05
GC_4_616 b_4 NI_4 NS_616 0 -1.8413322119209303e-06
GC_4_617 b_4 NI_4 NS_617 0 3.3050164038153076e-03
GC_4_618 b_4 NI_4 NS_618 0 -4.8021178342928932e-05
GC_4_619 b_4 NI_4 NS_619 0 -3.2253134973447741e-04
GC_4_620 b_4 NI_4 NS_620 0 -9.0109417998021166e-05
GC_4_621 b_4 NI_4 NS_621 0 1.7432495012061172e-04
GC_4_622 b_4 NI_4 NS_622 0 -2.5189239076991093e-04
GC_4_623 b_4 NI_4 NS_623 0 1.1631586436919605e-03
GC_4_624 b_4 NI_4 NS_624 0 -5.8183704093182009e-04
GC_4_625 b_4 NI_4 NS_625 0 3.6968073870633866e-04
GC_4_626 b_4 NI_4 NS_626 0 1.8752666597975395e-03
GC_4_627 b_4 NI_4 NS_627 0 -4.4996178209183717e-04
GC_4_628 b_4 NI_4 NS_628 0 9.0295454406442733e-05
GC_4_629 b_4 NI_4 NS_629 0 -4.5856193887274795e-04
GC_4_630 b_4 NI_4 NS_630 0 -4.6462764736873447e-04
GC_4_631 b_4 NI_4 NS_631 0 3.8048480039439209e-04
GC_4_632 b_4 NI_4 NS_632 0 -1.6482054443329327e-04
GC_4_633 b_4 NI_4 NS_633 0 4.1126070893005484e-04
GC_4_634 b_4 NI_4 NS_634 0 1.4706506396172066e-03
GC_4_635 b_4 NI_4 NS_635 0 -6.3405387300788396e-04
GC_4_636 b_4 NI_4 NS_636 0 -6.6990412337148309e-04
GC_4_637 b_4 NI_4 NS_637 0 7.1833917340243279e-05
GC_4_638 b_4 NI_4 NS_638 0 3.2018601183688705e-05
GC_4_639 b_4 NI_4 NS_639 0 1.4017862101918484e-03
GC_4_640 b_4 NI_4 NS_640 0 1.8753689565674181e-04
GC_4_641 b_4 NI_4 NS_641 0 -1.8068547188373617e-04
GC_4_642 b_4 NI_4 NS_642 0 1.6922299123871986e-04
GC_4_643 b_4 NI_4 NS_643 0 -3.1914150012934300e-04
GC_4_644 b_4 NI_4 NS_644 0 2.3487755375656153e-04
GC_4_645 b_4 NI_4 NS_645 0 1.0396678937707721e-05
GC_4_646 b_4 NI_4 NS_646 0 -2.7177462186975894e-04
GC_4_647 b_4 NI_4 NS_647 0 1.1072171978498116e-04
GC_4_648 b_4 NI_4 NS_648 0 1.2352429771196485e-05
GC_4_649 b_4 NI_4 NS_649 0 -1.7674768436029490e-03
GC_4_650 b_4 NI_4 NS_650 0 2.0872659921670530e-03
GC_4_651 b_4 NI_4 NS_651 0 -8.4304222663080951e-05
GC_4_652 b_4 NI_4 NS_652 0 3.0455192690586410e-05
GC_4_653 b_4 NI_4 NS_653 0 1.2855562465060645e-03
GC_4_654 b_4 NI_4 NS_654 0 2.4229830543293107e-04
GC_4_655 b_4 NI_4 NS_655 0 -8.0060001840199201e-04
GC_4_656 b_4 NI_4 NS_656 0 -1.4584233187646526e-03
GC_4_657 b_4 NI_4 NS_657 0 -2.8962714168134909e-04
GC_4_658 b_4 NI_4 NS_658 0 2.9537996650344571e-04
GC_4_659 b_4 NI_4 NS_659 0 2.9394604000572733e-06
GC_4_660 b_4 NI_4 NS_660 0 -5.7075544580254599e-07
GC_4_661 b_4 NI_4 NS_661 0 -9.2653446333004354e-06
GC_4_662 b_4 NI_4 NS_662 0 2.2410213796722903e-05
GC_4_663 b_4 NI_4 NS_663 0 1.1949593111108726e-04
GC_4_664 b_4 NI_4 NS_664 0 -2.3498513873235340e-05
GC_4_665 b_4 NI_4 NS_665 0 1.1983411701725668e-05
GC_4_666 b_4 NI_4 NS_666 0 3.5313486883429372e-05
GC_4_667 b_4 NI_4 NS_667 0 -7.4874820594826929e-06
GC_4_668 b_4 NI_4 NS_668 0 1.7522848921826836e-05
GC_4_669 b_4 NI_4 NS_669 0 1.5235210457751735e-04
GC_4_670 b_4 NI_4 NS_670 0 -7.2559658131728498e-05
GC_4_671 b_4 NI_4 NS_671 0 -2.4512172561037447e-04
GC_4_672 b_4 NI_4 NS_672 0 4.6970785578714322e-05
GD_4_1 b_4 NI_4 NA_1 0 -6.0404051628895707e-02
GD_4_2 b_4 NI_4 NA_2 0 1.1471403074301860e-02
GD_4_3 b_4 NI_4 NA_3 0 3.7780276852621718e-02
GD_4_4 b_4 NI_4 NA_4 0 9.4552368489063676e-02
GD_4_5 b_4 NI_4 NA_5 0 -2.1846663069441136e-02
GD_4_6 b_4 NI_4 NA_6 0 -1.8815260441414329e-02
GD_4_7 b_4 NI_4 NA_7 0 6.2067249436076940e-03
GD_4_8 b_4 NI_4 NA_8 0 -1.4753932160993802e-02
GD_4_9 b_4 NI_4 NA_9 0 -3.1807006864975206e-03
GD_4_10 b_4 NI_4 NA_10 0 3.0061871428493400e-03
GD_4_11 b_4 NI_4 NA_11 0 8.5494315936181621e-04
GD_4_12 b_4 NI_4 NA_12 0 -5.4585833604299918e-03
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 3.9255922856509952e-02
GC_5_2 b_5 NI_5 NS_2 0 8.4906406420566028e-05
GC_5_3 b_5 NI_5 NS_3 0 5.3213037231657238e-03
GC_5_4 b_5 NI_5 NS_4 0 7.7864468082119098e-05
GC_5_5 b_5 NI_5 NS_5 0 -3.9292101639275545e-03
GC_5_6 b_5 NI_5 NS_6 0 3.0866355596593335e-03
GC_5_7 b_5 NI_5 NS_7 0 -1.7463966475110596e-03
GC_5_8 b_5 NI_5 NS_8 0 7.6522113254428956e-03
GC_5_9 b_5 NI_5 NS_9 0 -9.4884937240854502e-03
GC_5_10 b_5 NI_5 NS_10 0 -5.9785944858851076e-03
GC_5_11 b_5 NI_5 NS_11 0 -2.6382611878225350e-04
GC_5_12 b_5 NI_5 NS_12 0 -1.1882059360947652e-04
GC_5_13 b_5 NI_5 NS_13 0 7.6099315043891488e-03
GC_5_14 b_5 NI_5 NS_14 0 2.6309735783813456e-04
GC_5_15 b_5 NI_5 NS_15 0 7.0235856597317242e-05
GC_5_16 b_5 NI_5 NS_16 0 2.2030319256351330e-03
GC_5_17 b_5 NI_5 NS_17 0 -1.1519151613016176e-03
GC_5_18 b_5 NI_5 NS_18 0 1.6540954058437076e-03
GC_5_19 b_5 NI_5 NS_19 0 1.1223345824188432e-03
GC_5_20 b_5 NI_5 NS_20 0 5.4039141023009326e-03
GC_5_21 b_5 NI_5 NS_21 0 2.9250243053733927e-04
GC_5_22 b_5 NI_5 NS_22 0 9.8879282896870046e-05
GC_5_23 b_5 NI_5 NS_23 0 -9.7263860482746083e-03
GC_5_24 b_5 NI_5 NS_24 0 4.0457099531868998e-03
GC_5_25 b_5 NI_5 NS_25 0 1.1626125657071566e-03
GC_5_26 b_5 NI_5 NS_26 0 3.4034004408279981e-04
GC_5_27 b_5 NI_5 NS_27 0 -3.7366477906818199e-04
GC_5_28 b_5 NI_5 NS_28 0 6.2673808995403654e-05
GC_5_29 b_5 NI_5 NS_29 0 -1.9765313112290659e-04
GC_5_30 b_5 NI_5 NS_30 0 2.5834166597401138e-04
GC_5_31 b_5 NI_5 NS_31 0 -8.3960394057362223e-05
GC_5_32 b_5 NI_5 NS_32 0 7.4307383211988963e-06
GC_5_33 b_5 NI_5 NS_33 0 -8.7301582356081459e-03
GC_5_34 b_5 NI_5 NS_34 0 -9.8459004977735042e-03
GC_5_35 b_5 NI_5 NS_35 0 1.0100869528499695e-04
GC_5_36 b_5 NI_5 NS_36 0 -5.6669580292478067e-05
GC_5_37 b_5 NI_5 NS_37 0 -4.8209041000187291e-04
GC_5_38 b_5 NI_5 NS_38 0 2.3272483731547446e-03
GC_5_39 b_5 NI_5 NS_39 0 5.9199581255972421e-03
GC_5_40 b_5 NI_5 NS_40 0 -1.5671446125624481e-04
GC_5_41 b_5 NI_5 NS_41 0 4.4812749839583024e-04
GC_5_42 b_5 NI_5 NS_42 0 4.0248478939143350e-04
GC_5_43 b_5 NI_5 NS_43 0 2.5527359346437796e-06
GC_5_44 b_5 NI_5 NS_44 0 3.5557784946793501e-06
GC_5_45 b_5 NI_5 NS_45 0 5.6281754698116808e-06
GC_5_46 b_5 NI_5 NS_46 0 -1.6198824868771408e-05
GC_5_47 b_5 NI_5 NS_47 0 -3.1726559552697789e-04
GC_5_48 b_5 NI_5 NS_48 0 -1.2513953714793065e-05
GC_5_49 b_5 NI_5 NS_49 0 1.9844323073000690e-05
GC_5_50 b_5 NI_5 NS_50 0 -2.8636864359057990e-05
GC_5_51 b_5 NI_5 NS_51 0 -1.7002672156305354e-05
GC_5_52 b_5 NI_5 NS_52 0 1.0656877360022343e-07
GC_5_53 b_5 NI_5 NS_53 0 5.0687603539202452e-05
GC_5_54 b_5 NI_5 NS_54 0 -3.5673429346612884e-05
GC_5_55 b_5 NI_5 NS_55 0 -8.7190713155115633e-05
GC_5_56 b_5 NI_5 NS_56 0 2.8753954698185322e-05
GC_5_57 b_5 NI_5 NS_57 0 -5.8437431343360486e-03
GC_5_58 b_5 NI_5 NS_58 0 -2.5992688754314245e-04
GC_5_59 b_5 NI_5 NS_59 0 -1.3292982173812582e-03
GC_5_60 b_5 NI_5 NS_60 0 3.0355052147258794e-03
GC_5_61 b_5 NI_5 NS_61 0 -9.5126401772885360e-04
GC_5_62 b_5 NI_5 NS_62 0 -2.2008466563582570e-03
GC_5_63 b_5 NI_5 NS_63 0 -5.0103479130262233e-03
GC_5_64 b_5 NI_5 NS_64 0 -5.7005805576151010e-03
GC_5_65 b_5 NI_5 NS_65 0 7.2765678784788455e-03
GC_5_66 b_5 NI_5 NS_66 0 -1.0999239210182389e-03
GC_5_67 b_5 NI_5 NS_67 0 -9.0613370146775706e-05
GC_5_68 b_5 NI_5 NS_68 0 -3.3558464459312651e-05
GC_5_69 b_5 NI_5 NS_69 0 4.0156481686963435e-03
GC_5_70 b_5 NI_5 NS_70 0 -2.3759595544820588e-03
GC_5_71 b_5 NI_5 NS_71 0 7.9215622525375339e-04
GC_5_72 b_5 NI_5 NS_72 0 1.1360894362744429e-03
GC_5_73 b_5 NI_5 NS_73 0 3.0544221532314393e-04
GC_5_74 b_5 NI_5 NS_74 0 2.2186151797783890e-03
GC_5_75 b_5 NI_5 NS_75 0 -3.3756750504002589e-03
GC_5_76 b_5 NI_5 NS_76 0 1.0898686606650575e-03
GC_5_77 b_5 NI_5 NS_77 0 -2.1849272191893724e-04
GC_5_78 b_5 NI_5 NS_78 0 5.6866315100970726e-06
GC_5_79 b_5 NI_5 NS_79 0 2.9342657956888695e-03
GC_5_80 b_5 NI_5 NS_80 0 -4.5477697113873551e-04
GC_5_81 b_5 NI_5 NS_81 0 -1.0827613662089343e-03
GC_5_82 b_5 NI_5 NS_82 0 -1.8172426413046785e-04
GC_5_83 b_5 NI_5 NS_83 0 -1.5170823785680925e-04
GC_5_84 b_5 NI_5 NS_84 0 8.3132763297223689e-05
GC_5_85 b_5 NI_5 NS_85 0 -3.1767124285321681e-04
GC_5_86 b_5 NI_5 NS_86 0 2.8571134671269080e-04
GC_5_87 b_5 NI_5 NS_87 0 -2.0423523715241740e-04
GC_5_88 b_5 NI_5 NS_88 0 -8.7120834806874039e-05
GC_5_89 b_5 NI_5 NS_89 0 2.1318505270864641e-03
GC_5_90 b_5 NI_5 NS_90 0 4.0851511747707985e-07
GC_5_91 b_5 NI_5 NS_91 0 -2.6501039890323157e-05
GC_5_92 b_5 NI_5 NS_92 0 1.2289428691585879e-04
GC_5_93 b_5 NI_5 NS_93 0 -4.6833155305197195e-04
GC_5_94 b_5 NI_5 NS_94 0 -7.2111847405685744e-04
GC_5_95 b_5 NI_5 NS_95 0 -7.0385127645895232e-04
GC_5_96 b_5 NI_5 NS_96 0 1.0700920481882131e-03
GC_5_97 b_5 NI_5 NS_97 0 8.2099507453705888e-05
GC_5_98 b_5 NI_5 NS_98 0 -6.0920722711648894e-05
GC_5_99 b_5 NI_5 NS_99 0 1.0117574893070006e-06
GC_5_100 b_5 NI_5 NS_100 0 -4.8294358437161441e-07
GC_5_101 b_5 NI_5 NS_101 0 -1.0041469975087210e-06
GC_5_102 b_5 NI_5 NS_102 0 2.5545879802911533e-06
GC_5_103 b_5 NI_5 NS_103 0 1.0881026975632944e-04
GC_5_104 b_5 NI_5 NS_104 0 -3.9564429649373152e-06
GC_5_105 b_5 NI_5 NS_105 0 -5.4194295292888450e-06
GC_5_106 b_5 NI_5 NS_106 0 7.8767466564199083e-06
GC_5_107 b_5 NI_5 NS_107 0 -6.9514270064990430e-06
GC_5_108 b_5 NI_5 NS_108 0 -1.6376175821319076e-06
GC_5_109 b_5 NI_5 NS_109 0 -7.1184987483230251e-06
GC_5_110 b_5 NI_5 NS_110 0 7.1693213655993989e-07
GC_5_111 b_5 NI_5 NS_111 0 9.7273291413036255e-06
GC_5_112 b_5 NI_5 NS_112 0 4.0972988851781749e-06
GC_5_113 b_5 NI_5 NS_113 0 3.4757877230602578e-02
GC_5_114 b_5 NI_5 NS_114 0 1.4285908315958662e-03
GC_5_115 b_5 NI_5 NS_115 0 5.8246829355904448e-03
GC_5_116 b_5 NI_5 NS_116 0 1.1407472833036352e-03
GC_5_117 b_5 NI_5 NS_117 0 -4.4989329353638859e-03
GC_5_118 b_5 NI_5 NS_118 0 -3.3622288087821334e-03
GC_5_119 b_5 NI_5 NS_119 0 4.1888735887329800e-03
GC_5_120 b_5 NI_5 NS_120 0 9.8493817124306726e-03
GC_5_121 b_5 NI_5 NS_121 0 4.6730983945963734e-04
GC_5_122 b_5 NI_5 NS_122 0 -4.9714329890086905e-03
GC_5_123 b_5 NI_5 NS_123 0 -3.4611869273765090e-04
GC_5_124 b_5 NI_5 NS_124 0 3.9560643956741757e-04
GC_5_125 b_5 NI_5 NS_125 0 9.6488309528021086e-03
GC_5_126 b_5 NI_5 NS_126 0 3.5231083082196408e-03
GC_5_127 b_5 NI_5 NS_127 0 5.3910614606855051e-04
GC_5_128 b_5 NI_5 NS_128 0 3.3158879071446463e-03
GC_5_129 b_5 NI_5 NS_129 0 2.4550411785959334e-03
GC_5_130 b_5 NI_5 NS_130 0 4.4743865182008550e-03
GC_5_131 b_5 NI_5 NS_131 0 3.0647654859365494e-03
GC_5_132 b_5 NI_5 NS_132 0 7.6251244386686739e-03
GC_5_133 b_5 NI_5 NS_133 0 4.3958183871924171e-04
GC_5_134 b_5 NI_5 NS_134 0 1.1146693101677806e-04
GC_5_135 b_5 NI_5 NS_135 0 -1.5839669244082148e-02
GC_5_136 b_5 NI_5 NS_136 0 1.3005523545564938e-02
GC_5_137 b_5 NI_5 NS_137 0 1.9133503178610973e-03
GC_5_138 b_5 NI_5 NS_138 0 3.9897100396051282e-04
GC_5_139 b_5 NI_5 NS_139 0 -7.3988404221756073e-04
GC_5_140 b_5 NI_5 NS_140 0 -4.3012283622233922e-07
GC_5_141 b_5 NI_5 NS_141 0 -4.0116847401094473e-04
GC_5_142 b_5 NI_5 NS_142 0 4.6161814261150465e-04
GC_5_143 b_5 NI_5 NS_143 0 -1.8700759973487409e-04
GC_5_144 b_5 NI_5 NS_144 0 4.4962329795423183e-05
GC_5_145 b_5 NI_5 NS_145 0 -8.4930949933557306e-03
GC_5_146 b_5 NI_5 NS_146 0 -1.1959306376016715e-02
GC_5_147 b_5 NI_5 NS_147 0 2.3586608241741655e-04
GC_5_148 b_5 NI_5 NS_148 0 -7.3130540340740860e-05
GC_5_149 b_5 NI_5 NS_149 0 -1.6032663930509823e-03
GC_5_150 b_5 NI_5 NS_150 0 3.5605087776960660e-03
GC_5_151 b_5 NI_5 NS_151 0 3.8194174490047547e-03
GC_5_152 b_5 NI_5 NS_152 0 -1.1618800347848134e-03
GC_5_153 b_5 NI_5 NS_153 0 9.7128552001649382e-05
GC_5_154 b_5 NI_5 NS_154 0 4.4580671647217741e-04
GC_5_155 b_5 NI_5 NS_155 0 -1.4552407116684348e-06
GC_5_156 b_5 NI_5 NS_156 0 3.2419541331341692e-06
GC_5_157 b_5 NI_5 NS_157 0 5.0113612610870148e-06
GC_5_158 b_5 NI_5 NS_158 0 -1.0945075609611899e-05
GC_5_159 b_5 NI_5 NS_159 0 -2.2221420917043809e-04
GC_5_160 b_5 NI_5 NS_160 0 -1.4552022294952967e-05
GC_5_161 b_5 NI_5 NS_161 0 1.6328445474177969e-05
GC_5_162 b_5 NI_5 NS_162 0 -1.8600795521773870e-05
GC_5_163 b_5 NI_5 NS_163 0 -8.0767790051412252e-06
GC_5_164 b_5 NI_5 NS_164 0 -9.2024029862728300e-06
GC_5_165 b_5 NI_5 NS_165 0 4.9664954267575066e-05
GC_5_166 b_5 NI_5 NS_166 0 -1.0182248542118506e-05
GC_5_167 b_5 NI_5 NS_167 0 -7.6913548773778359e-05
GC_5_168 b_5 NI_5 NS_168 0 -9.5243839757651823e-06
GC_5_169 b_5 NI_5 NS_169 0 2.6989211300599669e-02
GC_5_170 b_5 NI_5 NS_170 0 -8.4386319150128915e-04
GC_5_171 b_5 NI_5 NS_171 0 -1.9460633039193515e-03
GC_5_172 b_5 NI_5 NS_172 0 3.7443949577554408e-03
GC_5_173 b_5 NI_5 NS_173 0 1.0569242403260883e-03
GC_5_174 b_5 NI_5 NS_174 0 -3.7916553289368306e-04
GC_5_175 b_5 NI_5 NS_175 0 -9.3446228957583654e-03
GC_5_176 b_5 NI_5 NS_176 0 -3.7940206932850829e-03
GC_5_177 b_5 NI_5 NS_177 0 -1.3066320561298669e-03
GC_5_178 b_5 NI_5 NS_178 0 2.7861828183243786e-03
GC_5_179 b_5 NI_5 NS_179 0 -2.9107677086379421e-04
GC_5_180 b_5 NI_5 NS_180 0 2.3487895642491989e-04
GC_5_181 b_5 NI_5 NS_181 0 5.2061840433471540e-03
GC_5_182 b_5 NI_5 NS_182 0 -5.5271193144102500e-03
GC_5_183 b_5 NI_5 NS_183 0 8.5166089350565603e-04
GC_5_184 b_5 NI_5 NS_184 0 1.5028430640699857e-03
GC_5_185 b_5 NI_5 NS_185 0 2.8189484599676980e-04
GC_5_186 b_5 NI_5 NS_186 0 1.3819754804220272e-03
GC_5_187 b_5 NI_5 NS_187 0 -4.8241587449018904e-03
GC_5_188 b_5 NI_5 NS_188 0 -1.6647652561535260e-04
GC_5_189 b_5 NI_5 NS_189 0 -1.8588142242725319e-04
GC_5_190 b_5 NI_5 NS_190 0 -4.5725509491527699e-06
GC_5_191 b_5 NI_5 NS_191 0 2.1097177417388055e-03
GC_5_192 b_5 NI_5 NS_192 0 1.9641640314407207e-03
GC_5_193 b_5 NI_5 NS_193 0 -9.6364450439285468e-04
GC_5_194 b_5 NI_5 NS_194 0 -1.4031939445776438e-04
GC_5_195 b_5 NI_5 NS_195 0 -2.4112531614852093e-04
GC_5_196 b_5 NI_5 NS_196 0 -8.4638617696260557e-06
GC_5_197 b_5 NI_5 NS_197 0 -4.1669281871295732e-04
GC_5_198 b_5 NI_5 NS_198 0 3.2033563921010026e-04
GC_5_199 b_5 NI_5 NS_199 0 -2.1999514476152095e-04
GC_5_200 b_5 NI_5 NS_200 0 -9.5169664529712965e-05
GC_5_201 b_5 NI_5 NS_201 0 8.3068316002030118e-04
GC_5_202 b_5 NI_5 NS_202 0 -4.0393455624040324e-04
GC_5_203 b_5 NI_5 NS_203 0 -1.7883384735970385e-05
GC_5_204 b_5 NI_5 NS_204 0 1.0993220563728425e-04
GC_5_205 b_5 NI_5 NS_205 0 -5.5298481693348675e-04
GC_5_206 b_5 NI_5 NS_206 0 -4.2752852314615421e-04
GC_5_207 b_5 NI_5 NS_207 0 -2.0470058215717101e-03
GC_5_208 b_5 NI_5 NS_208 0 1.3332881980227616e-04
GC_5_209 b_5 NI_5 NS_209 0 -2.9643042165442816e-05
GC_5_210 b_5 NI_5 NS_210 0 -3.3649383177950486e-05
GC_5_211 b_5 NI_5 NS_211 0 1.3157909568449433e-06
GC_5_212 b_5 NI_5 NS_212 0 -9.2372066178027789e-07
GC_5_213 b_5 NI_5 NS_213 0 1.1669231170229968e-06
GC_5_214 b_5 NI_5 NS_214 0 1.8590746820617220e-06
GC_5_215 b_5 NI_5 NS_215 0 6.5307997703284074e-05
GC_5_216 b_5 NI_5 NS_216 0 -3.7685260909943962e-05
GC_5_217 b_5 NI_5 NS_217 0 -4.5025443447022134e-08
GC_5_218 b_5 NI_5 NS_218 0 7.2192038473696964e-06
GC_5_219 b_5 NI_5 NS_219 0 -8.0829895930168623e-07
GC_5_220 b_5 NI_5 NS_220 0 -6.0596552948207313e-07
GC_5_221 b_5 NI_5 NS_221 0 -7.8439897250288488e-06
GC_5_222 b_5 NI_5 NS_222 0 1.8834634144709982e-05
GC_5_223 b_5 NI_5 NS_223 0 2.1496455210699974e-05
GC_5_224 b_5 NI_5 NS_224 0 -2.4033905025778042e-05
GC_5_225 b_5 NI_5 NS_225 0 -1.2106205601191293e-02
GC_5_226 b_5 NI_5 NS_226 0 1.4909982959097168e-02
GC_5_227 b_5 NI_5 NS_227 0 8.0947304821390453e-03
GC_5_228 b_5 NI_5 NS_228 0 1.4158931219103890e-03
GC_5_229 b_5 NI_5 NS_229 0 1.0211747219819104e-02
GC_5_230 b_5 NI_5 NS_230 0 4.8709367374593247e-03
GC_5_231 b_5 NI_5 NS_231 0 -2.6890782796853813e-03
GC_5_232 b_5 NI_5 NS_232 0 9.0328960939674539e-03
GC_5_233 b_5 NI_5 NS_233 0 -2.6210843216404054e-03
GC_5_234 b_5 NI_5 NS_234 0 6.0127802046638663e-03
GC_5_235 b_5 NI_5 NS_235 0 2.4339527160985557e-04
GC_5_236 b_5 NI_5 NS_236 0 5.1806471772531792e-04
GC_5_237 b_5 NI_5 NS_237 0 1.0625102454481367e-02
GC_5_238 b_5 NI_5 NS_238 0 -2.3388602245150440e-03
GC_5_239 b_5 NI_5 NS_239 0 3.2969954400414439e-04
GC_5_240 b_5 NI_5 NS_240 0 3.0040780317189893e-03
GC_5_241 b_5 NI_5 NS_241 0 3.8281348454611576e-03
GC_5_242 b_5 NI_5 NS_242 0 1.9772686860660502e-03
GC_5_243 b_5 NI_5 NS_243 0 4.3258043780649647e-03
GC_5_244 b_5 NI_5 NS_244 0 7.8191526399162253e-03
GC_5_245 b_5 NI_5 NS_245 0 4.3700421889912577e-04
GC_5_246 b_5 NI_5 NS_246 0 1.9597685507233224e-04
GC_5_247 b_5 NI_5 NS_247 0 -8.5107127704808893e-03
GC_5_248 b_5 NI_5 NS_248 0 5.4135617494588048e-03
GC_5_249 b_5 NI_5 NS_249 0 1.4259872332751139e-03
GC_5_250 b_5 NI_5 NS_250 0 5.9823375683146370e-04
GC_5_251 b_5 NI_5 NS_251 0 -4.4119694723025488e-04
GC_5_252 b_5 NI_5 NS_252 0 -1.1397971188984709e-04
GC_5_253 b_5 NI_5 NS_253 0 -2.9715571277859121e-04
GC_5_254 b_5 NI_5 NS_254 0 5.9506149626159162e-05
GC_5_255 b_5 NI_5 NS_255 0 -6.0786291128760378e-05
GC_5_256 b_5 NI_5 NS_256 0 -7.2377899325126876e-05
GC_5_257 b_5 NI_5 NS_257 0 -2.6667419419627836e-03
GC_5_258 b_5 NI_5 NS_258 0 -4.1240002534539454e-03
GC_5_259 b_5 NI_5 NS_259 0 1.0482030560150569e-04
GC_5_260 b_5 NI_5 NS_260 0 1.6198733007778088e-05
GC_5_261 b_5 NI_5 NS_261 0 -8.3888696252179290e-04
GC_5_262 b_5 NI_5 NS_262 0 1.3838773290205848e-03
GC_5_263 b_5 NI_5 NS_263 0 3.3878601398016012e-03
GC_5_264 b_5 NI_5 NS_264 0 3.1238289642205792e-03
GC_5_265 b_5 NI_5 NS_265 0 1.3956060335376010e-04
GC_5_266 b_5 NI_5 NS_266 0 -9.5855602565912419e-05
GC_5_267 b_5 NI_5 NS_267 0 -1.1369184950210381e-06
GC_5_268 b_5 NI_5 NS_268 0 5.5410919633964626e-07
GC_5_269 b_5 NI_5 NS_269 0 5.7695693489375901e-06
GC_5_270 b_5 NI_5 NS_270 0 1.8571337379067113e-07
GC_5_271 b_5 NI_5 NS_271 0 -6.9920537162807800e-05
GC_5_272 b_5 NI_5 NS_272 0 -2.8351562945778284e-05
GC_5_273 b_5 NI_5 NS_273 0 1.0932919355900739e-05
GC_5_274 b_5 NI_5 NS_274 0 2.7634844674920470e-07
GC_5_275 b_5 NI_5 NS_275 0 2.3285970336293139e-06
GC_5_276 b_5 NI_5 NS_276 0 -1.4762226144958691e-05
GC_5_277 b_5 NI_5 NS_277 0 4.1567358343126321e-05
GC_5_278 b_5 NI_5 NS_278 0 2.0285600062793074e-05
GC_5_279 b_5 NI_5 NS_279 0 -5.4306150961600674e-05
GC_5_280 b_5 NI_5 NS_280 0 -5.0516505908263831e-05
GC_5_281 b_5 NI_5 NS_281 0 -4.5241116662553163e-02
GC_5_282 b_5 NI_5 NS_282 0 1.2126658278099183e-02
GC_5_283 b_5 NI_5 NS_283 0 -2.9182380150429795e-03
GC_5_284 b_5 NI_5 NS_284 0 3.7386200421143769e-03
GC_5_285 b_5 NI_5 NS_285 0 -4.3699494200614948e-03
GC_5_286 b_5 NI_5 NS_286 0 2.1341984242377317e-03
GC_5_287 b_5 NI_5 NS_287 0 -4.8443222586378480e-03
GC_5_288 b_5 NI_5 NS_288 0 -9.2083972724348317e-03
GC_5_289 b_5 NI_5 NS_289 0 -2.5373822466291259e-03
GC_5_290 b_5 NI_5 NS_290 0 -9.1021251796630145e-03
GC_5_291 b_5 NI_5 NS_291 0 6.2227033388843314e-04
GC_5_292 b_5 NI_5 NS_292 0 -1.4884668504702248e-04
GC_5_293 b_5 NI_5 NS_293 0 7.1329857603956038e-03
GC_5_294 b_5 NI_5 NS_294 0 -1.5514971393663856e-03
GC_5_295 b_5 NI_5 NS_295 0 1.5062842471312487e-03
GC_5_296 b_5 NI_5 NS_296 0 1.2893696660305353e-03
GC_5_297 b_5 NI_5 NS_297 0 5.4266406598106479e-03
GC_5_298 b_5 NI_5 NS_298 0 8.8710843935266607e-04
GC_5_299 b_5 NI_5 NS_299 0 -2.4576939074674479e-03
GC_5_300 b_5 NI_5 NS_300 0 1.1536036147651310e-03
GC_5_301 b_5 NI_5 NS_301 0 -3.6616848217801214e-04
GC_5_302 b_5 NI_5 NS_302 0 6.6445525464088506e-05
GC_5_303 b_5 NI_5 NS_303 0 7.7434764618249325e-03
GC_5_304 b_5 NI_5 NS_304 0 -2.6957583583778412e-03
GC_5_305 b_5 NI_5 NS_305 0 -1.7229508288891023e-03
GC_5_306 b_5 NI_5 NS_306 0 -2.1719262819729609e-05
GC_5_307 b_5 NI_5 NS_307 0 -2.7488932855731049e-04
GC_5_308 b_5 NI_5 NS_308 0 1.1878239739605731e-04
GC_5_309 b_5 NI_5 NS_309 0 -4.4658033831632257e-04
GC_5_310 b_5 NI_5 NS_310 0 4.1411167515916793e-04
GC_5_311 b_5 NI_5 NS_311 0 -3.0504463051359509e-04
GC_5_312 b_5 NI_5 NS_312 0 -1.1496658241061419e-04
GC_5_313 b_5 NI_5 NS_313 0 2.5842525410587056e-03
GC_5_314 b_5 NI_5 NS_314 0 -9.3118434286257724e-04
GC_5_315 b_5 NI_5 NS_315 0 -2.1793291717748532e-05
GC_5_316 b_5 NI_5 NS_316 0 1.7615227736192854e-04
GC_5_317 b_5 NI_5 NS_317 0 -9.5410186382213855e-04
GC_5_318 b_5 NI_5 NS_318 0 -8.8012865131547561e-04
GC_5_319 b_5 NI_5 NS_319 0 2.0326240592918898e-03
GC_5_320 b_5 NI_5 NS_320 0 1.2709729702076948e-03
GC_5_321 b_5 NI_5 NS_321 0 -1.2196516446975780e-04
GC_5_322 b_5 NI_5 NS_322 0 -1.5991032327953051e-04
GC_5_323 b_5 NI_5 NS_323 0 1.5547146297026832e-06
GC_5_324 b_5 NI_5 NS_324 0 -2.0148889242635988e-06
GC_5_325 b_5 NI_5 NS_325 0 2.5672981643010530e-06
GC_5_326 b_5 NI_5 NS_326 0 -2.5943822856299262e-06
GC_5_327 b_5 NI_5 NS_327 0 -7.1253127114650325e-05
GC_5_328 b_5 NI_5 NS_328 0 -6.3391827173071727e-05
GC_5_329 b_5 NI_5 NS_329 0 8.9353398906067046e-06
GC_5_330 b_5 NI_5 NS_330 0 1.7795412370628795e-06
GC_5_331 b_5 NI_5 NS_331 0 1.1846592981998867e-06
GC_5_332 b_5 NI_5 NS_332 0 -9.5678934487106601e-06
GC_5_333 b_5 NI_5 NS_333 0 2.3925003922085356e-05
GC_5_334 b_5 NI_5 NS_334 0 5.1828102197222885e-05
GC_5_335 b_5 NI_5 NS_335 0 -9.3275785468834632e-06
GC_5_336 b_5 NI_5 NS_336 0 -9.0459409327946764e-05
GC_5_337 b_5 NI_5 NS_337 0 -2.1720294406718275e-02
GC_5_338 b_5 NI_5 NS_338 0 1.6798521860743587e-03
GC_5_339 b_5 NI_5 NS_339 0 3.6043974572229028e-03
GC_5_340 b_5 NI_5 NS_340 0 2.4430212331954105e-03
GC_5_341 b_5 NI_5 NS_341 0 -5.3181847674778722e-03
GC_5_342 b_5 NI_5 NS_342 0 -6.5605009252241824e-03
GC_5_343 b_5 NI_5 NS_343 0 4.1121300400230867e-03
GC_5_344 b_5 NI_5 NS_344 0 2.0573913982215408e-03
GC_5_345 b_5 NI_5 NS_345 0 1.0332343411193885e-02
GC_5_346 b_5 NI_5 NS_346 0 -1.0197213546175712e-02
GC_5_347 b_5 NI_5 NS_347 0 -3.5358494178652241e-04
GC_5_348 b_5 NI_5 NS_348 0 1.5625094353726007e-04
GC_5_349 b_5 NI_5 NS_349 0 8.6981608579302649e-03
GC_5_350 b_5 NI_5 NS_350 0 3.0601460457480140e-03
GC_5_351 b_5 NI_5 NS_351 0 7.1707804375456628e-04
GC_5_352 b_5 NI_5 NS_352 0 2.0876809031375081e-03
GC_5_353 b_5 NI_5 NS_353 0 6.9603586024996750e-03
GC_5_354 b_5 NI_5 NS_354 0 1.0490131780615476e-03
GC_5_355 b_5 NI_5 NS_355 0 2.6266710926344423e-03
GC_5_356 b_5 NI_5 NS_356 0 3.9523114505835358e-03
GC_5_357 b_5 NI_5 NS_357 0 3.5523277622726343e-04
GC_5_358 b_5 NI_5 NS_358 0 1.3295437534013299e-04
GC_5_359 b_5 NI_5 NS_359 0 -4.1321520522758070e-03
GC_5_360 b_5 NI_5 NS_360 0 1.2930625152287066e-02
GC_5_361 b_5 NI_5 NS_361 0 9.9518265438490005e-04
GC_5_362 b_5 NI_5 NS_362 0 8.3432592184089753e-05
GC_5_363 b_5 NI_5 NS_363 0 -5.2970110635694966e-04
GC_5_364 b_5 NI_5 NS_364 0 7.2766756532874799e-05
GC_5_365 b_5 NI_5 NS_365 0 -1.6781578797079493e-04
GC_5_366 b_5 NI_5 NS_366 0 1.5339793186668050e-04
GC_5_367 b_5 NI_5 NS_367 0 -6.3877336420180571e-05
GC_5_368 b_5 NI_5 NS_368 0 2.5805606966206884e-05
GC_5_369 b_5 NI_5 NS_369 0 -4.3870371139444813e-03
GC_5_370 b_5 NI_5 NS_370 0 -3.1395911155158497e-03
GC_5_371 b_5 NI_5 NS_371 0 7.7194609924731536e-05
GC_5_372 b_5 NI_5 NS_372 0 -4.6487787916782550e-05
GC_5_373 b_5 NI_5 NS_373 0 -9.9880808214365048e-05
GC_5_374 b_5 NI_5 NS_374 0 1.6396446303191777e-03
GC_5_375 b_5 NI_5 NS_375 0 -2.4070897667531467e-04
GC_5_376 b_5 NI_5 NS_376 0 -5.4000804431157971e-04
GC_5_377 b_5 NI_5 NS_377 0 2.0123268353777957e-05
GC_5_378 b_5 NI_5 NS_378 0 2.4720901330126121e-04
GC_5_379 b_5 NI_5 NS_379 0 -5.7246384480495410e-07
GC_5_380 b_5 NI_5 NS_380 0 9.1028936054684004e-08
GC_5_381 b_5 NI_5 NS_381 0 -3.2764029084836441e-07
GC_5_382 b_5 NI_5 NS_382 0 1.1927936044744610e-06
GC_5_383 b_5 NI_5 NS_383 0 3.9302493573392963e-05
GC_5_384 b_5 NI_5 NS_384 0 6.1838636505175755e-05
GC_5_385 b_5 NI_5 NS_385 0 -2.8571316684170865e-06
GC_5_386 b_5 NI_5 NS_386 0 9.9821837589917490e-07
GC_5_387 b_5 NI_5 NS_387 0 -2.8073786932378614e-06
GC_5_388 b_5 NI_5 NS_388 0 -5.0432166161873116e-06
GC_5_389 b_5 NI_5 NS_389 0 1.4787343033818938e-05
GC_5_390 b_5 NI_5 NS_390 0 -9.2576157850498022e-06
GC_5_391 b_5 NI_5 NS_391 0 -2.9553523855348490e-05
GC_5_392 b_5 NI_5 NS_392 0 7.2103030241012901e-06
GC_5_393 b_5 NI_5 NS_393 0 5.8838610799422569e-02
GC_5_394 b_5 NI_5 NS_394 0 -8.1662674123075406e-04
GC_5_395 b_5 NI_5 NS_395 0 -1.7986335138458986e-03
GC_5_396 b_5 NI_5 NS_396 0 2.2781721099495557e-03
GC_5_397 b_5 NI_5 NS_397 0 2.8558879260481384e-03
GC_5_398 b_5 NI_5 NS_398 0 2.8094880422961481e-04
GC_5_399 b_5 NI_5 NS_399 0 -5.2690031174308103e-03
GC_5_400 b_5 NI_5 NS_400 0 6.4726576748678241e-04
GC_5_401 b_5 NI_5 NS_401 0 -6.1537719448901788e-03
GC_5_402 b_5 NI_5 NS_402 0 1.0731209688454828e-02
GC_5_403 b_5 NI_5 NS_403 0 -7.4197931662440359e-04
GC_5_404 b_5 NI_5 NS_404 0 -5.4346936213210781e-04
GC_5_405 b_5 NI_5 NS_405 0 1.5109443784985159e-03
GC_5_406 b_5 NI_5 NS_406 0 -3.9740441007757839e-03
GC_5_407 b_5 NI_5 NS_407 0 8.5127714743117090e-04
GC_5_408 b_5 NI_5 NS_408 0 1.2312434319921566e-03
GC_5_409 b_5 NI_5 NS_409 0 -1.5871471212555643e-04
GC_5_410 b_5 NI_5 NS_410 0 1.0935051819159214e-03
GC_5_411 b_5 NI_5 NS_411 0 -5.6242380321901587e-03
GC_5_412 b_5 NI_5 NS_412 0 9.6414810205926616e-04
GC_5_413 b_5 NI_5 NS_413 0 -1.0923918850305183e-04
GC_5_414 b_5 NI_5 NS_414 0 -7.3884098569328968e-05
GC_5_415 b_5 NI_5 NS_415 0 4.2412489849972472e-04
GC_5_416 b_5 NI_5 NS_416 0 5.3175006912769759e-03
GC_5_417 b_5 NI_5 NS_417 0 -3.6122808488653579e-04
GC_5_418 b_5 NI_5 NS_418 0 -1.6429755977220593e-04
GC_5_419 b_5 NI_5 NS_419 0 -4.3820101474811802e-04
GC_5_420 b_5 NI_5 NS_420 0 2.3869634296605828e-05
GC_5_421 b_5 NI_5 NS_421 0 -3.8853000698072746e-04
GC_5_422 b_5 NI_5 NS_422 0 3.6937540517281752e-04
GC_5_423 b_5 NI_5 NS_423 0 -2.0278482547937863e-04
GC_5_424 b_5 NI_5 NS_424 0 -3.0057326435520718e-05
GC_5_425 b_5 NI_5 NS_425 0 -7.2113834808548152e-03
GC_5_426 b_5 NI_5 NS_426 0 -1.0833815285636707e-03
GC_5_427 b_5 NI_5 NS_427 0 -1.0528095963081946e-06
GC_5_428 b_5 NI_5 NS_428 0 1.4310261402898141e-05
GC_5_429 b_5 NI_5 NS_429 0 -1.4062030232272110e-04
GC_5_430 b_5 NI_5 NS_430 0 8.0115417023036994e-04
GC_5_431 b_5 NI_5 NS_431 0 -1.0811712831981311e-03
GC_5_432 b_5 NI_5 NS_432 0 -2.8405401409620072e-03
GC_5_433 b_5 NI_5 NS_433 0 9.3874344259207271e-05
GC_5_434 b_5 NI_5 NS_434 0 2.1385118282154258e-04
GC_5_435 b_5 NI_5 NS_435 0 2.5547663097333727e-06
GC_5_436 b_5 NI_5 NS_436 0 -2.2362643826538031e-08
GC_5_437 b_5 NI_5 NS_437 0 -3.1766791373625915e-06
GC_5_438 b_5 NI_5 NS_438 0 -7.5027545806033233e-06
GC_5_439 b_5 NI_5 NS_439 0 -5.0754389283518150e-05
GC_5_440 b_5 NI_5 NS_440 0 7.5517330247909398e-05
GC_5_441 b_5 NI_5 NS_441 0 -2.5399134499401888e-06
GC_5_442 b_5 NI_5 NS_442 0 -1.1442734859512302e-05
GC_5_443 b_5 NI_5 NS_443 0 -2.9960486805044498e-06
GC_5_444 b_5 NI_5 NS_444 0 3.2800228740531214e-06
GC_5_445 b_5 NI_5 NS_445 0 2.2093981750129802e-06
GC_5_446 b_5 NI_5 NS_446 0 3.0645253087532553e-06
GC_5_447 b_5 NI_5 NS_447 0 4.6849575726335579e-07
GC_5_448 b_5 NI_5 NS_448 0 -8.2754733376323880e-06
GC_5_449 b_5 NI_5 NS_449 0 1.6594667329140951e-02
GC_5_450 b_5 NI_5 NS_450 0 7.0318859551580181e-05
GC_5_451 b_5 NI_5 NS_451 0 3.4521977071539126e-04
GC_5_452 b_5 NI_5 NS_452 0 -5.9571325588329610e-04
GC_5_453 b_5 NI_5 NS_453 0 5.5723014782172136e-04
GC_5_454 b_5 NI_5 NS_454 0 5.9051322702696307e-04
GC_5_455 b_5 NI_5 NS_455 0 9.6860272631444939e-04
GC_5_456 b_5 NI_5 NS_456 0 1.5952511360161209e-03
GC_5_457 b_5 NI_5 NS_457 0 -1.8403884151855566e-03
GC_5_458 b_5 NI_5 NS_458 0 2.0946128963686577e-03
GC_5_459 b_5 NI_5 NS_459 0 -5.2514714555208265e-04
GC_5_460 b_5 NI_5 NS_460 0 9.7683221468350054e-05
GC_5_461 b_5 NI_5 NS_461 0 1.0907044888765966e-03
GC_5_462 b_5 NI_5 NS_462 0 -1.4801753050581474e-03
GC_5_463 b_5 NI_5 NS_463 0 1.7808080112936694e-03
GC_5_464 b_5 NI_5 NS_464 0 2.3823357199193509e-04
GC_5_465 b_5 NI_5 NS_465 0 -1.7801516805619544e-03
GC_5_466 b_5 NI_5 NS_466 0 2.2762580253603689e-03
GC_5_467 b_5 NI_5 NS_467 0 3.1635955106169792e-03
GC_5_468 b_5 NI_5 NS_468 0 3.2254516397142962e-04
GC_5_469 b_5 NI_5 NS_469 0 6.6354827695972612e-04
GC_5_470 b_5 NI_5 NS_470 0 2.3564052648415452e-04
GC_5_471 b_5 NI_5 NS_471 0 -2.0617957575215480e-03
GC_5_472 b_5 NI_5 NS_472 0 9.8864751025473860e-03
GC_5_473 b_5 NI_5 NS_473 0 -6.7550175779437229e-04
GC_5_474 b_5 NI_5 NS_474 0 -1.1182329437895598e-03
GC_5_475 b_5 NI_5 NS_475 0 -1.3538842882976189e-03
GC_5_476 b_5 NI_5 NS_476 0 -7.6675928359321173e-05
GC_5_477 b_5 NI_5 NS_477 0 -4.3685064029532823e-04
GC_5_478 b_5 NI_5 NS_478 0 -4.4075101080811772e-04
GC_5_479 b_5 NI_5 NS_479 0 -1.4473566013818991e-04
GC_5_480 b_5 NI_5 NS_480 0 6.2679330690239759e-05
GC_5_481 b_5 NI_5 NS_481 0 -6.6117468612336095e-03
GC_5_482 b_5 NI_5 NS_482 0 -1.9570618735265050e-03
GC_5_483 b_5 NI_5 NS_483 0 4.4554872793219487e-05
GC_5_484 b_5 NI_5 NS_484 0 -4.4973188765054068e-05
GC_5_485 b_5 NI_5 NS_485 0 1.5725340361862436e-04
GC_5_486 b_5 NI_5 NS_486 0 8.0303519934894600e-04
GC_5_487 b_5 NI_5 NS_487 0 1.9112785606036201e-03
GC_5_488 b_5 NI_5 NS_488 0 -3.3766263260940369e-03
GC_5_489 b_5 NI_5 NS_489 0 1.7647765384315659e-04
GC_5_490 b_5 NI_5 NS_490 0 -7.0996282362690923e-05
GC_5_491 b_5 NI_5 NS_491 0 8.5063809165218610e-07
GC_5_492 b_5 NI_5 NS_492 0 1.0260547196361037e-06
GC_5_493 b_5 NI_5 NS_493 0 -9.2011063650423895e-07
GC_5_494 b_5 NI_5 NS_494 0 -4.4139528966129162e-06
GC_5_495 b_5 NI_5 NS_495 0 -7.0792848735296097e-05
GC_5_496 b_5 NI_5 NS_496 0 8.2935389400451748e-05
GC_5_497 b_5 NI_5 NS_497 0 -1.2442848322465373e-06
GC_5_498 b_5 NI_5 NS_498 0 -1.0140729101522833e-05
GC_5_499 b_5 NI_5 NS_499 0 -8.8664765604989586e-06
GC_5_500 b_5 NI_5 NS_500 0 3.3726463339194504e-06
GC_5_501 b_5 NI_5 NS_501 0 3.5762710489386950e-06
GC_5_502 b_5 NI_5 NS_502 0 -3.0691973680875193e-05
GC_5_503 b_5 NI_5 NS_503 0 -1.8496310141822279e-05
GC_5_504 b_5 NI_5 NS_504 0 4.4777898608903890e-05
GC_5_505 b_5 NI_5 NS_505 0 4.2544668957221676e-03
GC_5_506 b_5 NI_5 NS_506 0 -1.5443046706469695e-04
GC_5_507 b_5 NI_5 NS_507 0 2.7491875380055293e-04
GC_5_508 b_5 NI_5 NS_508 0 4.0106081381718022e-04
GC_5_509 b_5 NI_5 NS_509 0 -4.0779553367950946e-04
GC_5_510 b_5 NI_5 NS_510 0 2.2118047267543400e-04
GC_5_511 b_5 NI_5 NS_511 0 -1.4752092672482217e-03
GC_5_512 b_5 NI_5 NS_512 0 2.6979182414053334e-04
GC_5_513 b_5 NI_5 NS_513 0 -2.0291881528263243e-04
GC_5_514 b_5 NI_5 NS_514 0 -1.5814109058515170e-03
GC_5_515 b_5 NI_5 NS_515 0 2.1029624196141440e-04
GC_5_516 b_5 NI_5 NS_516 0 -2.8561516050730831e-04
GC_5_517 b_5 NI_5 NS_517 0 7.6273789845756799e-04
GC_5_518 b_5 NI_5 NS_518 0 -1.3190960804604700e-03
GC_5_519 b_5 NI_5 NS_519 0 1.0559651510436705e-03
GC_5_520 b_5 NI_5 NS_520 0 -6.1186043302756551e-04
GC_5_521 b_5 NI_5 NS_521 0 1.8188896722731540e-03
GC_5_522 b_5 NI_5 NS_522 0 2.1969489463263686e-03
GC_5_523 b_5 NI_5 NS_523 0 2.8228820553045119e-05
GC_5_524 b_5 NI_5 NS_524 0 3.0156984663805000e-03
GC_5_525 b_5 NI_5 NS_525 0 -3.6209655729794652e-04
GC_5_526 b_5 NI_5 NS_526 0 -2.8807158249168076e-05
GC_5_527 b_5 NI_5 NS_527 0 -2.9489487948157656e-03
GC_5_528 b_5 NI_5 NS_528 0 2.7203785654785991e-03
GC_5_529 b_5 NI_5 NS_529 0 3.0308276310638216e-04
GC_5_530 b_5 NI_5 NS_530 0 1.2537071708775672e-04
GC_5_531 b_5 NI_5 NS_531 0 -1.1205660743597295e-03
GC_5_532 b_5 NI_5 NS_532 0 2.2777945632469578e-04
GC_5_533 b_5 NI_5 NS_533 0 -6.5935645526805334e-04
GC_5_534 b_5 NI_5 NS_534 0 -2.4125327041803612e-05
GC_5_535 b_5 NI_5 NS_535 0 -1.4276108105348612e-04
GC_5_536 b_5 NI_5 NS_536 0 -5.0736650302146710e-05
GC_5_537 b_5 NI_5 NS_537 0 -9.6744724006084828e-05
GC_5_538 b_5 NI_5 NS_538 0 -4.7231635945829444e-03
GC_5_539 b_5 NI_5 NS_539 0 4.2607035722510576e-05
GC_5_540 b_5 NI_5 NS_540 0 -3.7792238035515479e-05
GC_5_541 b_5 NI_5 NS_541 0 -1.3105691515021270e-03
GC_5_542 b_5 NI_5 NS_542 0 5.5786216832441539e-04
GC_5_543 b_5 NI_5 NS_543 0 1.3155187617922483e-03
GC_5_544 b_5 NI_5 NS_544 0 -9.1643286886804144e-04
GC_5_545 b_5 NI_5 NS_545 0 -2.0428730230646506e-04
GC_5_546 b_5 NI_5 NS_546 0 8.0900192290243300e-05
GC_5_547 b_5 NI_5 NS_547 0 -7.7688516862456611e-07
GC_5_548 b_5 NI_5 NS_548 0 4.5650177089736916e-07
GC_5_549 b_5 NI_5 NS_549 0 -3.7809858369717807e-06
GC_5_550 b_5 NI_5 NS_550 0 -3.8835458510548324e-06
GC_5_551 b_5 NI_5 NS_551 0 -1.4841467840580382e-05
GC_5_552 b_5 NI_5 NS_552 0 6.4721694250394890e-05
GC_5_553 b_5 NI_5 NS_553 0 -9.0379234276820138e-06
GC_5_554 b_5 NI_5 NS_554 0 -5.8936089068786346e-06
GC_5_555 b_5 NI_5 NS_555 0 -4.7958612919862203e-06
GC_5_556 b_5 NI_5 NS_556 0 -4.4997406697481998e-06
GC_5_557 b_5 NI_5 NS_557 0 2.5692452596784524e-05
GC_5_558 b_5 NI_5 NS_558 0 -4.7797270674116811e-06
GC_5_559 b_5 NI_5 NS_559 0 -3.9493385349338664e-05
GC_5_560 b_5 NI_5 NS_560 0 -5.0474370656716838e-06
GC_5_561 b_5 NI_5 NS_561 0 6.9540425455901205e-04
GC_5_562 b_5 NI_5 NS_562 0 3.7827142030631311e-05
GC_5_563 b_5 NI_5 NS_563 0 1.2320224963636272e-03
GC_5_564 b_5 NI_5 NS_564 0 -1.3867989218284174e-04
GC_5_565 b_5 NI_5 NS_565 0 -1.1142250211358408e-03
GC_5_566 b_5 NI_5 NS_566 0 1.2983303305713295e-03
GC_5_567 b_5 NI_5 NS_567 0 -9.6308678339309696e-04
GC_5_568 b_5 NI_5 NS_568 0 7.1189469755260511e-04
GC_5_569 b_5 NI_5 NS_569 0 -2.7560385552192089e-03
GC_5_570 b_5 NI_5 NS_570 0 -3.0180073072404792e-03
GC_5_571 b_5 NI_5 NS_571 0 7.1991113399852180e-05
GC_5_572 b_5 NI_5 NS_572 0 -3.2740676926037830e-04
GC_5_573 b_5 NI_5 NS_573 0 2.8165679566524975e-03
GC_5_574 b_5 NI_5 NS_574 0 -1.5940867371301239e-03
GC_5_575 b_5 NI_5 NS_575 0 1.2681648474038912e-03
GC_5_576 b_5 NI_5 NS_576 0 5.1741972193926973e-04
GC_5_577 b_5 NI_5 NS_577 0 -1.3086168403006633e-03
GC_5_578 b_5 NI_5 NS_578 0 4.1156243806505614e-05
GC_5_579 b_5 NI_5 NS_579 0 1.6315819060569998e-03
GC_5_580 b_5 NI_5 NS_580 0 2.4417841598107565e-04
GC_5_581 b_5 NI_5 NS_581 0 4.8154138423239491e-04
GC_5_582 b_5 NI_5 NS_582 0 2.3802634626408098e-04
GC_5_583 b_5 NI_5 NS_583 0 2.1978262805187975e-04
GC_5_584 b_5 NI_5 NS_584 0 5.1342982039368880e-03
GC_5_585 b_5 NI_5 NS_585 0 -3.5469528466659502e-04
GC_5_586 b_5 NI_5 NS_586 0 -6.9365270423736418e-04
GC_5_587 b_5 NI_5 NS_587 0 -8.5901182367213432e-04
GC_5_588 b_5 NI_5 NS_588 0 4.5141393768456806e-05
GC_5_589 b_5 NI_5 NS_589 0 -3.3081418827198927e-04
GC_5_590 b_5 NI_5 NS_590 0 -2.7724700131748946e-04
GC_5_591 b_5 NI_5 NS_591 0 -8.3390310497796419e-05
GC_5_592 b_5 NI_5 NS_592 0 1.0532477204682679e-05
GC_5_593 b_5 NI_5 NS_593 0 -3.4380354148340611e-03
GC_5_594 b_5 NI_5 NS_594 0 -4.7631109611792786e-03
GC_5_595 b_5 NI_5 NS_595 0 2.7475111373256263e-05
GC_5_596 b_5 NI_5 NS_596 0 -5.1795565347348093e-05
GC_5_597 b_5 NI_5 NS_597 0 8.5947956264086927e-05
GC_5_598 b_5 NI_5 NS_598 0 7.8708984805025972e-04
GC_5_599 b_5 NI_5 NS_599 0 2.4790519629053036e-03
GC_5_600 b_5 NI_5 NS_600 0 6.8932619862987186e-04
GC_5_601 b_5 NI_5 NS_601 0 6.0240482963489692e-06
GC_5_602 b_5 NI_5 NS_602 0 3.2036882985159252e-04
GC_5_603 b_5 NI_5 NS_603 0 -8.7571341875527261e-07
GC_5_604 b_5 NI_5 NS_604 0 1.3609419016381165e-06
GC_5_605 b_5 NI_5 NS_605 0 3.2215924590736161e-06
GC_5_606 b_5 NI_5 NS_606 0 -3.3715884641142035e-06
GC_5_607 b_5 NI_5 NS_607 0 -1.0089361858062486e-04
GC_5_608 b_5 NI_5 NS_608 0 1.0649943054181901e-05
GC_5_609 b_5 NI_5 NS_609 0 7.1766640123985999e-06
GC_5_610 b_5 NI_5 NS_610 0 -5.2838506003107712e-06
GC_5_611 b_5 NI_5 NS_611 0 -6.8823445024146955e-06
GC_5_612 b_5 NI_5 NS_612 0 -5.4896806309357456e-06
GC_5_613 b_5 NI_5 NS_613 0 2.1866444239374423e-05
GC_5_614 b_5 NI_5 NS_614 0 -6.6659371105809843e-06
GC_5_615 b_5 NI_5 NS_615 0 -3.5631842337854163e-05
GC_5_616 b_5 NI_5 NS_616 0 7.4023037366239351e-07
GC_5_617 b_5 NI_5 NS_617 0 6.3396374328870330e-03
GC_5_618 b_5 NI_5 NS_618 0 -8.1728957910187817e-05
GC_5_619 b_5 NI_5 NS_619 0 -2.0144037165731476e-04
GC_5_620 b_5 NI_5 NS_620 0 7.0102362090007132e-04
GC_5_621 b_5 NI_5 NS_621 0 -3.1311903075118762e-04
GC_5_622 b_5 NI_5 NS_622 0 -6.9060723758360197e-04
GC_5_623 b_5 NI_5 NS_623 0 -5.2943903449673580e-04
GC_5_624 b_5 NI_5 NS_624 0 -8.6696463104387960e-04
GC_5_625 b_5 NI_5 NS_625 0 2.3194356980047459e-03
GC_5_626 b_5 NI_5 NS_626 0 6.6953672877149745e-04
GC_5_627 b_5 NI_5 NS_627 0 -6.5911680172538840e-04
GC_5_628 b_5 NI_5 NS_628 0 1.9484605949642610e-05
GC_5_629 b_5 NI_5 NS_629 0 4.5461546906664909e-04
GC_5_630 b_5 NI_5 NS_630 0 -4.8104261053511958e-04
GC_5_631 b_5 NI_5 NS_631 0 8.5903802954767541e-04
GC_5_632 b_5 NI_5 NS_632 0 -1.1629004717215304e-04
GC_5_633 b_5 NI_5 NS_633 0 6.7811457395313107e-04
GC_5_634 b_5 NI_5 NS_634 0 1.8218282808837177e-03
GC_5_635 b_5 NI_5 NS_635 0 -1.1267491850531872e-03
GC_5_636 b_5 NI_5 NS_636 0 2.5099798084032344e-03
GC_5_637 b_5 NI_5 NS_637 0 -2.0588961261730940e-04
GC_5_638 b_5 NI_5 NS_638 0 -5.3756855947519431e-05
GC_5_639 b_5 NI_5 NS_639 0 -6.4914850498560867e-04
GC_5_640 b_5 NI_5 NS_640 0 1.2846365322563915e-03
GC_5_641 b_5 NI_5 NS_641 0 3.0226115599134904e-05
GC_5_642 b_5 NI_5 NS_642 0 -2.2046284521170108e-05
GC_5_643 b_5 NI_5 NS_643 0 -6.6066231870579950e-04
GC_5_644 b_5 NI_5 NS_644 0 1.0574583008083859e-04
GC_5_645 b_5 NI_5 NS_645 0 -3.8210948574545460e-04
GC_5_646 b_5 NI_5 NS_646 0 4.5381661684520589e-05
GC_5_647 b_5 NI_5 NS_647 0 -1.0256425862845390e-04
GC_5_648 b_5 NI_5 NS_648 0 -3.9347875639281930e-05
GC_5_649 b_5 NI_5 NS_649 0 -5.7161204691478337e-05
GC_5_650 b_5 NI_5 NS_650 0 -2.6254042120012191e-03
GC_5_651 b_5 NI_5 NS_651 0 3.0917671705266979e-05
GC_5_652 b_5 NI_5 NS_652 0 -1.2756421451882390e-05
GC_5_653 b_5 NI_5 NS_653 0 -8.0844593578417213e-04
GC_5_654 b_5 NI_5 NS_654 0 3.6289713315849036e-04
GC_5_655 b_5 NI_5 NS_655 0 6.7660733409605038e-04
GC_5_656 b_5 NI_5 NS_656 0 4.6428108230074557e-04
GC_5_657 b_5 NI_5 NS_657 0 -1.5657969409611086e-04
GC_5_658 b_5 NI_5 NS_658 0 2.6270286674298096e-04
GC_5_659 b_5 NI_5 NS_659 0 -1.1175792809272251e-06
GC_5_660 b_5 NI_5 NS_660 0 4.9603348190359781e-07
GC_5_661 b_5 NI_5 NS_661 0 -6.1675786960312475e-07
GC_5_662 b_5 NI_5 NS_662 0 -5.0943520818239234e-06
GC_5_663 b_5 NI_5 NS_663 0 -1.6473284937289038e-06
GC_5_664 b_5 NI_5 NS_664 0 4.5927091941165784e-05
GC_5_665 b_5 NI_5 NS_665 0 -2.1796196280801462e-06
GC_5_666 b_5 NI_5 NS_666 0 -8.7083990521288370e-06
GC_5_667 b_5 NI_5 NS_667 0 -6.3290605740792056e-06
GC_5_668 b_5 NI_5 NS_668 0 -5.0551545479281091e-06
GC_5_669 b_5 NI_5 NS_669 0 2.2071775737077811e-05
GC_5_670 b_5 NI_5 NS_670 0 -1.1128590064090202e-05
GC_5_671 b_5 NI_5 NS_671 0 -3.8275351949699075e-05
GC_5_672 b_5 NI_5 NS_672 0 5.6072180722648661e-06
GD_5_1 b_5 NI_5 NA_1 0 -4.3599531985789163e-02
GD_5_2 b_5 NI_5 NA_2 0 2.9162948474715008e-03
GD_5_3 b_5 NI_5 NA_3 0 -6.6182539289799391e-02
GD_5_4 b_5 NI_5 NA_4 0 -2.1846663069386183e-02
GD_5_5 b_5 NI_5 NA_5 0 -1.6004991397018645e-01
GD_5_6 b_5 NI_5 NA_6 0 4.3724307229779942e-02
GD_5_7 b_5 NI_5 NA_7 0 -8.8798903932904502e-03
GD_5_8 b_5 NI_5 NA_8 0 -5.3666768120784872e-02
GD_5_9 b_5 NI_5 NA_9 0 -1.8740733839903729e-02
GD_5_10 b_5 NI_5 NA_10 0 -9.6464049561319665e-05
GD_5_11 b_5 NI_5 NA_11 0 1.9851491321819863e-04
GD_5_12 b_5 NI_5 NA_12 0 -9.3557202206627377e-03
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 -6.3897974355501107e-03
GC_6_2 b_6 NI_6 NS_2 0 -2.5326893473829042e-04
GC_6_3 b_6 NI_6 NS_3 0 -1.3426740229845514e-03
GC_6_4 b_6 NI_6 NS_4 0 3.0615288795078355e-03
GC_6_5 b_6 NI_6 NS_5 0 -9.8183977847637362e-04
GC_6_6 b_6 NI_6 NS_6 0 -2.2450650996153820e-03
GC_6_7 b_6 NI_6 NS_7 0 -5.0728768600043312e-03
GC_6_8 b_6 NI_6 NS_8 0 -5.7632622973405696e-03
GC_6_9 b_6 NI_6 NS_9 0 7.2881496558383904e-03
GC_6_10 b_6 NI_6 NS_10 0 -1.4230082272110793e-03
GC_6_11 b_6 NI_6 NS_11 0 -3.1156989322414849e-04
GC_6_12 b_6 NI_6 NS_12 0 4.3384388254709324e-04
GC_6_13 b_6 NI_6 NS_13 0 4.2215432821102730e-03
GC_6_14 b_6 NI_6 NS_14 0 -2.5833428306951600e-03
GC_6_15 b_6 NI_6 NS_15 0 8.0837411603049754e-04
GC_6_16 b_6 NI_6 NS_16 0 1.1386264035179170e-03
GC_6_17 b_6 NI_6 NS_17 0 4.4334332003116868e-04
GC_6_18 b_6 NI_6 NS_18 0 2.1270323315511182e-03
GC_6_19 b_6 NI_6 NS_19 0 -3.1835499923505480e-03
GC_6_20 b_6 NI_6 NS_20 0 1.1322991748361532e-03
GC_6_21 b_6 NI_6 NS_21 0 -2.3049875329692892e-04
GC_6_22 b_6 NI_6 NS_22 0 3.3301933494867572e-05
GC_6_23 b_6 NI_6 NS_23 0 3.3068057230811378e-03
GC_6_24 b_6 NI_6 NS_24 0 -8.6570998081726203e-04
GC_6_25 b_6 NI_6 NS_25 0 -1.1627426536230860e-03
GC_6_26 b_6 NI_6 NS_26 0 -8.8280599746901273e-05
GC_6_27 b_6 NI_6 NS_27 0 -1.5568734989224810e-04
GC_6_28 b_6 NI_6 NS_28 0 8.3490840879550440e-05
GC_6_29 b_6 NI_6 NS_29 0 -3.1787777221402460e-04
GC_6_30 b_6 NI_6 NS_30 0 2.4792683837216009e-04
GC_6_31 b_6 NI_6 NS_31 0 -2.0513994572316212e-04
GC_6_32 b_6 NI_6 NS_32 0 -1.0639250177406126e-04
GC_6_33 b_6 NI_6 NS_33 0 2.5969343421769430e-03
GC_6_34 b_6 NI_6 NS_34 0 1.2344002523842356e-03
GC_6_35 b_6 NI_6 NS_35 0 -6.1292942481195608e-05
GC_6_36 b_6 NI_6 NS_36 0 1.4455674590553631e-04
GC_6_37 b_6 NI_6 NS_37 0 -3.7073854381347755e-04
GC_6_38 b_6 NI_6 NS_38 0 -1.0402169006620140e-03
GC_6_39 b_6 NI_6 NS_39 0 -7.5674654860357867e-04
GC_6_40 b_6 NI_6 NS_40 0 1.0343240174487344e-03
GC_6_41 b_6 NI_6 NS_41 0 -7.8345589653925949e-07
GC_6_42 b_6 NI_6 NS_42 0 -2.2586606462677558e-04
GC_6_43 b_6 NI_6 NS_43 0 2.1316300591049575e-06
GC_6_44 b_6 NI_6 NS_44 0 1.1252689307393486e-06
GC_6_45 b_6 NI_6 NS_45 0 2.5045368743098642e-06
GC_6_46 b_6 NI_6 NS_46 0 1.6565171746260310e-06
GC_6_47 b_6 NI_6 NS_47 0 1.1025839531438946e-04
GC_6_48 b_6 NI_6 NS_48 0 -2.9691556780891948e-05
GC_6_49 b_6 NI_6 NS_49 0 -4.9179546928250589e-06
GC_6_50 b_6 NI_6 NS_50 0 1.9215066764768035e-06
GC_6_51 b_6 NI_6 NS_51 0 1.1896375179735152e-05
GC_6_52 b_6 NI_6 NS_52 0 -1.0032959266300238e-06
GC_6_53 b_6 NI_6 NS_53 0 -2.2105309166194161e-05
GC_6_54 b_6 NI_6 NS_54 0 1.6304046014973890e-05
GC_6_55 b_6 NI_6 NS_55 0 3.8049426923109821e-05
GC_6_56 b_6 NI_6 NS_56 0 -6.5227122792226786e-06
GC_6_57 b_6 NI_6 NS_57 0 1.2032637891320740e-02
GC_6_58 b_6 NI_6 NS_58 0 -7.2270226862494041e-04
GC_6_59 b_6 NI_6 NS_59 0 -1.1910284465165759e-03
GC_6_60 b_6 NI_6 NS_60 0 -1.1286308443558650e-03
GC_6_61 b_6 NI_6 NS_61 0 9.9826007770340182e-04
GC_6_62 b_6 NI_6 NS_62 0 3.4854179319756889e-04
GC_6_63 b_6 NI_6 NS_63 0 4.5306469299303334e-03
GC_6_64 b_6 NI_6 NS_64 0 1.2211091454242095e-03
GC_6_65 b_6 NI_6 NS_65 0 -6.6820236634058464e-03
GC_6_66 b_6 NI_6 NS_66 0 3.5747103329925420e-03
GC_6_67 b_6 NI_6 NS_67 0 -1.6137197653010897e-04
GC_6_68 b_6 NI_6 NS_68 0 6.3875543864629146e-04
GC_6_69 b_6 NI_6 NS_69 0 3.8026641850379613e-05
GC_6_70 b_6 NI_6 NS_70 0 -3.6917289180751168e-03
GC_6_71 b_6 NI_6 NS_71 0 8.0985043945402979e-04
GC_6_72 b_6 NI_6 NS_72 0 4.8595397565351134e-04
GC_6_73 b_6 NI_6 NS_73 0 1.5118653123384826e-04
GC_6_74 b_6 NI_6 NS_74 0 1.5726199271828389e-03
GC_6_75 b_6 NI_6 NS_75 0 1.2904708773205037e-03
GC_6_76 b_6 NI_6 NS_76 0 -1.5030878472648938e-03
GC_6_77 b_6 NI_6 NS_77 0 9.3449949980510007e-05
GC_6_78 b_6 NI_6 NS_78 0 -1.9605129454013796e-05
GC_6_79 b_6 NI_6 NS_79 0 5.6161683856409167e-04
GC_6_80 b_6 NI_6 NS_80 0 2.5506483565828761e-03
GC_6_81 b_6 NI_6 NS_81 0 3.2641404145840189e-04
GC_6_82 b_6 NI_6 NS_82 0 1.0814512994659079e-04
GC_6_83 b_6 NI_6 NS_83 0 -1.7961350877259682e-04
GC_6_84 b_6 NI_6 NS_84 0 -4.0826359738068434e-05
GC_6_85 b_6 NI_6 NS_85 0 1.2862152786597734e-04
GC_6_86 b_6 NI_6 NS_86 0 -2.6556661984781079e-04
GC_6_87 b_6 NI_6 NS_87 0 3.4747760964606416e-04
GC_6_88 b_6 NI_6 NS_88 0 -1.4933843406635878e-04
GC_6_89 b_6 NI_6 NS_89 0 -1.5144877905476153e-02
GC_6_90 b_6 NI_6 NS_90 0 2.3793619515202783e-03
GC_6_91 b_6 NI_6 NS_91 0 -2.1725120545996147e-04
GC_6_92 b_6 NI_6 NS_92 0 -2.8037863194058712e-04
GC_6_93 b_6 NI_6 NS_93 0 4.4112449348023882e-03
GC_6_94 b_6 NI_6 NS_94 0 1.4099792854984283e-03
GC_6_95 b_6 NI_6 NS_95 0 6.8708671874466694e-03
GC_6_96 b_6 NI_6 NS_96 0 -5.2392284240832055e-03
GC_6_97 b_6 NI_6 NS_97 0 1.1178129382874915e-03
GC_6_98 b_6 NI_6 NS_98 0 1.3642544628398548e-04
GC_6_99 b_6 NI_6 NS_99 0 -1.8415218408556629e-07
GC_6_100 b_6 NI_6 NS_100 0 -4.9394087234017859e-06
GC_6_101 b_6 NI_6 NS_101 0 -4.1493492266969074e-05
GC_6_102 b_6 NI_6 NS_102 0 -3.9763491122351126e-05
GC_6_103 b_6 NI_6 NS_103 0 -3.7080463241743848e-04
GC_6_104 b_6 NI_6 NS_104 0 3.3286600653242317e-04
GC_6_105 b_6 NI_6 NS_105 0 -5.4693408707160976e-05
GC_6_106 b_6 NI_6 NS_106 0 -5.5405343873106804e-05
GC_6_107 b_6 NI_6 NS_107 0 -4.9200192694162740e-05
GC_6_108 b_6 NI_6 NS_108 0 -1.0547459974037342e-05
GC_6_109 b_6 NI_6 NS_109 0 3.0569263639514138e-04
GC_6_110 b_6 NI_6 NS_110 0 -2.8722204617331334e-04
GC_6_111 b_6 NI_6 NS_111 0 -5.6334344393858620e-04
GC_6_112 b_6 NI_6 NS_112 0 2.8088331574917762e-04
GC_6_113 b_6 NI_6 NS_113 0 2.6597972873199240e-02
GC_6_114 b_6 NI_6 NS_114 0 -8.3746175878914768e-04
GC_6_115 b_6 NI_6 NS_115 0 -1.8272418774961214e-03
GC_6_116 b_6 NI_6 NS_116 0 3.8984134861736381e-03
GC_6_117 b_6 NI_6 NS_117 0 1.0402788885111791e-03
GC_6_118 b_6 NI_6 NS_118 0 -3.2871410829326820e-04
GC_6_119 b_6 NI_6 NS_119 0 -9.8877834306805527e-03
GC_6_120 b_6 NI_6 NS_120 0 -3.7811999428784600e-03
GC_6_121 b_6 NI_6 NS_121 0 -1.5496381115084636e-03
GC_6_122 b_6 NI_6 NS_122 0 2.3303385167877159e-03
GC_6_123 b_6 NI_6 NS_123 0 -4.1464690174630167e-04
GC_6_124 b_6 NI_6 NS_124 0 -2.4631858875464708e-05
GC_6_125 b_6 NI_6 NS_125 0 5.6562834173213006e-03
GC_6_126 b_6 NI_6 NS_126 0 -6.1506372459045697e-03
GC_6_127 b_6 NI_6 NS_127 0 1.1720249732532118e-03
GC_6_128 b_6 NI_6 NS_128 0 1.7308458933909870e-03
GC_6_129 b_6 NI_6 NS_129 0 4.7278939376157217e-04
GC_6_130 b_6 NI_6 NS_130 0 1.8533894887244630e-03
GC_6_131 b_6 NI_6 NS_131 0 -5.0851002786954647e-03
GC_6_132 b_6 NI_6 NS_132 0 1.5509155084316638e-04
GC_6_133 b_6 NI_6 NS_133 0 -2.3040988039788488e-04
GC_6_134 b_6 NI_6 NS_134 0 -2.7503614059939287e-05
GC_6_135 b_6 NI_6 NS_135 0 2.4868171775595999e-03
GC_6_136 b_6 NI_6 NS_136 0 2.8878410974216896e-03
GC_6_137 b_6 NI_6 NS_137 0 -1.1638277521313219e-03
GC_6_138 b_6 NI_6 NS_138 0 -1.4323730973363750e-04
GC_6_139 b_6 NI_6 NS_139 0 -3.9402696983477115e-04
GC_6_140 b_6 NI_6 NS_140 0 6.4033254267449938e-05
GC_6_141 b_6 NI_6 NS_141 0 -5.7285674020416321e-04
GC_6_142 b_6 NI_6 NS_142 0 5.0309144512027300e-04
GC_6_143 b_6 NI_6 NS_143 0 -3.5340939021313286e-04
GC_6_144 b_6 NI_6 NS_144 0 -1.2701656279973252e-04
GC_6_145 b_6 NI_6 NS_145 0 -6.1998991961537662e-04
GC_6_146 b_6 NI_6 NS_146 0 -8.3127016707978572e-04
GC_6_147 b_6 NI_6 NS_147 0 -3.7576784602017946e-05
GC_6_148 b_6 NI_6 NS_148 0 1.6148703380106154e-04
GC_6_149 b_6 NI_6 NS_149 0 -7.1504344039808763e-04
GC_6_150 b_6 NI_6 NS_150 0 -5.5142715209515641e-04
GC_6_151 b_6 NI_6 NS_151 0 -1.0252926936768062e-03
GC_6_152 b_6 NI_6 NS_152 0 -9.6717133989675404e-04
GC_6_153 b_6 NI_6 NS_153 0 5.6909722820694839e-05
GC_6_154 b_6 NI_6 NS_154 0 -7.7398421223092532e-05
GC_6_155 b_6 NI_6 NS_155 0 1.4545001979742871e-06
GC_6_156 b_6 NI_6 NS_156 0 1.8107271753119784e-07
GC_6_157 b_6 NI_6 NS_157 0 -3.1829227494648007e-06
GC_6_158 b_6 NI_6 NS_158 0 4.6012058864503603e-06
GC_6_159 b_6 NI_6 NS_159 0 6.1819659496273292e-05
GC_6_160 b_6 NI_6 NS_160 0 1.3721932439979825e-05
GC_6_161 b_6 NI_6 NS_161 0 -5.1515587828568870e-06
GC_6_162 b_6 NI_6 NS_162 0 5.3360972908134910e-06
GC_6_163 b_6 NI_6 NS_163 0 1.0608991544031773e-06
GC_6_164 b_6 NI_6 NS_164 0 2.1639646630718277e-06
GC_6_165 b_6 NI_6 NS_165 0 -2.5173884000866439e-05
GC_6_166 b_6 NI_6 NS_166 0 -1.9972854348854508e-05
GC_6_167 b_6 NI_6 NS_167 0 2.2885449489094574e-05
GC_6_168 b_6 NI_6 NS_168 0 3.8354284660467587e-05
GC_6_169 b_6 NI_6 NS_169 0 5.2611173123535988e-03
GC_6_170 b_6 NI_6 NS_170 0 -1.4446755189502954e-03
GC_6_171 b_6 NI_6 NS_171 0 -1.5058079172474142e-03
GC_6_172 b_6 NI_6 NS_172 0 -1.4352623017342204e-03
GC_6_173 b_6 NI_6 NS_173 0 -3.9263870268664200e-04
GC_6_174 b_6 NI_6 NS_174 0 8.0826351442854190e-04
GC_6_175 b_6 NI_6 NS_175 0 4.7945383371966388e-03
GC_6_176 b_6 NI_6 NS_176 0 -4.7617583962480335e-04
GC_6_177 b_6 NI_6 NS_177 0 -3.9753895549601848e-03
GC_6_178 b_6 NI_6 NS_178 0 -1.7587520754717050e-03
GC_6_179 b_6 NI_6 NS_179 0 -1.3886792395772699e-04
GC_6_180 b_6 NI_6 NS_180 0 7.2685637820553916e-04
GC_6_181 b_6 NI_6 NS_181 0 9.1338579209281339e-04
GC_6_182 b_6 NI_6 NS_182 0 -2.7491081364146974e-03
GC_6_183 b_6 NI_6 NS_183 0 1.0979251236180288e-03
GC_6_184 b_6 NI_6 NS_184 0 6.0131867554968910e-04
GC_6_185 b_6 NI_6 NS_185 0 9.0939266746659152e-04
GC_6_186 b_6 NI_6 NS_186 0 1.1361251319718540e-03
GC_6_187 b_6 NI_6 NS_187 0 1.7045646241883384e-03
GC_6_188 b_6 NI_6 NS_188 0 -2.4860657744294511e-03
GC_6_189 b_6 NI_6 NS_189 0 9.7859251360304966e-05
GC_6_190 b_6 NI_6 NS_190 0 -5.8372778425853063e-05
GC_6_191 b_6 NI_6 NS_191 0 3.5051835049566462e-03
GC_6_192 b_6 NI_6 NS_192 0 5.0803000828510214e-03
GC_6_193 b_6 NI_6 NS_193 0 3.3688937898263926e-04
GC_6_194 b_6 NI_6 NS_194 0 -1.5566461415075354e-05
GC_6_195 b_6 NI_6 NS_195 0 -2.3857886335995967e-04
GC_6_196 b_6 NI_6 NS_196 0 -1.6350139985961006e-07
GC_6_197 b_6 NI_6 NS_197 0 1.9882301834673764e-04
GC_6_198 b_6 NI_6 NS_198 0 -1.9992883678408588e-04
GC_6_199 b_6 NI_6 NS_199 0 3.6454801651637981e-04
GC_6_200 b_6 NI_6 NS_200 0 -9.7169942370140192e-05
GC_6_201 b_6 NI_6 NS_201 0 -1.5278548446071927e-02
GC_6_202 b_6 NI_6 NS_202 0 1.8372239903478144e-03
GC_6_203 b_6 NI_6 NS_203 0 -2.2191141534569288e-04
GC_6_204 b_6 NI_6 NS_204 0 -3.1094019685644076e-04
GC_6_205 b_6 NI_6 NS_205 0 4.7744086698173665e-03
GC_6_206 b_6 NI_6 NS_206 0 1.9067385497160863e-03
GC_6_207 b_6 NI_6 NS_207 0 5.4014192378224451e-03
GC_6_208 b_6 NI_6 NS_208 0 -4.1644053390039355e-03
GC_6_209 b_6 NI_6 NS_209 0 1.1613846415989976e-03
GC_6_210 b_6 NI_6 NS_210 0 3.7782698335562587e-04
GC_6_211 b_6 NI_6 NS_211 0 -3.3728978004512149e-06
GC_6_212 b_6 NI_6 NS_212 0 -2.8875224737233763e-06
GC_6_213 b_6 NI_6 NS_213 0 -3.7912087523907256e-05
GC_6_214 b_6 NI_6 NS_214 0 -3.3743935094598493e-05
GC_6_215 b_6 NI_6 NS_215 0 -2.3296012894840978e-04
GC_6_216 b_6 NI_6 NS_216 0 2.1070988092934887e-04
GC_6_217 b_6 NI_6 NS_217 0 -5.5623602755966605e-05
GC_6_218 b_6 NI_6 NS_218 0 -4.1523025595025220e-05
GC_6_219 b_6 NI_6 NS_219 0 -3.6381468076485655e-05
GC_6_220 b_6 NI_6 NS_220 0 -1.2374187497496625e-05
GC_6_221 b_6 NI_6 NS_221 0 2.9572101839388010e-04
GC_6_222 b_6 NI_6 NS_222 0 -2.2809499656841763e-04
GC_6_223 b_6 NI_6 NS_223 0 -5.2276230576959212e-04
GC_6_224 b_6 NI_6 NS_224 0 1.9857930666271730e-04
GC_6_225 b_6 NI_6 NS_225 0 -4.5241116662555293e-02
GC_6_226 b_6 NI_6 NS_226 0 1.2126658278099084e-02
GC_6_227 b_6 NI_6 NS_227 0 -2.9182380150428971e-03
GC_6_228 b_6 NI_6 NS_228 0 3.7386200421144749e-03
GC_6_229 b_6 NI_6 NS_229 0 -4.3699494200615538e-03
GC_6_230 b_6 NI_6 NS_230 0 2.1341984242379004e-03
GC_6_231 b_6 NI_6 NS_231 0 -4.8443222586382027e-03
GC_6_232 b_6 NI_6 NS_232 0 -9.2083972724343547e-03
GC_6_233 b_6 NI_6 NS_233 0 -2.5373822466301706e-03
GC_6_234 b_6 NI_6 NS_234 0 -9.1021251796622529e-03
GC_6_235 b_6 NI_6 NS_235 0 6.2227033389343728e-04
GC_6_236 b_6 NI_6 NS_236 0 -1.4884668504813606e-04
GC_6_237 b_6 NI_6 NS_237 0 7.1329857603946219e-03
GC_6_238 b_6 NI_6 NS_238 0 -1.5514971393661820e-03
GC_6_239 b_6 NI_6 NS_239 0 1.5062842471312370e-03
GC_6_240 b_6 NI_6 NS_240 0 1.2893696660307705e-03
GC_6_241 b_6 NI_6 NS_241 0 5.4266406598088551e-03
GC_6_242 b_6 NI_6 NS_242 0 8.8710843935299643e-04
GC_6_243 b_6 NI_6 NS_243 0 -2.4576939074685100e-03
GC_6_244 b_6 NI_6 NS_244 0 1.1536036147647912e-03
GC_6_245 b_6 NI_6 NS_245 0 -3.6616848217794167e-04
GC_6_246 b_6 NI_6 NS_246 0 6.6445525464088167e-05
GC_6_247 b_6 NI_6 NS_247 0 7.7434764618211256e-03
GC_6_248 b_6 NI_6 NS_248 0 -2.6957583583794697e-03
GC_6_249 b_6 NI_6 NS_249 0 -1.7229508288888460e-03
GC_6_250 b_6 NI_6 NS_250 0 -2.1719262819543259e-05
GC_6_251 b_6 NI_6 NS_251 0 -2.7488932855736784e-04
GC_6_252 b_6 NI_6 NS_252 0 1.1878239739588959e-04
GC_6_253 b_6 NI_6 NS_253 0 -4.4658033831650710e-04
GC_6_254 b_6 NI_6 NS_254 0 4.1411167515914684e-04
GC_6_255 b_6 NI_6 NS_255 0 -3.0504463051364821e-04
GC_6_256 b_6 NI_6 NS_256 0 -1.1496658241065375e-04
GC_6_257 b_6 NI_6 NS_257 0 2.5842525410578582e-03
GC_6_258 b_6 NI_6 NS_258 0 -9.3118434286859056e-04
GC_6_259 b_6 NI_6 NS_259 0 -2.1793291717698655e-05
GC_6_260 b_6 NI_6 NS_260 0 1.7615227736194150e-04
GC_6_261 b_6 NI_6 NS_261 0 -9.5410186382302239e-04
GC_6_262 b_6 NI_6 NS_262 0 -8.8012865131508594e-04
GC_6_263 b_6 NI_6 NS_263 0 2.0326240592959486e-03
GC_6_264 b_6 NI_6 NS_264 0 1.2709729702061305e-03
GC_6_265 b_6 NI_6 NS_265 0 -1.2196516446979658e-04
GC_6_266 b_6 NI_6 NS_266 0 -1.5991032327936029e-04
GC_6_267 b_6 NI_6 NS_267 0 1.5547146297027715e-06
GC_6_268 b_6 NI_6 NS_268 0 -2.0148889242618869e-06
GC_6_269 b_6 NI_6 NS_269 0 2.5672981642926102e-06
GC_6_270 b_6 NI_6 NS_270 0 -2.5943822856504625e-06
GC_6_271 b_6 NI_6 NS_271 0 -7.1253127114792166e-05
GC_6_272 b_6 NI_6 NS_272 0 -6.3391827172810854e-05
GC_6_273 b_6 NI_6 NS_273 0 8.9353398905816426e-06
GC_6_274 b_6 NI_6 NS_274 0 1.7795412370263578e-06
GC_6_275 b_6 NI_6 NS_275 0 1.1846592981844321e-06
GC_6_276 b_6 NI_6 NS_276 0 -9.5678934487099452e-06
GC_6_277 b_6 NI_6 NS_277 0 2.3925003922109865e-05
GC_6_278 b_6 NI_6 NS_278 0 5.1828102197169150e-05
GC_6_279 b_6 NI_6 NS_279 0 -9.3275785469453220e-06
GC_6_280 b_6 NI_6 NS_280 0 -9.0459409327877917e-05
GC_6_281 b_6 NI_6 NS_281 0 -7.0221195990799470e-02
GC_6_282 b_6 NI_6 NS_282 0 7.7287865068711168e-03
GC_6_283 b_6 NI_6 NS_283 0 -1.1468598097740387e-03
GC_6_284 b_6 NI_6 NS_284 0 -1.9281462042801322e-03
GC_6_285 b_6 NI_6 NS_285 0 5.4000021940564103e-05
GC_6_286 b_6 NI_6 NS_286 0 -1.5107805040825695e-03
GC_6_287 b_6 NI_6 NS_287 0 6.0382734312435706e-03
GC_6_288 b_6 NI_6 NS_288 0 3.9066645447778181e-03
GC_6_289 b_6 NI_6 NS_289 0 3.4392357304708679e-03
GC_6_290 b_6 NI_6 NS_290 0 6.4176255080952167e-03
GC_6_291 b_6 NI_6 NS_291 0 6.3580842807799663e-04
GC_6_292 b_6 NI_6 NS_292 0 -4.6029903631664409e-04
GC_6_293 b_6 NI_6 NS_293 0 -1.7345318767350377e-03
GC_6_294 b_6 NI_6 NS_294 0 -5.5162055281232775e-03
GC_6_295 b_6 NI_6 NS_295 0 1.2128264263384099e-03
GC_6_296 b_6 NI_6 NS_296 0 6.2243912379950886e-04
GC_6_297 b_6 NI_6 NS_297 0 5.5680794663752454e-04
GC_6_298 b_6 NI_6 NS_298 0 7.0796176372456840e-04
GC_6_299 b_6 NI_6 NS_299 0 2.1434657025631984e-03
GC_6_300 b_6 NI_6 NS_300 0 -2.5831012900761042e-03
GC_6_301 b_6 NI_6 NS_301 0 1.5037744397198086e-04
GC_6_302 b_6 NI_6 NS_302 0 -7.1427707694032030e-05
GC_6_303 b_6 NI_6 NS_303 0 1.7330574023106363e-03
GC_6_304 b_6 NI_6 NS_304 0 5.4700212002679162e-03
GC_6_305 b_6 NI_6 NS_305 0 4.9894535029470545e-04
GC_6_306 b_6 NI_6 NS_306 0 9.9456208593305001e-06
GC_6_307 b_6 NI_6 NS_307 0 -4.1163406850591678e-04
GC_6_308 b_6 NI_6 NS_308 0 6.1096096365317418e-05
GC_6_309 b_6 NI_6 NS_309 0 1.0368867691638526e-04
GC_6_310 b_6 NI_6 NS_310 0 -2.9710034241006527e-04
GC_6_311 b_6 NI_6 NS_311 0 4.4277362839301225e-04
GC_6_312 b_6 NI_6 NS_312 0 -2.1028889162985604e-04
GC_6_313 b_6 NI_6 NS_313 0 -2.0499550123340361e-02
GC_6_314 b_6 NI_6 NS_314 0 1.9724831832668242e-03
GC_6_315 b_6 NI_6 NS_315 0 -2.9696788428571104e-04
GC_6_316 b_6 NI_6 NS_316 0 -3.8682747195160964e-04
GC_6_317 b_6 NI_6 NS_317 0 6.2209716601193052e-03
GC_6_318 b_6 NI_6 NS_318 0 2.1929631495115295e-03
GC_6_319 b_6 NI_6 NS_319 0 9.5415143774320484e-03
GC_6_320 b_6 NI_6 NS_320 0 -6.1346210356371528e-03
GC_6_321 b_6 NI_6 NS_321 0 1.5228725641527341e-03
GC_6_322 b_6 NI_6 NS_322 0 5.1721805341494224e-04
GC_6_323 b_6 NI_6 NS_323 0 -3.4453009419638390e-06
GC_6_324 b_6 NI_6 NS_324 0 -5.1893156461268684e-06
GC_6_325 b_6 NI_6 NS_325 0 -5.8966569205838467e-05
GC_6_326 b_6 NI_6 NS_326 0 -3.3885179162401832e-05
GC_6_327 b_6 NI_6 NS_327 0 -3.9058862712342999e-04
GC_6_328 b_6 NI_6 NS_328 0 2.2036006450497288e-04
GC_6_329 b_6 NI_6 NS_329 0 -6.7038391325446484e-05
GC_6_330 b_6 NI_6 NS_330 0 -3.8464342003035053e-05
GC_6_331 b_6 NI_6 NS_331 0 -6.7968322123646046e-05
GC_6_332 b_6 NI_6 NS_332 0 -2.8017396877024774e-05
GC_6_333 b_6 NI_6 NS_333 0 4.3673068514262181e-04
GC_6_334 b_6 NI_6 NS_334 0 -4.1536320568485638e-04
GC_6_335 b_6 NI_6 NS_335 0 -8.0801209502633423e-04
GC_6_336 b_6 NI_6 NS_336 0 4.0256071189161336e-04
GC_6_337 b_6 NI_6 NS_337 0 5.7573995023942726e-02
GC_6_338 b_6 NI_6 NS_338 0 -7.8908432183411004e-04
GC_6_339 b_6 NI_6 NS_339 0 -1.7550542069091327e-03
GC_6_340 b_6 NI_6 NS_340 0 2.3937903761521552e-03
GC_6_341 b_6 NI_6 NS_341 0 2.8923399177407357e-03
GC_6_342 b_6 NI_6 NS_342 0 2.8225286742782871e-04
GC_6_343 b_6 NI_6 NS_343 0 -5.6229684162300694e-03
GC_6_344 b_6 NI_6 NS_344 0 5.6045715252262007e-04
GC_6_345 b_6 NI_6 NS_345 0 -6.4091422020177711e-03
GC_6_346 b_6 NI_6 NS_346 0 1.0277525061076086e-02
GC_6_347 b_6 NI_6 NS_347 0 -5.3710528181329412e-04
GC_6_348 b_6 NI_6 NS_348 0 -2.6664432400759188e-04
GC_6_349 b_6 NI_6 NS_349 0 1.8473492048460588e-03
GC_6_350 b_6 NI_6 NS_350 0 -4.4300295537771303e-03
GC_6_351 b_6 NI_6 NS_351 0 1.0620724899402293e-03
GC_6_352 b_6 NI_6 NS_352 0 1.3769930609840006e-03
GC_6_353 b_6 NI_6 NS_353 0 -1.0672661250876091e-04
GC_6_354 b_6 NI_6 NS_354 0 1.2707692528954322e-03
GC_6_355 b_6 NI_6 NS_355 0 -5.9327847793131973e-03
GC_6_356 b_6 NI_6 NS_356 0 9.8778558334581602e-04
GC_6_357 b_6 NI_6 NS_357 0 -1.4813178555228470e-04
GC_6_358 b_6 NI_6 NS_358 0 -8.4416546535572536e-05
GC_6_359 b_6 NI_6 NS_359 0 1.0332063175602002e-03
GC_6_360 b_6 NI_6 NS_360 0 5.3252605127526069e-03
GC_6_361 b_6 NI_6 NS_361 0 -4.7987269228076207e-04
GC_6_362 b_6 NI_6 NS_362 0 -1.7923478726856177e-04
GC_6_363 b_6 NI_6 NS_363 0 -5.0274838507825619e-04
GC_6_364 b_6 NI_6 NS_364 0 7.2378405314032693e-05
GC_6_365 b_6 NI_6 NS_365 0 -4.4711456784797136e-04
GC_6_366 b_6 NI_6 NS_366 0 4.6474053763787075e-04
GC_6_367 b_6 NI_6 NS_367 0 -2.5256704698739844e-04
GC_6_368 b_6 NI_6 NS_368 0 -3.9026797580889770e-05
GC_6_369 b_6 NI_6 NS_369 0 -8.1484255062545131e-03
GC_6_370 b_6 NI_6 NS_370 0 -1.9148405400463144e-03
GC_6_371 b_6 NI_6 NS_371 0 -1.5473165649173515e-05
GC_6_372 b_6 NI_6 NS_372 0 3.6747395338755709e-05
GC_6_373 b_6 NI_6 NS_373 0 -8.7894504029356957e-05
GC_6_374 b_6 NI_6 NS_374 0 7.6916528992207239e-04
GC_6_375 b_6 NI_6 NS_375 0 9.0364342352851449e-05
GC_6_376 b_6 NI_6 NS_376 0 -2.9101782588587663e-03
GC_6_377 b_6 NI_6 NS_377 0 3.3469560357641165e-04
GC_6_378 b_6 NI_6 NS_378 0 2.3824812517143074e-04
GC_6_379 b_6 NI_6 NS_379 0 -4.7633284126463947e-07
GC_6_380 b_6 NI_6 NS_380 0 1.1738497303080073e-06
GC_6_381 b_6 NI_6 NS_381 0 -3.5728064173385826e-06
GC_6_382 b_6 NI_6 NS_382 0 -5.8905708512987411e-06
GC_6_383 b_6 NI_6 NS_383 0 -1.0067177299003648e-04
GC_6_384 b_6 NI_6 NS_384 0 1.3975659954970626e-04
GC_6_385 b_6 NI_6 NS_385 0 -8.4457507687535872e-06
GC_6_386 b_6 NI_6 NS_386 0 -1.6314926647700301e-05
GC_6_387 b_6 NI_6 NS_387 0 -1.3114897652128513e-05
GC_6_388 b_6 NI_6 NS_388 0 6.4495574226803021e-06
GC_6_389 b_6 NI_6 NS_389 0 2.2592176650883798e-05
GC_6_390 b_6 NI_6 NS_390 0 -4.4891236453262563e-05
GC_6_391 b_6 NI_6 NS_391 0 -4.7049414974223146e-05
GC_6_392 b_6 NI_6 NS_392 0 6.2087849185503806e-05
GC_6_393 b_6 NI_6 NS_393 0 -1.5074112611669547e-02
GC_6_394 b_6 NI_6 NS_394 0 -1.3247136509706382e-03
GC_6_395 b_6 NI_6 NS_395 0 -8.4916649294436398e-04
GC_6_396 b_6 NI_6 NS_396 0 -1.0111910962236606e-03
GC_6_397 b_6 NI_6 NS_397 0 -1.1790192022934978e-03
GC_6_398 b_6 NI_6 NS_398 0 1.3800284987719072e-03
GC_6_399 b_6 NI_6 NS_399 0 8.5020681007498371e-04
GC_6_400 b_6 NI_6 NS_400 0 -7.4005573565451906e-04
GC_6_401 b_6 NI_6 NS_401 0 -3.1906880525983234e-03
GC_6_402 b_6 NI_6 NS_402 0 -8.5706095281366142e-03
GC_6_403 b_6 NI_6 NS_403 0 3.1831922393774866e-05
GC_6_404 b_6 NI_6 NS_404 0 1.8335857851780563e-04
GC_6_405 b_6 NI_6 NS_405 0 1.9449516362423599e-03
GC_6_406 b_6 NI_6 NS_406 0 -2.3077120784840066e-03
GC_6_407 b_6 NI_6 NS_407 0 7.4376387219267988e-04
GC_6_408 b_6 NI_6 NS_408 0 1.7762228561358798e-04
GC_6_409 b_6 NI_6 NS_409 0 9.5984305028983636e-04
GC_6_410 b_6 NI_6 NS_410 0 -1.9577709839496819e-03
GC_6_411 b_6 NI_6 NS_411 0 1.2352236853775903e-03
GC_6_412 b_6 NI_6 NS_412 0 -2.2346515268515032e-03
GC_6_413 b_6 NI_6 NS_413 0 3.7411300779960107e-05
GC_6_414 b_6 NI_6 NS_414 0 7.0984910278763069e-06
GC_6_415 b_6 NI_6 NS_415 0 7.4412934126063118e-03
GC_6_416 b_6 NI_6 NS_416 0 1.1498965242843140e-03
GC_6_417 b_6 NI_6 NS_417 0 -1.1913406468304412e-04
GC_6_418 b_6 NI_6 NS_418 0 3.1478848249251722e-05
GC_6_419 b_6 NI_6 NS_419 0 -1.3213190232659635e-04
GC_6_420 b_6 NI_6 NS_420 0 1.2295628807027515e-04
GC_6_421 b_6 NI_6 NS_421 0 1.9358902555498668e-04
GC_6_422 b_6 NI_6 NS_422 0 -3.5776762458411088e-04
GC_6_423 b_6 NI_6 NS_423 0 3.4607944821244806e-04
GC_6_424 b_6 NI_6 NS_424 0 -1.0717382421495076e-04
GC_6_425 b_6 NI_6 NS_425 0 -7.7708114292729833e-03
GC_6_426 b_6 NI_6 NS_426 0 3.0732171071050376e-03
GC_6_427 b_6 NI_6 NS_427 0 -2.1447016470920057e-04
GC_6_428 b_6 NI_6 NS_428 0 -1.6643308406975228e-04
GC_6_429 b_6 NI_6 NS_429 0 3.8500278684386242e-03
GC_6_430 b_6 NI_6 NS_430 0 5.0804070178390233e-04
GC_6_431 b_6 NI_6 NS_431 0 2.3161102807572912e-03
GC_6_432 b_6 NI_6 NS_432 0 -1.0753088856177279e-03
GC_6_433 b_6 NI_6 NS_433 0 7.6279979155452666e-04
GC_6_434 b_6 NI_6 NS_434 0 3.3799073269589330e-04
GC_6_435 b_6 NI_6 NS_435 0 -2.6770843380316565e-06
GC_6_436 b_6 NI_6 NS_436 0 -4.3129783381924086e-06
GC_6_437 b_6 NI_6 NS_437 0 -2.0059599544932234e-05
GC_6_438 b_6 NI_6 NS_438 0 -5.6038610948406577e-06
GC_6_439 b_6 NI_6 NS_439 0 -3.3886610269537352e-05
GC_6_440 b_6 NI_6 NS_440 0 -6.9192244312858353e-05
GC_6_441 b_6 NI_6 NS_441 0 -2.7013065716494706e-05
GC_6_442 b_6 NI_6 NS_442 0 1.6625666886667365e-06
GC_6_443 b_6 NI_6 NS_443 0 -1.4439314177669654e-05
GC_6_444 b_6 NI_6 NS_444 0 -8.9562218876720209e-06
GC_6_445 b_6 NI_6 NS_445 0 2.3636326284917123e-04
GC_6_446 b_6 NI_6 NS_446 0 -1.3182694890300287e-04
GC_6_447 b_6 NI_6 NS_447 0 -3.9255774461582460e-04
GC_6_448 b_6 NI_6 NS_448 0 9.5573920238566380e-05
GC_6_449 b_6 NI_6 NS_449 0 4.1248735162764810e-03
GC_6_450 b_6 NI_6 NS_450 0 -1.5392334138855340e-04
GC_6_451 b_6 NI_6 NS_451 0 2.7446041455701309e-04
GC_6_452 b_6 NI_6 NS_452 0 4.0117508684405390e-04
GC_6_453 b_6 NI_6 NS_453 0 -4.0838844077429801e-04
GC_6_454 b_6 NI_6 NS_454 0 2.2079773903083732e-04
GC_6_455 b_6 NI_6 NS_455 0 -1.4768738065859084e-03
GC_6_456 b_6 NI_6 NS_456 0 2.6789300943580078e-04
GC_6_457 b_6 NI_6 NS_457 0 -2.0974100046736773e-04
GC_6_458 b_6 NI_6 NS_458 0 -1.5836128807355163e-03
GC_6_459 b_6 NI_6 NS_459 0 2.4930988362040788e-04
GC_6_460 b_6 NI_6 NS_460 0 -3.0220887383720728e-04
GC_6_461 b_6 NI_6 NS_461 0 7.5794081165339946e-04
GC_6_462 b_6 NI_6 NS_462 0 -1.3224230678526938e-03
GC_6_463 b_6 NI_6 NS_463 0 1.0549633435392666e-03
GC_6_464 b_6 NI_6 NS_464 0 -6.1054241004261786e-04
GC_6_465 b_6 NI_6 NS_465 0 1.8024077582086784e-03
GC_6_466 b_6 NI_6 NS_466 0 2.1958211206104770e-03
GC_6_467 b_6 NI_6 NS_467 0 2.1552121217345443e-05
GC_6_468 b_6 NI_6 NS_468 0 3.0033475850761203e-03
GC_6_469 b_6 NI_6 NS_469 0 -3.6056586731095605e-04
GC_6_470 b_6 NI_6 NS_470 0 -3.0601841440734669e-05
GC_6_471 b_6 NI_6 NS_471 0 -2.9682062250617394e-03
GC_6_472 b_6 NI_6 NS_472 0 2.6848353164432627e-03
GC_6_473 b_6 NI_6 NS_473 0 3.0309159413286770e-04
GC_6_474 b_6 NI_6 NS_474 0 1.3050530604736380e-04
GC_6_475 b_6 NI_6 NS_475 0 -1.1219286661006515e-03
GC_6_476 b_6 NI_6 NS_476 0 2.1765067958349267e-04
GC_6_477 b_6 NI_6 NS_477 0 -6.5007171853895924e-04
GC_6_478 b_6 NI_6 NS_478 0 -3.8175466618938976e-05
GC_6_479 b_6 NI_6 NS_479 0 -1.3739808880823678e-04
GC_6_480 b_6 NI_6 NS_480 0 -4.8361442042399443e-05
GC_6_481 b_6 NI_6 NS_481 0 -1.1893402914425454e-04
GC_6_482 b_6 NI_6 NS_482 0 -4.7085156800219033e-03
GC_6_483 b_6 NI_6 NS_483 0 4.2051358884184206e-05
GC_6_484 b_6 NI_6 NS_484 0 -4.1593807455531568e-05
GC_6_485 b_6 NI_6 NS_485 0 -1.2917437469166537e-03
GC_6_486 b_6 NI_6 NS_486 0 5.7009472433763983e-04
GC_6_487 b_6 NI_6 NS_487 0 1.3332622966487366e-03
GC_6_488 b_6 NI_6 NS_488 0 -9.4753626799196381e-04
GC_6_489 b_6 NI_6 NS_489 0 -2.0495660229746432e-04
GC_6_490 b_6 NI_6 NS_490 0 7.9387880350116242e-05
GC_6_491 b_6 NI_6 NS_491 0 -5.8380314157202833e-07
GC_6_492 b_6 NI_6 NS_492 0 5.5713215026827839e-07
GC_6_493 b_6 NI_6 NS_493 0 -4.5690054010163056e-06
GC_6_494 b_6 NI_6 NS_494 0 -3.8528124466534184e-06
GC_6_495 b_6 NI_6 NS_495 0 -1.3739069078403906e-05
GC_6_496 b_6 NI_6 NS_496 0 6.6748953827505198e-05
GC_6_497 b_6 NI_6 NS_497 0 -9.0077353996205181e-06
GC_6_498 b_6 NI_6 NS_498 0 -5.2421504971679114e-06
GC_6_499 b_6 NI_6 NS_499 0 -5.1694465983000774e-06
GC_6_500 b_6 NI_6 NS_500 0 -4.0149249769916971e-06
GC_6_501 b_6 NI_6 NS_501 0 2.7231027217142593e-05
GC_6_502 b_6 NI_6 NS_502 0 -2.8880396130925465e-06
GC_6_503 b_6 NI_6 NS_503 0 -4.2303480978834104e-05
GC_6_504 b_6 NI_6 NS_504 0 -7.2877499946991101e-06
GC_6_505 b_6 NI_6 NS_505 0 3.2475988588530737e-04
GC_6_506 b_6 NI_6 NS_506 0 -3.0980755351632355e-05
GC_6_507 b_6 NI_6 NS_507 0 -2.7049335834402997e-04
GC_6_508 b_6 NI_6 NS_508 0 3.0755494883873486e-07
GC_6_509 b_6 NI_6 NS_509 0 5.7804873432713563e-05
GC_6_510 b_6 NI_6 NS_510 0 -2.5250137170588171e-04
GC_6_511 b_6 NI_6 NS_511 0 7.7777544805279493e-04
GC_6_512 b_6 NI_6 NS_512 0 -7.3612716011832674e-04
GC_6_513 b_6 NI_6 NS_513 0 6.0068956357490089e-04
GC_6_514 b_6 NI_6 NS_514 0 1.5362306355449814e-03
GC_6_515 b_6 NI_6 NS_515 0 -4.4887833616709741e-04
GC_6_516 b_6 NI_6 NS_516 0 4.9316877858891263e-04
GC_6_517 b_6 NI_6 NS_517 0 -9.5111009758652655e-04
GC_6_518 b_6 NI_6 NS_518 0 -4.1093769778040296e-04
GC_6_519 b_6 NI_6 NS_519 0 4.4685531535597047e-04
GC_6_520 b_6 NI_6 NS_520 0 -5.0679412967350281e-04
GC_6_521 b_6 NI_6 NS_521 0 -1.6899424812091807e-04
GC_6_522 b_6 NI_6 NS_522 0 1.7756182987460907e-03
GC_6_523 b_6 NI_6 NS_523 0 -1.5595263523983200e-03
GC_6_524 b_6 NI_6 NS_524 0 -1.6134266411175280e-03
GC_6_525 b_6 NI_6 NS_525 0 1.9758872463832827e-04
GC_6_526 b_6 NI_6 NS_526 0 2.2939891003050673e-05
GC_6_527 b_6 NI_6 NS_527 0 3.0621028333172890e-03
GC_6_528 b_6 NI_6 NS_528 0 -2.6507979605404873e-03
GC_6_529 b_6 NI_6 NS_529 0 -4.6323500928077823e-04
GC_6_530 b_6 NI_6 NS_530 0 4.3061304152824736e-04
GC_6_531 b_6 NI_6 NS_531 0 -5.2546504666810343e-04
GC_6_532 b_6 NI_6 NS_532 0 6.0746583774064905e-04
GC_6_533 b_6 NI_6 NS_533 0 -2.1664565743844403e-04
GC_6_534 b_6 NI_6 NS_534 0 -7.3814588941002366e-04
GC_6_535 b_6 NI_6 NS_535 0 2.6808936304540358e-04
GC_6_536 b_6 NI_6 NS_536 0 -8.4522447808610859e-05
GC_6_537 b_6 NI_6 NS_537 0 1.7585085945280596e-03
GC_6_538 b_6 NI_6 NS_538 0 4.3790216031835442e-03
GC_6_539 b_6 NI_6 NS_539 0 -1.2295043446657205e-04
GC_6_540 b_6 NI_6 NS_540 0 2.5274194493526460e-04
GC_6_541 b_6 NI_6 NS_541 0 1.9986443681628066e-03
GC_6_542 b_6 NI_6 NS_542 0 -1.1613514529612795e-03
GC_6_543 b_6 NI_6 NS_543 0 -2.3427737692966501e-03
GC_6_544 b_6 NI_6 NS_544 0 -1.0191935613952268e-03
GC_6_545 b_6 NI_6 NS_545 0 -8.3276574332181888e-04
GC_6_546 b_6 NI_6 NS_546 0 7.8983909183181610e-04
GC_6_547 b_6 NI_6 NS_547 0 4.1005859113034898e-06
GC_6_548 b_6 NI_6 NS_548 0 -1.0082129638830073e-05
GC_6_549 b_6 NI_6 NS_549 0 1.1896386455800313e-05
GC_6_550 b_6 NI_6 NS_550 0 7.5866838301214451e-05
GC_6_551 b_6 NI_6 NS_551 0 1.7878025274318225e-04
GC_6_552 b_6 NI_6 NS_552 0 -2.5847034722376901e-04
GC_6_553 b_6 NI_6 NS_553 0 9.2186020446343567e-05
GC_6_554 b_6 NI_6 NS_554 0 8.6736325376870403e-05
GC_6_555 b_6 NI_6 NS_555 0 1.5660615008568634e-05
GC_6_556 b_6 NI_6 NS_556 0 5.3836253128689956e-05
GC_6_557 b_6 NI_6 NS_557 0 3.2767425826198452e-04
GC_6_558 b_6 NI_6 NS_558 0 -3.1004316323483177e-04
GC_6_559 b_6 NI_6 NS_559 0 -5.8095040744610181e-04
GC_6_560 b_6 NI_6 NS_560 0 2.9966114667718537e-04
GC_6_561 b_6 NI_6 NS_561 0 7.8306304411304081e-03
GC_6_562 b_6 NI_6 NS_562 0 -9.1683925925114531e-05
GC_6_563 b_6 NI_6 NS_563 0 -1.7746160872506806e-04
GC_6_564 b_6 NI_6 NS_564 0 7.1868147592501466e-04
GC_6_565 b_6 NI_6 NS_565 0 -3.1687559950458149e-04
GC_6_566 b_6 NI_6 NS_566 0 -6.9173339832620041e-04
GC_6_567 b_6 NI_6 NS_567 0 -5.4972304468600566e-04
GC_6_568 b_6 NI_6 NS_568 0 -7.7045896933784319e-04
GC_6_569 b_6 NI_6 NS_569 0 2.2332214597009111e-03
GC_6_570 b_6 NI_6 NS_570 0 7.1014888290253165e-04
GC_6_571 b_6 NI_6 NS_571 0 -5.9311172812271144e-04
GC_6_572 b_6 NI_6 NS_572 0 3.0662366387872674e-04
GC_6_573 b_6 NI_6 NS_573 0 5.1812684369175984e-04
GC_6_574 b_6 NI_6 NS_574 0 -6.3159516210462333e-04
GC_6_575 b_6 NI_6 NS_575 0 9.9893440500923377e-04
GC_6_576 b_6 NI_6 NS_576 0 -1.8583036461284092e-04
GC_6_577 b_6 NI_6 NS_577 0 8.3923943504146117e-04
GC_6_578 b_6 NI_6 NS_578 0 2.2099106605655301e-03
GC_6_579 b_6 NI_6 NS_579 0 -1.3060481659055707e-03
GC_6_580 b_6 NI_6 NS_580 0 2.6968060309998949e-03
GC_6_581 b_6 NI_6 NS_581 0 -2.7300723073428869e-04
GC_6_582 b_6 NI_6 NS_582 0 -6.8984088293617320e-05
GC_6_583 b_6 NI_6 NS_583 0 -5.1686945231735706e-04
GC_6_584 b_6 NI_6 NS_584 0 1.3705710614126049e-03
GC_6_585 b_6 NI_6 NS_585 0 5.5089905865154061e-05
GC_6_586 b_6 NI_6 NS_586 0 -1.2475501631719770e-06
GC_6_587 b_6 NI_6 NS_587 0 -7.3218037447717456e-04
GC_6_588 b_6 NI_6 NS_588 0 2.4700416215009044e-04
GC_6_589 b_6 NI_6 NS_589 0 -4.8231904909167863e-04
GC_6_590 b_6 NI_6 NS_590 0 6.0035738308550890e-05
GC_6_591 b_6 NI_6 NS_591 0 -1.1685653964179025e-04
GC_6_592 b_6 NI_6 NS_592 0 -4.0207276257792016e-05
GC_6_593 b_6 NI_6 NS_593 0 -4.7116972504774907e-04
GC_6_594 b_6 NI_6 NS_594 0 -2.7219927014738472e-03
GC_6_595 b_6 NI_6 NS_595 0 2.7566797171434813e-05
GC_6_596 b_6 NI_6 NS_596 0 -2.4079029042196973e-05
GC_6_597 b_6 NI_6 NS_597 0 -8.6665643406788140e-04
GC_6_598 b_6 NI_6 NS_598 0 4.0256217825814411e-04
GC_6_599 b_6 NI_6 NS_599 0 1.0381717063385474e-03
GC_6_600 b_6 NI_6 NS_600 0 2.5633695602200822e-04
GC_6_601 b_6 NI_6 NS_601 0 -1.3608131901578926e-04
GC_6_602 b_6 NI_6 NS_602 0 1.3811464717459644e-04
GC_6_603 b_6 NI_6 NS_603 0 -2.2894717286716935e-06
GC_6_604 b_6 NI_6 NS_604 0 2.5428301028417049e-06
GC_6_605 b_6 NI_6 NS_605 0 3.2788243194813181e-07
GC_6_606 b_6 NI_6 NS_606 0 -3.3797397164999160e-06
GC_6_607 b_6 NI_6 NS_607 0 -5.6560745901816103e-05
GC_6_608 b_6 NI_6 NS_608 0 3.6649605506612936e-05
GC_6_609 b_6 NI_6 NS_609 0 5.6224632493187334e-06
GC_6_610 b_6 NI_6 NS_610 0 -9.4040692107749236e-06
GC_6_611 b_6 NI_6 NS_611 0 -7.7875081786996801e-07
GC_6_612 b_6 NI_6 NS_612 0 -6.4072670726654406e-06
GC_6_613 b_6 NI_6 NS_613 0 2.7637026871309909e-05
GC_6_614 b_6 NI_6 NS_614 0 -3.7206385895770900e-05
GC_6_615 b_6 NI_6 NS_615 0 -5.0132657712728133e-05
GC_6_616 b_6 NI_6 NS_616 0 4.6877754415077757e-05
GC_6_617 b_6 NI_6 NS_617 0 -2.3410134868431338e-03
GC_6_618 b_6 NI_6 NS_618 0 -1.4592120124547753e-04
GC_6_619 b_6 NI_6 NS_619 0 -2.9574812599215413e-04
GC_6_620 b_6 NI_6 NS_620 0 -2.2219333376224284e-04
GC_6_621 b_6 NI_6 NS_621 0 3.4396351331089712e-04
GC_6_622 b_6 NI_6 NS_622 0 9.8879390522643845e-05
GC_6_623 b_6 NI_6 NS_623 0 6.5727150602835503e-04
GC_6_624 b_6 NI_6 NS_624 0 3.5060643253915884e-04
GC_6_625 b_6 NI_6 NS_625 0 -2.3804550581438687e-03
GC_6_626 b_6 NI_6 NS_626 0 8.6613055194374299e-04
GC_6_627 b_6 NI_6 NS_627 0 4.2805024028761661e-05
GC_6_628 b_6 NI_6 NS_628 0 -1.3746500195885148e-04
GC_6_629 b_6 NI_6 NS_629 0 -4.6578060797313858e-04
GC_6_630 b_6 NI_6 NS_630 0 -1.4216440208705094e-03
GC_6_631 b_6 NI_6 NS_631 0 3.5578243272977434e-04
GC_6_632 b_6 NI_6 NS_632 0 -2.4250780211550855e-04
GC_6_633 b_6 NI_6 NS_633 0 -8.1205697688913514e-04
GC_6_634 b_6 NI_6 NS_634 0 7.9176137443731100e-04
GC_6_635 b_6 NI_6 NS_635 0 -1.0272272853189095e-03
GC_6_636 b_6 NI_6 NS_636 0 -1.2913300692369233e-03
GC_6_637 b_6 NI_6 NS_637 0 1.1282428361610281e-04
GC_6_638 b_6 NI_6 NS_638 0 4.6795616690125644e-05
GC_6_639 b_6 NI_6 NS_639 0 2.1446308426480076e-03
GC_6_640 b_6 NI_6 NS_640 0 -3.3902611692299164e-03
GC_6_641 b_6 NI_6 NS_641 0 -3.1125597857620447e-04
GC_6_642 b_6 NI_6 NS_642 0 3.2872412443047880e-04
GC_6_643 b_6 NI_6 NS_643 0 -2.7674281534997326e-04
GC_6_644 b_6 NI_6 NS_644 0 2.8375751743664869e-04
GC_6_645 b_6 NI_6 NS_645 0 -4.5507978257578489e-05
GC_6_646 b_6 NI_6 NS_646 0 -5.1070189586881144e-04
GC_6_647 b_6 NI_6 NS_647 0 1.9193616919434324e-04
GC_6_648 b_6 NI_6 NS_648 0 -5.1968389223120261e-05
GC_6_649 b_6 NI_6 NS_649 0 5.0559147052699985e-04
GC_6_650 b_6 NI_6 NS_650 0 2.0558406489625770e-03
GC_6_651 b_6 NI_6 NS_651 0 -1.0539427332937972e-04
GC_6_652 b_6 NI_6 NS_652 0 1.0218758455390171e-04
GC_6_653 b_6 NI_6 NS_653 0 1.3877274826662757e-03
GC_6_654 b_6 NI_6 NS_654 0 -5.7087677839179286e-04
GC_6_655 b_6 NI_6 NS_655 0 -8.9845490945242567e-05
GC_6_656 b_6 NI_6 NS_656 0 -8.0107204918809024e-05
GC_6_657 b_6 NI_6 NS_657 0 -4.6426038117269213e-04
GC_6_658 b_6 NI_6 NS_658 0 3.8565921154690516e-04
GC_6_659 b_6 NI_6 NS_659 0 1.1023303886345413e-06
GC_6_660 b_6 NI_6 NS_660 0 -4.6245681066646056e-06
GC_6_661 b_6 NI_6 NS_661 0 -1.5055318432106766e-06
GC_6_662 b_6 NI_6 NS_662 0 3.3036193134451506e-05
GC_6_663 b_6 NI_6 NS_663 0 4.8184089445316061e-05
GC_6_664 b_6 NI_6 NS_664 0 -1.4853572942141456e-04
GC_6_665 b_6 NI_6 NS_665 0 4.1107244786259592e-05
GC_6_666 b_6 NI_6 NS_666 0 4.8683867301209557e-05
GC_6_667 b_6 NI_6 NS_667 0 3.7451952049515895e-06
GC_6_668 b_6 NI_6 NS_668 0 1.9133957983795259e-05
GC_6_669 b_6 NI_6 NS_669 0 2.3198471715609915e-04
GC_6_670 b_6 NI_6 NS_670 0 -1.1083300977560067e-04
GC_6_671 b_6 NI_6 NS_671 0 -3.7076854327114579e-04
GC_6_672 b_6 NI_6 NS_672 0 6.4778805290101104e-05
GD_6_1 b_6 NI_6 NA_1 0 2.3305025613390463e-03
GD_6_2 b_6 NI_6 NA_2 0 -2.0018996693931462e-02
GD_6_3 b_6 NI_6 NA_3 0 -1.8764971022868782e-02
GD_6_4 b_6 NI_6 NA_4 0 -1.8815260441502397e-02
GD_6_5 b_6 NI_6 NA_5 0 4.3724307229775994e-02
GD_6_6 b_6 NI_6 NA_6 0 9.3943293126935001e-02
GD_6_7 b_6 NI_6 NA_7 0 -5.3950200966531130e-02
GD_6_8 b_6 NI_6 NA_8 0 1.1454479886740563e-02
GD_6_9 b_6 NI_6 NA_9 0 5.6753650763431353e-05
GD_6_10 b_6 NI_6 NA_10 0 -3.1486186037215699e-03
GD_6_11 b_6 NI_6 NA_11 0 -1.2049855159344423e-02
GD_6_12 b_6 NI_6 NA_12 0 5.0915336871031943e-03
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 8.7304398110413670e-02
GC_7_2 b_7 NI_7 NS_2 0 -6.0122120129970941e-04
GC_7_3 b_7 NI_7 NS_3 0 4.0530896420450596e-03
GC_7_4 b_7 NI_7 NS_4 0 -1.5490071474414846e-03
GC_7_5 b_7 NI_7 NS_5 0 7.8453436218839739e-05
GC_7_6 b_7 NI_7 NS_6 0 5.5038400272796380e-03
GC_7_7 b_7 NI_7 NS_7 0 -1.2061496917185495e-03
GC_7_8 b_7 NI_7 NS_8 0 1.1589545008593634e-02
GC_7_9 b_7 NI_7 NS_9 0 -1.5625989539396291e-02
GC_7_10 b_7 NI_7 NS_10 0 5.5669629573582551e-03
GC_7_11 b_7 NI_7 NS_11 0 1.0316180314501646e-04
GC_7_12 b_7 NI_7 NS_12 0 6.3074953738341571e-05
GC_7_13 b_7 NI_7 NS_13 0 2.9428163021877115e-03
GC_7_14 b_7 NI_7 NS_14 0 6.1115288388197630e-04
GC_7_15 b_7 NI_7 NS_15 0 2.5123131252852084e-04
GC_7_16 b_7 NI_7 NS_16 0 2.0083417416855505e-03
GC_7_17 b_7 NI_7 NS_17 0 -6.7042076153026302e-03
GC_7_18 b_7 NI_7 NS_18 0 6.5997323108334238e-03
GC_7_19 b_7 NI_7 NS_19 0 -1.7608760307172573e-04
GC_7_20 b_7 NI_7 NS_20 0 6.1387843672513868e-03
GC_7_21 b_7 NI_7 NS_21 0 3.5322564792489416e-04
GC_7_22 b_7 NI_7 NS_22 0 8.5689308268441439e-05
GC_7_23 b_7 NI_7 NS_23 0 -1.9433940848689175e-02
GC_7_24 b_7 NI_7 NS_24 0 9.2620152802493614e-04
GC_7_25 b_7 NI_7 NS_25 0 1.2635821915308511e-03
GC_7_26 b_7 NI_7 NS_26 0 5.8042423561609181e-04
GC_7_27 b_7 NI_7 NS_27 0 -5.2180237914950381e-04
GC_7_28 b_7 NI_7 NS_28 0 -2.3816938882796813e-04
GC_7_29 b_7 NI_7 NS_29 0 -4.6673986766791080e-04
GC_7_30 b_7 NI_7 NS_30 0 2.2032709024447352e-04
GC_7_31 b_7 NI_7 NS_31 0 -1.9651045295060175e-04
GC_7_32 b_7 NI_7 NS_32 0 -7.9602561659266277e-06
GC_7_33 b_7 NI_7 NS_33 0 -7.8911477550939954e-03
GC_7_34 b_7 NI_7 NS_34 0 -1.4291063158345248e-02
GC_7_35 b_7 NI_7 NS_35 0 2.0902396211503149e-04
GC_7_36 b_7 NI_7 NS_36 0 -3.7711964779295488e-05
GC_7_37 b_7 NI_7 NS_37 0 -2.1997658538199590e-03
GC_7_38 b_7 NI_7 NS_38 0 2.7833234031218353e-03
GC_7_39 b_7 NI_7 NS_39 0 8.0639162651206363e-03
GC_7_40 b_7 NI_7 NS_40 0 -2.7509416758489764e-03
GC_7_41 b_7 NI_7 NS_41 0 -2.3262065734184006e-04
GC_7_42 b_7 NI_7 NS_42 0 4.2506571793002313e-04
GC_7_43 b_7 NI_7 NS_43 0 1.2389195699588522e-06
GC_7_44 b_7 NI_7 NS_44 0 5.6803064886268140e-06
GC_7_45 b_7 NI_7 NS_45 0 2.0723810303613784e-06
GC_7_46 b_7 NI_7 NS_46 0 -2.5087260721120609e-05
GC_7_47 b_7 NI_7 NS_47 0 -5.1687721697926605e-04
GC_7_48 b_7 NI_7 NS_48 0 1.0480751537451303e-04
GC_7_49 b_7 NI_7 NS_49 0 2.2190710886336585e-05
GC_7_50 b_7 NI_7 NS_50 0 -4.9175704823575178e-05
GC_7_51 b_7 NI_7 NS_51 0 -3.0195695432547267e-05
GC_7_52 b_7 NI_7 NS_52 0 -1.3421877435324565e-05
GC_7_53 b_7 NI_7 NS_53 0 1.1106904931526395e-04
GC_7_54 b_7 NI_7 NS_54 0 -5.2454594377881233e-05
GC_7_55 b_7 NI_7 NS_55 0 -1.8572327369162088e-04
GC_7_56 b_7 NI_7 NS_56 0 2.4900950676778824e-05
GC_7_57 b_7 NI_7 NS_57 0 -3.7744081428270092e-02
GC_7_58 b_7 NI_7 NS_58 0 -9.0932264974805284e-05
GC_7_59 b_7 NI_7 NS_59 0 -3.0858689607549323e-04
GC_7_60 b_7 NI_7 NS_60 0 2.4212140736379613e-03
GC_7_61 b_7 NI_7 NS_61 0 -2.5417475313663320e-03
GC_7_62 b_7 NI_7 NS_62 0 -1.4090481662047591e-03
GC_7_63 b_7 NI_7 NS_63 0 -5.7681344956309792e-03
GC_7_64 b_7 NI_7 NS_64 0 -6.2456448782983835e-03
GC_7_65 b_7 NI_7 NS_65 0 8.1080997461518475e-03
GC_7_66 b_7 NI_7 NS_66 0 -9.8242341333005991e-03
GC_7_67 b_7 NI_7 NS_67 0 3.5721824755533574e-04
GC_7_68 b_7 NI_7 NS_68 0 4.3932322268337508e-04
GC_7_69 b_7 NI_7 NS_69 0 5.3359142992845596e-03
GC_7_70 b_7 NI_7 NS_70 0 -2.2773339839630190e-03
GC_7_71 b_7 NI_7 NS_71 0 5.2666382728496538e-04
GC_7_72 b_7 NI_7 NS_72 0 5.6600073516327443e-04
GC_7_73 b_7 NI_7 NS_73 0 1.0159074818504297e-03
GC_7_74 b_7 NI_7 NS_74 0 2.3597400573463676e-03
GC_7_75 b_7 NI_7 NS_75 0 -1.6045620963018079e-04
GC_7_76 b_7 NI_7 NS_76 0 6.9411562634617420e-05
GC_7_77 b_7 NI_7 NS_77 0 -1.7845474784796174e-04
GC_7_78 b_7 NI_7 NS_78 0 7.8033621587364523e-05
GC_7_79 b_7 NI_7 NS_79 0 1.0261232391483371e-03
GC_7_80 b_7 NI_7 NS_80 0 -3.4202526036688280e-03
GC_7_81 b_7 NI_7 NS_81 0 -8.9230910426287523e-04
GC_7_82 b_7 NI_7 NS_82 0 1.7320729742644272e-04
GC_7_83 b_7 NI_7 NS_83 0 -3.2388660654319983e-05
GC_7_84 b_7 NI_7 NS_84 0 3.6437987106879414e-05
GC_7_85 b_7 NI_7 NS_85 0 -2.3531942786668880e-04
GC_7_86 b_7 NI_7 NS_86 0 -2.8014087548466039e-05
GC_7_87 b_7 NI_7 NS_87 0 -9.9213685850908889e-05
GC_7_88 b_7 NI_7 NS_88 0 -1.3351814042990515e-04
GC_7_89 b_7 NI_7 NS_89 0 8.0871988385318640e-03
GC_7_90 b_7 NI_7 NS_90 0 -3.6638662887031450e-05
GC_7_91 b_7 NI_7 NS_91 0 -5.7313388012101221e-05
GC_7_92 b_7 NI_7 NS_92 0 1.2753681639939484e-04
GC_7_93 b_7 NI_7 NS_93 0 -4.6378670170234856e-04
GC_7_94 b_7 NI_7 NS_94 0 -1.4512536239903531e-03
GC_7_95 b_7 NI_7 NS_95 0 -2.0239529926139888e-04
GC_7_96 b_7 NI_7 NS_96 0 2.0288549986224374e-03
GC_7_97 b_7 NI_7 NS_97 0 -3.9067901948646632e-04
GC_7_98 b_7 NI_7 NS_98 0 -6.7787755302215283e-05
GC_7_99 b_7 NI_7 NS_99 0 -2.1470203941051075e-06
GC_7_100 b_7 NI_7 NS_100 0 -2.3909737711461923e-06
GC_7_101 b_7 NI_7 NS_101 0 5.7483737560034770e-06
GC_7_102 b_7 NI_7 NS_102 0 1.4820634674224101e-05
GC_7_103 b_7 NI_7 NS_103 0 1.7966600367736200e-04
GC_7_104 b_7 NI_7 NS_104 0 -1.6573033964355750e-04
GC_7_105 b_7 NI_7 NS_105 0 -8.1028247260549806e-07
GC_7_106 b_7 NI_7 NS_106 0 2.7997753219445724e-05
GC_7_107 b_7 NI_7 NS_107 0 5.2009873171056939e-06
GC_7_108 b_7 NI_7 NS_108 0 4.7376995607246434e-07
GC_7_109 b_7 NI_7 NS_109 0 -1.9362264172321905e-05
GC_7_110 b_7 NI_7 NS_110 0 1.8911107066334327e-05
GC_7_111 b_7 NI_7 NS_111 0 4.0892770381326488e-05
GC_7_112 b_7 NI_7 NS_112 0 -1.0329265962825315e-05
GC_7_113 b_7 NI_7 NS_113 0 3.8795067795017950e-02
GC_7_114 b_7 NI_7 NS_114 0 1.9750542861029304e-04
GC_7_115 b_7 NI_7 NS_115 0 5.2441381790850243e-03
GC_7_116 b_7 NI_7 NS_116 0 -5.0639849259712143e-05
GC_7_117 b_7 NI_7 NS_117 0 -3.8439901486907874e-03
GC_7_118 b_7 NI_7 NS_118 0 2.9963247926830111e-03
GC_7_119 b_7 NI_7 NS_119 0 -1.1812884697322771e-03
GC_7_120 b_7 NI_7 NS_120 0 7.1585111778305040e-03
GC_7_121 b_7 NI_7 NS_121 0 -8.4626749362283309e-03
GC_7_122 b_7 NI_7 NS_122 0 -5.6478453618065546e-03
GC_7_123 b_7 NI_7 NS_123 0 -1.6913173611970002e-04
GC_7_124 b_7 NI_7 NS_124 0 -1.8144928396625668e-04
GC_7_125 b_7 NI_7 NS_125 0 8.2792212334501167e-03
GC_7_126 b_7 NI_7 NS_126 0 5.1720878020842923e-04
GC_7_127 b_7 NI_7 NS_127 0 2.7691025390390333e-04
GC_7_128 b_7 NI_7 NS_128 0 2.3814244004107085e-03
GC_7_129 b_7 NI_7 NS_129 0 -7.2951634884521664e-04
GC_7_130 b_7 NI_7 NS_130 0 3.1567003907469401e-03
GC_7_131 b_7 NI_7 NS_131 0 6.1194599778299839e-04
GC_7_132 b_7 NI_7 NS_132 0 5.3578776252239087e-03
GC_7_133 b_7 NI_7 NS_133 0 3.3841060791703646e-04
GC_7_134 b_7 NI_7 NS_134 0 1.7577813560604177e-04
GC_7_135 b_7 NI_7 NS_135 0 -1.0819859358058943e-02
GC_7_136 b_7 NI_7 NS_136 0 5.3913820168409107e-03
GC_7_137 b_7 NI_7 NS_137 0 9.9973975282443292e-04
GC_7_138 b_7 NI_7 NS_138 0 4.5517616987618631e-04
GC_7_139 b_7 NI_7 NS_139 0 -5.4244451223313449e-04
GC_7_140 b_7 NI_7 NS_140 0 1.8787830252739710e-06
GC_7_141 b_7 NI_7 NS_141 0 -2.7958400500440031e-04
GC_7_142 b_7 NI_7 NS_142 0 2.1243215299802159e-04
GC_7_143 b_7 NI_7 NS_143 0 -1.3207582852797835e-04
GC_7_144 b_7 NI_7 NS_144 0 1.2753242153247739e-05
GC_7_145 b_7 NI_7 NS_145 0 -8.0524317465783379e-03
GC_7_146 b_7 NI_7 NS_146 0 -1.1297655016081086e-02
GC_7_147 b_7 NI_7 NS_147 0 1.4347883842292291e-04
GC_7_148 b_7 NI_7 NS_148 0 -4.5514726057819185e-05
GC_7_149 b_7 NI_7 NS_149 0 -1.1618775368556940e-03
GC_7_150 b_7 NI_7 NS_150 0 2.3711141662536837e-03
GC_7_151 b_7 NI_7 NS_151 0 6.1320464700320102e-03
GC_7_152 b_7 NI_7 NS_152 0 -2.1279855865388687e-04
GC_7_153 b_7 NI_7 NS_153 0 1.3792545076917709e-04
GC_7_154 b_7 NI_7 NS_154 0 3.3187763860138472e-04
GC_7_155 b_7 NI_7 NS_155 0 -2.2625934400794294e-08
GC_7_156 b_7 NI_7 NS_156 0 4.3694038747229684e-06
GC_7_157 b_7 NI_7 NS_157 0 4.1984813915157843e-06
GC_7_158 b_7 NI_7 NS_158 0 -1.9601858204855516e-05
GC_7_159 b_7 NI_7 NS_159 0 -3.6146939135671337e-04
GC_7_160 b_7 NI_7 NS_160 0 7.4582472430135633e-05
GC_7_161 b_7 NI_7 NS_161 0 1.8606664139732309e-05
GC_7_162 b_7 NI_7 NS_162 0 -3.6500753531045666e-05
GC_7_163 b_7 NI_7 NS_163 0 -2.0254702025645061e-05
GC_7_164 b_7 NI_7 NS_164 0 -1.2254882260334200e-05
GC_7_165 b_7 NI_7 NS_165 0 8.2425155540443262e-05
GC_7_166 b_7 NI_7 NS_166 0 -3.4698500511977674e-05
GC_7_167 b_7 NI_7 NS_167 0 -1.3711722737260002e-04
GC_7_168 b_7 NI_7 NS_168 0 1.1500336898521128e-05
GC_7_169 b_7 NI_7 NS_169 0 -8.2280834145318574e-03
GC_7_170 b_7 NI_7 NS_170 0 -2.3837370115176060e-04
GC_7_171 b_7 NI_7 NS_171 0 -1.3510034806754323e-03
GC_7_172 b_7 NI_7 NS_172 0 2.9662468753484808e-03
GC_7_173 b_7 NI_7 NS_173 0 -9.2138232963066477e-04
GC_7_174 b_7 NI_7 NS_174 0 -2.2289397577289912e-03
GC_7_175 b_7 NI_7 NS_175 0 -4.8028512757118469e-03
GC_7_176 b_7 NI_7 NS_176 0 -5.4465581545335611e-03
GC_7_177 b_7 NI_7 NS_177 0 6.6780373885692275e-03
GC_7_178 b_7 NI_7 NS_178 0 -1.5237086673296517e-03
GC_7_179 b_7 NI_7 NS_179 0 1.6747671394221251e-04
GC_7_180 b_7 NI_7 NS_180 0 -3.0856848391990196e-05
GC_7_181 b_7 NI_7 NS_181 0 4.0263033397161434e-03
GC_7_182 b_7 NI_7 NS_182 0 -2.6519574755876443e-03
GC_7_183 b_7 NI_7 NS_183 0 6.9140887688269256e-04
GC_7_184 b_7 NI_7 NS_184 0 1.0151562673966067e-03
GC_7_185 b_7 NI_7 NS_185 0 7.1352989709970189e-04
GC_7_186 b_7 NI_7 NS_186 0 2.1040188619635062e-03
GC_7_187 b_7 NI_7 NS_187 0 -3.0951634400913368e-03
GC_7_188 b_7 NI_7 NS_188 0 8.4633238507332315e-04
GC_7_189 b_7 NI_7 NS_189 0 -1.9656287550761257e-04
GC_7_190 b_7 NI_7 NS_190 0 -3.6504364566705176e-06
GC_7_191 b_7 NI_7 NS_191 0 2.5992903858731036e-03
GC_7_192 b_7 NI_7 NS_192 0 5.4805897879403621e-05
GC_7_193 b_7 NI_7 NS_193 0 -7.9285856059706737e-04
GC_7_194 b_7 NI_7 NS_194 0 -1.2485858719601963e-04
GC_7_195 b_7 NI_7 NS_195 0 -2.1064989308799796e-04
GC_7_196 b_7 NI_7 NS_196 0 5.0355621137776984e-05
GC_7_197 b_7 NI_7 NS_197 0 -2.6612980420956107e-04
GC_7_198 b_7 NI_7 NS_198 0 1.3769874454978680e-04
GC_7_199 b_7 NI_7 NS_199 0 -1.2376747751928843e-04
GC_7_200 b_7 NI_7 NS_200 0 -8.5167744465343816e-05
GC_7_201 b_7 NI_7 NS_201 0 7.8164186085514121e-04
GC_7_202 b_7 NI_7 NS_202 0 -7.9134408292485582e-04
GC_7_203 b_7 NI_7 NS_203 0 -3.9438199385837136e-05
GC_7_204 b_7 NI_7 NS_204 0 6.8819462196090394e-05
GC_7_205 b_7 NI_7 NS_205 0 -1.9211240642398106e-04
GC_7_206 b_7 NI_7 NS_206 0 -4.7540070049875580e-04
GC_7_207 b_7 NI_7 NS_207 0 4.9724636543148663e-04
GC_7_208 b_7 NI_7 NS_208 0 1.2130326488450970e-03
GC_7_209 b_7 NI_7 NS_209 0 8.9668980481192065e-06
GC_7_210 b_7 NI_7 NS_210 0 2.0842974946515924e-07
GC_7_211 b_7 NI_7 NS_211 0 -1.6851757960187553e-06
GC_7_212 b_7 NI_7 NS_212 0 -3.7129175061898191e-07
GC_7_213 b_7 NI_7 NS_213 0 4.4123157210272904e-06
GC_7_214 b_7 NI_7 NS_214 0 4.5135015225271191e-06
GC_7_215 b_7 NI_7 NS_215 0 1.6767756936053080e-05
GC_7_216 b_7 NI_7 NS_216 0 -8.8235344594474467e-05
GC_7_217 b_7 NI_7 NS_217 0 3.9265157875156934e-06
GC_7_218 b_7 NI_7 NS_218 0 8.3148982085170756e-06
GC_7_219 b_7 NI_7 NS_219 0 -4.7725574127819770e-08
GC_7_220 b_7 NI_7 NS_220 0 -2.8866313194389458e-06
GC_7_221 b_7 NI_7 NS_221 0 1.1959584208648860e-05
GC_7_222 b_7 NI_7 NS_222 0 1.1578073844319966e-05
GC_7_223 b_7 NI_7 NS_223 0 -8.7168575127440477e-06
GC_7_224 b_7 NI_7 NS_224 0 -1.6252124349234261e-05
GC_7_225 b_7 NI_7 NS_225 0 -2.1720294406733967e-02
GC_7_226 b_7 NI_7 NS_226 0 1.6798521860743418e-03
GC_7_227 b_7 NI_7 NS_227 0 3.6043974572228586e-03
GC_7_228 b_7 NI_7 NS_228 0 2.4430212331954981e-03
GC_7_229 b_7 NI_7 NS_229 0 -5.3181847674780751e-03
GC_7_230 b_7 NI_7 NS_230 0 -6.5605009252241494e-03
GC_7_231 b_7 NI_7 NS_231 0 4.1121300400224587e-03
GC_7_232 b_7 NI_7 NS_232 0 2.0573913982210668e-03
GC_7_233 b_7 NI_7 NS_233 0 1.0332343411193564e-02
GC_7_234 b_7 NI_7 NS_234 0 -1.0197213546177038e-02
GC_7_235 b_7 NI_7 NS_235 0 -3.5358494178708532e-04
GC_7_236 b_7 NI_7 NS_236 0 1.5625094353297135e-04
GC_7_237 b_7 NI_7 NS_237 0 8.6981608579305095e-03
GC_7_238 b_7 NI_7 NS_238 0 3.0601460457475348e-03
GC_7_239 b_7 NI_7 NS_239 0 7.1707804375454665e-04
GC_7_240 b_7 NI_7 NS_240 0 2.0876809031374478e-03
GC_7_241 b_7 NI_7 NS_241 0 6.9603586024997851e-03
GC_7_242 b_7 NI_7 NS_242 0 1.0490131780613104e-03
GC_7_243 b_7 NI_7 NS_243 0 2.6266710926345273e-03
GC_7_244 b_7 NI_7 NS_244 0 3.9523114505835982e-03
GC_7_245 b_7 NI_7 NS_245 0 3.5523277622726609e-04
GC_7_246 b_7 NI_7 NS_246 0 1.3295437534011230e-04
GC_7_247 b_7 NI_7 NS_247 0 -4.1321520522764020e-03
GC_7_248 b_7 NI_7 NS_248 0 1.2930625152287758e-02
GC_7_249 b_7 NI_7 NS_249 0 9.9518265438494949e-04
GC_7_250 b_7 NI_7 NS_250 0 8.3432592184031653e-05
GC_7_251 b_7 NI_7 NS_251 0 -5.2970110635698836e-04
GC_7_252 b_7 NI_7 NS_252 0 7.2766756532889192e-05
GC_7_253 b_7 NI_7 NS_253 0 -1.6781578797079008e-04
GC_7_254 b_7 NI_7 NS_254 0 1.5339793186673598e-04
GC_7_255 b_7 NI_7 NS_255 0 -6.3877336420185016e-05
GC_7_256 b_7 NI_7 NS_256 0 2.5805606966230360e-05
GC_7_257 b_7 NI_7 NS_257 0 -4.3870371139475405e-03
GC_7_258 b_7 NI_7 NS_258 0 -3.1395911155164421e-03
GC_7_259 b_7 NI_7 NS_259 0 7.7194609924733813e-05
GC_7_260 b_7 NI_7 NS_260 0 -4.6487787916813931e-05
GC_7_261 b_7 NI_7 NS_261 0 -9.9880808214146906e-05
GC_7_262 b_7 NI_7 NS_262 0 1.6396446303196519e-03
GC_7_263 b_7 NI_7 NS_263 0 -2.4070897667517765e-04
GC_7_264 b_7 NI_7 NS_264 0 -5.4000804431366604e-04
GC_7_265 b_7 NI_7 NS_265 0 2.0123268353895678e-05
GC_7_266 b_7 NI_7 NS_266 0 2.4720901330132697e-04
GC_7_267 b_7 NI_7 NS_267 0 -5.7246384480366195e-07
GC_7_268 b_7 NI_7 NS_268 0 9.1028936055968278e-08
GC_7_269 b_7 NI_7 NS_269 0 -3.2764029085354502e-07
GC_7_270 b_7 NI_7 NS_270 0 1.1927936044754459e-06
GC_7_271 b_7 NI_7 NS_271 0 3.9302493573440187e-05
GC_7_272 b_7 NI_7 NS_272 0 6.1838636505258453e-05
GC_7_273 b_7 NI_7 NS_273 0 -2.8571316684267265e-06
GC_7_274 b_7 NI_7 NS_274 0 9.9821837589841744e-07
GC_7_275 b_7 NI_7 NS_275 0 -2.8073786932446491e-06
GC_7_276 b_7 NI_7 NS_276 0 -5.0432166161818940e-06
GC_7_277 b_7 NI_7 NS_277 0 1.4787343033813460e-05
GC_7_278 b_7 NI_7 NS_278 0 -9.2576157850699802e-06
GC_7_279 b_7 NI_7 NS_279 0 -2.9553523855349937e-05
GC_7_280 b_7 NI_7 NS_280 0 7.2103030241356102e-06
GC_7_281 b_7 NI_7 NS_281 0 5.7573995023942177e-02
GC_7_282 b_7 NI_7 NS_282 0 -7.8908432183426595e-04
GC_7_283 b_7 NI_7 NS_283 0 -1.7550542069091760e-03
GC_7_284 b_7 NI_7 NS_284 0 2.3937903761522875e-03
GC_7_285 b_7 NI_7 NS_285 0 2.8923399177405739e-03
GC_7_286 b_7 NI_7 NS_286 0 2.8225286742789848e-04
GC_7_287 b_7 NI_7 NS_287 0 -5.6229684162306393e-03
GC_7_288 b_7 NI_7 NS_288 0 5.6045715252253496e-04
GC_7_289 b_7 NI_7 NS_289 0 -6.4091422020186367e-03
GC_7_290 b_7 NI_7 NS_290 0 1.0277525061075699e-02
GC_7_291 b_7 NI_7 NS_291 0 -5.3710528180944109e-04
GC_7_292 b_7 NI_7 NS_292 0 -2.6664432400433233e-04
GC_7_293 b_7 NI_7 NS_293 0 1.8473492048455659e-03
GC_7_294 b_7 NI_7 NS_294 0 -4.4300295537775466e-03
GC_7_295 b_7 NI_7 NS_295 0 1.0620724899400834e-03
GC_7_296 b_7 NI_7 NS_296 0 1.3769930609841129e-03
GC_7_297 b_7 NI_7 NS_297 0 -1.0672661251000725e-04
GC_7_298 b_7 NI_7 NS_298 0 1.2707692528946587e-03
GC_7_299 b_7 NI_7 NS_299 0 -5.9327847793137429e-03
GC_7_300 b_7 NI_7 NS_300 0 9.8778558334483351e-04
GC_7_301 b_7 NI_7 NS_301 0 -1.4813178555224025e-04
GC_7_302 b_7 NI_7 NS_302 0 -8.4416546535512322e-05
GC_7_303 b_7 NI_7 NS_303 0 1.0332063175590501e-03
GC_7_304 b_7 NI_7 NS_304 0 5.3252605127487021e-03
GC_7_305 b_7 NI_7 NS_305 0 -4.7987269228077215e-04
GC_7_306 b_7 NI_7 NS_306 0 -1.7923478726825621e-04
GC_7_307 b_7 NI_7 NS_307 0 -5.0274838507819157e-04
GC_7_308 b_7 NI_7 NS_308 0 7.2378405313898401e-05
GC_7_309 b_7 NI_7 NS_309 0 -4.4711456784811730e-04
GC_7_310 b_7 NI_7 NS_310 0 4.6474053763776645e-04
GC_7_311 b_7 NI_7 NS_311 0 -2.5256704698743785e-04
GC_7_312 b_7 NI_7 NS_312 0 -3.9026797580952016e-05
GC_7_313 b_7 NI_7 NS_313 0 -8.1484255062484849e-03
GC_7_314 b_7 NI_7 NS_314 0 -1.9148405400521806e-03
GC_7_315 b_7 NI_7 NS_315 0 -1.5473165649112963e-05
GC_7_316 b_7 NI_7 NS_316 0 3.6747395338811911e-05
GC_7_317 b_7 NI_7 NS_317 0 -8.7894504030742025e-05
GC_7_318 b_7 NI_7 NS_318 0 7.6916528992173228e-04
GC_7_319 b_7 NI_7 NS_319 0 9.0364342356141677e-05
GC_7_320 b_7 NI_7 NS_320 0 -2.9101782588543314e-03
GC_7_321 b_7 NI_7 NS_321 0 3.3469560357612553e-04
GC_7_322 b_7 NI_7 NS_322 0 2.3824812517159061e-04
GC_7_323 b_7 NI_7 NS_323 0 -4.7633284126767397e-07
GC_7_324 b_7 NI_7 NS_324 0 1.1738497303107371e-06
GC_7_325 b_7 NI_7 NS_325 0 -3.5728064172987708e-06
GC_7_326 b_7 NI_7 NS_326 0 -5.8905708512529666e-06
GC_7_327 b_7 NI_7 NS_327 0 -1.0067177299038797e-04
GC_7_328 b_7 NI_7 NS_328 0 1.3975659954929394e-04
GC_7_329 b_7 NI_7 NS_329 0 -8.4457507686533307e-06
GC_7_330 b_7 NI_7 NS_330 0 -1.6314926647700877e-05
GC_7_331 b_7 NI_7 NS_331 0 -1.3114897652135895e-05
GC_7_332 b_7 NI_7 NS_332 0 6.4495574226490991e-06
GC_7_333 b_7 NI_7 NS_333 0 2.2592176651009304e-05
GC_7_334 b_7 NI_7 NS_334 0 -4.4891236453239490e-05
GC_7_335 b_7 NI_7 NS_335 0 -4.7049414974394910e-05
GC_7_336 b_7 NI_7 NS_336 0 6.2087849185408329e-05
GC_7_337 b_7 NI_7 NS_337 0 -6.1752887316885940e-02
GC_7_338 b_7 NI_7 NS_338 0 1.5398314481293992e-02
GC_7_339 b_7 NI_7 NS_339 0 4.0794377955196076e-03
GC_7_340 b_7 NI_7 NS_340 0 2.2311526676195357e-03
GC_7_341 b_7 NI_7 NS_341 0 1.2091801295770163e-02
GC_7_342 b_7 NI_7 NS_342 0 -1.7196203301661871e-04
GC_7_343 b_7 NI_7 NS_343 0 -1.6782750564553827e-05
GC_7_344 b_7 NI_7 NS_344 0 1.7468346860453129e-03
GC_7_345 b_7 NI_7 NS_345 0 1.0065207572285613e-02
GC_7_346 b_7 NI_7 NS_346 0 7.3687457331607946e-03
GC_7_347 b_7 NI_7 NS_347 0 7.8777605130315152e-04
GC_7_348 b_7 NI_7 NS_348 0 9.3595939680525759e-04
GC_7_349 b_7 NI_7 NS_349 0 6.2907520265543726e-03
GC_7_350 b_7 NI_7 NS_350 0 -1.6717997343726752e-03
GC_7_351 b_7 NI_7 NS_351 0 4.9605856960055852e-04
GC_7_352 b_7 NI_7 NS_352 0 1.6144853279210895e-03
GC_7_353 b_7 NI_7 NS_353 0 7.1433858213407310e-03
GC_7_354 b_7 NI_7 NS_354 0 -4.4376869358747260e-04
GC_7_355 b_7 NI_7 NS_355 0 3.7540745338271219e-03
GC_7_356 b_7 NI_7 NS_356 0 3.4883092898264586e-03
GC_7_357 b_7 NI_7 NS_357 0 2.3809645203201070e-04
GC_7_358 b_7 NI_7 NS_358 0 1.7052332770383212e-04
GC_7_359 b_7 NI_7 NS_359 0 3.6246271583005173e-03
GC_7_360 b_7 NI_7 NS_360 0 4.9259439606099695e-03
GC_7_361 b_7 NI_7 NS_361 0 3.2034007782027725e-04
GC_7_362 b_7 NI_7 NS_362 0 8.6325662171038688e-05
GC_7_363 b_7 NI_7 NS_363 0 -2.7097214054292622e-04
GC_7_364 b_7 NI_7 NS_364 0 1.3177145378624676e-04
GC_7_365 b_7 NI_7 NS_365 0 4.6209451715555922e-05
GC_7_366 b_7 NI_7 NS_366 0 -9.5191797977918800e-05
GC_7_367 b_7 NI_7 NS_367 0 2.9383875036579589e-05
GC_7_368 b_7 NI_7 NS_368 0 -4.6271911233844458e-06
GC_7_369 b_7 NI_7 NS_369 0 3.8484347604193873e-04
GC_7_370 b_7 NI_7 NS_370 0 6.1407271774723280e-03
GC_7_371 b_7 NI_7 NS_371 0 -2.7488556055175529e-05
GC_7_372 b_7 NI_7 NS_372 0 -1.0967158125727395e-05
GC_7_373 b_7 NI_7 NS_373 0 8.8257550668104730e-04
GC_7_374 b_7 NI_7 NS_374 0 1.8206378541206196e-04
GC_7_375 b_7 NI_7 NS_375 0 -1.9210381674425790e-03
GC_7_376 b_7 NI_7 NS_376 0 2.0539697222589828e-03
GC_7_377 b_7 NI_7 NS_377 0 2.3693991432986638e-04
GC_7_378 b_7 NI_7 NS_378 0 -3.3235096270397435e-04
GC_7_379 b_7 NI_7 NS_379 0 -5.4037696935484395e-08
GC_7_380 b_7 NI_7 NS_380 0 -1.2770268807552219e-06
GC_7_381 b_7 NI_7 NS_381 0 4.7147854534190380e-06
GC_7_382 b_7 NI_7 NS_382 0 1.4450271788978095e-05
GC_7_383 b_7 NI_7 NS_383 0 2.4165860384830291e-04
GC_7_384 b_7 NI_7 NS_384 0 -9.4762146277973633e-05
GC_7_385 b_7 NI_7 NS_385 0 -1.3235134592024867e-06
GC_7_386 b_7 NI_7 NS_386 0 2.7791046861496300e-05
GC_7_387 b_7 NI_7 NS_387 0 6.7997207648331516e-06
GC_7_388 b_7 NI_7 NS_388 0 2.0215011245197359e-06
GC_7_389 b_7 NI_7 NS_389 0 -2.5764229378091695e-05
GC_7_390 b_7 NI_7 NS_390 0 1.1164290363121390e-05
GC_7_391 b_7 NI_7 NS_391 0 4.2259168241590537e-05
GC_7_392 b_7 NI_7 NS_392 0 -1.5704088767566514e-06
GC_7_393 b_7 NI_7 NS_393 0 -1.3219958273246015e-02
GC_7_394 b_7 NI_7 NS_394 0 1.2044449083902765e-02
GC_7_395 b_7 NI_7 NS_395 0 -2.2023344575709397e-03
GC_7_396 b_7 NI_7 NS_396 0 1.4394743987853136e-03
GC_7_397 b_7 NI_7 NS_397 0 -2.4020460292128142e-03
GC_7_398 b_7 NI_7 NS_398 0 4.3204556206904816e-03
GC_7_399 b_7 NI_7 NS_399 0 -9.8944804927672656e-04
GC_7_400 b_7 NI_7 NS_400 0 -2.9570758796023701e-03
GC_7_401 b_7 NI_7 NS_401 0 -1.1571807928308451e-02
GC_7_402 b_7 NI_7 NS_402 0 -3.3375374356219793e-03
GC_7_403 b_7 NI_7 NS_403 0 3.3294280737468780e-04
GC_7_404 b_7 NI_7 NS_404 0 -3.8181711718840005e-04
GC_7_405 b_7 NI_7 NS_405 0 3.0706477843229023e-03
GC_7_406 b_7 NI_7 NS_406 0 2.7298466753090158e-04
GC_7_407 b_7 NI_7 NS_407 0 9.7712036860211579e-04
GC_7_408 b_7 NI_7 NS_408 0 6.3661363947187905e-04
GC_7_409 b_7 NI_7 NS_409 0 4.2160893262319522e-03
GC_7_410 b_7 NI_7 NS_410 0 -6.9945736704659799e-04
GC_7_411 b_7 NI_7 NS_411 0 -1.0010219503949281e-03
GC_7_412 b_7 NI_7 NS_412 0 5.8035147746363384e-04
GC_7_413 b_7 NI_7 NS_413 0 -1.4614069636603540e-04
GC_7_414 b_7 NI_7 NS_414 0 -4.2750998104374631e-05
GC_7_415 b_7 NI_7 NS_415 0 4.1349476973865842e-03
GC_7_416 b_7 NI_7 NS_416 0 -3.9764447797501276e-04
GC_7_417 b_7 NI_7 NS_417 0 -4.7548246833205169e-04
GC_7_418 b_7 NI_7 NS_418 0 -1.4229995897005934e-04
GC_7_419 b_7 NI_7 NS_419 0 -2.8838813921668759e-04
GC_7_420 b_7 NI_7 NS_420 0 3.6416699210840484e-05
GC_7_421 b_7 NI_7 NS_421 0 -3.0280954547604928e-04
GC_7_422 b_7 NI_7 NS_422 0 1.4279920494428153e-04
GC_7_423 b_7 NI_7 NS_423 0 -1.2864878741512231e-04
GC_7_424 b_7 NI_7 NS_424 0 -6.9474722913984215e-05
GC_7_425 b_7 NI_7 NS_425 0 -2.0656948235934416e-03
GC_7_426 b_7 NI_7 NS_426 0 1.0998431088655470e-04
GC_7_427 b_7 NI_7 NS_427 0 -1.2583815430837339e-05
GC_7_428 b_7 NI_7 NS_428 0 4.3597938609654304e-05
GC_7_429 b_7 NI_7 NS_429 0 -3.1386874931827819e-04
GC_7_430 b_7 NI_7 NS_430 0 4.5855053122625330e-06
GC_7_431 b_7 NI_7 NS_431 0 1.7956689939263842e-03
GC_7_432 b_7 NI_7 NS_432 0 -1.6189845445517979e-03
GC_7_433 b_7 NI_7 NS_433 0 1.6420192561298345e-04
GC_7_434 b_7 NI_7 NS_434 0 -1.0933660562329580e-04
GC_7_435 b_7 NI_7 NS_435 0 -9.1430453361306615e-07
GC_7_436 b_7 NI_7 NS_436 0 5.7008151200381833e-07
GC_7_437 b_7 NI_7 NS_437 0 -3.3604341693647267e-06
GC_7_438 b_7 NI_7 NS_438 0 -8.5252954626182258e-06
GC_7_439 b_7 NI_7 NS_439 0 -1.3595339613434789e-04
GC_7_440 b_7 NI_7 NS_440 0 1.3045759120776374e-04
GC_7_441 b_7 NI_7 NS_441 0 -2.8519312401497478e-07
GC_7_442 b_7 NI_7 NS_442 0 -2.0711806879558494e-05
GC_7_443 b_7 NI_7 NS_443 0 -4.5062864523304360e-06
GC_7_444 b_7 NI_7 NS_444 0 -4.1284726552457513e-06
GC_7_445 b_7 NI_7 NS_445 0 4.7744941253621739e-05
GC_7_446 b_7 NI_7 NS_446 0 -1.4665627501920916e-05
GC_7_447 b_7 NI_7 NS_447 0 -7.3836531193764989e-05
GC_7_448 b_7 NI_7 NS_448 0 3.5158644673219927e-07
GC_7_449 b_7 NI_7 NS_449 0 1.9416340477248037e-03
GC_7_450 b_7 NI_7 NS_450 0 3.2031069121061846e-05
GC_7_451 b_7 NI_7 NS_451 0 1.2362677810949087e-03
GC_7_452 b_7 NI_7 NS_452 0 -1.4019328443516641e-04
GC_7_453 b_7 NI_7 NS_453 0 -1.1064620981862752e-03
GC_7_454 b_7 NI_7 NS_454 0 1.3027347410189706e-03
GC_7_455 b_7 NI_7 NS_455 0 -9.4255987248407841e-04
GC_7_456 b_7 NI_7 NS_456 0 7.3844347527987143e-04
GC_7_457 b_7 NI_7 NS_457 0 -2.7176362442539702e-03
GC_7_458 b_7 NI_7 NS_458 0 -2.9728876614769292e-03
GC_7_459 b_7 NI_7 NS_459 0 -4.2741186297398469e-04
GC_7_460 b_7 NI_7 NS_460 0 -2.8669292556414937e-04
GC_7_461 b_7 NI_7 NS_461 0 2.8452512812607179e-03
GC_7_462 b_7 NI_7 NS_462 0 -1.5783737902452875e-03
GC_7_463 b_7 NI_7 NS_463 0 1.2720878519667789e-03
GC_7_464 b_7 NI_7 NS_464 0 5.0811948482776443e-04
GC_7_465 b_7 NI_7 NS_465 0 -1.2121712727414741e-03
GC_7_466 b_7 NI_7 NS_466 0 3.9743192887015566e-05
GC_7_467 b_7 NI_7 NS_467 0 1.7014784482072124e-03
GC_7_468 b_7 NI_7 NS_468 0 2.6297830655008575e-04
GC_7_469 b_7 NI_7 NS_469 0 4.7531370668388057e-04
GC_7_470 b_7 NI_7 NS_470 0 2.3895384275885101e-04
GC_7_471 b_7 NI_7 NS_471 0 5.6138880223451462e-04
GC_7_472 b_7 NI_7 NS_472 0 5.2959347769498738e-03
GC_7_473 b_7 NI_7 NS_473 0 -3.8315521011859227e-04
GC_7_474 b_7 NI_7 NS_474 0 -7.1333702535724243e-04
GC_7_475 b_7 NI_7 NS_475 0 -8.5783890823391904e-04
GC_7_476 b_7 NI_7 NS_476 0 5.5285626863937674e-05
GC_7_477 b_7 NI_7 NS_477 0 -3.1464640976360052e-04
GC_7_478 b_7 NI_7 NS_478 0 -2.8183841873436957e-04
GC_7_479 b_7 NI_7 NS_479 0 -7.7628730691232763e-05
GC_7_480 b_7 NI_7 NS_480 0 1.2030353622625843e-05
GC_7_481 b_7 NI_7 NS_481 0 -3.3267425705263858e-03
GC_7_482 b_7 NI_7 NS_482 0 -3.9758477081037946e-03
GC_7_483 b_7 NI_7 NS_483 0 2.1321771538213565e-05
GC_7_484 b_7 NI_7 NS_484 0 -4.9501045425208177e-05
GC_7_485 b_7 NI_7 NS_485 0 1.7771430906501565e-04
GC_7_486 b_7 NI_7 NS_486 0 7.0102832119618231e-04
GC_7_487 b_7 NI_7 NS_487 0 1.9353827545452115e-03
GC_7_488 b_7 NI_7 NS_488 0 7.4141649333171744e-04
GC_7_489 b_7 NI_7 NS_489 0 9.7630824368022689e-06
GC_7_490 b_7 NI_7 NS_490 0 2.8783995955702181e-04
GC_7_491 b_7 NI_7 NS_491 0 -7.9279169472216695e-07
GC_7_492 b_7 NI_7 NS_492 0 8.8023398284171155e-07
GC_7_493 b_7 NI_7 NS_493 0 3.0800025171703479e-06
GC_7_494 b_7 NI_7 NS_494 0 -1.3996584621727187e-06
GC_7_495 b_7 NI_7 NS_495 0 -6.9636293523275532e-05
GC_7_496 b_7 NI_7 NS_496 0 -4.4378253013111257e-06
GC_7_497 b_7 NI_7 NS_497 0 6.0845856910755715e-06
GC_7_498 b_7 NI_7 NS_498 0 -1.4896805142121222e-06
GC_7_499 b_7 NI_7 NS_499 0 -4.2626239907210441e-06
GC_7_500 b_7 NI_7 NS_500 0 -4.5033614261094362e-06
GC_7_501 b_7 NI_7 NS_501 0 1.4125508773382949e-05
GC_7_502 b_7 NI_7 NS_502 0 -4.5832129628627790e-07
GC_7_503 b_7 NI_7 NS_503 0 -2.1253532751351136e-05
GC_7_504 b_7 NI_7 NS_504 0 -4.8241592713713076e-06
GC_7_505 b_7 NI_7 NS_505 0 9.1985770989384159e-03
GC_7_506 b_7 NI_7 NS_506 0 -1.0820501378984417e-04
GC_7_507 b_7 NI_7 NS_507 0 -1.6063129023330595e-04
GC_7_508 b_7 NI_7 NS_508 0 7.1864938050028809e-04
GC_7_509 b_7 NI_7 NS_509 0 -3.0035343932253522e-04
GC_7_510 b_7 NI_7 NS_510 0 -6.6812393559640142e-04
GC_7_511 b_7 NI_7 NS_511 0 -5.3910156607360124e-04
GC_7_512 b_7 NI_7 NS_512 0 -6.6289476589820220e-04
GC_7_513 b_7 NI_7 NS_513 0 2.2077767129615755e-03
GC_7_514 b_7 NI_7 NS_514 0 8.7822518735310422e-04
GC_7_515 b_7 NI_7 NS_515 0 -5.8618430119382228e-04
GC_7_516 b_7 NI_7 NS_516 0 -6.0962253889866748e-05
GC_7_517 b_7 NI_7 NS_517 0 5.0516146836935931e-04
GC_7_518 b_7 NI_7 NS_518 0 -5.4384456051354045e-04
GC_7_519 b_7 NI_7 NS_519 0 1.0216386658711374e-03
GC_7_520 b_7 NI_7 NS_520 0 -1.8622408191131201e-04
GC_7_521 b_7 NI_7 NS_521 0 9.0450363067691691e-04
GC_7_522 b_7 NI_7 NS_522 0 2.4153264421862878e-03
GC_7_523 b_7 NI_7 NS_523 0 -1.3445721143413418e-03
GC_7_524 b_7 NI_7 NS_524 0 2.8634763232446513e-03
GC_7_525 b_7 NI_7 NS_525 0 -2.7446836934943758e-04
GC_7_526 b_7 NI_7 NS_526 0 -7.7418457258273166e-05
GC_7_527 b_7 NI_7 NS_527 0 -7.8717474944824378e-04
GC_7_528 b_7 NI_7 NS_528 0 1.9332009858710972e-03
GC_7_529 b_7 NI_7 NS_529 0 8.3349822201380741e-05
GC_7_530 b_7 NI_7 NS_530 0 -4.1723557272405908e-05
GC_7_531 b_7 NI_7 NS_531 0 -7.6069469408923229e-04
GC_7_532 b_7 NI_7 NS_532 0 2.5886898945016925e-04
GC_7_533 b_7 NI_7 NS_533 0 -4.9253576842020832e-04
GC_7_534 b_7 NI_7 NS_534 0 9.6951372476714186e-05
GC_7_535 b_7 NI_7 NS_535 0 -1.2771378812152242e-04
GC_7_536 b_7 NI_7 NS_536 0 -3.2309038683280210e-05
GC_7_537 b_7 NI_7 NS_537 0 -1.4100993532129660e-03
GC_7_538 b_7 NI_7 NS_538 0 -2.8958206540548479e-03
GC_7_539 b_7 NI_7 NS_539 0 3.0377894405012113e-05
GC_7_540 b_7 NI_7 NS_540 0 -2.9095056493627517e-05
GC_7_541 b_7 NI_7 NS_541 0 -8.3607874690853792e-04
GC_7_542 b_7 NI_7 NS_542 0 5.5527328898710140e-04
GC_7_543 b_7 NI_7 NS_543 0 1.1176247829539827e-03
GC_7_544 b_7 NI_7 NS_544 0 -2.8919811407196092e-04
GC_7_545 b_7 NI_7 NS_545 0 -1.0514581613633885e-04
GC_7_546 b_7 NI_7 NS_546 0 1.5838089721766319e-04
GC_7_547 b_7 NI_7 NS_547 0 -1.9868375409852420e-06
GC_7_548 b_7 NI_7 NS_548 0 2.5378489837198238e-06
GC_7_549 b_7 NI_7 NS_549 0 -2.0655322968377255e-06
GC_7_550 b_7 NI_7 NS_550 0 -3.9515092409119731e-06
GC_7_551 b_7 NI_7 NS_551 0 -4.8380755288607008e-05
GC_7_552 b_7 NI_7 NS_552 0 7.0574630662485551e-05
GC_7_553 b_7 NI_7 NS_553 0 2.3995859699995955e-06
GC_7_554 b_7 NI_7 NS_554 0 -1.0993444398806265e-05
GC_7_555 b_7 NI_7 NS_555 0 -1.9735405225411254e-06
GC_7_556 b_7 NI_7 NS_556 0 -4.9972427498075156e-06
GC_7_557 b_7 NI_7 NS_557 0 2.4599797672495279e-05
GC_7_558 b_7 NI_7 NS_558 0 -4.1451023789745232e-05
GC_7_559 b_7 NI_7 NS_559 0 -4.9294270682901142e-05
GC_7_560 b_7 NI_7 NS_560 0 5.5827426882182847e-05
GC_7_561 b_7 NI_7 NS_561 0 -1.7513274191163383e-02
GC_7_562 b_7 NI_7 NS_562 0 6.2692913950541745e-04
GC_7_563 b_7 NI_7 NS_563 0 8.0498192394194441e-04
GC_7_564 b_7 NI_7 NS_564 0 8.1000824932674802e-04
GC_7_565 b_7 NI_7 NS_565 0 -1.6184484045361671e-03
GC_7_566 b_7 NI_7 NS_566 0 -2.4432493191596343e-03
GC_7_567 b_7 NI_7 NS_567 0 1.2162876038703263e-03
GC_7_568 b_7 NI_7 NS_568 0 -3.6566454443763048e-04
GC_7_569 b_7 NI_7 NS_569 0 4.0419266586423702e-03
GC_7_570 b_7 NI_7 NS_570 0 -4.0562196170569427e-03
GC_7_571 b_7 NI_7 NS_571 0 -3.1815896679466643e-04
GC_7_572 b_7 NI_7 NS_572 0 1.6430966133070441e-04
GC_7_573 b_7 NI_7 NS_573 0 2.5152980162466893e-03
GC_7_574 b_7 NI_7 NS_574 0 -1.6564678125002689e-04
GC_7_575 b_7 NI_7 NS_575 0 1.0452547707196630e-03
GC_7_576 b_7 NI_7 NS_576 0 6.4452650446861659e-04
GC_7_577 b_7 NI_7 NS_577 0 1.0876289110995235e-03
GC_7_578 b_7 NI_7 NS_578 0 -1.5186341414447522e-03
GC_7_579 b_7 NI_7 NS_579 0 2.5713168007455559e-03
GC_7_580 b_7 NI_7 NS_580 0 -1.7437366641275516e-04
GC_7_581 b_7 NI_7 NS_581 0 3.5079276319887638e-04
GC_7_582 b_7 NI_7 NS_582 0 1.7554417196054457e-04
GC_7_583 b_7 NI_7 NS_583 0 2.4325350531634485e-03
GC_7_584 b_7 NI_7 NS_584 0 5.7447965226383986e-03
GC_7_585 b_7 NI_7 NS_585 0 -5.9984672812242640e-05
GC_7_586 b_7 NI_7 NS_586 0 -6.7719109870962495e-04
GC_7_587 b_7 NI_7 NS_587 0 -6.0503983355215528e-04
GC_7_588 b_7 NI_7 NS_588 0 1.8785373372793475e-04
GC_7_589 b_7 NI_7 NS_589 0 -1.6670827904258323e-04
GC_7_590 b_7 NI_7 NS_590 0 -1.0491864427533381e-04
GC_7_591 b_7 NI_7 NS_591 0 -6.3607770944085687e-05
GC_7_592 b_7 NI_7 NS_592 0 2.4854902125176369e-05
GC_7_593 b_7 NI_7 NS_593 0 8.3313264989172669e-04
GC_7_594 b_7 NI_7 NS_594 0 1.0473768561850142e-03
GC_7_595 b_7 NI_7 NS_595 0 1.4736836908016978e-05
GC_7_596 b_7 NI_7 NS_596 0 -3.1671095305039369e-05
GC_7_597 b_7 NI_7 NS_597 0 3.7319105064010017e-04
GC_7_598 b_7 NI_7 NS_598 0 4.1477653696333079e-04
GC_7_599 b_7 NI_7 NS_599 0 -2.2355184734368680e-03
GC_7_600 b_7 NI_7 NS_600 0 5.8076485757799440e-04
GC_7_601 b_7 NI_7 NS_601 0 -1.6288533290259409e-04
GC_7_602 b_7 NI_7 NS_602 0 -2.2751855138467616e-04
GC_7_603 b_7 NI_7 NS_603 0 1.3468051966644361e-06
GC_7_604 b_7 NI_7 NS_604 0 -5.0923232848472253e-07
GC_7_605 b_7 NI_7 NS_605 0 7.3044406817345779e-06
GC_7_606 b_7 NI_7 NS_606 0 9.0616786473065354e-06
GC_7_607 b_7 NI_7 NS_607 0 1.3378574547620809e-04
GC_7_608 b_7 NI_7 NS_608 0 -1.5806843204310811e-04
GC_7_609 b_7 NI_7 NS_609 0 5.9660815146600699e-06
GC_7_610 b_7 NI_7 NS_610 0 2.2325765582574377e-05
GC_7_611 b_7 NI_7 NS_611 0 6.0023983387604992e-06
GC_7_612 b_7 NI_7 NS_612 0 6.8479528775348272e-06
GC_7_613 b_7 NI_7 NS_613 0 -3.7525102279885913e-05
GC_7_614 b_7 NI_7 NS_614 0 2.0239371137867120e-05
GC_7_615 b_7 NI_7 NS_615 0 6.7721926180459364e-05
GC_7_616 b_7 NI_7 NS_616 0 -9.5876283356738320e-06
GC_7_617 b_7 NI_7 NS_617 0 2.6113910399560666e-02
GC_7_618 b_7 NI_7 NS_618 0 -2.8081568320264681e-04
GC_7_619 b_7 NI_7 NS_619 0 -4.7191378253243741e-04
GC_7_620 b_7 NI_7 NS_620 0 5.6101976288284094e-04
GC_7_621 b_7 NI_7 NS_621 0 1.0796920309497724e-03
GC_7_622 b_7 NI_7 NS_622 0 2.3879991424983056e-04
GC_7_623 b_7 NI_7 NS_623 0 -1.1434196351042161e-03
GC_7_624 b_7 NI_7 NS_624 0 9.1466303617375986e-04
GC_7_625 b_7 NI_7 NS_625 0 -2.7851048566760669e-03
GC_7_626 b_7 NI_7 NS_626 0 4.4659259725283529e-03
GC_7_627 b_7 NI_7 NS_627 0 -3.7630184465256941e-04
GC_7_628 b_7 NI_7 NS_628 0 1.1957781522193980e-04
GC_7_629 b_7 NI_7 NS_629 0 5.7688607417266991e-05
GC_7_630 b_7 NI_7 NS_630 0 -1.2281864553706902e-03
GC_7_631 b_7 NI_7 NS_631 0 7.6765881944232492e-04
GC_7_632 b_7 NI_7 NS_632 0 1.3467173557900770e-04
GC_7_633 b_7 NI_7 NS_633 0 -4.5904687874349221e-04
GC_7_634 b_7 NI_7 NS_634 0 6.9709949778156593e-04
GC_7_635 b_7 NI_7 NS_635 0 -1.6687602019109322e-03
GC_7_636 b_7 NI_7 NS_636 0 9.5919841623389986e-04
GC_7_637 b_7 NI_7 NS_637 0 -1.2970759022220090e-04
GC_7_638 b_7 NI_7 NS_638 0 -8.9930709460930055e-05
GC_7_639 b_7 NI_7 NS_639 0 1.3907437472162256e-04
GC_7_640 b_7 NI_7 NS_640 0 2.1918276102541453e-03
GC_7_641 b_7 NI_7 NS_641 0 5.7125449278527534e-05
GC_7_642 b_7 NI_7 NS_642 0 -1.8310638396010779e-04
GC_7_643 b_7 NI_7 NS_643 0 -5.0642899256663539e-04
GC_7_644 b_7 NI_7 NS_644 0 1.5579893701996999e-04
GC_7_645 b_7 NI_7 NS_645 0 -3.0540480418361266e-04
GC_7_646 b_7 NI_7 NS_646 0 1.2386945641429417e-04
GC_7_647 b_7 NI_7 NS_647 0 -9.8125158265736887e-05
GC_7_648 b_7 NI_7 NS_648 0 -1.7925822106694510e-05
GC_7_649 b_7 NI_7 NS_649 0 -1.0666344494805024e-03
GC_7_650 b_7 NI_7 NS_650 0 4.9152476372507008e-04
GC_7_651 b_7 NI_7 NS_651 0 2.7611644512680409e-05
GC_7_652 b_7 NI_7 NS_652 0 -1.8833014962130707e-05
GC_7_653 b_7 NI_7 NS_653 0 -5.0002447538430111e-04
GC_7_654 b_7 NI_7 NS_654 0 4.8131757480364152e-04
GC_7_655 b_7 NI_7 NS_655 0 -1.7105298186980756e-03
GC_7_656 b_7 NI_7 NS_656 0 -1.7722953190643545e-03
GC_7_657 b_7 NI_7 NS_657 0 -1.9516320925264954e-04
GC_7_658 b_7 NI_7 NS_658 0 -6.8472775576559536e-05
GC_7_659 b_7 NI_7 NS_659 0 -8.5581324188424492e-08
GC_7_660 b_7 NI_7 NS_660 0 1.0152563601776208e-06
GC_7_661 b_7 NI_7 NS_661 0 -6.1146546546799872e-06
GC_7_662 b_7 NI_7 NS_662 0 -3.2297373997504695e-06
GC_7_663 b_7 NI_7 NS_663 0 7.4821653403485012e-05
GC_7_664 b_7 NI_7 NS_664 0 1.2540044745888398e-04
GC_7_665 b_7 NI_7 NS_665 0 -8.7626478164731640e-06
GC_7_666 b_7 NI_7 NS_666 0 -1.0173665950323262e-05
GC_7_667 b_7 NI_7 NS_667 0 -3.7344315344775170e-06
GC_7_668 b_7 NI_7 NS_668 0 3.8930408997456101e-06
GC_7_669 b_7 NI_7 NS_669 0 8.0137038748085305e-06
GC_7_670 b_7 NI_7 NS_670 0 -4.3991496038594260e-05
GC_7_671 b_7 NI_7 NS_671 0 -2.9717983490859048e-05
GC_7_672 b_7 NI_7 NS_672 0 6.4752625915261874e-05
GD_7_1 b_7 NI_7 NA_1 0 -8.1417525917316158e-02
GD_7_2 b_7 NI_7 NA_2 0 4.0311334785615174e-02
GD_7_3 b_7 NI_7 NA_3 0 -4.4479508840142540e-02
GD_7_4 b_7 NI_7 NA_4 0 6.2067249436090670e-03
GD_7_5 b_7 NI_7 NA_5 0 -8.8798903932468653e-03
GD_7_6 b_7 NI_7 NA_6 0 -5.3950200966555152e-02
GD_7_7 b_7 NI_7 NA_7 0 -1.1840012451103814e-01
GD_7_8 b_7 NI_7 NA_8 0 1.1794143850451896e-02
GD_7_9 b_7 NI_7 NA_9 0 -7.4585849631141554e-04
GD_7_10 b_7 NI_7 NA_10 0 -1.2216992980849823e-02
GD_7_11 b_7 NI_7 NA_11 0 5.8730314809384929e-03
GD_7_12 b_7 NI_7 NA_12 0 -2.7059768597431776e-02
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 -3.7701362339117923e-02
GC_8_2 b_8 NI_8 NS_2 0 -9.0949517691875411e-05
GC_8_3 b_8 NI_8 NS_3 0 -3.4758651154012714e-04
GC_8_4 b_8 NI_8 NS_4 0 2.3768057867345283e-03
GC_8_5 b_8 NI_8 NS_5 0 -2.4923580644024292e-03
GC_8_6 b_8 NI_8 NS_6 0 -1.4025237067786145e-03
GC_8_7 b_8 NI_8 NS_7 0 -5.5894393074068750e-03
GC_8_8 b_8 NI_8 NS_8 0 -6.1963786255550624e-03
GC_8_9 b_8 NI_8 NS_9 0 7.9811227553672533e-03
GC_8_10 b_8 NI_8 NS_10 0 -9.6907931229274717e-03
GC_8_11 b_8 NI_8 NS_11 0 3.0169147987239801e-05
GC_8_12 b_8 NI_8 NS_12 0 5.5634538323658816e-04
GC_8_13 b_8 NI_8 NS_13 0 5.1817747285672578e-03
GC_8_14 b_8 NI_8 NS_14 0 -2.0646373902258107e-03
GC_8_15 b_8 NI_8 NS_15 0 4.0474550878685106e-04
GC_8_16 b_8 NI_8 NS_16 0 4.6321923703225500e-04
GC_8_17 b_8 NI_8 NS_17 0 8.7973404643514237e-04
GC_8_18 b_8 NI_8 NS_18 0 2.1873013167598714e-03
GC_8_19 b_8 NI_8 NS_19 0 -1.4206434911967045e-06
GC_8_20 b_8 NI_8 NS_20 0 7.6879833360049351e-05
GC_8_21 b_8 NI_8 NS_21 0 -1.5187627701662986e-04
GC_8_22 b_8 NI_8 NS_22 0 1.0322612231400896e-04
GC_8_23 b_8 NI_8 NS_23 0 6.5162768212875929e-04
GC_8_24 b_8 NI_8 NS_24 0 -4.1065977893939712e-03
GC_8_25 b_8 NI_8 NS_25 0 -8.1744060234879335e-04
GC_8_26 b_8 NI_8 NS_26 0 2.7486033359995634e-04
GC_8_27 b_8 NI_8 NS_27 0 -2.9096148470728116e-06
GC_8_28 b_8 NI_8 NS_28 0 -3.0287635173485761e-05
GC_8_29 b_8 NI_8 NS_29 0 -2.2523373499274495e-04
GC_8_30 b_8 NI_8 NS_30 0 -8.7724037906983341e-05
GC_8_31 b_8 NI_8 NS_31 0 -7.0284200181654083e-05
GC_8_32 b_8 NI_8 NS_32 0 -1.4317018525544168e-04
GC_8_33 b_8 NI_8 NS_33 0 9.2805573395963528e-03
GC_8_34 b_8 NI_8 NS_34 0 8.0023686719944221e-04
GC_8_35 b_8 NI_8 NS_35 0 -5.9514575065484083e-05
GC_8_36 b_8 NI_8 NS_36 0 1.3298812055321960e-04
GC_8_37 b_8 NI_8 NS_37 0 -5.7895331746050623e-04
GC_8_38 b_8 NI_8 NS_38 0 -1.7065018604394365e-03
GC_8_39 b_8 NI_8 NS_39 0 -5.2353237640212220e-04
GC_8_40 b_8 NI_8 NS_40 0 2.3359122362103767e-03
GC_8_41 b_8 NI_8 NS_41 0 -4.6952452662645341e-04
GC_8_42 b_8 NI_8 NS_42 0 -2.9728910195324923e-04
GC_8_43 b_8 NI_8 NS_43 0 -1.2103061999836554e-07
GC_8_44 b_8 NI_8 NS_44 0 -1.3562405209713885e-06
GC_8_45 b_8 NI_8 NS_45 0 5.3033514290090266e-06
GC_8_46 b_8 NI_8 NS_46 0 1.3704186934945203e-05
GC_8_47 b_8 NI_8 NS_47 0 1.6474620008079973e-04
GC_8_48 b_8 NI_8 NS_48 0 -1.4824621166130493e-04
GC_8_49 b_8 NI_8 NS_49 0 -4.9275000630012078e-08
GC_8_50 b_8 NI_8 NS_50 0 2.5780093194347015e-05
GC_8_51 b_8 NI_8 NS_51 0 1.3619426543821471e-05
GC_8_52 b_8 NI_8 NS_52 0 -7.5222429831532371e-07
GC_8_53 b_8 NI_8 NS_53 0 -3.5922423279747189e-05
GC_8_54 b_8 NI_8 NS_54 0 3.8364746744645178e-05
GC_8_55 b_8 NI_8 NS_55 0 6.8212066014245587e-05
GC_8_56 b_8 NI_8 NS_56 0 -3.3336323581681639e-05
GC_8_57 b_8 NI_8 NS_57 0 3.5910367315377334e-02
GC_8_58 b_8 NI_8 NS_58 0 -3.1429226743136620e-04
GC_8_59 b_8 NI_8 NS_59 0 -9.8606758519918748e-04
GC_8_60 b_8 NI_8 NS_60 0 -7.4407239656676231e-04
GC_8_61 b_8 NI_8 NS_61 0 1.3776247464893981e-03
GC_8_62 b_8 NI_8 NS_62 0 -5.8709030361661695e-04
GC_8_63 b_8 NI_8 NS_63 0 5.8524960557292784e-03
GC_8_64 b_8 NI_8 NS_64 0 1.0117589782781267e-03
GC_8_65 b_8 NI_8 NS_65 0 -2.3683178004469257e-03
GC_8_66 b_8 NI_8 NS_66 0 1.0272689602108722e-02
GC_8_67 b_8 NI_8 NS_67 0 -6.2157140847982409e-04
GC_8_68 b_8 NI_8 NS_68 0 5.6000171216566473e-04
GC_8_69 b_8 NI_8 NS_69 0 -1.2606988330545394e-03
GC_8_70 b_8 NI_8 NS_70 0 -1.0364921425743199e-03
GC_8_71 b_8 NI_8 NS_71 0 7.4875507557971743e-04
GC_8_72 b_8 NI_8 NS_72 0 4.8267935796434514e-04
GC_8_73 b_8 NI_8 NS_73 0 4.9234937065061231e-04
GC_8_74 b_8 NI_8 NS_74 0 5.3901312214271113e-03
GC_8_75 b_8 NI_8 NS_75 0 3.5274397044036569e-04
GC_8_76 b_8 NI_8 NS_76 0 1.7455762014535698e-04
GC_8_77 b_8 NI_8 NS_77 0 1.2493285449657830e-04
GC_8_78 b_8 NI_8 NS_78 0 -9.6936990730190278e-05
GC_8_79 b_8 NI_8 NS_79 0 -5.3911521061958071e-03
GC_8_80 b_8 NI_8 NS_80 0 6.9711323626783272e-03
GC_8_81 b_8 NI_8 NS_81 0 6.0619714866488991e-04
GC_8_82 b_8 NI_8 NS_82 0 -9.4366346682388266e-05
GC_8_83 b_8 NI_8 NS_83 0 -3.9814487410868183e-04
GC_8_84 b_8 NI_8 NS_84 0 8.4054051878379632e-06
GC_8_85 b_8 NI_8 NS_85 0 -2.3339141158918872e-05
GC_8_86 b_8 NI_8 NS_86 0 9.1540846724593849e-05
GC_8_87 b_8 NI_8 NS_87 0 1.1974575860350826e-04
GC_8_88 b_8 NI_8 NS_88 0 2.7722550734265016e-05
GC_8_89 b_8 NI_8 NS_89 0 -1.4763940327449938e-02
GC_8_90 b_8 NI_8 NS_90 0 -2.3762289663730499e-03
GC_8_91 b_8 NI_8 NS_91 0 -4.2613218751471486e-05
GC_8_92 b_8 NI_8 NS_92 0 -2.3098353251976766e-04
GC_8_93 b_8 NI_8 NS_93 0 2.2834434537554282e-03
GC_8_94 b_8 NI_8 NS_94 0 2.8685343114617039e-03
GC_8_95 b_8 NI_8 NS_95 0 5.0342847802211941e-03
GC_8_96 b_8 NI_8 NS_96 0 -5.9581456547065205e-03
GC_8_97 b_8 NI_8 NS_97 0 5.1150303657498150e-04
GC_8_98 b_8 NI_8 NS_98 0 5.9032712986205088e-04
GC_8_99 b_8 NI_8 NS_99 0 1.4572920346562476e-06
GC_8_100 b_8 NI_8 NS_100 0 1.6908306902622924e-06
GC_8_101 b_8 NI_8 NS_101 0 -2.7054273301181821e-05
GC_8_102 b_8 NI_8 NS_102 0 -2.9496064331023846e-05
GC_8_103 b_8 NI_8 NS_103 0 -2.5735080158102291e-04
GC_8_104 b_8 NI_8 NS_104 0 4.3914125023765513e-04
GC_8_105 b_8 NI_8 NS_105 0 -3.6131219803846711e-05
GC_8_106 b_8 NI_8 NS_106 0 -5.5776953002320738e-05
GC_8_107 b_8 NI_8 NS_107 0 -4.1377972421387506e-05
GC_8_108 b_8 NI_8 NS_108 0 -8.0878654924007422e-06
GC_8_109 b_8 NI_8 NS_109 0 2.2984231418618752e-04
GC_8_110 b_8 NI_8 NS_110 0 -1.7204653426360682e-04
GC_8_111 b_8 NI_8 NS_111 0 -4.1222525109969616e-04
GC_8_112 b_8 NI_8 NS_112 0 1.5602551283216843e-04
GC_8_113 b_8 NI_8 NS_113 0 -4.7108844398643258e-03
GC_8_114 b_8 NI_8 NS_114 0 -2.7057613611124881e-04
GC_8_115 b_8 NI_8 NS_115 0 -1.2981495452324512e-03
GC_8_116 b_8 NI_8 NS_116 0 2.9646937939682154e-03
GC_8_117 b_8 NI_8 NS_117 0 -9.0101273618577377e-04
GC_8_118 b_8 NI_8 NS_118 0 -2.1585934591388206e-03
GC_8_119 b_8 NI_8 NS_119 0 -4.8241010355927864e-03
GC_8_120 b_8 NI_8 NS_120 0 -5.2327791563066490e-03
GC_8_121 b_8 NI_8 NS_121 0 6.6113530061501181e-03
GC_8_122 b_8 NI_8 NS_122 0 -1.2399264939466589e-03
GC_8_123 b_8 NI_8 NS_123 0 -2.7231652954970269e-04
GC_8_124 b_8 NI_8 NS_124 0 -5.8239358577085053e-05
GC_8_125 b_8 NI_8 NS_125 0 3.9896801950792182e-03
GC_8_126 b_8 NI_8 NS_126 0 -2.5678389338233518e-03
GC_8_127 b_8 NI_8 NS_127 0 7.3641777279517470e-04
GC_8_128 b_8 NI_8 NS_128 0 1.0236524976485945e-03
GC_8_129 b_8 NI_8 NS_129 0 7.3404456570490327e-04
GC_8_130 b_8 NI_8 NS_130 0 2.3515104468547878e-03
GC_8_131 b_8 NI_8 NS_131 0 -3.0485347367965477e-03
GC_8_132 b_8 NI_8 NS_132 0 1.0842577934802597e-03
GC_8_133 b_8 NI_8 NS_133 0 -1.9783189680264729e-04
GC_8_134 b_8 NI_8 NS_134 0 -8.6295389435328291e-06
GC_8_135 b_8 NI_8 NS_135 0 2.3282267874790564e-03
GC_8_136 b_8 NI_8 NS_136 0 5.7151092053213056e-04
GC_8_137 b_8 NI_8 NS_137 0 -7.9255932660440343e-04
GC_8_138 b_8 NI_8 NS_138 0 -1.0153501657687751e-04
GC_8_139 b_8 NI_8 NS_139 0 -2.7113352381955415e-04
GC_8_140 b_8 NI_8 NS_140 0 6.1973332087672544e-05
GC_8_141 b_8 NI_8 NS_141 0 -3.4873616518592011e-04
GC_8_142 b_8 NI_8 NS_142 0 1.9196022250065958e-04
GC_8_143 b_8 NI_8 NS_143 0 -1.6152454343230097e-04
GC_8_144 b_8 NI_8 NS_144 0 -1.0442915857276137e-04
GC_8_145 b_8 NI_8 NS_145 0 7.8243403053790731e-04
GC_8_146 b_8 NI_8 NS_146 0 -4.3737885597535140e-04
GC_8_147 b_8 NI_8 NS_147 0 -4.1987216208936425e-05
GC_8_148 b_8 NI_8 NS_148 0 8.3393285725287552e-05
GC_8_149 b_8 NI_8 NS_149 0 -2.9876630299346398e-04
GC_8_150 b_8 NI_8 NS_150 0 -6.1646384841066034e-04
GC_8_151 b_8 NI_8 NS_151 0 2.0354368494853941e-04
GC_8_152 b_8 NI_8 NS_152 0 9.6545422649131044e-04
GC_8_153 b_8 NI_8 NS_153 0 -3.6004383185213625e-06
GC_8_154 b_8 NI_8 NS_154 0 -1.0300740019439410e-04
GC_8_155 b_8 NI_8 NS_155 0 2.2385732610214035e-07
GC_8_156 b_8 NI_8 NS_156 0 -1.3347125161928656e-08
GC_8_157 b_8 NI_8 NS_157 0 7.6529026012833897e-07
GC_8_158 b_8 NI_8 NS_158 0 4.8152492440183336e-06
GC_8_159 b_8 NI_8 NS_159 0 3.3833487260139727e-05
GC_8_160 b_8 NI_8 NS_160 0 -6.0533840475718263e-05
GC_8_161 b_8 NI_8 NS_161 0 -2.4540247746433256e-07
GC_8_162 b_8 NI_8 NS_162 0 9.1689172101014618e-06
GC_8_163 b_8 NI_8 NS_163 0 1.7848319040184138e-06
GC_8_164 b_8 NI_8 NS_164 0 4.1267889074732776e-07
GC_8_165 b_8 NI_8 NS_165 0 -1.7052453410798780e-05
GC_8_166 b_8 NI_8 NS_166 0 -3.6587089270224698e-06
GC_8_167 b_8 NI_8 NS_167 0 2.0952939396572112e-05
GC_8_168 b_8 NI_8 NS_168 0 1.2817498122600194e-05
GC_8_169 b_8 NI_8 NS_169 0 1.1842650810292668e-02
GC_8_170 b_8 NI_8 NS_170 0 -7.2521038553269984e-04
GC_8_171 b_8 NI_8 NS_171 0 -1.1313545394730366e-03
GC_8_172 b_8 NI_8 NS_172 0 -1.1311517575342746e-03
GC_8_173 b_8 NI_8 NS_173 0 9.5330693731836454e-04
GC_8_174 b_8 NI_8 NS_174 0 3.3415515629529023e-04
GC_8_175 b_8 NI_8 NS_175 0 4.1690772209938094e-03
GC_8_176 b_8 NI_8 NS_176 0 1.0302037479530395e-03
GC_8_177 b_8 NI_8 NS_177 0 -5.8912814116800528e-03
GC_8_178 b_8 NI_8 NS_178 0 3.3053768409968941e-03
GC_8_179 b_8 NI_8 NS_179 0 -4.9250640759443366e-04
GC_8_180 b_8 NI_8 NS_180 0 3.5152937801968581e-04
GC_8_181 b_8 NI_8 NS_181 0 2.6535154767815764e-04
GC_8_182 b_8 NI_8 NS_182 0 -3.2422231045397638e-03
GC_8_183 b_8 NI_8 NS_183 0 6.2509022745122790e-04
GC_8_184 b_8 NI_8 NS_184 0 4.1636414722856480e-04
GC_8_185 b_8 NI_8 NS_185 0 2.4331667145777487e-04
GC_8_186 b_8 NI_8 NS_186 0 1.5777783061692423e-03
GC_8_187 b_8 NI_8 NS_187 0 9.3434572320551126e-04
GC_8_188 b_8 NI_8 NS_188 0 -1.1539185529056088e-03
GC_8_189 b_8 NI_8 NS_189 0 5.9006497812733951e-05
GC_8_190 b_8 NI_8 NS_190 0 -9.8351545604651395e-06
GC_8_191 b_8 NI_8 NS_191 0 8.5116331058316948e-04
GC_8_192 b_8 NI_8 NS_192 0 2.4042279701405470e-03
GC_8_193 b_8 NI_8 NS_193 0 1.2560314525198431e-04
GC_8_194 b_8 NI_8 NS_194 0 5.7032581258312694e-05
GC_8_195 b_8 NI_8 NS_195 0 -2.0477979791696152e-04
GC_8_196 b_8 NI_8 NS_196 0 1.7448236318041321e-05
GC_8_197 b_8 NI_8 NS_197 0 1.0462875316985923e-04
GC_8_198 b_8 NI_8 NS_198 0 -1.3838927664821214e-04
GC_8_199 b_8 NI_8 NS_199 0 2.0754026954036340e-04
GC_8_200 b_8 NI_8 NS_200 0 -2.2819396009709907e-05
GC_8_201 b_8 NI_8 NS_201 0 -9.4772238826387814e-03
GC_8_202 b_8 NI_8 NS_202 0 5.7440921416854261e-04
GC_8_203 b_8 NI_8 NS_203 0 -1.1239263406409420e-04
GC_8_204 b_8 NI_8 NS_204 0 -1.6637232888435023e-04
GC_8_205 b_8 NI_8 NS_205 0 2.5983750767696930e-03
GC_8_206 b_8 NI_8 NS_206 0 1.4392307009514183e-03
GC_8_207 b_8 NI_8 NS_207 0 2.8563323868143792e-03
GC_8_208 b_8 NI_8 NS_208 0 -2.4036037360849393e-03
GC_8_209 b_8 NI_8 NS_209 0 5.7602435479317581e-04
GC_8_210 b_8 NI_8 NS_210 0 3.3119793354134675e-04
GC_8_211 b_8 NI_8 NS_211 0 -9.6470845240197665e-07
GC_8_212 b_8 NI_8 NS_212 0 -9.6680916382231768e-07
GC_8_213 b_8 NI_8 NS_213 0 -1.5589765477559549e-05
GC_8_214 b_8 NI_8 NS_214 0 -1.2977505443485080e-05
GC_8_215 b_8 NI_8 NS_215 0 -7.9312499640541101e-05
GC_8_216 b_8 NI_8 NS_216 0 1.0143600172926782e-04
GC_8_217 b_8 NI_8 NS_217 0 -2.4181462017808656e-05
GC_8_218 b_8 NI_8 NS_218 0 -1.9458132785035099e-05
GC_8_219 b_8 NI_8 NS_219 0 -1.7406629508539774e-05
GC_8_220 b_8 NI_8 NS_220 0 -7.7274045355829043e-06
GC_8_221 b_8 NI_8 NS_221 0 1.8336965072920494e-04
GC_8_222 b_8 NI_8 NS_222 0 -8.5640317900223737e-05
GC_8_223 b_8 NI_8 NS_223 0 -3.0286086554602256e-04
GC_8_224 b_8 NI_8 NS_224 0 4.9418538354988681e-05
GC_8_225 b_8 NI_8 NS_225 0 5.8838610799363013e-02
GC_8_226 b_8 NI_8 NS_226 0 -8.1662674122995630e-04
GC_8_227 b_8 NI_8 NS_227 0 -1.7986335138466018e-03
GC_8_228 b_8 NI_8 NS_228 0 2.2781721099493940e-03
GC_8_229 b_8 NI_8 NS_229 0 2.8558879260476865e-03
GC_8_230 b_8 NI_8 NS_230 0 2.8094880422853690e-04
GC_8_231 b_8 NI_8 NS_231 0 -5.2690031174306142e-03
GC_8_232 b_8 NI_8 NS_232 0 6.4726576748248528e-04
GC_8_233 b_8 NI_8 NS_233 0 -6.1537719448878560e-03
GC_8_234 b_8 NI_8 NS_234 0 1.0731209688448437e-02
GC_8_235 b_8 NI_8 NS_235 0 -7.4197931662514215e-04
GC_8_236 b_8 NI_8 NS_236 0 -5.4346936212871242e-04
GC_8_237 b_8 NI_8 NS_237 0 1.5109443785001611e-03
GC_8_238 b_8 NI_8 NS_238 0 -3.9740441007787659e-03
GC_8_239 b_8 NI_8 NS_239 0 8.5127714743056645e-04
GC_8_240 b_8 NI_8 NS_240 0 1.2312434319917721e-03
GC_8_241 b_8 NI_8 NS_241 0 -1.5871471212427642e-04
GC_8_242 b_8 NI_8 NS_242 0 1.0935051819098976e-03
GC_8_243 b_8 NI_8 NS_243 0 -5.6242380321875557e-03
GC_8_244 b_8 NI_8 NS_244 0 9.6414810205618128e-04
GC_8_245 b_8 NI_8 NS_245 0 -1.0923918850320045e-04
GC_8_246 b_8 NI_8 NS_246 0 -7.3884098569136237e-05
GC_8_247 b_8 NI_8 NS_247 0 4.2412489850930413e-04
GC_8_248 b_8 NI_8 NS_248 0 5.3175006912689416e-03
GC_8_249 b_8 NI_8 NS_249 0 -3.6122808488746186e-04
GC_8_250 b_8 NI_8 NS_250 0 -1.6429755977192181e-04
GC_8_251 b_8 NI_8 NS_251 0 -4.3820101474770874e-04
GC_8_252 b_8 NI_8 NS_252 0 2.3869634296652852e-05
GC_8_253 b_8 NI_8 NS_253 0 -3.8853000698057318e-04
GC_8_254 b_8 NI_8 NS_254 0 3.6937540517236698e-04
GC_8_255 b_8 NI_8 NS_255 0 -2.0278482547925032e-04
GC_8_256 b_8 NI_8 NS_256 0 -3.0057326435664270e-05
GC_8_257 b_8 NI_8 NS_257 0 -7.2113834808388132e-03
GC_8_258 b_8 NI_8 NS_258 0 -1.0833815285557118e-03
GC_8_259 b_8 NI_8 NS_259 0 -1.0528095964133737e-06
GC_8_260 b_8 NI_8 NS_260 0 1.4310261403075042e-05
GC_8_261 b_8 NI_8 NS_261 0 -1.4062030232278060e-04
GC_8_262 b_8 NI_8 NS_262 0 8.0115417022692532e-04
GC_8_263 b_8 NI_8 NS_263 0 -1.0811712832026704e-03
GC_8_264 b_8 NI_8 NS_264 0 -2.8405401409544433e-03
GC_8_265 b_8 NI_8 NS_265 0 9.3874344258759509e-05
GC_8_266 b_8 NI_8 NS_266 0 2.1385118282095806e-04
GC_8_267 b_8 NI_8 NS_267 0 2.5547663097286497e-06
GC_8_268 b_8 NI_8 NS_268 0 -2.2362643834537344e-08
GC_8_269 b_8 NI_8 NS_269 0 -3.1766791373595134e-06
GC_8_270 b_8 NI_8 NS_270 0 -7.5027545805439302e-06
GC_8_271 b_8 NI_8 NS_271 0 -5.0754389283158208e-05
GC_8_272 b_8 NI_8 NS_272 0 7.5517330247385091e-05
GC_8_273 b_8 NI_8 NS_273 0 -2.5399134499214016e-06
GC_8_274 b_8 NI_8 NS_274 0 -1.1442734859423478e-05
GC_8_275 b_8 NI_8 NS_275 0 -2.9960486804561185e-06
GC_8_276 b_8 NI_8 NS_276 0 3.2800228740388069e-06
GC_8_277 b_8 NI_8 NS_277 0 2.2093981749824921e-06
GC_8_278 b_8 NI_8 NS_278 0 3.0645253089288681e-06
GC_8_279 b_8 NI_8 NS_279 0 4.6849575739329720e-07
GC_8_280 b_8 NI_8 NS_280 0 -8.2754733378780529e-06
GC_8_281 b_8 NI_8 NS_281 0 -1.5074112611669558e-02
GC_8_282 b_8 NI_8 NS_282 0 -1.3247136509707228e-03
GC_8_283 b_8 NI_8 NS_283 0 -8.4916649294427226e-04
GC_8_284 b_8 NI_8 NS_284 0 -1.0111910962236302e-03
GC_8_285 b_8 NI_8 NS_285 0 -1.1790192022934686e-03
GC_8_286 b_8 NI_8 NS_286 0 1.3800284987720661e-03
GC_8_287 b_8 NI_8 NS_287 0 8.5020681007478064e-04
GC_8_288 b_8 NI_8 NS_288 0 -7.4005573565397197e-04
GC_8_289 b_8 NI_8 NS_289 0 -3.1906880525988763e-03
GC_8_290 b_8 NI_8 NS_290 0 -8.5706095281360885e-03
GC_8_291 b_8 NI_8 NS_291 0 3.1831922393934501e-05
GC_8_292 b_8 NI_8 NS_292 0 1.8335857851359554e-04
GC_8_293 b_8 NI_8 NS_293 0 1.9449516362421960e-03
GC_8_294 b_8 NI_8 NS_294 0 -2.3077120784836900e-03
GC_8_295 b_8 NI_8 NS_295 0 7.4376387219276022e-04
GC_8_296 b_8 NI_8 NS_296 0 1.7762228561363260e-04
GC_8_297 b_8 NI_8 NS_297 0 9.5984305028980936e-04
GC_8_298 b_8 NI_8 NS_298 0 -1.9577709839487959e-03
GC_8_299 b_8 NI_8 NS_299 0 1.2352236853773930e-03
GC_8_300 b_8 NI_8 NS_300 0 -2.2346515268508245e-03
GC_8_301 b_8 NI_8 NS_301 0 3.7411300779965067e-05
GC_8_302 b_8 NI_8 NS_302 0 7.0984910278038644e-06
GC_8_303 b_8 NI_8 NS_303 0 7.4412934126043924e-03
GC_8_304 b_8 NI_8 NS_304 0 1.1498965242875720e-03
GC_8_305 b_8 NI_8 NS_305 0 -1.1913406468282949e-04
GC_8_306 b_8 NI_8 NS_306 0 3.1478848249002566e-05
GC_8_307 b_8 NI_8 NS_307 0 -1.3213190232674158e-04
GC_8_308 b_8 NI_8 NS_308 0 1.2295628807032253e-04
GC_8_309 b_8 NI_8 NS_309 0 1.9358902555497321e-04
GC_8_310 b_8 NI_8 NS_310 0 -3.5776762458390688e-04
GC_8_311 b_8 NI_8 NS_311 0 3.4607944821240708e-04
GC_8_312 b_8 NI_8 NS_312 0 -1.0717382421487860e-04
GC_8_313 b_8 NI_8 NS_313 0 -7.7708114292799049e-03
GC_8_314 b_8 NI_8 NS_314 0 3.0732171071030322e-03
GC_8_315 b_8 NI_8 NS_315 0 -2.1447016470917170e-04
GC_8_316 b_8 NI_8 NS_316 0 -1.6643308406983119e-04
GC_8_317 b_8 NI_8 NS_317 0 3.8500278684389048e-03
GC_8_318 b_8 NI_8 NS_318 0 5.0804070178527103e-04
GC_8_319 b_8 NI_8 NS_319 0 2.3161102807582241e-03
GC_8_320 b_8 NI_8 NS_320 0 -1.0753088856217360e-03
GC_8_321 b_8 NI_8 NS_321 0 7.6279979155473700e-04
GC_8_322 b_8 NI_8 NS_322 0 3.3799073269609312e-04
GC_8_323 b_8 NI_8 NS_323 0 -2.6770843380295609e-06
GC_8_324 b_8 NI_8 NS_324 0 -4.3129783381894432e-06
GC_8_325 b_8 NI_8 NS_325 0 -2.0059599544944133e-05
GC_8_326 b_8 NI_8 NS_326 0 -5.6038610948449140e-06
GC_8_327 b_8 NI_8 NS_327 0 -3.3886610269498490e-05
GC_8_328 b_8 NI_8 NS_328 0 -6.9192244312633720e-05
GC_8_329 b_8 NI_8 NS_329 0 -2.7013065716516596e-05
GC_8_330 b_8 NI_8 NS_330 0 1.6625666886538100e-06
GC_8_331 b_8 NI_8 NS_331 0 -1.4439314177683642e-05
GC_8_332 b_8 NI_8 NS_332 0 -8.9562218876626341e-06
GC_8_333 b_8 NI_8 NS_333 0 2.3636326284915934e-04
GC_8_334 b_8 NI_8 NS_334 0 -1.3182694890305445e-04
GC_8_335 b_8 NI_8 NS_335 0 -3.9255774461583213e-04
GC_8_336 b_8 NI_8 NS_336 0 9.5573920238650487e-05
GC_8_337 b_8 NI_8 NS_337 0 -1.3219958273245893e-02
GC_8_338 b_8 NI_8 NS_338 0 1.2044449083902896e-02
GC_8_339 b_8 NI_8 NS_339 0 -2.2023344575709688e-03
GC_8_340 b_8 NI_8 NS_340 0 1.4394743987854676e-03
GC_8_341 b_8 NI_8 NS_341 0 -2.4020460292130644e-03
GC_8_342 b_8 NI_8 NS_342 0 4.3204556206903177e-03
GC_8_343 b_8 NI_8 NS_343 0 -9.8944804927660946e-04
GC_8_344 b_8 NI_8 NS_344 0 -2.9570758796032283e-03
GC_8_345 b_8 NI_8 NS_345 0 -1.1571807928307381e-02
GC_8_346 b_8 NI_8 NS_346 0 -3.3375374356228154e-03
GC_8_347 b_8 NI_8 NS_347 0 3.3294280737056827e-04
GC_8_348 b_8 NI_8 NS_348 0 -3.8181711718655111e-04
GC_8_349 b_8 NI_8 NS_349 0 3.0706477843235589e-03
GC_8_350 b_8 NI_8 NS_350 0 2.7298466753063731e-04
GC_8_351 b_8 NI_8 NS_351 0 9.7712036860207849e-04
GC_8_352 b_8 NI_8 NS_352 0 6.3661363947170092e-04
GC_8_353 b_8 NI_8 NS_353 0 4.2160893262332636e-03
GC_8_354 b_8 NI_8 NS_354 0 -6.9945736704739986e-04
GC_8_355 b_8 NI_8 NS_355 0 -1.0010219503938298e-03
GC_8_356 b_8 NI_8 NS_356 0 5.8035147746360956e-04
GC_8_357 b_8 NI_8 NS_357 0 -1.4614069636611072e-04
GC_8_358 b_8 NI_8 NS_358 0 -4.2750998104355915e-05
GC_8_359 b_8 NI_8 NS_359 0 4.1349476973905359e-03
GC_8_360 b_8 NI_8 NS_360 0 -3.9764447797403568e-04
GC_8_361 b_8 NI_8 NS_361 0 -4.7548246833235781e-04
GC_8_362 b_8 NI_8 NS_362 0 -1.4229995897022051e-04
GC_8_363 b_8 NI_8 NS_363 0 -2.8838813921661175e-04
GC_8_364 b_8 NI_8 NS_364 0 3.6416699211002572e-05
GC_8_365 b_8 NI_8 NS_365 0 -3.0280954547585667e-04
GC_8_366 b_8 NI_8 NS_366 0 1.4279920494428706e-04
GC_8_367 b_8 NI_8 NS_367 0 -1.2864878741505642e-04
GC_8_368 b_8 NI_8 NS_368 0 -6.9474722913941294e-05
GC_8_369 b_8 NI_8 NS_369 0 -2.0656948235928218e-03
GC_8_370 b_8 NI_8 NS_370 0 1.0998431089140485e-04
GC_8_371 b_8 NI_8 NS_371 0 -1.2583815430886603e-05
GC_8_372 b_8 NI_8 NS_372 0 4.3597938609623973e-05
GC_8_373 b_8 NI_8 NS_373 0 -3.1386874931739142e-04
GC_8_374 b_8 NI_8 NS_374 0 4.5855053120460093e-06
GC_8_375 b_8 NI_8 NS_375 0 1.7956689939236424e-03
GC_8_376 b_8 NI_8 NS_376 0 -1.6189845445503631e-03
GC_8_377 b_8 NI_8 NS_377 0 1.6420192561303901e-04
GC_8_378 b_8 NI_8 NS_378 0 -1.0933660562340007e-04
GC_8_379 b_8 NI_8 NS_379 0 -9.1430453361256163e-07
GC_8_380 b_8 NI_8 NS_380 0 5.7008151200426080e-07
GC_8_381 b_8 NI_8 NS_381 0 -3.3604341693534599e-06
GC_8_382 b_8 NI_8 NS_382 0 -8.5252954626387088e-06
GC_8_383 b_8 NI_8 NS_383 0 -1.3595339613429869e-04
GC_8_384 b_8 NI_8 NS_384 0 1.3045759120769597e-04
GC_8_385 b_8 NI_8 NS_385 0 -2.8519312402597430e-07
GC_8_386 b_8 NI_8 NS_386 0 -2.0711806879561618e-05
GC_8_387 b_8 NI_8 NS_387 0 -4.5062864523150233e-06
GC_8_388 b_8 NI_8 NS_388 0 -4.1284726552468033e-06
GC_8_389 b_8 NI_8 NS_389 0 4.7744941253586041e-05
GC_8_390 b_8 NI_8 NS_390 0 -1.4665627501880328e-05
GC_8_391 b_8 NI_8 NS_391 0 -7.3836531193694570e-05
GC_8_392 b_8 NI_8 NS_392 0 3.5158644668853118e-07
GC_8_393 b_8 NI_8 NS_393 0 -8.9831662039037280e-02
GC_8_394 b_8 NI_8 NS_394 0 8.1182576345562724e-03
GC_8_395 b_8 NI_8 NS_395 0 -1.6302047095767650e-04
GC_8_396 b_8 NI_8 NS_396 0 -1.2312486582295292e-03
GC_8_397 b_8 NI_8 NS_397 0 -1.1820419976382942e-03
GC_8_398 b_8 NI_8 NS_398 0 -1.4322565865959550e-03
GC_8_399 b_8 NI_8 NS_399 0 1.7020210857515861e-03
GC_8_400 b_8 NI_8 NS_400 0 2.6344280177284410e-03
GC_8_401 b_8 NI_8 NS_401 0 8.9198451063080067e-03
GC_8_402 b_8 NI_8 NS_402 0 2.6151858326569946e-05
GC_8_403 b_8 NI_8 NS_403 0 4.0839437176639736e-04
GC_8_404 b_8 NI_8 NS_404 0 -5.1067903011279886e-04
GC_8_405 b_8 NI_8 NS_405 0 -9.1398532921717443e-04
GC_8_406 b_8 NI_8 NS_406 0 -2.4837353908558949e-03
GC_8_407 b_8 NI_8 NS_407 0 5.0902955113272532e-04
GC_8_408 b_8 NI_8 NS_408 0 1.6853201321361428e-04
GC_8_409 b_8 NI_8 NS_409 0 1.9367213188890598e-04
GC_8_410 b_8 NI_8 NS_410 0 -1.5543542481506463e-03
GC_8_411 b_8 NI_8 NS_411 0 1.1059204987755751e-03
GC_8_412 b_8 NI_8 NS_412 0 -1.7748306112879792e-03
GC_8_413 b_8 NI_8 NS_413 0 3.2922375116739687e-05
GC_8_414 b_8 NI_8 NS_414 0 -7.0299199333421975e-06
GC_8_415 b_8 NI_8 NS_415 0 3.5597358386459869e-03
GC_8_416 b_8 NI_8 NS_416 0 1.2747699215571312e-03
GC_8_417 b_8 NI_8 NS_417 0 -5.3974662882680925e-05
GC_8_418 b_8 NI_8 NS_418 0 -1.8920482526242861e-05
GC_8_419 b_8 NI_8 NS_419 0 -1.4196466364502222e-04
GC_8_420 b_8 NI_8 NS_420 0 1.0940145121616458e-04
GC_8_421 b_8 NI_8 NS_421 0 1.6324790100073834e-04
GC_8_422 b_8 NI_8 NS_422 0 -2.0264263830581053e-04
GC_8_423 b_8 NI_8 NS_423 0 2.1656152418501266e-04
GC_8_424 b_8 NI_8 NS_424 0 -1.7379037273173213e-05
GC_8_425 b_8 NI_8 NS_425 0 -4.9616176283164646e-03
GC_8_426 b_8 NI_8 NS_426 0 2.3813642763591573e-03
GC_8_427 b_8 NI_8 NS_427 0 -1.2869769443119456e-04
GC_8_428 b_8 NI_8 NS_428 0 -1.0590539895066958e-04
GC_8_429 b_8 NI_8 NS_429 0 2.4510447348120219e-03
GC_8_430 b_8 NI_8 NS_430 0 5.2897555801877875e-04
GC_8_431 b_8 NI_8 NS_431 0 1.4384377500757967e-03
GC_8_432 b_8 NI_8 NS_432 0 -4.9026164698968847e-04
GC_8_433 b_8 NI_8 NS_433 0 4.6980769477506385e-04
GC_8_434 b_8 NI_8 NS_434 0 5.8544353493171875e-05
GC_8_435 b_8 NI_8 NS_435 0 -3.9956618809661566e-07
GC_8_436 b_8 NI_8 NS_436 0 -1.8447855246339831e-06
GC_8_437 b_8 NI_8 NS_437 0 -7.2809999897697955e-06
GC_8_438 b_8 NI_8 NS_438 0 2.0657345225447104e-06
GC_8_439 b_8 NI_8 NS_439 0 -5.6723196978261363e-06
GC_8_440 b_8 NI_8 NS_440 0 -1.4548575033896866e-04
GC_8_441 b_8 NI_8 NS_441 0 -1.0952659485793752e-05
GC_8_442 b_8 NI_8 NS_442 0 9.6733234625462481e-06
GC_8_443 b_8 NI_8 NS_443 0 -6.5463127281775253e-06
GC_8_444 b_8 NI_8 NS_444 0 5.8580225782437329e-06
GC_8_445 b_8 NI_8 NS_445 0 1.0916903903397294e-04
GC_8_446 b_8 NI_8 NS_446 0 -4.1670552841557912e-05
GC_8_447 b_8 NI_8 NS_447 0 -1.7207234302517606e-04
GC_8_448 b_8 NI_8 NS_448 0 2.7289506334373191e-05
GC_8_449 b_8 NI_8 NS_449 0 6.5575966872793495e-03
GC_8_450 b_8 NI_8 NS_450 0 -8.5830992450166248e-05
GC_8_451 b_8 NI_8 NS_451 0 -1.9560044582087296e-04
GC_8_452 b_8 NI_8 NS_452 0 7.0113140806893912e-04
GC_8_453 b_8 NI_8 NS_453 0 -3.0825255711977513e-04
GC_8_454 b_8 NI_8 NS_454 0 -6.8120270407258940e-04
GC_8_455 b_8 NI_8 NS_455 0 -5.3653208588292853e-04
GC_8_456 b_8 NI_8 NS_456 0 -8.2810383287276203e-04
GC_8_457 b_8 NI_8 NS_457 0 2.2767881748169253e-03
GC_8_458 b_8 NI_8 NS_458 0 7.1800469727908013e-04
GC_8_459 b_8 NI_8 NS_459 0 -1.3373192929670342e-04
GC_8_460 b_8 NI_8 NS_460 0 9.7607751780677359e-05
GC_8_461 b_8 NI_8 NS_461 0 4.3128990319371492e-04
GC_8_462 b_8 NI_8 NS_462 0 -4.5673399573489500e-04
GC_8_463 b_8 NI_8 NS_463 0 8.6764235192738389e-04
GC_8_464 b_8 NI_8 NS_464 0 -1.0956052484965504e-04
GC_8_465 b_8 NI_8 NS_465 0 6.2746489213366056e-04
GC_8_466 b_8 NI_8 NS_466 0 1.9121310627720539e-03
GC_8_467 b_8 NI_8 NS_467 0 -1.2033475633369149e-03
GC_8_468 b_8 NI_8 NS_468 0 2.5524455117089707e-03
GC_8_469 b_8 NI_8 NS_469 0 -2.0076716642376333e-04
GC_8_470 b_8 NI_8 NS_470 0 -5.8802109304380533e-05
GC_8_471 b_8 NI_8 NS_471 0 -1.0135002201420214e-03
GC_8_472 b_8 NI_8 NS_472 0 1.3388406714337096e-03
GC_8_473 b_8 NI_8 NS_473 0 5.9371646448839064e-05
GC_8_474 b_8 NI_8 NS_474 0 -2.0587236093817637e-05
GC_8_475 b_8 NI_8 NS_475 0 -6.7535725235467884e-04
GC_8_476 b_8 NI_8 NS_476 0 9.0745627408502931e-05
GC_8_477 b_8 NI_8 NS_477 0 -3.9092414423361611e-04
GC_8_478 b_8 NI_8 NS_478 0 5.0439706941557888e-05
GC_8_479 b_8 NI_8 NS_479 0 -1.0766422471414869e-04
GC_8_480 b_8 NI_8 NS_480 0 -3.4998175636262423e-05
GC_8_481 b_8 NI_8 NS_481 0 -4.0384742239682730e-04
GC_8_482 b_8 NI_8 NS_482 0 -3.3770410101010657e-03
GC_8_483 b_8 NI_8 NS_483 0 3.7921578629109889e-05
GC_8_484 b_8 NI_8 NS_484 0 -1.9107425996638272e-05
GC_8_485 b_8 NI_8 NS_485 0 -8.7697648881110131e-04
GC_8_486 b_8 NI_8 NS_486 0 4.9605543421912010e-04
GC_8_487 b_8 NI_8 NS_487 0 1.2288554237786663e-03
GC_8_488 b_8 NI_8 NS_488 0 2.8811119889896020e-04
GC_8_489 b_8 NI_8 NS_489 0 -1.5361158018475986e-04
GC_8_490 b_8 NI_8 NS_490 0 2.9714120241646001e-04
GC_8_491 b_8 NI_8 NS_491 0 -1.0363969700615352e-06
GC_8_492 b_8 NI_8 NS_492 0 1.0092114316843305e-06
GC_8_493 b_8 NI_8 NS_493 0 -1.3461347410100946e-06
GC_8_494 b_8 NI_8 NS_494 0 -7.7025207375511750e-06
GC_8_495 b_8 NI_8 NS_495 0 -3.2445933987941964e-05
GC_8_496 b_8 NI_8 NS_496 0 7.4271488501924398e-05
GC_8_497 b_8 NI_8 NS_497 0 -2.2469475903780322e-06
GC_8_498 b_8 NI_8 NS_498 0 -1.3260175990159059e-05
GC_8_499 b_8 NI_8 NS_499 0 -9.0686502764242929e-06
GC_8_500 b_8 NI_8 NS_500 0 -5.2684078249294194e-06
GC_8_501 b_8 NI_8 NS_501 0 2.7479714462166694e-05
GC_8_502 b_8 NI_8 NS_502 0 -1.8543638352156872e-05
GC_8_503 b_8 NI_8 NS_503 0 -5.0924396634151740e-05
GC_8_504 b_8 NI_8 NS_504 0 1.4311934486344560e-05
GC_8_505 b_8 NI_8 NS_505 0 -3.3963333878717977e-03
GC_8_506 b_8 NI_8 NS_506 0 -1.3409448314773996e-04
GC_8_507 b_8 NI_8 NS_507 0 -3.0684957325257051e-04
GC_8_508 b_8 NI_8 NS_508 0 -2.2206889072041869e-04
GC_8_509 b_8 NI_8 NS_509 0 3.3254355225319655e-04
GC_8_510 b_8 NI_8 NS_510 0 8.2569294914034940e-05
GC_8_511 b_8 NI_8 NS_511 0 6.5238648451365362e-04
GC_8_512 b_8 NI_8 NS_512 0 2.7949118117238215e-04
GC_8_513 b_8 NI_8 NS_513 0 -2.3645459689356470e-03
GC_8_514 b_8 NI_8 NS_514 0 7.6659522928249231e-04
GC_8_515 b_8 NI_8 NS_515 0 2.3459978023479490e-04
GC_8_516 b_8 NI_8 NS_516 0 1.5568595333369299e-04
GC_8_517 b_8 NI_8 NS_517 0 -4.6490198111633107e-04
GC_8_518 b_8 NI_8 NS_518 0 -1.4673840308627041e-03
GC_8_519 b_8 NI_8 NS_519 0 3.4673195161808536e-04
GC_8_520 b_8 NI_8 NS_520 0 -2.4201800443309453e-04
GC_8_521 b_8 NI_8 NS_521 0 -8.6843612685098153e-04
GC_8_522 b_8 NI_8 NS_522 0 7.1309991645854189e-04
GC_8_523 b_8 NI_8 NS_523 0 -1.0605230007730776e-03
GC_8_524 b_8 NI_8 NS_524 0 -1.3650763921787719e-03
GC_8_525 b_8 NI_8 NS_525 0 1.1836651280649094e-04
GC_8_526 b_8 NI_8 NS_526 0 5.2362338727428835e-05
GC_8_527 b_8 NI_8 NS_527 0 2.0728416496434599e-03
GC_8_528 b_8 NI_8 NS_528 0 -3.7917014302665925e-03
GC_8_529 b_8 NI_8 NS_529 0 -3.1234729205297564e-04
GC_8_530 b_8 NI_8 NS_530 0 3.6359294260357385e-04
GC_8_531 b_8 NI_8 NS_531 0 -2.6722982926298241e-04
GC_8_532 b_8 NI_8 NS_532 0 2.7061718008933484e-04
GC_8_533 b_8 NI_8 NS_533 0 -5.8007784594822064e-05
GC_8_534 b_8 NI_8 NS_534 0 -5.2675396282647103e-04
GC_8_535 b_8 NI_8 NS_535 0 1.9021966028286296e-04
GC_8_536 b_8 NI_8 NS_536 0 -6.0137246334175128e-05
GC_8_537 b_8 NI_8 NS_537 0 1.2205496797727652e-03
GC_8_538 b_8 NI_8 NS_538 0 1.6796172339909178e-03
GC_8_539 b_8 NI_8 NS_539 0 -1.0133682474315056e-04
GC_8_540 b_8 NI_8 NS_540 0 1.0806259809562085e-04
GC_8_541 b_8 NI_8 NS_541 0 1.2612841702435232e-03
GC_8_542 b_8 NI_8 NS_542 0 -6.3848484973783092e-04
GC_8_543 b_8 NI_8 NS_543 0 1.0559170600090376e-04
GC_8_544 b_8 NI_8 NS_544 0 3.4003695713278801e-04
GC_8_545 b_8 NI_8 NS_545 0 -5.0106875083968114e-04
GC_8_546 b_8 NI_8 NS_546 0 3.8825309279335533e-04
GC_8_547 b_8 NI_8 NS_547 0 6.5613236486776359e-07
GC_8_548 b_8 NI_8 NS_548 0 -4.6184345407637282e-06
GC_8_549 b_8 NI_8 NS_549 0 -1.1951247215611575e-07
GC_8_550 b_8 NI_8 NS_550 0 3.3216378748150168e-05
GC_8_551 b_8 NI_8 NS_551 0 2.6899497867666725e-05
GC_8_552 b_8 NI_8 NS_552 0 -1.6963389710647351e-04
GC_8_553 b_8 NI_8 NS_553 0 4.5553460775706770e-05
GC_8_554 b_8 NI_8 NS_554 0 4.8639987449224296e-05
GC_8_555 b_8 NI_8 NS_555 0 4.6997769517136263e-06
GC_8_556 b_8 NI_8 NS_556 0 1.7341739637796108e-05
GC_8_557 b_8 NI_8 NS_557 0 2.3750597745190712e-04
GC_8_558 b_8 NI_8 NS_558 0 -1.0737598510310003e-04
GC_8_559 b_8 NI_8 NS_559 0 -3.7730814788135346e-04
GC_8_560 b_8 NI_8 NS_560 0 5.7521953639564811e-05
GC_8_561 b_8 NI_8 NS_561 0 2.6509271169464815e-02
GC_8_562 b_8 NI_8 NS_562 0 -2.8560267373162136e-04
GC_8_563 b_8 NI_8 NS_563 0 -4.6672448184517429e-04
GC_8_564 b_8 NI_8 NS_564 0 5.6166547167501918e-04
GC_8_565 b_8 NI_8 NS_565 0 1.0830866259422826e-03
GC_8_566 b_8 NI_8 NS_566 0 2.4769511767044682e-04
GC_8_567 b_8 NI_8 NS_567 0 -1.1485844227287010e-03
GC_8_568 b_8 NI_8 NS_568 0 9.4539014346843662e-04
GC_8_569 b_8 NI_8 NS_569 0 -2.8069487227108795e-03
GC_8_570 b_8 NI_8 NS_570 0 4.5021822344547963e-03
GC_8_571 b_8 NI_8 NS_571 0 -2.3787033187878964e-04
GC_8_572 b_8 NI_8 NS_572 0 1.4291726896386304e-04
GC_8_573 b_8 NI_8 NS_573 0 4.7113619346268534e-05
GC_8_574 b_8 NI_8 NS_574 0 -1.2076189545108572e-03
GC_8_575 b_8 NI_8 NS_575 0 7.7334494509442679e-04
GC_8_576 b_8 NI_8 NS_576 0 1.3893067117181002e-04
GC_8_577 b_8 NI_8 NS_577 0 -4.8497811809194297e-04
GC_8_578 b_8 NI_8 NS_578 0 7.4306481863431657e-04
GC_8_579 b_8 NI_8 NS_579 0 -1.6970850942715145e-03
GC_8_580 b_8 NI_8 NS_580 0 9.7327851358419086e-04
GC_8_581 b_8 NI_8 NS_581 0 -1.2707743894692879e-04
GC_8_582 b_8 NI_8 NS_582 0 -9.1179174914762947e-05
GC_8_583 b_8 NI_8 NS_583 0 3.3113896436750317e-05
GC_8_584 b_8 NI_8 NS_584 0 2.2189855260750166e-03
GC_8_585 b_8 NI_8 NS_585 0 6.4554428098657210e-05
GC_8_586 b_8 NI_8 NS_586 0 -1.8152559370240748e-04
GC_8_587 b_8 NI_8 NS_587 0 -5.0940186686729044e-04
GC_8_588 b_8 NI_8 NS_588 0 1.5196497028021952e-04
GC_8_589 b_8 NI_8 NS_589 0 -3.0484838175635643e-04
GC_8_590 b_8 NI_8 NS_590 0 1.2518113152991552e-04
GC_8_591 b_8 NI_8 NS_591 0 -9.8987499009759030e-05
GC_8_592 b_8 NI_8 NS_592 0 -1.5066502203259927e-05
GC_8_593 b_8 NI_8 NS_593 0 -1.1915552964821496e-03
GC_8_594 b_8 NI_8 NS_594 0 3.3027167186815750e-04
GC_8_595 b_8 NI_8 NS_595 0 3.0081174530165801e-05
GC_8_596 b_8 NI_8 NS_596 0 -2.1064678215533579e-05
GC_8_597 b_8 NI_8 NS_597 0 -5.1575977597390597e-04
GC_8_598 b_8 NI_8 NS_598 0 5.2073917480604474e-04
GC_8_599 b_8 NI_8 NS_599 0 -1.5817023723736165e-03
GC_8_600 b_8 NI_8 NS_600 0 -1.8552751220749818e-03
GC_8_601 b_8 NI_8 NS_601 0 -1.9381343302395519e-04
GC_8_602 b_8 NI_8 NS_602 0 -6.2506513491215898e-05
GC_8_603 b_8 NI_8 NS_603 0 -3.5796024728632278e-09
GC_8_604 b_8 NI_8 NS_604 0 1.2054900528434939e-06
GC_8_605 b_8 NI_8 NS_605 0 -6.1440954896463143e-06
GC_8_606 b_8 NI_8 NS_606 0 -3.8983646880151463e-06
GC_8_607 b_8 NI_8 NS_607 0 6.7383185378896263e-05
GC_8_608 b_8 NI_8 NS_608 0 1.3609504520200328e-04
GC_8_609 b_8 NI_8 NS_609 0 -9.1000076740467679e-06
GC_8_610 b_8 NI_8 NS_610 0 -1.1808584822006427e-05
GC_8_611 b_8 NI_8 NS_611 0 -4.6496437462680050e-06
GC_8_612 b_8 NI_8 NS_612 0 4.1895675167047390e-06
GC_8_613 b_8 NI_8 NS_613 0 8.5648152681988957e-06
GC_8_614 b_8 NI_8 NS_614 0 -4.9521760414303914e-05
GC_8_615 b_8 NI_8 NS_615 0 -3.2055345758357767e-05
GC_8_616 b_8 NI_8 NS_616 0 7.2202900640065860e-05
GC_8_617 b_8 NI_8 NS_617 0 -9.1923781034170520e-03
GC_8_618 b_8 NI_8 NS_618 0 -3.8938211451324477e-04
GC_8_619 b_8 NI_8 NS_619 0 -2.0088073306993973e-04
GC_8_620 b_8 NI_8 NS_620 0 -2.5626596970543730e-04
GC_8_621 b_8 NI_8 NS_621 0 -4.5221635030302755e-04
GC_8_622 b_8 NI_8 NS_622 0 4.5388850062803669e-04
GC_8_623 b_8 NI_8 NS_623 0 -2.6344463725557529e-04
GC_8_624 b_8 NI_8 NS_624 0 -2.7046631190547592e-04
GC_8_625 b_8 NI_8 NS_625 0 -8.1399467283976249e-04
GC_8_626 b_8 NI_8 NS_626 0 -3.4082571711312694e-03
GC_8_627 b_8 NI_8 NS_627 0 1.6788045223697700e-04
GC_8_628 b_8 NI_8 NS_628 0 1.7526250150448126e-04
GC_8_629 b_8 NI_8 NS_629 0 3.2045654769394119e-04
GC_8_630 b_8 NI_8 NS_630 0 -5.4830393196626890e-04
GC_8_631 b_8 NI_8 NS_631 0 3.3513751138635525e-04
GC_8_632 b_8 NI_8 NS_632 0 -1.7527674756684719e-04
GC_8_633 b_8 NI_8 NS_633 0 -7.2668002061238262e-04
GC_8_634 b_8 NI_8 NS_634 0 -3.5729647473673289e-04
GC_8_635 b_8 NI_8 NS_635 0 -5.4064369337252166e-04
GC_8_636 b_8 NI_8 NS_636 0 -1.6464202148030263e-03
GC_8_637 b_8 NI_8 NS_637 0 3.9572703324286465e-05
GC_8_638 b_8 NI_8 NS_638 0 3.0058013462048214e-05
GC_8_639 b_8 NI_8 NS_639 0 3.8188818093275955e-03
GC_8_640 b_8 NI_8 NS_640 0 -2.4089955777632367e-03
GC_8_641 b_8 NI_8 NS_641 0 -3.0411111979548368e-04
GC_8_642 b_8 NI_8 NS_642 0 1.0299526214439775e-04
GC_8_643 b_8 NI_8 NS_643 0 -1.2627382383429886e-04
GC_8_644 b_8 NI_8 NS_644 0 1.9055209170985838e-04
GC_8_645 b_8 NI_8 NS_645 0 6.8673979440144302e-05
GC_8_646 b_8 NI_8 NS_646 0 -3.5983483095626832e-04
GC_8_647 b_8 NI_8 NS_647 0 1.5424281531754296e-04
GC_8_648 b_8 NI_8 NS_648 0 -3.1182372873486882e-05
GC_8_649 b_8 NI_8 NS_649 0 1.2365757055137600e-03
GC_8_650 b_8 NI_8 NS_650 0 2.0564199013048999e-03
GC_8_651 b_8 NI_8 NS_651 0 -1.0111765128609580e-04
GC_8_652 b_8 NI_8 NS_652 0 4.2923810169033012e-05
GC_8_653 b_8 NI_8 NS_653 0 1.1568680958842616e-03
GC_8_654 b_8 NI_8 NS_654 0 -5.7811228241794221e-04
GC_8_655 b_8 NI_8 NS_655 0 -5.1286801854374447e-05
GC_8_656 b_8 NI_8 NS_656 0 9.0047981688393987e-04
GC_8_657 b_8 NI_8 NS_657 0 -3.6517973885834629e-04
GC_8_658 b_8 NI_8 NS_658 0 -2.3174511402499231e-05
GC_8_659 b_8 NI_8 NS_659 0 1.3099471393420952e-06
GC_8_660 b_8 NI_8 NS_660 0 -2.6250987448442553e-06
GC_8_661 b_8 NI_8 NS_661 0 -5.4500961227497421e-07
GC_8_662 b_8 NI_8 NS_662 0 1.4278614618032664e-05
GC_8_663 b_8 NI_8 NS_663 0 -8.7080612547193808e-05
GC_8_664 b_8 NI_8 NS_664 0 -1.9499223684521678e-04
GC_8_665 b_8 NI_8 NS_665 0 2.4925786637137105e-05
GC_8_666 b_8 NI_8 NS_666 0 3.0063957453142614e-05
GC_8_667 b_8 NI_8 NS_667 0 3.6416934071107764e-06
GC_8_668 b_8 NI_8 NS_668 0 6.3643839087499105e-06
GC_8_669 b_8 NI_8 NS_669 0 1.4328613965147781e-04
GC_8_670 b_8 NI_8 NS_670 0 -3.4079664259897528e-06
GC_8_671 b_8 NI_8 NS_671 0 -2.0326020729257585e-04
GC_8_672 b_8 NI_8 NS_672 0 -4.8355957809548004e-05
GD_8_1 b_8 NI_8 NA_1 0 4.0846446920752434e-02
GD_8_2 b_8 NI_8 NA_2 0 -4.7215764370710719e-02
GD_8_3 b_8 NI_8 NA_3 0 3.0795733089672493e-03
GD_8_4 b_8 NI_8 NA_4 0 -1.4753932160989892e-02
GD_8_5 b_8 NI_8 NA_5 0 -5.3666768120727466e-02
GD_8_6 b_8 NI_8 NA_6 0 1.1454479886759988e-02
GD_8_7 b_8 NI_8 NA_7 0 1.1794143850457886e-02
GD_8_8 b_8 NI_8 NA_8 0 1.2860800167683892e-01
GD_8_9 b_8 NI_8 NA_9 0 -1.1065509962177342e-02
GD_8_10 b_8 NI_8 NA_10 0 4.9507838724109779e-03
GD_8_11 b_8 NI_8 NA_11 0 -2.8015666332153334e-02
GD_8_12 b_8 NI_8 NA_12 0 8.8545031458919388e-03
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 4.6820193733009777e-03
GC_9_2 b_9 NI_9 NS_2 0 1.3455451164569191e-04
GC_9_3 b_9 NI_9 NS_3 0 -1.7937763128366191e-04
GC_9_4 b_9 NI_9 NS_4 0 -1.8179982547134464e-04
GC_9_5 b_9 NI_9 NS_5 0 1.1938773449187453e-04
GC_9_6 b_9 NI_9 NS_6 0 -2.8494641304710813e-04
GC_9_7 b_9 NI_9 NS_7 0 1.1086842889318381e-03
GC_9_8 b_9 NI_9 NS_8 0 -7.6331996237358028e-04
GC_9_9 b_9 NI_9 NS_9 0 1.6985078722223522e-03
GC_9_10 b_9 NI_9 NS_10 0 5.0716159345861320e-04
GC_9_11 b_9 NI_9 NS_11 0 -3.8893313591794161e-04
GC_9_12 b_9 NI_9 NS_12 0 2.1793810144571835e-04
GC_9_13 b_9 NI_9 NS_13 0 1.3070139610573839e-03
GC_9_14 b_9 NI_9 NS_14 0 -6.5820893135271139e-04
GC_9_15 b_9 NI_9 NS_15 0 1.2840784158057467e-03
GC_9_16 b_9 NI_9 NS_16 0 -5.6987637296982583e-05
GC_9_17 b_9 NI_9 NS_17 0 1.1039119511465022e-03
GC_9_18 b_9 NI_9 NS_18 0 2.3356345754331959e-03
GC_9_19 b_9 NI_9 NS_19 0 1.4822839493117796e-03
GC_9_20 b_9 NI_9 NS_20 0 8.8246726382791517e-05
GC_9_21 b_9 NI_9 NS_21 0 4.2063044098893375e-04
GC_9_22 b_9 NI_9 NS_22 0 1.9173293128909403e-04
GC_9_23 b_9 NI_9 NS_23 0 -1.2679167005112782e-04
GC_9_24 b_9 NI_9 NS_24 0 9.1803020593417481e-03
GC_9_25 b_9 NI_9 NS_25 0 -7.3660576921357769e-04
GC_9_26 b_9 NI_9 NS_26 0 -7.3117782619629406e-04
GC_9_27 b_9 NI_9 NS_27 0 -9.6407865161816312e-04
GC_9_28 b_9 NI_9 NS_28 0 -9.3676360295974956e-05
GC_9_29 b_9 NI_9 NS_29 0 -4.0627976559064113e-04
GC_9_30 b_9 NI_9 NS_30 0 -4.1332466723879749e-04
GC_9_31 b_9 NI_9 NS_31 0 -8.3705885274028345e-05
GC_9_32 b_9 NI_9 NS_32 0 -3.0450248696298647e-06
GC_9_33 b_9 NI_9 NS_33 0 -5.0694599385429509e-03
GC_9_34 b_9 NI_9 NS_34 0 -1.3984832079220544e-03
GC_9_35 b_9 NI_9 NS_35 0 1.2594835051516269e-05
GC_9_36 b_9 NI_9 NS_36 0 -2.2330847104459686e-05
GC_9_37 b_9 NI_9 NS_37 0 2.6398337714938995e-05
GC_9_38 b_9 NI_9 NS_38 0 2.9797190786075821e-04
GC_9_39 b_9 NI_9 NS_39 0 1.3575794346306147e-03
GC_9_40 b_9 NI_9 NS_40 0 -2.1416889199587642e-03
GC_9_41 b_9 NI_9 NS_41 0 6.4852876908834644e-05
GC_9_42 b_9 NI_9 NS_42 0 1.4315027374501684e-04
GC_9_43 b_9 NI_9 NS_43 0 -1.9190585948826536e-06
GC_9_44 b_9 NI_9 NS_44 0 1.8204297699309113e-06
GC_9_45 b_9 NI_9 NS_45 0 -1.3029505583412322e-06
GC_9_46 b_9 NI_9 NS_46 0 -7.5787941748140525e-06
GC_9_47 b_9 NI_9 NS_47 0 -1.1522831343385523e-04
GC_9_48 b_9 NI_9 NS_48 0 8.3892111363659236e-05
GC_9_49 b_9 NI_9 NS_49 0 2.6508552589837500e-06
GC_9_50 b_9 NI_9 NS_50 0 -1.7725512114260788e-05
GC_9_51 b_9 NI_9 NS_51 0 -1.1609215501782093e-05
GC_9_52 b_9 NI_9 NS_52 0 -1.4127494152208948e-05
GC_9_53 b_9 NI_9 NS_53 0 5.3961300645250788e-05
GC_9_54 b_9 NI_9 NS_54 0 -2.0720651495250077e-05
GC_9_55 b_9 NI_9 NS_55 0 -9.3365193214066015e-05
GC_9_56 b_9 NI_9 NS_56 0 5.0058813621006560e-06
GC_9_57 b_9 NI_9 NS_57 0 6.8933819317371975e-03
GC_9_58 b_9 NI_9 NS_58 0 -1.0644520660841122e-04
GC_9_59 b_9 NI_9 NS_59 0 2.0352845610878479e-04
GC_9_60 b_9 NI_9 NS_60 0 1.3318975982351267e-05
GC_9_61 b_9 NI_9 NS_61 0 1.1210497364423441e-04
GC_9_62 b_9 NI_9 NS_62 0 2.4840970216945138e-04
GC_9_63 b_9 NI_9 NS_63 0 -2.9209880167959399e-04
GC_9_64 b_9 NI_9 NS_64 0 1.2655702757035381e-03
GC_9_65 b_9 NI_9 NS_65 0 -1.6527243209261983e-03
GC_9_66 b_9 NI_9 NS_66 0 6.1720321042234977e-04
GC_9_67 b_9 NI_9 NS_67 0 2.2969805698756112e-05
GC_9_68 b_9 NI_9 NS_68 0 -6.7241150208200752e-04
GC_9_69 b_9 NI_9 NS_69 0 -5.0508664300454465e-04
GC_9_70 b_9 NI_9 NS_70 0 -9.5467609399883476e-04
GC_9_71 b_9 NI_9 NS_71 0 5.8454731615151397e-04
GC_9_72 b_9 NI_9 NS_72 0 -3.7083277568562519e-04
GC_9_73 b_9 NI_9 NS_73 0 1.4122577837828887e-03
GC_9_74 b_9 NI_9 NS_74 0 1.0497249932318320e-03
GC_9_75 b_9 NI_9 NS_75 0 -7.0611981297373039e-04
GC_9_76 b_9 NI_9 NS_76 0 2.2659496003996837e-03
GC_9_77 b_9 NI_9 NS_77 0 -1.9643866248943300e-04
GC_9_78 b_9 NI_9 NS_78 0 -3.9496959101380790e-05
GC_9_79 b_9 NI_9 NS_79 0 -2.8171317767991689e-03
GC_9_80 b_9 NI_9 NS_80 0 1.8507465934603036e-03
GC_9_81 b_9 NI_9 NS_81 0 3.4238746154201477e-04
GC_9_82 b_9 NI_9 NS_82 0 3.9183739306527469e-04
GC_9_83 b_9 NI_9 NS_83 0 -7.2355628482087357e-04
GC_9_84 b_9 NI_9 NS_84 0 6.4083023709937838e-05
GC_9_85 b_9 NI_9 NS_85 0 -4.8192077080356382e-04
GC_9_86 b_9 NI_9 NS_86 0 -8.8720984606139423e-06
GC_9_87 b_9 NI_9 NS_87 0 -1.0675296667507107e-04
GC_9_88 b_9 NI_9 NS_88 0 -3.9732297252253097e-05
GC_9_89 b_9 NI_9 NS_89 0 -1.2492284417949349e-03
GC_9_90 b_9 NI_9 NS_90 0 -5.7938783285366151e-03
GC_9_91 b_9 NI_9 NS_91 0 5.3639413470012642e-05
GC_9_92 b_9 NI_9 NS_92 0 -2.3815449607107405e-05
GC_9_93 b_9 NI_9 NS_93 0 -1.1841675076438498e-03
GC_9_94 b_9 NI_9 NS_94 0 4.7077786491127733e-04
GC_9_95 b_9 NI_9 NS_95 0 2.2133158999136514e-03
GC_9_96 b_9 NI_9 NS_96 0 9.0375708430026288e-04
GC_9_97 b_9 NI_9 NS_97 0 -5.5571860225965378e-05
GC_9_98 b_9 NI_9 NS_98 0 8.5588308608973684e-05
GC_9_99 b_9 NI_9 NS_99 0 -1.8478033189094941e-06
GC_9_100 b_9 NI_9 NS_100 0 6.1298819363270878e-07
GC_9_101 b_9 NI_9 NS_101 0 4.5507247071036966e-06
GC_9_102 b_9 NI_9 NS_102 0 -3.6783055166380175e-06
GC_9_103 b_9 NI_9 NS_103 0 -1.4969050344469165e-04
GC_9_104 b_9 NI_9 NS_104 0 -7.6982179370288942e-05
GC_9_105 b_9 NI_9 NS_105 0 1.1121307654498568e-05
GC_9_106 b_9 NI_9 NS_106 0 -2.1018406954294489e-06
GC_9_107 b_9 NI_9 NS_107 0 6.6808464656234170e-06
GC_9_108 b_9 NI_9 NS_108 0 -1.1074127821092204e-05
GC_9_109 b_9 NI_9 NS_109 0 3.3025178294554193e-05
GC_9_110 b_9 NI_9 NS_110 0 4.5271129853257535e-05
GC_9_111 b_9 NI_9 NS_111 0 -2.7214012701548313e-05
GC_9_112 b_9 NI_9 NS_112 0 -8.3981291251004116e-05
GC_9_113 b_9 NI_9 NS_113 0 1.1882631102822000e-02
GC_9_114 b_9 NI_9 NS_114 0 1.4764342989833561e-04
GC_9_115 b_9 NI_9 NS_115 0 -5.3398686662380099e-05
GC_9_116 b_9 NI_9 NS_116 0 -4.2102087572420678e-04
GC_9_117 b_9 NI_9 NS_117 0 3.8317487005453928e-04
GC_9_118 b_9 NI_9 NS_118 0 -3.7460189626586755e-05
GC_9_119 b_9 NI_9 NS_119 0 1.4796056176766233e-03
GC_9_120 b_9 NI_9 NS_120 0 -6.7680496518397434e-06
GC_9_121 b_9 NI_9 NS_121 0 7.6812323413617790e-04
GC_9_122 b_9 NI_9 NS_122 0 1.4996449982156196e-03
GC_9_123 b_9 NI_9 NS_123 0 -6.6989975854509019e-04
GC_9_124 b_9 NI_9 NS_124 0 2.0341095115673433e-04
GC_9_125 b_9 NI_9 NS_125 0 1.5028186362214245e-03
GC_9_126 b_9 NI_9 NS_126 0 -1.1499122455179605e-03
GC_9_127 b_9 NI_9 NS_127 0 1.8186828969276815e-03
GC_9_128 b_9 NI_9 NS_128 0 5.9667258851469708e-05
GC_9_129 b_9 NI_9 NS_129 0 8.4398209847270692e-05
GC_9_130 b_9 NI_9 NS_130 0 2.7198332830253771e-03
GC_9_131 b_9 NI_9 NS_131 0 2.9815000925641935e-03
GC_9_132 b_9 NI_9 NS_132 0 2.1941592178053096e-04
GC_9_133 b_9 NI_9 NS_133 0 6.0527599184139608e-04
GC_9_134 b_9 NI_9 NS_134 0 2.8814940486919830e-04
GC_9_135 b_9 NI_9 NS_135 0 -7.2197180975616324e-04
GC_9_136 b_9 NI_9 NS_136 0 1.1775135480021529e-02
GC_9_137 b_9 NI_9 NS_137 0 -8.4249396361468819e-04
GC_9_138 b_9 NI_9 NS_138 0 -1.0914240584642518e-03
GC_9_139 b_9 NI_9 NS_139 0 -1.3554585215734979e-03
GC_9_140 b_9 NI_9 NS_140 0 -1.1284117148347986e-05
GC_9_141 b_9 NI_9 NS_141 0 -5.1981516851299769e-04
GC_9_142 b_9 NI_9 NS_142 0 -4.4011104029951424e-04
GC_9_143 b_9 NI_9 NS_143 0 -1.3884847390258011e-04
GC_9_144 b_9 NI_9 NS_144 0 3.8054941468428748e-05
GC_9_145 b_9 NI_9 NS_145 0 -6.2717937526371604e-03
GC_9_146 b_9 NI_9 NS_146 0 -1.5195153023896844e-03
GC_9_147 b_9 NI_9 NS_147 0 3.3755317058809882e-05
GC_9_148 b_9 NI_9 NS_148 0 -4.5268963100435592e-05
GC_9_149 b_9 NI_9 NS_149 0 1.0857337633124402e-04
GC_9_150 b_9 NI_9 NS_150 0 7.5451808166348254e-04
GC_9_151 b_9 NI_9 NS_151 0 9.3791498970179185e-04
GC_9_152 b_9 NI_9 NS_152 0 -3.1098494944524274e-03
GC_9_153 b_9 NI_9 NS_153 0 1.9400010602378744e-05
GC_9_154 b_9 NI_9 NS_154 0 8.1218386611998906e-05
GC_9_155 b_9 NI_9 NS_155 0 -2.1435995808330310e-07
GC_9_156 b_9 NI_9 NS_156 0 1.4075854966144826e-06
GC_9_157 b_9 NI_9 NS_157 0 -1.6694584153990589e-06
GC_9_158 b_9 NI_9 NS_158 0 -9.7022253062794245e-06
GC_9_159 b_9 NI_9 NS_159 0 -1.2083548515405254e-04
GC_9_160 b_9 NI_9 NS_160 0 1.1974123843556082e-04
GC_9_161 b_9 NI_9 NS_161 0 1.1021616179431005e-06
GC_9_162 b_9 NI_9 NS_162 0 -2.0671068150308007e-05
GC_9_163 b_9 NI_9 NS_163 0 -1.5485134567533730e-05
GC_9_164 b_9 NI_9 NS_164 0 -4.9914990418443104e-06
GC_9_165 b_9 NI_9 NS_165 0 4.0908954193444895e-05
GC_9_166 b_9 NI_9 NS_166 0 -4.3805200845320286e-05
GC_9_167 b_9 NI_9 NS_167 0 -8.1823357208872852e-05
GC_9_168 b_9 NI_9 NS_168 0 4.5837541201366886e-05
GC_9_169 b_9 NI_9 NS_169 0 8.3541258382938393e-03
GC_9_170 b_9 NI_9 NS_170 0 -1.5596779753314320e-04
GC_9_171 b_9 NI_9 NS_171 0 2.9992008258203877e-04
GC_9_172 b_9 NI_9 NS_172 0 1.6281321917315317e-04
GC_9_173 b_9 NI_9 NS_173 0 -7.2501531760112996e-05
GC_9_174 b_9 NI_9 NS_174 0 3.3259414805536823e-04
GC_9_175 b_9 NI_9 NS_175 0 -8.9291454119769015e-04
GC_9_176 b_9 NI_9 NS_176 0 1.2037554243242861e-03
GC_9_177 b_9 NI_9 NS_177 0 -1.5304361208722716e-03
GC_9_178 b_9 NI_9 NS_178 0 -2.8040310377854352e-04
GC_9_179 b_9 NI_9 NS_179 0 -7.1976696993412913e-05
GC_9_180 b_9 NI_9 NS_180 0 -4.3687741543247917e-04
GC_9_181 b_9 NI_9 NS_181 0 -1.3282069440057968e-05
GC_9_182 b_9 NI_9 NS_182 0 -1.3372988690780240e-03
GC_9_183 b_9 NI_9 NS_183 0 8.4212323447791382e-04
GC_9_184 b_9 NI_9 NS_184 0 -4.9874178830061568e-04
GC_9_185 b_9 NI_9 NS_185 0 1.7715174851964887e-03
GC_9_186 b_9 NI_9 NS_186 0 1.6514170984605065e-03
GC_9_187 b_9 NI_9 NS_187 0 -4.2767996000196143e-04
GC_9_188 b_9 NI_9 NS_188 0 2.6322706769468553e-03
GC_9_189 b_9 NI_9 NS_189 0 -2.2164509615892915e-04
GC_9_190 b_9 NI_9 NS_190 0 -3.6807200594334724e-05
GC_9_191 b_9 NI_9 NS_191 0 -2.7962257153364019e-03
GC_9_192 b_9 NI_9 NS_192 0 2.2968638823893175e-03
GC_9_193 b_9 NI_9 NS_193 0 2.5995171705698770e-04
GC_9_194 b_9 NI_9 NS_194 0 3.1486733049412039e-04
GC_9_195 b_9 NI_9 NS_195 0 -8.7293648607055842e-04
GC_9_196 b_9 NI_9 NS_196 0 5.9799869603462516e-05
GC_9_197 b_9 NI_9 NS_197 0 -4.4767132611169198e-04
GC_9_198 b_9 NI_9 NS_198 0 -4.9558419342296026e-06
GC_9_199 b_9 NI_9 NS_199 0 -1.0010037658396160e-04
GC_9_200 b_9 NI_9 NS_200 0 -2.7372519025515961e-05
GC_9_201 b_9 NI_9 NS_201 0 -9.3885194285238513e-04
GC_9_202 b_9 NI_9 NS_202 0 -4.9262550703032346e-03
GC_9_203 b_9 NI_9 NS_203 0 4.9795896337529949e-05
GC_9_204 b_9 NI_9 NS_204 0 -3.2849116563780163e-05
GC_9_205 b_9 NI_9 NS_205 0 -1.0385789816069601e-03
GC_9_206 b_9 NI_9 NS_206 0 6.1131235076372495e-04
GC_9_207 b_9 NI_9 NS_207 0 1.3134074791239722e-03
GC_9_208 b_9 NI_9 NS_208 0 -3.7140542410153305e-05
GC_9_209 b_9 NI_9 NS_209 0 -1.1646922975173986e-04
GC_9_210 b_9 NI_9 NS_210 0 1.1464536013113547e-04
GC_9_211 b_9 NI_9 NS_211 0 -8.6928792501424128e-07
GC_9_212 b_9 NI_9 NS_212 0 7.0669456043002657e-07
GC_9_213 b_9 NI_9 NS_213 0 -6.8625981140867011e-07
GC_9_214 b_9 NI_9 NS_214 0 -3.6740313875643924e-06
GC_9_215 b_9 NI_9 NS_215 0 -5.5523096424088058e-05
GC_9_216 b_9 NI_9 NS_216 0 9.0751851989141830e-06
GC_9_217 b_9 NI_9 NS_217 0 -4.6765968021492481e-07
GC_9_218 b_9 NI_9 NS_218 0 -4.3128747410621659e-06
GC_9_219 b_9 NI_9 NS_219 0 -8.7701489183284435e-07
GC_9_220 b_9 NI_9 NS_220 0 -4.6204918300469818e-06
GC_9_221 b_9 NI_9 NS_221 0 1.9695804147523425e-05
GC_9_222 b_9 NI_9 NS_222 0 1.2629825504410162e-05
GC_9_223 b_9 NI_9 NS_223 0 -2.3089587112919471e-05
GC_9_224 b_9 NI_9 NS_224 0 -2.7862051852016453e-05
GC_9_225 b_9 NI_9 NS_225 0 1.6594667329139692e-02
GC_9_226 b_9 NI_9 NS_226 0 7.0318859551569312e-05
GC_9_227 b_9 NI_9 NS_227 0 3.4521977071536746e-04
GC_9_228 b_9 NI_9 NS_228 0 -5.9571325588324764e-04
GC_9_229 b_9 NI_9 NS_229 0 5.5723014782166661e-04
GC_9_230 b_9 NI_9 NS_230 0 5.9051322702690886e-04
GC_9_231 b_9 NI_9 NS_231 0 9.6860272631444603e-04
GC_9_232 b_9 NI_9 NS_232 0 1.5952511360160658e-03
GC_9_233 b_9 NI_9 NS_233 0 -1.8403884151855716e-03
GC_9_234 b_9 NI_9 NS_234 0 2.0946128963686104e-03
GC_9_235 b_9 NI_9 NS_235 0 -5.2514714555220246e-04
GC_9_236 b_9 NI_9 NS_236 0 9.7683221468087257e-05
GC_9_237 b_9 NI_9 NS_237 0 1.0907044888765528e-03
GC_9_238 b_9 NI_9 NS_238 0 -1.4801753050581214e-03
GC_9_239 b_9 NI_9 NS_239 0 1.7808080112936536e-03
GC_9_240 b_9 NI_9 NS_240 0 2.3823357199195946e-04
GC_9_241 b_9 NI_9 NS_241 0 -1.7801516805620770e-03
GC_9_242 b_9 NI_9 NS_242 0 2.2762580253603702e-03
GC_9_243 b_9 NI_9 NS_243 0 3.1635955106168300e-03
GC_9_244 b_9 NI_9 NS_244 0 3.2254516397133421e-04
GC_9_245 b_9 NI_9 NS_245 0 6.6354827695973425e-04
GC_9_246 b_9 NI_9 NS_246 0 2.3564052648416184e-04
GC_9_247 b_9 NI_9 NS_247 0 -2.0617957575215702e-03
GC_9_248 b_9 NI_9 NS_248 0 9.8864751025469957e-03
GC_9_249 b_9 NI_9 NS_249 0 -6.7550175779439929e-04
GC_9_250 b_9 NI_9 NS_250 0 -1.1182329437895210e-03
GC_9_251 b_9 NI_9 NS_251 0 -1.3538842882976131e-03
GC_9_252 b_9 NI_9 NS_252 0 -7.6675928359332354e-05
GC_9_253 b_9 NI_9 NS_253 0 -4.3685064029532936e-04
GC_9_254 b_9 NI_9 NS_254 0 -4.4075101080813127e-04
GC_9_255 b_9 NI_9 NS_255 0 -1.4473566013819080e-04
GC_9_256 b_9 NI_9 NS_256 0 6.2679330690234027e-05
GC_9_257 b_9 NI_9 NS_257 0 -6.6117468612332669e-03
GC_9_258 b_9 NI_9 NS_258 0 -1.9570618735265306e-03
GC_9_259 b_9 NI_9 NS_259 0 4.4554872793218802e-05
GC_9_260 b_9 NI_9 NS_260 0 -4.4973188765047184e-05
GC_9_261 b_9 NI_9 NS_261 0 1.5725340361858218e-04
GC_9_262 b_9 NI_9 NS_262 0 8.0303519934886165e-04
GC_9_263 b_9 NI_9 NS_263 0 1.9112785606035635e-03
GC_9_264 b_9 NI_9 NS_264 0 -3.3766263260939021e-03
GC_9_265 b_9 NI_9 NS_265 0 1.7647765384314553e-04
GC_9_266 b_9 NI_9 NS_266 0 -7.0996282362700423e-05
GC_9_267 b_9 NI_9 NS_267 0 8.5063809165205915e-07
GC_9_268 b_9 NI_9 NS_268 0 1.0260547196360690e-06
GC_9_269 b_9 NI_9 NS_269 0 -9.2011063650338917e-07
GC_9_270 b_9 NI_9 NS_270 0 -4.4139528966115161e-06
GC_9_271 b_9 NI_9 NS_271 0 -7.0792848735291638e-05
GC_9_272 b_9 NI_9 NS_272 0 8.2935389400432165e-05
GC_9_273 b_9 NI_9 NS_273 0 -1.2442848322446925e-06
GC_9_274 b_9 NI_9 NS_274 0 -1.0140729101520384e-05
GC_9_275 b_9 NI_9 NS_275 0 -8.8664765604982487e-06
GC_9_276 b_9 NI_9 NS_276 0 3.3726463339187262e-06
GC_9_277 b_9 NI_9 NS_277 0 3.5762710489409879e-06
GC_9_278 b_9 NI_9 NS_278 0 -3.0691973680872618e-05
GC_9_279 b_9 NI_9 NS_279 0 -1.8496310141823543e-05
GC_9_280 b_9 NI_9 NS_280 0 4.4777898608898780e-05
GC_9_281 b_9 NI_9 NS_281 0 4.1248735162779694e-03
GC_9_282 b_9 NI_9 NS_282 0 -1.5392334138853949e-04
GC_9_283 b_9 NI_9 NS_283 0 2.7446041455699965e-04
GC_9_284 b_9 NI_9 NS_284 0 4.0117508684404588e-04
GC_9_285 b_9 NI_9 NS_285 0 -4.0838844077429329e-04
GC_9_286 b_9 NI_9 NS_286 0 2.2079773903080536e-04
GC_9_287 b_9 NI_9 NS_287 0 -1.4768738065858121e-03
GC_9_288 b_9 NI_9 NS_288 0 2.6789300943573383e-04
GC_9_289 b_9 NI_9 NS_289 0 -2.0974100046716539e-04
GC_9_290 b_9 NI_9 NS_290 0 -1.5836128807354864e-03
GC_9_291 b_9 NI_9 NS_291 0 2.4930988362045276e-04
GC_9_292 b_9 NI_9 NS_292 0 -3.0220887383606209e-04
GC_9_293 b_9 NI_9 NS_293 0 7.5794081165343752e-04
GC_9_294 b_9 NI_9 NS_294 0 -1.3224230678526132e-03
GC_9_295 b_9 NI_9 NS_295 0 1.0549633435392796e-03
GC_9_296 b_9 NI_9 NS_296 0 -6.1054241004260799e-04
GC_9_297 b_9 NI_9 NS_297 0 1.8024077582086168e-03
GC_9_298 b_9 NI_9 NS_298 0 2.1958211206105113e-03
GC_9_299 b_9 NI_9 NS_299 0 2.1552121217277606e-05
GC_9_300 b_9 NI_9 NS_300 0 3.0033475850760735e-03
GC_9_301 b_9 NI_9 NS_301 0 -3.6056586731093995e-04
GC_9_302 b_9 NI_9 NS_302 0 -3.0601841440729404e-05
GC_9_303 b_9 NI_9 NS_303 0 -2.9682062250619263e-03
GC_9_304 b_9 NI_9 NS_304 0 2.6848353164425926e-03
GC_9_305 b_9 NI_9 NS_305 0 3.0309159413288982e-04
GC_9_306 b_9 NI_9 NS_306 0 1.3050530604742777e-04
GC_9_307 b_9 NI_9 NS_307 0 -1.1219286661006283e-03
GC_9_308 b_9 NI_9 NS_308 0 2.1765067958345541e-04
GC_9_309 b_9 NI_9 NS_309 0 -6.5007171853898081e-04
GC_9_310 b_9 NI_9 NS_310 0 -3.8175466618986309e-05
GC_9_311 b_9 NI_9 NS_311 0 -1.3739808880823339e-04
GC_9_312 b_9 NI_9 NS_312 0 -4.8361442042419351e-05
GC_9_313 b_9 NI_9 NS_313 0 -1.1893402914246730e-04
GC_9_314 b_9 NI_9 NS_314 0 -4.7085156800225746e-03
GC_9_315 b_9 NI_9 NS_315 0 4.2051358884187370e-05
GC_9_316 b_9 NI_9 NS_316 0 -4.1593807455516627e-05
GC_9_317 b_9 NI_9 NS_317 0 -1.2917437469168664e-03
GC_9_318 b_9 NI_9 NS_318 0 5.7009472433745248e-04
GC_9_319 b_9 NI_9 NS_319 0 1.3332622966488949e-03
GC_9_320 b_9 NI_9 NS_320 0 -9.4753626799040256e-04
GC_9_321 b_9 NI_9 NS_321 0 -2.0495660229751932e-04
GC_9_322 b_9 NI_9 NS_322 0 7.9387880350139715e-05
GC_9_323 b_9 NI_9 NS_323 0 -5.8380314157147257e-07
GC_9_324 b_9 NI_9 NS_324 0 5.5713215027144534e-07
GC_9_325 b_9 NI_9 NS_325 0 -4.5690054010003060e-06
GC_9_326 b_9 NI_9 NS_326 0 -3.8528124466517836e-06
GC_9_327 b_9 NI_9 NS_327 0 -1.3739069078470229e-05
GC_9_328 b_9 NI_9 NS_328 0 6.6748953827353206e-05
GC_9_329 b_9 NI_9 NS_329 0 -9.0077353995985325e-06
GC_9_330 b_9 NI_9 NS_330 0 -5.2421504971637313e-06
GC_9_331 b_9 NI_9 NS_331 0 -5.1694465982979259e-06
GC_9_332 b_9 NI_9 NS_332 0 -4.0149249770027653e-06
GC_9_333 b_9 NI_9 NS_333 0 2.7231027217172198e-05
GC_9_334 b_9 NI_9 NS_334 0 -2.8880396130673914e-06
GC_9_335 b_9 NI_9 NS_335 0 -4.2303480978865634e-05
GC_9_336 b_9 NI_9 NS_336 0 -7.2877499947508316e-06
GC_9_337 b_9 NI_9 NS_337 0 1.9416340477204470e-03
GC_9_338 b_9 NI_9 NS_338 0 3.2031069121110730e-05
GC_9_339 b_9 NI_9 NS_339 0 1.2362677810948688e-03
GC_9_340 b_9 NI_9 NS_340 0 -1.4019328443518687e-04
GC_9_341 b_9 NI_9 NS_341 0 -1.1064620981862683e-03
GC_9_342 b_9 NI_9 NS_342 0 1.3027347410189054e-03
GC_9_343 b_9 NI_9 NS_343 0 -9.4255987248396500e-04
GC_9_344 b_9 NI_9 NS_344 0 7.3844347527969741e-04
GC_9_345 b_9 NI_9 NS_345 0 -2.7176362442537334e-03
GC_9_346 b_9 NI_9 NS_346 0 -2.9728876614770238e-03
GC_9_347 b_9 NI_9 NS_347 0 -4.2741186297786207e-04
GC_9_348 b_9 NI_9 NS_348 0 -2.8669292556651472e-04
GC_9_349 b_9 NI_9 NS_349 0 2.8452512812607864e-03
GC_9_350 b_9 NI_9 NS_350 0 -1.5783737902453155e-03
GC_9_351 b_9 NI_9 NS_351 0 1.2720878519667559e-03
GC_9_352 b_9 NI_9 NS_352 0 5.0811948482773137e-04
GC_9_353 b_9 NI_9 NS_353 0 -1.2121712727412204e-03
GC_9_354 b_9 NI_9 NS_354 0 3.9743192886841897e-05
GC_9_355 b_9 NI_9 NS_355 0 1.7014784482074642e-03
GC_9_356 b_9 NI_9 NS_356 0 2.6297830655009176e-04
GC_9_357 b_9 NI_9 NS_357 0 4.7531370668385157e-04
GC_9_358 b_9 NI_9 NS_358 0 2.3895384275884345e-04
GC_9_359 b_9 NI_9 NS_359 0 5.6138880223526955e-04
GC_9_360 b_9 NI_9 NS_360 0 5.2959347769502034e-03
GC_9_361 b_9 NI_9 NS_361 0 -3.8315521011862805e-04
GC_9_362 b_9 NI_9 NS_362 0 -7.1333702535733221e-04
GC_9_363 b_9 NI_9 NS_363 0 -8.5783890823397336e-04
GC_9_364 b_9 NI_9 NS_364 0 5.5285626863899930e-05
GC_9_365 b_9 NI_9 NS_365 0 -3.1464640976369305e-04
GC_9_366 b_9 NI_9 NS_366 0 -2.8183841873458023e-04
GC_9_367 b_9 NI_9 NS_367 0 -7.7628730691169621e-05
GC_9_368 b_9 NI_9 NS_368 0 1.2030353622552723e-05
GC_9_369 b_9 NI_9 NS_369 0 -3.3267425705240353e-03
GC_9_370 b_9 NI_9 NS_370 0 -3.9758477080991221e-03
GC_9_371 b_9 NI_9 NS_371 0 2.1321771538154930e-05
GC_9_372 b_9 NI_9 NS_372 0 -4.9501045425165453e-05
GC_9_373 b_9 NI_9 NS_373 0 1.7771430906535186e-04
GC_9_374 b_9 NI_9 NS_374 0 7.0102832119513638e-04
GC_9_375 b_9 NI_9 NS_375 0 1.9353827545411338e-03
GC_9_376 b_9 NI_9 NS_376 0 7.4141649333222615e-04
GC_9_377 b_9 NI_9 NS_377 0 9.7630824367461496e-06
GC_9_378 b_9 NI_9 NS_378 0 2.8783995955676653e-04
GC_9_379 b_9 NI_9 NS_379 0 -7.9279169472333861e-07
GC_9_380 b_9 NI_9 NS_380 0 8.8023398283821129e-07
GC_9_381 b_9 NI_9 NS_381 0 3.0800025171700536e-06
GC_9_382 b_9 NI_9 NS_382 0 -1.3996584621532602e-06
GC_9_383 b_9 NI_9 NS_383 0 -6.9636293522993151e-05
GC_9_384 b_9 NI_9 NS_384 0 -4.4378253014710921e-06
GC_9_385 b_9 NI_9 NS_385 0 6.0845856910682362e-06
GC_9_386 b_9 NI_9 NS_386 0 -1.4896805141753180e-06
GC_9_387 b_9 NI_9 NS_387 0 -4.2626239906972602e-06
GC_9_388 b_9 NI_9 NS_388 0 -4.5033614261040847e-06
GC_9_389 b_9 NI_9 NS_389 0 1.4125508773321784e-05
GC_9_390 b_9 NI_9 NS_390 0 -4.5832129622218000e-07
GC_9_391 b_9 NI_9 NS_391 0 -2.1253532751230519e-05
GC_9_392 b_9 NI_9 NS_392 0 -4.8241592714370949e-06
GC_9_393 b_9 NI_9 NS_393 0 6.5575966872878097e-03
GC_9_394 b_9 NI_9 NS_394 0 -8.5830992450280360e-05
GC_9_395 b_9 NI_9 NS_395 0 -1.9560044582076560e-04
GC_9_396 b_9 NI_9 NS_396 0 7.0113140806892893e-04
GC_9_397 b_9 NI_9 NS_397 0 -3.0825255711964286e-04
GC_9_398 b_9 NI_9 NS_398 0 -6.8120270407243111e-04
GC_9_399 b_9 NI_9 NS_399 0 -5.3653208588290825e-04
GC_9_400 b_9 NI_9 NS_400 0 -8.2810383287203941e-04
GC_9_401 b_9 NI_9 NS_401 0 2.2767881748167206e-03
GC_9_402 b_9 NI_9 NS_402 0 7.1800469728009657e-04
GC_9_403 b_9 NI_9 NS_403 0 -1.3373192929660131e-04
GC_9_404 b_9 NI_9 NS_404 0 9.7607751778178706e-05
GC_9_405 b_9 NI_9 NS_405 0 4.3128990319366088e-04
GC_9_406 b_9 NI_9 NS_406 0 -4.5673399573435106e-04
GC_9_407 b_9 NI_9 NS_407 0 8.6764235192750131e-04
GC_9_408 b_9 NI_9 NS_408 0 -1.0956052484965418e-04
GC_9_409 b_9 NI_9 NS_409 0 6.2746489213409760e-04
GC_9_410 b_9 NI_9 NS_410 0 1.9121310627733259e-03
GC_9_411 b_9 NI_9 NS_411 0 -1.2033475633371159e-03
GC_9_412 b_9 NI_9 NS_412 0 2.5524455117099938e-03
GC_9_413 b_9 NI_9 NS_413 0 -2.0076716642375943e-04
GC_9_414 b_9 NI_9 NS_414 0 -5.8802109304449291e-05
GC_9_415 b_9 NI_9 NS_415 0 -1.0135002201435649e-03
GC_9_416 b_9 NI_9 NS_416 0 1.3388406714373875e-03
GC_9_417 b_9 NI_9 NS_417 0 5.9371646449022728e-05
GC_9_418 b_9 NI_9 NS_418 0 -2.0587236094056162e-05
GC_9_419 b_9 NI_9 NS_419 0 -6.7535725235482607e-04
GC_9_420 b_9 NI_9 NS_420 0 9.0745627408578866e-05
GC_9_421 b_9 NI_9 NS_421 0 -3.9092414423357903e-04
GC_9_422 b_9 NI_9 NS_422 0 5.0439706941769043e-05
GC_9_423 b_9 NI_9 NS_423 0 -1.0766422471417303e-04
GC_9_424 b_9 NI_9 NS_424 0 -3.4998175636169162e-05
GC_9_425 b_9 NI_9 NS_425 0 -4.0384742240385043e-04
GC_9_426 b_9 NI_9 NS_426 0 -3.3770410101022471e-03
GC_9_427 b_9 NI_9 NS_427 0 3.7921578629147301e-05
GC_9_428 b_9 NI_9 NS_428 0 -1.9107425996722373e-05
GC_9_429 b_9 NI_9 NS_429 0 -8.7697648881071891e-04
GC_9_430 b_9 NI_9 NS_430 0 4.9605543422051547e-04
GC_9_431 b_9 NI_9 NS_431 0 1.2288554237793903e-03
GC_9_432 b_9 NI_9 NS_432 0 2.8811119889508548e-04
GC_9_433 b_9 NI_9 NS_433 0 -1.5361158018453752e-04
GC_9_434 b_9 NI_9 NS_434 0 2.9714120241663197e-04
GC_9_435 b_9 NI_9 NS_435 0 -1.0363969700598619e-06
GC_9_436 b_9 NI_9 NS_436 0 1.0092114316872981e-06
GC_9_437 b_9 NI_9 NS_437 0 -1.3461347410236005e-06
GC_9_438 b_9 NI_9 NS_438 0 -7.7025207375585053e-06
GC_9_439 b_9 NI_9 NS_439 0 -3.2445933987915198e-05
GC_9_440 b_9 NI_9 NS_440 0 7.4271488502179213e-05
GC_9_441 b_9 NI_9 NS_441 0 -2.2469475904022281e-06
GC_9_442 b_9 NI_9 NS_442 0 -1.3260175990176927e-05
GC_9_443 b_9 NI_9 NS_443 0 -9.0686502764366003e-06
GC_9_444 b_9 NI_9 NS_444 0 -5.2684078249172450e-06
GC_9_445 b_9 NI_9 NS_445 0 2.7479714462143472e-05
GC_9_446 b_9 NI_9 NS_446 0 -1.8543638352216629e-05
GC_9_447 b_9 NI_9 NS_447 0 -5.0924396634146231e-05
GC_9_448 b_9 NI_9 NS_448 0 1.4311934486445154e-05
GC_9_449 b_9 NI_9 NS_449 0 2.5247980355020002e-03
GC_9_450 b_9 NI_9 NS_450 0 1.4710313368974031e-02
GC_9_451 b_9 NI_9 NS_451 0 8.2619352647212690e-03
GC_9_452 b_9 NI_9 NS_452 0 1.4985133862097987e-03
GC_9_453 b_9 NI_9 NS_453 0 1.0249904836596329e-02
GC_9_454 b_9 NI_9 NS_454 0 5.1619435267735566e-03
GC_9_455 b_9 NI_9 NS_455 0 -2.9918828077657904e-03
GC_9_456 b_9 NI_9 NS_456 0 9.8656148851220659e-03
GC_9_457 b_9 NI_9 NS_457 0 -3.1687870787734406e-03
GC_9_458 b_9 NI_9 NS_458 0 6.9153751696843027e-03
GC_9_459 b_9 NI_9 NS_459 0 2.6996266456174754e-04
GC_9_460 b_9 NI_9 NS_460 0 6.5327873026185758e-04
GC_9_461 b_9 NI_9 NS_461 0 1.0467854392101527e-02
GC_9_462 b_9 NI_9 NS_462 0 -1.9132729995608290e-03
GC_9_463 b_9 NI_9 NS_463 0 4.2702129557944756e-04
GC_9_464 b_9 NI_9 NS_464 0 3.0437028297275086e-03
GC_9_465 b_9 NI_9 NS_465 0 3.8753930220827258e-03
GC_9_466 b_9 NI_9 NS_466 0 2.8320447973731373e-03
GC_9_467 b_9 NI_9 NS_467 0 4.1982933499541851e-03
GC_9_468 b_9 NI_9 NS_468 0 8.3505196172775943e-03
GC_9_469 b_9 NI_9 NS_469 0 4.3191378120000878e-04
GC_9_470 b_9 NI_9 NS_470 0 1.6169645700237867e-04
GC_9_471 b_9 NI_9 NS_471 0 -9.2116590205516130e-03
GC_9_472 b_9 NI_9 NS_472 0 7.6270852077894935e-03
GC_9_473 b_9 NI_9 NS_473 0 1.4948087492136395e-03
GC_9_474 b_9 NI_9 NS_474 0 4.3106164413618818e-04
GC_9_475 b_9 NI_9 NS_475 0 -5.5000633834982214e-04
GC_9_476 b_9 NI_9 NS_476 0 -7.5624040852503285e-05
GC_9_477 b_9 NI_9 NS_477 0 -3.1239027731875103e-04
GC_9_478 b_9 NI_9 NS_478 0 1.7054545264081171e-04
GC_9_479 b_9 NI_9 NS_479 0 -8.1310243618824216e-05
GC_9_480 b_9 NI_9 NS_480 0 -3.6915557234246350e-05
GC_9_481 b_9 NI_9 NS_481 0 -5.8766089881410787e-03
GC_9_482 b_9 NI_9 NS_482 0 -4.6187889613036734e-03
GC_9_483 b_9 NI_9 NS_483 0 1.2095613407326467e-04
GC_9_484 b_9 NI_9 NS_484 0 -1.8938624479076750e-05
GC_9_485 b_9 NI_9 NS_485 0 -7.0347298269695193e-04
GC_9_486 b_9 NI_9 NS_486 0 2.0182410115955596e-03
GC_9_487 b_9 NI_9 NS_487 0 3.7763291076257474e-03
GC_9_488 b_9 NI_9 NS_488 0 1.5535528692815317e-03
GC_9_489 b_9 NI_9 NS_489 0 2.4040298979492711e-04
GC_9_490 b_9 NI_9 NS_490 0 -2.6460403844141431e-05
GC_9_491 b_9 NI_9 NS_491 0 2.0886624939318416e-07
GC_9_492 b_9 NI_9 NS_492 0 1.3233540831239346e-06
GC_9_493 b_9 NI_9 NS_493 0 7.8881668842725300e-07
GC_9_494 b_9 NI_9 NS_494 0 -3.9964493828097052e-06
GC_9_495 b_9 NI_9 NS_495 0 -8.2043881397486816e-05
GC_9_496 b_9 NI_9 NS_496 0 8.2305498286765899e-05
GC_9_497 b_9 NI_9 NS_497 0 2.3851863508574594e-06
GC_9_498 b_9 NI_9 NS_498 0 -9.5805462424077242e-06
GC_9_499 b_9 NI_9 NS_499 0 -4.9096478199199823e-06
GC_9_500 b_9 NI_9 NS_500 0 -9.2238988223816164e-06
GC_9_501 b_9 NI_9 NS_501 0 3.6031056303510595e-05
GC_9_502 b_9 NI_9 NS_502 0 -1.0748204840069785e-05
GC_9_503 b_9 NI_9 NS_503 0 -6.0747891294564730e-05
GC_9_504 b_9 NI_9 NS_504 0 -1.9761997652449887e-06
GC_9_505 b_9 NI_9 NS_505 0 -4.5487796352564662e-02
GC_9_506 b_9 NI_9 NS_506 0 1.2148228660640269e-02
GC_9_507 b_9 NI_9 NS_507 0 -2.9338491313858480e-03
GC_9_508 b_9 NI_9 NS_508 0 3.7223078412582664e-03
GC_9_509 b_9 NI_9 NS_509 0 -4.3639025693567009e-03
GC_9_510 b_9 NI_9 NS_510 0 2.1017782713831771e-03
GC_9_511 b_9 NI_9 NS_511 0 -4.7808389670069102e-03
GC_9_512 b_9 NI_9 NS_512 0 -9.2825516534754144e-03
GC_9_513 b_9 NI_9 NS_513 0 -2.4143535033857555e-03
GC_9_514 b_9 NI_9 NS_514 0 -9.2045340358129796e-03
GC_9_515 b_9 NI_9 NS_515 0 4.6184473684348688e-04
GC_9_516 b_9 NI_9 NS_516 0 1.6663514010241144e-04
GC_9_517 b_9 NI_9 NS_517 0 7.2088874857577220e-03
GC_9_518 b_9 NI_9 NS_518 0 -1.5917336433331104e-03
GC_9_519 b_9 NI_9 NS_519 0 1.5076664056013192e-03
GC_9_520 b_9 NI_9 NS_520 0 1.2646463673084253e-03
GC_9_521 b_9 NI_9 NS_521 0 5.5694862594700672e-03
GC_9_522 b_9 NI_9 NS_522 0 8.2374936308816558e-04
GC_9_523 b_9 NI_9 NS_523 0 -2.3798214792863539e-03
GC_9_524 b_9 NI_9 NS_524 0 1.1646685864850712e-03
GC_9_525 b_9 NI_9 NS_525 0 -3.7364946906555337e-04
GC_9_526 b_9 NI_9 NS_526 0 6.8805461772152772e-05
GC_9_527 b_9 NI_9 NS_527 0 7.9978305804422733e-03
GC_9_528 b_9 NI_9 NS_528 0 -2.7376528324723729e-03
GC_9_529 b_9 NI_9 NS_529 0 -1.7443061658780959e-03
GC_9_530 b_9 NI_9 NS_530 0 -2.4148591880055804e-05
GC_9_531 b_9 NI_9 NS_531 0 -2.8142285364360451e-04
GC_9_532 b_9 NI_9 NS_532 0 1.2194196255424714e-04
GC_9_533 b_9 NI_9 NS_533 0 -4.5359873834361421e-04
GC_9_534 b_9 NI_9 NS_534 0 3.9177316353462995e-04
GC_9_535 b_9 NI_9 NS_535 0 -2.9623790450574204e-04
GC_9_536 b_9 NI_9 NS_536 0 -1.2279932372062576e-04
GC_9_537 b_9 NI_9 NS_537 0 3.0255442046477469e-03
GC_9_538 b_9 NI_9 NS_538 0 -6.4864083202423946e-04
GC_9_539 b_9 NI_9 NS_539 0 -2.6897399974703586e-05
GC_9_540 b_9 NI_9 NS_540 0 1.7986425700643462e-04
GC_9_541 b_9 NI_9 NS_541 0 -9.3160705693087135e-04
GC_9_542 b_9 NI_9 NS_542 0 -9.7637406028100861e-04
GC_9_543 b_9 NI_9 NS_543 0 1.8590623756113394e-03
GC_9_544 b_9 NI_9 NS_544 0 1.6027031518645264e-03
GC_9_545 b_9 NI_9 NS_545 0 -1.2831012875595368e-04
GC_9_546 b_9 NI_9 NS_546 0 -1.7211462906121749e-04
GC_9_547 b_9 NI_9 NS_547 0 1.6045233974695179e-06
GC_9_548 b_9 NI_9 NS_548 0 -2.1324659601866400e-06
GC_9_549 b_9 NI_9 NS_549 0 3.7688557184548187e-06
GC_9_550 b_9 NI_9 NS_550 0 -1.9773669689776115e-06
GC_9_551 b_9 NI_9 NS_551 0 -6.8083975012310762e-05
GC_9_552 b_9 NI_9 NS_552 0 -8.9521503356574099e-05
GC_9_553 b_9 NI_9 NS_553 0 9.4196724112307239e-06
GC_9_554 b_9 NI_9 NS_554 0 4.0979500173543544e-06
GC_9_555 b_9 NI_9 NS_555 0 2.4615715259585929e-06
GC_9_556 b_9 NI_9 NS_556 0 -1.1024984342040940e-05
GC_9_557 b_9 NI_9 NS_557 0 2.6530205701223499e-05
GC_9_558 b_9 NI_9 NS_558 0 6.1448239003761022e-05
GC_9_559 b_9 NI_9 NS_559 0 -1.0121360653444262e-05
GC_9_560 b_9 NI_9 NS_560 0 -1.0469942576158123e-04
GC_9_561 b_9 NI_9 NS_561 0 -1.2339460024620904e-02
GC_9_562 b_9 NI_9 NS_562 0 1.5846354246809688e-03
GC_9_563 b_9 NI_9 NS_563 0 3.7051082345272131e-03
GC_9_564 b_9 NI_9 NS_564 0 2.4603662628618207e-03
GC_9_565 b_9 NI_9 NS_565 0 -5.2611608997405277e-03
GC_9_566 b_9 NI_9 NS_566 0 -6.3979683759242800e-03
GC_9_567 b_9 NI_9 NS_567 0 4.0078752075361082e-03
GC_9_568 b_9 NI_9 NS_568 0 2.5416635664440635e-03
GC_9_569 b_9 NI_9 NS_569 0 1.0136069275778857e-02
GC_9_570 b_9 NI_9 NS_570 0 -9.6415195120840031e-03
GC_9_571 b_9 NI_9 NS_571 0 -6.6842177128775566e-04
GC_9_572 b_9 NI_9 NS_572 0 5.3367257005240362e-04
GC_9_573 b_9 NI_9 NS_573 0 8.6833936288767590e-03
GC_9_574 b_9 NI_9 NS_574 0 3.3057946206562798e-03
GC_9_575 b_9 NI_9 NS_575 0 7.8724626817749076e-04
GC_9_576 b_9 NI_9 NS_576 0 2.0745267491033494e-03
GC_9_577 b_9 NI_9 NS_577 0 7.2191421889326460e-03
GC_9_578 b_9 NI_9 NS_578 0 1.6343651060941162e-03
GC_9_579 b_9 NI_9 NS_579 0 2.5992257205273784e-03
GC_9_580 b_9 NI_9 NS_580 0 4.3715633733231521e-03
GC_9_581 b_9 NI_9 NS_581 0 3.5240276956963255e-04
GC_9_582 b_9 NI_9 NS_582 0 1.0351618503230559e-04
GC_9_583 b_9 NI_9 NS_583 0 -4.5456942019812020e-03
GC_9_584 b_9 NI_9 NS_584 0 1.4407891628132205e-02
GC_9_585 b_9 NI_9 NS_585 0 1.0571347388658690e-03
GC_9_586 b_9 NI_9 NS_586 0 -2.4327580233868151e-05
GC_9_587 b_9 NI_9 NS_587 0 -5.9672236130086254e-04
GC_9_588 b_9 NI_9 NS_588 0 9.1789594268748968e-05
GC_9_589 b_9 NI_9 NS_589 0 -1.7944462537753617e-04
GC_9_590 b_9 NI_9 NS_590 0 2.1211104306915807e-04
GC_9_591 b_9 NI_9 NS_591 0 -7.5002204617271990e-05
GC_9_592 b_9 NI_9 NS_592 0 4.3474499455337071e-05
GC_9_593 b_9 NI_9 NS_593 0 -5.9431781270191638e-03
GC_9_594 b_9 NI_9 NS_594 0 -3.3187183759156498e-03
GC_9_595 b_9 NI_9 NS_595 0 8.5373790590596486e-05
GC_9_596 b_9 NI_9 NS_596 0 -6.5301450676977010e-05
GC_9_597 b_9 NI_9 NS_597 0 -3.4575409487594102e-05
GC_9_598 b_9 NI_9 NS_598 0 1.9728702383117959e-03
GC_9_599 b_9 NI_9 NS_599 0 -2.0814144959787413e-04
GC_9_600 b_9 NI_9 NS_600 0 -1.0923361934782405e-03
GC_9_601 b_9 NI_9 NS_601 0 6.7147092839219628e-05
GC_9_602 b_9 NI_9 NS_602 0 2.9052599824354683e-04
GC_9_603 b_9 NI_9 NS_603 0 -1.9245354080711748e-07
GC_9_604 b_9 NI_9 NS_604 0 7.2388099753888941e-07
GC_9_605 b_9 NI_9 NS_605 0 -1.4758363015917262e-06
GC_9_606 b_9 NI_9 NS_606 0 5.0749362455750604e-07
GC_9_607 b_9 NI_9 NS_607 0 3.5454796719600520e-05
GC_9_608 b_9 NI_9 NS_608 0 8.6835399351779311e-05
GC_9_609 b_9 NI_9 NS_609 0 -4.6804733072841924e-06
GC_9_610 b_9 NI_9 NS_610 0 -7.5284268064295607e-07
GC_9_611 b_9 NI_9 NS_611 0 -5.7916195433411756e-06
GC_9_612 b_9 NI_9 NS_612 0 -4.3944524610906531e-06
GC_9_613 b_9 NI_9 NS_613 0 1.7500238311531857e-05
GC_9_614 b_9 NI_9 NS_614 0 -1.6580121941438681e-05
GC_9_615 b_9 NI_9 NS_615 0 -3.6993400938359115e-05
GC_9_616 b_9 NI_9 NS_616 0 1.7379742673017344e-05
GC_9_617 b_9 NI_9 NS_617 0 5.6746496340041475e-02
GC_9_618 b_9 NI_9 NS_618 0 -7.8728806715615371e-04
GC_9_619 b_9 NI_9 NS_619 0 -1.8256131036097404e-03
GC_9_620 b_9 NI_9 NS_620 0 2.2759316103577914e-03
GC_9_621 b_9 NI_9 NS_621 0 2.8300063910071762e-03
GC_9_622 b_9 NI_9 NS_622 0 2.3731408861818126e-04
GC_9_623 b_9 NI_9 NS_623 0 -5.2608056493072706e-03
GC_9_624 b_9 NI_9 NS_624 0 4.7288411081683750e-04
GC_9_625 b_9 NI_9 NS_625 0 -6.0836554097264293e-03
GC_9_626 b_9 NI_9 NS_626 0 1.0464821360319227e-02
GC_9_627 b_9 NI_9 NS_627 0 -6.3081003831909430e-04
GC_9_628 b_9 NI_9 NS_628 0 -8.4396225363583856e-05
GC_9_629 b_9 NI_9 NS_629 0 1.5620587675221783e-03
GC_9_630 b_9 NI_9 NS_630 0 -4.1083484927387313e-03
GC_9_631 b_9 NI_9 NS_631 0 8.2241960170820259e-04
GC_9_632 b_9 NI_9 NS_632 0 1.2136134837888446e-03
GC_9_633 b_9 NI_9 NS_633 0 -1.2742833565008250e-04
GC_9_634 b_9 NI_9 NS_634 0 8.2893525537435658e-04
GC_9_635 b_9 NI_9 NS_635 0 -5.5432921628288225e-03
GC_9_636 b_9 NI_9 NS_636 0 8.0374405703384987e-04
GC_9_637 b_9 NI_9 NS_637 0 -1.1589360712551038e-04
GC_9_638 b_9 NI_9 NS_638 0 -6.4086897278720043e-05
GC_9_639 b_9 NI_9 NS_639 0 7.6761035015287388e-04
GC_9_640 b_9 NI_9 NS_640 0 4.8048080279888706e-03
GC_9_641 b_9 NI_9 NS_641 0 -3.9895006231018855e-04
GC_9_642 b_9 NI_9 NS_642 0 -1.3836698107608415e-04
GC_9_643 b_9 NI_9 NS_643 0 -4.2774098817720371e-04
GC_9_644 b_9 NI_9 NS_644 0 1.5423701391438644e-05
GC_9_645 b_9 NI_9 NS_645 0 -3.9811863573486350e-04
GC_9_646 b_9 NI_9 NS_646 0 3.3411242004319490e-04
GC_9_647 b_9 NI_9 NS_647 0 -1.9656248381826882e-04
GC_9_648 b_9 NI_9 NS_648 0 -4.3232910920465931e-05
GC_9_649 b_9 NI_9 NS_649 0 -6.1049046588483096e-03
GC_9_650 b_9 NI_9 NS_650 0 -1.0187971846443351e-03
GC_9_651 b_9 NI_9 NS_651 0 -3.9046165132329755e-06
GC_9_652 b_9 NI_9 NS_652 0 2.6099896198696751e-05
GC_9_653 b_9 NI_9 NS_653 0 -2.1995136571248506e-04
GC_9_654 b_9 NI_9 NS_654 0 6.0948943844317777e-04
GC_9_655 b_9 NI_9 NS_655 0 -1.1170299443558733e-03
GC_9_656 b_9 NI_9 NS_656 0 -2.2107386660610634e-03
GC_9_657 b_9 NI_9 NS_657 0 5.7628822107779684e-05
GC_9_658 b_9 NI_9 NS_658 0 1.9491593307818287e-04
GC_9_659 b_9 NI_9 NS_659 0 2.2139502980485369e-06
GC_9_660 b_9 NI_9 NS_660 0 -3.0163817874773194e-07
GC_9_661 b_9 NI_9 NS_661 0 -1.6298160766423781e-06
GC_9_662 b_9 NI_9 NS_662 0 -6.1592170160813568e-06
GC_9_663 b_9 NI_9 NS_663 0 -5.4196328521911126e-05
GC_9_664 b_9 NI_9 NS_664 0 3.8239461185968447e-05
GC_9_665 b_9 NI_9 NS_665 0 3.9962968135579465e-07
GC_9_666 b_9 NI_9 NS_666 0 -8.7100510485647145e-06
GC_9_667 b_9 NI_9 NS_667 0 -9.5715923892600592e-07
GC_9_668 b_9 NI_9 NS_668 0 1.1465102965116001e-06
GC_9_669 b_9 NI_9 NS_669 0 6.2297045956049642e-06
GC_9_670 b_9 NI_9 NS_670 0 1.3998296308067613e-05
GC_9_671 b_9 NI_9 NS_671 0 -1.1852031610343953e-06
GC_9_672 b_9 NI_9 NS_672 0 -2.5956778430169536e-05
GD_9_1 b_9 NI_9 NA_1 0 -1.1601535750909230e-02
GD_9_2 b_9 NI_9 NA_2 0 -5.2820242332787977e-04
GD_9_3 b_9 NI_9 NA_3 0 -2.0309520865218159e-02
GD_9_4 b_9 NI_9 NA_4 0 -3.1807006864988225e-03
GD_9_5 b_9 NI_9 NA_5 0 -1.8740733839900259e-02
GD_9_6 b_9 NI_9 NA_6 0 5.6753650755863215e-05
GD_9_7 b_9 NI_9 NA_7 0 -7.4585849628671980e-04
GD_9_8 b_9 NI_9 NA_8 0 -1.1065509962177301e-02
GD_9_9 b_9 NI_9 NA_9 0 -1.7891309399444710e-01
GD_9_10 b_9 NI_9 NA_10 0 4.2603485398233089e-02
GD_9_11 b_9 NI_9 NA_11 0 -2.1712256038430095e-02
GD_9_12 b_9 NI_9 NA_12 0 -5.3530411270550825e-02
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 5.5660533841491418e-03
GC_10_2 b_10 NI_10 NS_2 0 -1.0145321138742508e-04
GC_10_3 b_10 NI_10 NS_3 0 1.9992950229114022e-04
GC_10_4 b_10 NI_10 NS_4 0 1.6140516246590521e-05
GC_10_5 b_10 NI_10 NS_5 0 1.0372911734711688e-04
GC_10_6 b_10 NI_10 NS_6 0 2.4325577023124706e-04
GC_10_7 b_10 NI_10 NS_7 0 -3.1611090393750187e-04
GC_10_8 b_10 NI_10 NS_8 0 1.2476672671575153e-03
GC_10_9 b_10 NI_10 NS_9 0 -1.7128848404921206e-03
GC_10_10 b_10 NI_10 NS_10 0 5.6251575511910578e-04
GC_10_11 b_10 NI_10 NS_11 0 3.8290556158678435e-04
GC_10_12 b_10 NI_10 NS_12 0 -9.3814592350347891e-04
GC_10_13 b_10 NI_10 NS_13 0 -5.3111055563115860e-04
GC_10_14 b_10 NI_10 NS_14 0 -1.0183091500540061e-03
GC_10_15 b_10 NI_10 NS_15 0 5.9511083819849936e-04
GC_10_16 b_10 NI_10 NS_16 0 -3.8076081417925034e-04
GC_10_17 b_10 NI_10 NS_17 0 1.3702353233691279e-03
GC_10_18 b_10 NI_10 NS_18 0 1.0770191555470802e-03
GC_10_19 b_10 NI_10 NS_19 0 -7.6306369664619420e-04
GC_10_20 b_10 NI_10 NS_20 0 2.2130015074527973e-03
GC_10_21 b_10 NI_10 NS_21 0 -2.1002614300629155e-04
GC_10_22 b_10 NI_10 NS_22 0 -2.7445049667442537e-06
GC_10_23 b_10 NI_10 NS_23 0 -2.8947164745079298e-03
GC_10_24 b_10 NI_10 NS_24 0 1.8290981455364595e-03
GC_10_25 b_10 NI_10 NS_25 0 3.4458234987822314e-04
GC_10_26 b_10 NI_10 NS_26 0 3.5811355743310279e-04
GC_10_27 b_10 NI_10 NS_27 0 -8.0098250863451851e-04
GC_10_28 b_10 NI_10 NS_28 0 8.1147455517372493e-05
GC_10_29 b_10 NI_10 NS_29 0 -5.4047661649025383e-04
GC_10_30 b_10 NI_10 NS_30 0 -1.0269537315857403e-04
GC_10_31 b_10 NI_10 NS_31 0 -8.9800300916865875e-05
GC_10_32 b_10 NI_10 NS_32 0 -5.5939958532665852e-05
GC_10_33 b_10 NI_10 NS_33 0 -1.2217264407971822e-03
GC_10_34 b_10 NI_10 NS_34 0 -5.7137305867599264e-03
GC_10_35 b_10 NI_10 NS_35 0 5.1376449979174775e-05
GC_10_36 b_10 NI_10 NS_36 0 -2.2848655436044756e-05
GC_10_37 b_10 NI_10 NS_37 0 -1.1269313238583809e-03
GC_10_38 b_10 NI_10 NS_38 0 4.1506642029952604e-04
GC_10_39 b_10 NI_10 NS_39 0 2.1247866607427483e-03
GC_10_40 b_10 NI_10 NS_40 0 4.3545860347734351e-04
GC_10_41 b_10 NI_10 NS_41 0 -8.8815121691411636e-05
GC_10_42 b_10 NI_10 NS_42 0 1.6625290195647769e-04
GC_10_43 b_10 NI_10 NS_43 0 -1.0222119359361018e-06
GC_10_44 b_10 NI_10 NS_44 0 1.2395205604994968e-06
GC_10_45 b_10 NI_10 NS_45 0 5.6207858849467538e-06
GC_10_46 b_10 NI_10 NS_46 0 -1.9364294416772242e-06
GC_10_47 b_10 NI_10 NS_47 0 -1.3162829318799312e-04
GC_10_48 b_10 NI_10 NS_48 0 -7.4360257118877905e-05
GC_10_49 b_10 NI_10 NS_49 0 1.7462363966871331e-05
GC_10_50 b_10 NI_10 NS_50 0 -2.1723022339134512e-06
GC_10_51 b_10 NI_10 NS_51 0 -6.0489143191562036e-06
GC_10_52 b_10 NI_10 NS_52 0 -1.1046712097869805e-05
GC_10_53 b_10 NI_10 NS_53 0 4.1274347070401510e-05
GC_10_54 b_10 NI_10 NS_54 0 4.4225436589831017e-05
GC_10_55 b_10 NI_10 NS_55 0 -4.3629130832453214e-05
GC_10_56 b_10 NI_10 NS_56 0 -7.7747881122419330e-05
GC_10_57 b_10 NI_10 NS_57 0 -4.8613628801506721e-03
GC_10_58 b_10 NI_10 NS_58 0 1.2504095849440632e-05
GC_10_59 b_10 NI_10 NS_59 0 -8.5592895262754423e-05
GC_10_60 b_10 NI_10 NS_60 0 8.1985214466439611e-05
GC_10_61 b_10 NI_10 NS_61 0 -1.5105019694403078e-04
GC_10_62 b_10 NI_10 NS_62 0 -5.6342206206565790e-05
GC_10_63 b_10 NI_10 NS_63 0 -3.4950084920877403e-04
GC_10_64 b_10 NI_10 NS_64 0 -8.4344312354502180e-04
GC_10_65 b_10 NI_10 NS_65 0 8.4168984435071593e-04
GC_10_66 b_10 NI_10 NS_66 0 -8.5660294286592524e-04
GC_10_67 b_10 NI_10 NS_67 0 -8.3025956914738527e-05
GC_10_68 b_10 NI_10 NS_68 0 -3.0335263408532017e-04
GC_10_69 b_10 NI_10 NS_69 0 -5.2232730692931221e-05
GC_10_70 b_10 NI_10 NS_70 0 -3.6360763275076303e-04
GC_10_71 b_10 NI_10 NS_71 0 2.5710647125130567e-04
GC_10_72 b_10 NI_10 NS_72 0 -4.3842628548458319e-04
GC_10_73 b_10 NI_10 NS_73 0 7.1113824972579836e-04
GC_10_74 b_10 NI_10 NS_74 0 2.6094297775498810e-04
GC_10_75 b_10 NI_10 NS_75 0 -9.1662656257207251e-04
GC_10_76 b_10 NI_10 NS_76 0 -6.4155290721422170e-04
GC_10_77 b_10 NI_10 NS_77 0 1.1410892663373651e-04
GC_10_78 b_10 NI_10 NS_78 0 5.8382742747880837e-05
GC_10_79 b_10 NI_10 NS_79 0 3.8663637365452313e-03
GC_10_80 b_10 NI_10 NS_80 0 -1.7525553831205356e-03
GC_10_81 b_10 NI_10 NS_81 0 -4.3608719419681622e-04
GC_10_82 b_10 NI_10 NS_82 0 3.2550078920480226e-04
GC_10_83 b_10 NI_10 NS_83 0 -3.1011544371377478e-04
GC_10_84 b_10 NI_10 NS_84 0 4.5865175709280487e-04
GC_10_85 b_10 NI_10 NS_85 0 -4.7654157987919698e-05
GC_10_86 b_10 NI_10 NS_86 0 -4.6737828820803910e-04
GC_10_87 b_10 NI_10 NS_87 0 1.8169937734188016e-04
GC_10_88 b_10 NI_10 NS_88 0 -1.7472912262263646e-05
GC_10_89 b_10 NI_10 NS_89 0 7.9546172492063233e-04
GC_10_90 b_10 NI_10 NS_90 0 4.7628415835837632e-03
GC_10_91 b_10 NI_10 NS_91 0 -1.0855606152508781e-04
GC_10_92 b_10 NI_10 NS_92 0 1.8723149207925744e-04
GC_10_93 b_10 NI_10 NS_93 0 1.6604547346932563e-03
GC_10_94 b_10 NI_10 NS_94 0 -8.3590331480051057e-04
GC_10_95 b_10 NI_10 NS_95 0 -3.1566913070130410e-03
GC_10_96 b_10 NI_10 NS_96 0 -1.3331616079306483e-03
GC_10_97 b_10 NI_10 NS_97 0 -5.1394661386954302e-04
GC_10_98 b_10 NI_10 NS_98 0 4.8358058258140592e-04
GC_10_99 b_10 NI_10 NS_99 0 5.2981377580906157e-06
GC_10_100 b_10 NI_10 NS_100 0 -5.9206901969538221e-06
GC_10_101 b_10 NI_10 NS_101 0 1.0611129974103056e-06
GC_10_102 b_10 NI_10 NS_102 0 6.1285182886358910e-05
GC_10_103 b_10 NI_10 NS_103 0 3.0114607946986246e-04
GC_10_104 b_10 NI_10 NS_104 0 -1.6904585293545996e-04
GC_10_105 b_10 NI_10 NS_105 0 4.7392356731498849e-05
GC_10_106 b_10 NI_10 NS_106 0 7.3875693362907948e-05
GC_10_107 b_10 NI_10 NS_107 0 1.1853743967778757e-05
GC_10_108 b_10 NI_10 NS_108 0 4.5739162550081268e-05
GC_10_109 b_10 NI_10 NS_109 0 1.7738831963387566e-04
GC_10_110 b_10 NI_10 NS_110 0 -1.9777833066233225e-04
GC_10_111 b_10 NI_10 NS_111 0 -3.1917549713487194e-04
GC_10_112 b_10 NI_10 NS_112 0 2.1291102533672150e-04
GC_10_113 b_10 NI_10 NS_113 0 8.0622616758051213e-03
GC_10_114 b_10 NI_10 NS_114 0 -1.5147958968021583e-04
GC_10_115 b_10 NI_10 NS_115 0 3.0541915684601027e-04
GC_10_116 b_10 NI_10 NS_116 0 1.6335775894027850e-04
GC_10_117 b_10 NI_10 NS_117 0 -7.9987552419010606e-05
GC_10_118 b_10 NI_10 NS_118 0 3.3356406188098098e-04
GC_10_119 b_10 NI_10 NS_119 0 -9.2575855701834567e-04
GC_10_120 b_10 NI_10 NS_120 0 1.2090068577250868e-03
GC_10_121 b_10 NI_10 NS_121 0 -1.5895623139254402e-03
GC_10_122 b_10 NI_10 NS_122 0 -3.8700471426989256e-04
GC_10_123 b_10 NI_10 NS_123 0 1.1951301586374245e-04
GC_10_124 b_10 NI_10 NS_124 0 -3.3159016631891837e-04
GC_10_125 b_10 NI_10 NS_125 0 6.1336311600065895e-06
GC_10_126 b_10 NI_10 NS_126 0 -1.5464995924787033e-03
GC_10_127 b_10 NI_10 NS_127 0 9.7343882697011747e-04
GC_10_128 b_10 NI_10 NS_128 0 -6.1912788012127200e-04
GC_10_129 b_10 NI_10 NS_129 0 1.9281476701832523e-03
GC_10_130 b_10 NI_10 NS_130 0 1.8630683813437776e-03
GC_10_131 b_10 NI_10 NS_131 0 -4.4927500656012572e-04
GC_10_132 b_10 NI_10 NS_132 0 2.7060367652638052e-03
GC_10_133 b_10 NI_10 NS_133 0 -3.2995533555218515e-04
GC_10_134 b_10 NI_10 NS_134 0 -2.9811296601054575e-05
GC_10_135 b_10 NI_10 NS_135 0 -2.4211673695565075e-03
GC_10_136 b_10 NI_10 NS_136 0 2.7066650125579764e-03
GC_10_137 b_10 NI_10 NS_137 0 3.2268182754199257e-04
GC_10_138 b_10 NI_10 NS_138 0 3.1889536375297634e-04
GC_10_139 b_10 NI_10 NS_139 0 -1.0964657468359763e-03
GC_10_140 b_10 NI_10 NS_140 0 2.9468117661316445e-04
GC_10_141 b_10 NI_10 NS_141 0 -7.2148819670719909e-04
GC_10_142 b_10 NI_10 NS_142 0 -1.8717931940941966e-05
GC_10_143 b_10 NI_10 NS_143 0 -1.2988785710843257e-04
GC_10_144 b_10 NI_10 NS_144 0 -6.6050004640677483e-05
GC_10_145 b_10 NI_10 NS_145 0 -7.5857983994717377e-04
GC_10_146 b_10 NI_10 NS_146 0 -5.5940445553688822e-03
GC_10_147 b_10 NI_10 NS_147 0 5.8518715740409734e-05
GC_10_148 b_10 NI_10 NS_148 0 -3.8795707393012613e-05
GC_10_149 b_10 NI_10 NS_149 0 -1.2958630157924856e-03
GC_10_150 b_10 NI_10 NS_150 0 5.4380859927564322e-04
GC_10_151 b_10 NI_10 NS_151 0 1.5320740886250312e-03
GC_10_152 b_10 NI_10 NS_152 0 -6.5140497969666251e-05
GC_10_153 b_10 NI_10 NS_153 0 -1.4958657324600039e-04
GC_10_154 b_10 NI_10 NS_154 0 1.8029244868930818e-04
GC_10_155 b_10 NI_10 NS_155 0 -9.0707459757462009e-07
GC_10_156 b_10 NI_10 NS_156 0 4.2021229901378245e-07
GC_10_157 b_10 NI_10 NS_157 0 6.0058677843125302e-06
GC_10_158 b_10 NI_10 NS_158 0 -2.4411451994410255e-06
GC_10_159 b_10 NI_10 NS_159 0 -8.8381023001191507e-05
GC_10_160 b_10 NI_10 NS_160 0 -1.9622247308033257e-05
GC_10_161 b_10 NI_10 NS_161 0 1.3051385205870293e-05
GC_10_162 b_10 NI_10 NS_162 0 -6.5008808585585442e-06
GC_10_163 b_10 NI_10 NS_163 0 -4.8254306562329737e-06
GC_10_164 b_10 NI_10 NS_164 0 -5.1549035295421951e-06
GC_10_165 b_10 NI_10 NS_165 0 2.1021661776715161e-05
GC_10_166 b_10 NI_10 NS_166 0 -9.2628863185413231e-06
GC_10_167 b_10 NI_10 NS_167 0 -4.0870480982445407e-05
GC_10_168 b_10 NI_10 NS_168 0 1.2329322906523544e-06
GC_10_169 b_10 NI_10 NS_169 0 -4.8220290292311325e-03
GC_10_170 b_10 NI_10 NS_170 0 8.1014462567925299e-06
GC_10_171 b_10 NI_10 NS_171 0 -1.8579110550175575e-04
GC_10_172 b_10 NI_10 NS_172 0 7.5669461402399181e-05
GC_10_173 b_10 NI_10 NS_173 0 -1.1905336900617859e-04
GC_10_174 b_10 NI_10 NS_174 0 -1.7175623636045688e-04
GC_10_175 b_10 NI_10 NS_175 0 4.4306678526276878e-05
GC_10_176 b_10 NI_10 NS_176 0 -1.0739952950735738e-03
GC_10_177 b_10 NI_10 NS_177 0 1.0894129461492665e-03
GC_10_178 b_10 NI_10 NS_178 0 -5.0462019154268231e-05
GC_10_179 b_10 NI_10 NS_179 0 -1.4218737152122806e-04
GC_10_180 b_10 NI_10 NS_180 0 7.4389031959595298e-05
GC_10_181 b_10 NI_10 NS_181 0 -4.1158124747239008e-04
GC_10_182 b_10 NI_10 NS_182 0 -3.2487793677007210e-04
GC_10_183 b_10 NI_10 NS_183 0 3.8850714071462410e-04
GC_10_184 b_10 NI_10 NS_184 0 -4.6949377487965710e-04
GC_10_185 b_10 NI_10 NS_185 0 2.0966579713584344e-04
GC_10_186 b_10 NI_10 NS_186 0 1.0461961465596862e-03
GC_10_187 b_10 NI_10 NS_187 0 -1.4394810726187745e-03
GC_10_188 b_10 NI_10 NS_188 0 -1.3501915266898655e-03
GC_10_189 b_10 NI_10 NS_189 0 1.2089471799873410e-04
GC_10_190 b_10 NI_10 NS_190 0 5.9695122355758822e-05
GC_10_191 b_10 NI_10 NS_191 0 3.7622566574743712e-03
GC_10_192 b_10 NI_10 NS_192 0 -2.2908599282019390e-03
GC_10_193 b_10 NI_10 NS_193 0 -4.7923894773763809e-04
GC_10_194 b_10 NI_10 NS_194 0 3.2762336628890142e-04
GC_10_195 b_10 NI_10 NS_195 0 -4.3239448104813655e-04
GC_10_196 b_10 NI_10 NS_196 0 4.7632357880416954e-04
GC_10_197 b_10 NI_10 NS_197 0 -4.9976557412876507e-05
GC_10_198 b_10 NI_10 NS_198 0 -5.0453787232201345e-04
GC_10_199 b_10 NI_10 NS_199 0 1.6528289762705796e-04
GC_10_200 b_10 NI_10 NS_200 0 -1.5927763877052739e-05
GC_10_201 b_10 NI_10 NS_201 0 1.7151528197471210e-03
GC_10_202 b_10 NI_10 NS_202 0 3.6008122969167942e-03
GC_10_203 b_10 NI_10 NS_203 0 -1.1146193223273622e-04
GC_10_204 b_10 NI_10 NS_204 0 1.7564959984266314e-04
GC_10_205 b_10 NI_10 NS_205 0 1.5058143802232132e-03
GC_10_206 b_10 NI_10 NS_206 0 -7.2804425506086475e-04
GC_10_207 b_10 NI_10 NS_207 0 -2.3375350693142756e-03
GC_10_208 b_10 NI_10 NS_208 0 -5.8274616820572461e-04
GC_10_209 b_10 NI_10 NS_209 0 -7.2179203897093918e-04
GC_10_210 b_10 NI_10 NS_210 0 5.0053665904037630e-04
GC_10_211 b_10 NI_10 NS_211 0 4.8217365205917011e-06
GC_10_212 b_10 NI_10 NS_212 0 -4.3372150851098637e-06
GC_10_213 b_10 NI_10 NS_213 0 -1.1612599990639485e-06
GC_10_214 b_10 NI_10 NS_214 0 5.5955075002346411e-05
GC_10_215 b_10 NI_10 NS_215 0 2.2287175037153677e-04
GC_10_216 b_10 NI_10 NS_216 0 -1.5966784911227491e-04
GC_10_217 b_10 NI_10 NS_217 0 4.8453017270881900e-05
GC_10_218 b_10 NI_10 NS_218 0 7.3424305143455134e-05
GC_10_219 b_10 NI_10 NS_219 0 7.1263624059392596e-06
GC_10_220 b_10 NI_10 NS_220 0 3.8255164872392118e-05
GC_10_221 b_10 NI_10 NS_221 0 2.1947760902536899e-04
GC_10_222 b_10 NI_10 NS_222 0 -1.6130824447482692e-04
GC_10_223 b_10 NI_10 NS_223 0 -3.6770304792313403e-04
GC_10_224 b_10 NI_10 NS_224 0 1.3817210153535076e-04
GC_10_225 b_10 NI_10 NS_225 0 4.2544668957390647e-03
GC_10_226 b_10 NI_10 NS_226 0 -1.5443046706477525e-04
GC_10_227 b_10 NI_10 NS_227 0 2.7491875380062134e-04
GC_10_228 b_10 NI_10 NS_228 0 4.0106081381715685e-04
GC_10_229 b_10 NI_10 NS_229 0 -4.0779553367940218e-04
GC_10_230 b_10 NI_10 NS_230 0 2.2118047267551710e-04
GC_10_231 b_10 NI_10 NS_231 0 -1.4752092672480198e-03
GC_10_232 b_10 NI_10 NS_232 0 2.6979182414096171e-04
GC_10_233 b_10 NI_10 NS_233 0 -2.0291881528233444e-04
GC_10_234 b_10 NI_10 NS_234 0 -1.5814109058509610e-03
GC_10_235 b_10 NI_10 NS_235 0 2.1029624195738090e-04
GC_10_236 b_10 NI_10 NS_236 0 -2.8561516050463901e-04
GC_10_237 b_10 NI_10 NS_237 0 7.6273789845787763e-04
GC_10_238 b_10 NI_10 NS_238 0 -1.3190960804602687e-03
GC_10_239 b_10 NI_10 NS_239 0 1.0559651510437199e-03
GC_10_240 b_10 NI_10 NS_240 0 -6.1186043302765354e-04
GC_10_241 b_10 NI_10 NS_241 0 1.8188896722741326e-03
GC_10_242 b_10 NI_10 NS_242 0 2.1969489463265156e-03
GC_10_243 b_10 NI_10 NS_243 0 2.8228820553654495e-05
GC_10_244 b_10 NI_10 NS_244 0 3.0156984663808630e-03
GC_10_245 b_10 NI_10 NS_245 0 -3.6209655729798701e-04
GC_10_246 b_10 NI_10 NS_246 0 -2.8807158249186701e-05
GC_10_247 b_10 NI_10 NS_247 0 -2.9489487948136032e-03
GC_10_248 b_10 NI_10 NS_248 0 2.7203785654799592e-03
GC_10_249 b_10 NI_10 NS_249 0 3.0308276310628133e-04
GC_10_250 b_10 NI_10 NS_250 0 1.2537071708762024e-04
GC_10_251 b_10 NI_10 NS_251 0 -1.1205660743597004e-03
GC_10_252 b_10 NI_10 NS_252 0 2.2777945632477533e-04
GC_10_253 b_10 NI_10 NS_253 0 -6.5935645526795511e-04
GC_10_254 b_10 NI_10 NS_254 0 -2.4125327041817246e-05
GC_10_255 b_10 NI_10 NS_255 0 -1.4276108105344289e-04
GC_10_256 b_10 NI_10 NS_256 0 -5.0736650302135197e-05
GC_10_257 b_10 NI_10 NS_257 0 -9.6744724005030306e-05
GC_10_258 b_10 NI_10 NS_258 0 -4.7231635945798071e-03
GC_10_259 b_10 NI_10 NS_259 0 4.2607035722476789e-05
GC_10_260 b_10 NI_10 NS_260 0 -3.7792238035519721e-05
GC_10_261 b_10 NI_10 NS_261 0 -1.3105691515015614e-03
GC_10_262 b_10 NI_10 NS_262 0 5.5786216832412895e-04
GC_10_263 b_10 NI_10 NS_263 0 1.3155187617906023e-03
GC_10_264 b_10 NI_10 NS_264 0 -9.1643286886471575e-04
GC_10_265 b_10 NI_10 NS_265 0 -2.0428730230636889e-04
GC_10_266 b_10 NI_10 NS_266 0 8.0900192290151536e-05
GC_10_267 b_10 NI_10 NS_267 0 -7.7688516861417016e-07
GC_10_268 b_10 NI_10 NS_268 0 4.5650177089890340e-07
GC_10_269 b_10 NI_10 NS_269 0 -3.7809858369163979e-06
GC_10_270 b_10 NI_10 NS_270 0 -3.8835458510850266e-06
GC_10_271 b_10 NI_10 NS_271 0 -1.4841467840912970e-05
GC_10_272 b_10 NI_10 NS_272 0 6.4721694250020109e-05
GC_10_273 b_10 NI_10 NS_273 0 -9.0379234276162638e-06
GC_10_274 b_10 NI_10 NS_274 0 -5.8936089069025988e-06
GC_10_275 b_10 NI_10 NS_275 0 -4.7958612919943646e-06
GC_10_276 b_10 NI_10 NS_276 0 -4.4997406697654547e-06
GC_10_277 b_10 NI_10 NS_277 0 2.5692452596864863e-05
GC_10_278 b_10 NI_10 NS_278 0 -4.7797270673943372e-06
GC_10_279 b_10 NI_10 NS_279 0 -3.9493385349447003e-05
GC_10_280 b_10 NI_10 NS_280 0 -5.0474370657362582e-06
GC_10_281 b_10 NI_10 NS_281 0 3.2475988589142536e-04
GC_10_282 b_10 NI_10 NS_282 0 -3.0980755351694365e-05
GC_10_283 b_10 NI_10 NS_283 0 -2.7049335834396178e-04
GC_10_284 b_10 NI_10 NS_284 0 3.0755494882822207e-07
GC_10_285 b_10 NI_10 NS_285 0 5.7804873432796166e-05
GC_10_286 b_10 NI_10 NS_286 0 -2.5250137170579242e-04
GC_10_287 b_10 NI_10 NS_287 0 7.7777544805290031e-04
GC_10_288 b_10 NI_10 NS_288 0 -7.3612716011788721e-04
GC_10_289 b_10 NI_10 NS_289 0 6.0068956357493743e-04
GC_10_290 b_10 NI_10 NS_290 0 1.5362306355457273e-03
GC_10_291 b_10 NI_10 NS_291 0 -4.4887833616584564e-04
GC_10_292 b_10 NI_10 NS_292 0 4.9316877858661596e-04
GC_10_293 b_10 NI_10 NS_293 0 -9.5111009758647137e-04
GC_10_294 b_10 NI_10 NS_294 0 -4.1093769777995041e-04
GC_10_295 b_10 NI_10 NS_295 0 4.4685531535609033e-04
GC_10_296 b_10 NI_10 NS_296 0 -5.0679412967351138e-04
GC_10_297 b_10 NI_10 NS_297 0 -1.6899424812046789e-04
GC_10_298 b_10 NI_10 NS_298 0 1.7756182987470760e-03
GC_10_299 b_10 NI_10 NS_299 0 -1.5595263523983044e-03
GC_10_300 b_10 NI_10 NS_300 0 -1.6134266411166815e-03
GC_10_301 b_10 NI_10 NS_301 0 1.9758872463830182e-04
GC_10_302 b_10 NI_10 NS_302 0 2.2939891002988677e-05
GC_10_303 b_10 NI_10 NS_303 0 3.0621028333165305e-03
GC_10_304 b_10 NI_10 NS_304 0 -2.6507979605367624e-03
GC_10_305 b_10 NI_10 NS_305 0 -4.6323500928067236e-04
GC_10_306 b_10 NI_10 NS_306 0 4.3061304152795853e-04
GC_10_307 b_10 NI_10 NS_307 0 -5.2546504666825609e-04
GC_10_308 b_10 NI_10 NS_308 0 6.0746583774074934e-04
GC_10_309 b_10 NI_10 NS_309 0 -2.1664565743840443e-04
GC_10_310 b_10 NI_10 NS_310 0 -7.3814588940984455e-04
GC_10_311 b_10 NI_10 NS_311 0 2.6808936304539567e-04
GC_10_312 b_10 NI_10 NS_312 0 -8.4522447808540603e-05
GC_10_313 b_10 NI_10 NS_313 0 1.7585085945195384e-03
GC_10_314 b_10 NI_10 NS_314 0 4.3790216031834714e-03
GC_10_315 b_10 NI_10 NS_315 0 -1.2295043446659763e-04
GC_10_316 b_10 NI_10 NS_316 0 2.5274194493517466e-04
GC_10_317 b_10 NI_10 NS_317 0 1.9986443681637728e-03
GC_10_318 b_10 NI_10 NS_318 0 -1.1613514529600489e-03
GC_10_319 b_10 NI_10 NS_319 0 -2.3427737692953933e-03
GC_10_320 b_10 NI_10 NS_320 0 -1.0191935614002133e-03
GC_10_321 b_10 NI_10 NS_321 0 -8.3276574332143659e-04
GC_10_322 b_10 NI_10 NS_322 0 7.8983909183194599e-04
GC_10_323 b_10 NI_10 NS_323 0 4.1005859113086474e-06
GC_10_324 b_10 NI_10 NS_324 0 -1.0082129638827108e-05
GC_10_325 b_10 NI_10 NS_325 0 1.1896386455780984e-05
GC_10_326 b_10 NI_10 NS_326 0 7.5866838301205344e-05
GC_10_327 b_10 NI_10 NS_327 0 1.7878025274319177e-04
GC_10_328 b_10 NI_10 NS_328 0 -2.5847034722342532e-04
GC_10_329 b_10 NI_10 NS_329 0 9.2186020446311258e-05
GC_10_330 b_10 NI_10 NS_330 0 8.6736325376847404e-05
GC_10_331 b_10 NI_10 NS_331 0 1.5660615008542640e-05
GC_10_332 b_10 NI_10 NS_332 0 5.3836253128710996e-05
GC_10_333 b_10 NI_10 NS_333 0 3.2767425826198013e-04
GC_10_334 b_10 NI_10 NS_334 0 -3.1004316323493878e-04
GC_10_335 b_10 NI_10 NS_335 0 -5.8095040744614269e-04
GC_10_336 b_10 NI_10 NS_336 0 2.9966114667734811e-04
GC_10_337 b_10 NI_10 NS_337 0 9.1985770989343827e-03
GC_10_338 b_10 NI_10 NS_338 0 -1.0820501378981644e-04
GC_10_339 b_10 NI_10 NS_339 0 -1.6063129023330083e-04
GC_10_340 b_10 NI_10 NS_340 0 7.1864938050028853e-04
GC_10_341 b_10 NI_10 NS_341 0 -3.0035343932252628e-04
GC_10_342 b_10 NI_10 NS_342 0 -6.6812393559638364e-04
GC_10_343 b_10 NI_10 NS_343 0 -5.3910156607370934e-04
GC_10_344 b_10 NI_10 NS_344 0 -6.6289476589821272e-04
GC_10_345 b_10 NI_10 NS_345 0 2.2077767129614870e-03
GC_10_346 b_10 NI_10 NS_346 0 8.7822518735301966e-04
GC_10_347 b_10 NI_10 NS_347 0 -5.8618430119410363e-04
GC_10_348 b_10 NI_10 NS_348 0 -6.0962253891542498e-05
GC_10_349 b_10 NI_10 NS_349 0 5.0516146836935693e-04
GC_10_350 b_10 NI_10 NS_350 0 -5.4384456051354403e-04
GC_10_351 b_10 NI_10 NS_351 0 1.0216386658711484e-03
GC_10_352 b_10 NI_10 NS_352 0 -1.8622408191131131e-04
GC_10_353 b_10 NI_10 NS_353 0 9.0450363067688265e-04
GC_10_354 b_10 NI_10 NS_354 0 2.4153264421864760e-03
GC_10_355 b_10 NI_10 NS_355 0 -1.3445721143414773e-03
GC_10_356 b_10 NI_10 NS_356 0 2.8634763232447845e-03
GC_10_357 b_10 NI_10 NS_357 0 -2.7446836934943297e-04
GC_10_358 b_10 NI_10 NS_358 0 -7.7418457258289199e-05
GC_10_359 b_10 NI_10 NS_359 0 -7.8717474944907623e-04
GC_10_360 b_10 NI_10 NS_360 0 1.9332009858715807e-03
GC_10_361 b_10 NI_10 NS_361 0 8.3349822201453383e-05
GC_10_362 b_10 NI_10 NS_362 0 -4.1723557272445942e-05
GC_10_363 b_10 NI_10 NS_363 0 -7.6069469408929149e-04
GC_10_364 b_10 NI_10 NS_364 0 2.5886898945015537e-04
GC_10_365 b_10 NI_10 NS_365 0 -4.9253576842028313e-04
GC_10_366 b_10 NI_10 NS_366 0 9.6951372476780594e-05
GC_10_367 b_10 NI_10 NS_367 0 -1.2771378812158357e-04
GC_10_368 b_10 NI_10 NS_368 0 -3.2309038683276300e-05
GC_10_369 b_10 NI_10 NS_369 0 -1.4100993532130666e-03
GC_10_370 b_10 NI_10 NS_370 0 -2.8958206540550748e-03
GC_10_371 b_10 NI_10 NS_371 0 3.0377894405023122e-05
GC_10_372 b_10 NI_10 NS_372 0 -2.9095056493557884e-05
GC_10_373 b_10 NI_10 NS_373 0 -8.3607874690891826e-04
GC_10_374 b_10 NI_10 NS_374 0 5.5527328898686331e-04
GC_10_375 b_10 NI_10 NS_375 0 1.1176247829536605e-03
GC_10_376 b_10 NI_10 NS_376 0 -2.8919811407268072e-04
GC_10_377 b_10 NI_10 NS_377 0 -1.0514581613634938e-04
GC_10_378 b_10 NI_10 NS_378 0 1.5838089721760410e-04
GC_10_379 b_10 NI_10 NS_379 0 -1.9868375409847965e-06
GC_10_380 b_10 NI_10 NS_380 0 2.5378489837188006e-06
GC_10_381 b_10 NI_10 NS_381 0 -2.0655322968412818e-06
GC_10_382 b_10 NI_10 NS_382 0 -3.9515092409097319e-06
GC_10_383 b_10 NI_10 NS_383 0 -4.8380755288547059e-05
GC_10_384 b_10 NI_10 NS_384 0 7.0574630662517535e-05
GC_10_385 b_10 NI_10 NS_385 0 2.3995859699921501e-06
GC_10_386 b_10 NI_10 NS_386 0 -1.0993444398803190e-05
GC_10_387 b_10 NI_10 NS_387 0 -1.9735405225393076e-06
GC_10_388 b_10 NI_10 NS_388 0 -4.9972427498032381e-06
GC_10_389 b_10 NI_10 NS_389 0 2.4599797672478257e-05
GC_10_390 b_10 NI_10 NS_390 0 -4.1451023789747394e-05
GC_10_391 b_10 NI_10 NS_391 0 -4.9294270682877160e-05
GC_10_392 b_10 NI_10 NS_392 0 5.5827426882194116e-05
GC_10_393 b_10 NI_10 NS_393 0 -3.3963333878714850e-03
GC_10_394 b_10 NI_10 NS_394 0 -1.3409448314771256e-04
GC_10_395 b_10 NI_10 NS_395 0 -3.0684957325263258e-04
GC_10_396 b_10 NI_10 NS_396 0 -2.2206889072041389e-04
GC_10_397 b_10 NI_10 NS_397 0 3.3254355225314066e-04
GC_10_398 b_10 NI_10 NS_398 0 8.2569294913938812e-05
GC_10_399 b_10 NI_10 NS_399 0 6.5238648451375857e-04
GC_10_400 b_10 NI_10 NS_400 0 2.7949118117199303e-04
GC_10_401 b_10 NI_10 NS_401 0 -2.3645459689352164e-03
GC_10_402 b_10 NI_10 NS_402 0 7.6659522928217594e-04
GC_10_403 b_10 NI_10 NS_403 0 2.3459978023441039e-04
GC_10_404 b_10 NI_10 NS_404 0 1.5568595333633264e-04
GC_10_405 b_10 NI_10 NS_405 0 -4.6490198111620503e-04
GC_10_406 b_10 NI_10 NS_406 0 -1.4673840308627780e-03
GC_10_407 b_10 NI_10 NS_407 0 3.4673195161804898e-04
GC_10_408 b_10 NI_10 NS_408 0 -2.4201800443309914e-04
GC_10_409 b_10 NI_10 NS_409 0 -8.6843612685103975e-04
GC_10_410 b_10 NI_10 NS_410 0 7.1309991645816047e-04
GC_10_411 b_10 NI_10 NS_411 0 -1.0605230007730464e-03
GC_10_412 b_10 NI_10 NS_412 0 -1.3650763921791180e-03
GC_10_413 b_10 NI_10 NS_413 0 1.1836651280650772e-04
GC_10_414 b_10 NI_10 NS_414 0 5.2362338727465487e-05
GC_10_415 b_10 NI_10 NS_415 0 2.0728416496440306e-03
GC_10_416 b_10 NI_10 NS_416 0 -3.7917014302686234e-03
GC_10_417 b_10 NI_10 NS_417 0 -3.1234729205303549e-04
GC_10_418 b_10 NI_10 NS_418 0 3.6359294260374689e-04
GC_10_419 b_10 NI_10 NS_419 0 -2.6722982926290028e-04
GC_10_420 b_10 NI_10 NS_420 0 2.7061718008929131e-04
GC_10_421 b_10 NI_10 NS_421 0 -5.8007784594856229e-05
GC_10_422 b_10 NI_10 NS_422 0 -5.2675396282657870e-04
GC_10_423 b_10 NI_10 NS_423 0 1.9021966028286751e-04
GC_10_424 b_10 NI_10 NS_424 0 -6.0137246334221606e-05
GC_10_425 b_10 NI_10 NS_425 0 1.2205496797781609e-03
GC_10_426 b_10 NI_10 NS_426 0 1.6796172339911505e-03
GC_10_427 b_10 NI_10 NS_427 0 -1.0133682474313649e-04
GC_10_428 b_10 NI_10 NS_428 0 1.0806259809567410e-04
GC_10_429 b_10 NI_10 NS_429 0 1.2612841702429277e-03
GC_10_430 b_10 NI_10 NS_430 0 -6.3848484973859669e-04
GC_10_431 b_10 NI_10 NS_431 0 1.0559170600027212e-04
GC_10_432 b_10 NI_10 NS_432 0 3.4003695713591056e-04
GC_10_433 b_10 NI_10 NS_433 0 -5.0106875083994298e-04
GC_10_434 b_10 NI_10 NS_434 0 3.8825309279326127e-04
GC_10_435 b_10 NI_10 NS_435 0 6.5613236486231621e-07
GC_10_436 b_10 NI_10 NS_436 0 -4.6184345407669825e-06
GC_10_437 b_10 NI_10 NS_437 0 -1.1951247214626264e-07
GC_10_438 b_10 NI_10 NS_438 0 3.3216378748157079e-05
GC_10_439 b_10 NI_10 NS_439 0 2.6899497867644143e-05
GC_10_440 b_10 NI_10 NS_440 0 -1.6963389710666901e-04
GC_10_441 b_10 NI_10 NS_441 0 4.5553460775726618e-05
GC_10_442 b_10 NI_10 NS_442 0 4.8639987449238011e-05
GC_10_443 b_10 NI_10 NS_443 0 4.6997769517277625e-06
GC_10_444 b_10 NI_10 NS_444 0 1.7341739637790175e-05
GC_10_445 b_10 NI_10 NS_445 0 2.3750597745191807e-04
GC_10_446 b_10 NI_10 NS_446 0 -1.0737598510306202e-04
GC_10_447 b_10 NI_10 NS_447 0 -3.7730814788134863e-04
GC_10_448 b_10 NI_10 NS_448 0 5.7521953639500945e-05
GC_10_449 b_10 NI_10 NS_449 0 -4.5487796352469717e-02
GC_10_450 b_10 NI_10 NS_450 0 1.2148228660622947e-02
GC_10_451 b_10 NI_10 NS_451 0 -2.9338491313903262e-03
GC_10_452 b_10 NI_10 NS_452 0 3.7223078412648770e-03
GC_10_453 b_10 NI_10 NS_453 0 -4.3639025693651603e-03
GC_10_454 b_10 NI_10 NS_454 0 2.1017782713832504e-03
GC_10_455 b_10 NI_10 NS_455 0 -4.7808389670266948e-03
GC_10_456 b_10 NI_10 NS_456 0 -9.2825516534799177e-03
GC_10_457 b_10 NI_10 NS_457 0 -2.4143535034039910e-03
GC_10_458 b_10 NI_10 NS_458 0 -9.2045340358214607e-03
GC_10_459 b_10 NI_10 NS_459 0 4.6184473684863153e-04
GC_10_460 b_10 NI_10 NS_460 0 1.6663514009215927e-04
GC_10_461 b_10 NI_10 NS_461 0 7.2088874857509921e-03
GC_10_462 b_10 NI_10 NS_462 0 -1.5917336433372068e-03
GC_10_463 b_10 NI_10 NS_463 0 1.5076664056002829e-03
GC_10_464 b_10 NI_10 NS_464 0 1.2646463673094824e-03
GC_10_465 b_10 NI_10 NS_465 0 5.5694862594595964e-03
GC_10_466 b_10 NI_10 NS_466 0 8.2374936308513545e-04
GC_10_467 b_10 NI_10 NS_467 0 -2.3798214792909414e-03
GC_10_468 b_10 NI_10 NS_468 0 1.1646685864811872e-03
GC_10_469 b_10 NI_10 NS_469 0 -3.7364946906528362e-04
GC_10_470 b_10 NI_10 NS_470 0 6.8805461772328887e-05
GC_10_471 b_10 NI_10 NS_471 0 7.9978305804297156e-03
GC_10_472 b_10 NI_10 NS_472 0 -2.7376528324836724e-03
GC_10_473 b_10 NI_10 NS_473 0 -1.7443061658775809e-03
GC_10_474 b_10 NI_10 NS_474 0 -2.4148591878878221e-05
GC_10_475 b_10 NI_10 NS_475 0 -2.8142285364354352e-04
GC_10_476 b_10 NI_10 NS_476 0 1.2194196255368447e-04
GC_10_477 b_10 NI_10 NS_477 0 -4.5359873834408129e-04
GC_10_478 b_10 NI_10 NS_478 0 3.9177316353436876e-04
GC_10_479 b_10 NI_10 NS_479 0 -2.9623790450584081e-04
GC_10_480 b_10 NI_10 NS_480 0 -1.2279932372078259e-04
GC_10_481 b_10 NI_10 NS_481 0 3.0255442046472174e-03
GC_10_482 b_10 NI_10 NS_482 0 -6.4864083203891370e-04
GC_10_483 b_10 NI_10 NS_483 0 -2.6897399974606204e-05
GC_10_484 b_10 NI_10 NS_484 0 1.7986425700651577e-04
GC_10_485 b_10 NI_10 NS_485 0 -9.3160705693325551e-04
GC_10_486 b_10 NI_10 NS_486 0 -9.7637406028076976e-04
GC_10_487 b_10 NI_10 NS_487 0 1.8590623756186868e-03
GC_10_488 b_10 NI_10 NS_488 0 1.6027031518604153e-03
GC_10_489 b_10 NI_10 NS_489 0 -1.2831012875612403e-04
GC_10_490 b_10 NI_10 NS_490 0 -1.7211462906089873e-04
GC_10_491 b_10 NI_10 NS_491 0 1.6045233974689146e-06
GC_10_492 b_10 NI_10 NS_492 0 -2.1324659601838096e-06
GC_10_493 b_10 NI_10 NS_493 0 3.7688557184455496e-06
GC_10_494 b_10 NI_10 NS_494 0 -1.9773669689927742e-06
GC_10_495 b_10 NI_10 NS_495 0 -6.8083975012517696e-05
GC_10_496 b_10 NI_10 NS_496 0 -8.9521503356245193e-05
GC_10_497 b_10 NI_10 NS_497 0 9.4196724112200547e-06
GC_10_498 b_10 NI_10 NS_498 0 4.0979500173139212e-06
GC_10_499 b_10 NI_10 NS_499 0 2.4615715259327533e-06
GC_10_500 b_10 NI_10 NS_500 0 -1.1024984342044325e-05
GC_10_501 b_10 NI_10 NS_501 0 2.6530205701270414e-05
GC_10_502 b_10 NI_10 NS_502 0 6.1448239003678162e-05
GC_10_503 b_10 NI_10 NS_503 0 -1.0121360653554940e-05
GC_10_504 b_10 NI_10 NS_504 0 -1.0469942576147917e-04
GC_10_505 b_10 NI_10 NS_505 0 -7.0032339542678637e-02
GC_10_506 b_10 NI_10 NS_506 0 7.7264337451599394e-03
GC_10_507 b_10 NI_10 NS_507 0 -1.1547515523642263e-03
GC_10_508 b_10 NI_10 NS_508 0 -1.9316721952989057e-03
GC_10_509 b_10 NI_10 NS_509 0 5.4897070836686560e-05
GC_10_510 b_10 NI_10 NS_510 0 -1.5219944999826176e-03
GC_10_511 b_10 NI_10 NS_511 0 6.0551906648040220e-03
GC_10_512 b_10 NI_10 NS_512 0 3.8808489535665856e-03
GC_10_513 b_10 NI_10 NS_513 0 3.4825812148877753e-03
GC_10_514 b_10 NI_10 NS_514 0 6.4001220165893777e-03
GC_10_515 b_10 NI_10 NS_515 0 3.4976086349794791e-04
GC_10_516 b_10 NI_10 NS_516 0 -3.6871371666580293e-04
GC_10_517 b_10 NI_10 NS_517 0 -1.7150147931642172e-03
GC_10_518 b_10 NI_10 NS_518 0 -5.5367257063207624e-03
GC_10_519 b_10 NI_10 NS_519 0 1.2139242201110656e-03
GC_10_520 b_10 NI_10 NS_520 0 6.0894741863111999e-04
GC_10_521 b_10 NI_10 NS_521 0 6.1928415428136329e-04
GC_10_522 b_10 NI_10 NS_522 0 6.8970506338981009e-04
GC_10_523 b_10 NI_10 NS_523 0 2.1629083614137408e-03
GC_10_524 b_10 NI_10 NS_524 0 -2.5960251056557971e-03
GC_10_525 b_10 NI_10 NS_525 0 1.4848436502291242e-04
GC_10_526 b_10 NI_10 NS_526 0 -7.0479501048348428e-05
GC_10_527 b_10 NI_10 NS_527 0 1.9366952635722274e-03
GC_10_528 b_10 NI_10 NS_528 0 5.4205079645468154e-03
GC_10_529 b_10 NI_10 NS_529 0 4.8203131486403503e-04
GC_10_530 b_10 NI_10 NS_530 0 6.9304132430641971e-06
GC_10_531 b_10 NI_10 NS_531 0 -4.1745366339802681e-04
GC_10_532 b_10 NI_10 NS_532 0 6.6932707621063012e-05
GC_10_533 b_10 NI_10 NS_533 0 1.0578672007219452e-04
GC_10_534 b_10 NI_10 NS_534 0 -3.3411627256307999e-04
GC_10_535 b_10 NI_10 NS_535 0 4.5513092086648603e-04
GC_10_536 b_10 NI_10 NS_536 0 -2.0995874167543523e-04
GC_10_537 b_10 NI_10 NS_537 0 -2.0167511321573569e-02
GC_10_538 b_10 NI_10 NS_538 0 2.4864864043547693e-03
GC_10_539 b_10 NI_10 NS_539 0 -3.0109873114080737e-04
GC_10_540 b_10 NI_10 NS_540 0 -3.8039947574534716e-04
GC_10_541 b_10 NI_10 NS_541 0 6.2539489247624130e-03
GC_10_542 b_10 NI_10 NS_542 0 2.0711391879524510e-03
GC_10_543 b_10 NI_10 NS_543 0 9.2169888595222890e-03
GC_10_544 b_10 NI_10 NS_544 0 -5.9759043499543491e-03
GC_10_545 b_10 NI_10 NS_545 0 1.5247510664135216e-03
GC_10_546 b_10 NI_10 NS_546 0 4.8302720997836474e-04
GC_10_547 b_10 NI_10 NS_547 0 -3.7560224748666402e-06
GC_10_548 b_10 NI_10 NS_548 0 -5.6092195610710997e-06
GC_10_549 b_10 NI_10 NS_549 0 -5.8644457917325555e-05
GC_10_550 b_10 NI_10 NS_550 0 -3.1303239357249781e-05
GC_10_551 b_10 NI_10 NS_551 0 -3.7524376844588032e-04
GC_10_552 b_10 NI_10 NS_552 0 1.9811236300446128e-04
GC_10_553 b_10 NI_10 NS_553 0 -6.4557521438444668e-05
GC_10_554 b_10 NI_10 NS_554 0 -3.3901755313040594e-05
GC_10_555 b_10 NI_10 NS_555 0 -6.6099636867311212e-05
GC_10_556 b_10 NI_10 NS_556 0 -2.7599238201845731e-05
GC_10_557 b_10 NI_10 NS_557 0 4.3735307367133035e-04
GC_10_558 b_10 NI_10 NS_558 0 -4.1081737492961785e-04
GC_10_559 b_10 NI_10 NS_559 0 -8.0594051616109650e-04
GC_10_560 b_10 NI_10 NS_560 0 3.9693329043397654e-04
GC_10_561 b_10 NI_10 NS_561 0 5.7434285216554325e-02
GC_10_562 b_10 NI_10 NS_562 0 -7.8096423303067135e-04
GC_10_563 b_10 NI_10 NS_563 0 -1.7649582837868908e-03
GC_10_564 b_10 NI_10 NS_564 0 2.3941417913815517e-03
GC_10_565 b_10 NI_10 NS_565 0 2.8812338170611834e-03
GC_10_566 b_10 NI_10 NS_566 0 2.6566787309148033e-04
GC_10_567 b_10 NI_10 NS_567 0 -5.6069433122297894e-03
GC_10_568 b_10 NI_10 NS_568 0 4.9244666721707728e-04
GC_10_569 b_10 NI_10 NS_569 0 -6.3581741134312569e-03
GC_10_570 b_10 NI_10 NS_570 0 1.0169290054741247e-02
GC_10_571 b_10 NI_10 NS_571 0 -7.6138103010757344e-04
GC_10_572 b_10 NI_10 NS_572 0 3.0400926107607980e-05
GC_10_573 b_10 NI_10 NS_573 0 1.9032017236546908e-03
GC_10_574 b_10 NI_10 NS_574 0 -4.4859297146334666e-03
GC_10_575 b_10 NI_10 NS_575 0 1.0553095129953902e-03
GC_10_576 b_10 NI_10 NS_576 0 1.3589755216437936e-03
GC_10_577 b_10 NI_10 NS_577 0 -9.0134658970031209e-06
GC_10_578 b_10 NI_10 NS_578 0 1.1728772907548520e-03
GC_10_579 b_10 NI_10 NS_579 0 -5.8436637079250179e-03
GC_10_580 b_10 NI_10 NS_580 0 9.4976866331969705e-04
GC_10_581 b_10 NI_10 NS_581 0 -1.5340828563586628e-04
GC_10_582 b_10 NI_10 NS_582 0 -8.1534168087330251e-05
GC_10_583 b_10 NI_10 NS_583 0 1.2920501835578125e-03
GC_10_584 b_10 NI_10 NS_584 0 5.2330587846349703e-03
GC_10_585 b_10 NI_10 NS_585 0 -4.9894056287758213e-04
GC_10_586 b_10 NI_10 NS_586 0 -1.8074639022476227e-04
GC_10_587 b_10 NI_10 NS_587 0 -5.0411159345730891e-04
GC_10_588 b_10 NI_10 NS_588 0 7.6264330709567777e-05
GC_10_589 b_10 NI_10 NS_589 0 -4.5612509097745277e-04
GC_10_590 b_10 NI_10 NS_590 0 4.4236381567471102e-04
GC_10_591 b_10 NI_10 NS_591 0 -2.4602366516808028e-04
GC_10_592 b_10 NI_10 NS_592 0 -4.8690735916362865e-05
GC_10_593 b_10 NI_10 NS_593 0 -7.5535675398475059e-03
GC_10_594 b_10 NI_10 NS_594 0 -1.5776459721931612e-03
GC_10_595 b_10 NI_10 NS_595 0 -2.0328255694817244e-05
GC_10_596 b_10 NI_10 NS_596 0 4.2794299386370916e-05
GC_10_597 b_10 NI_10 NS_597 0 -9.0318469653142695e-05
GC_10_598 b_10 NI_10 NS_598 0 6.4024157100633200e-04
GC_10_599 b_10 NI_10 NS_599 0 -1.6179958643791574e-04
GC_10_600 b_10 NI_10 NS_600 0 -2.5374174946464147e-03
GC_10_601 b_10 NI_10 NS_601 0 3.1862102138714992e-04
GC_10_602 b_10 NI_10 NS_602 0 2.1875096644603405e-04
GC_10_603 b_10 NI_10 NS_603 0 -5.0195635069949873e-07
GC_10_604 b_10 NI_10 NS_604 0 1.2291285014520426e-06
GC_10_605 b_10 NI_10 NS_605 0 -2.3042430254065419e-06
GC_10_606 b_10 NI_10 NS_606 0 -4.7508742159655183e-06
GC_10_607 b_10 NI_10 NS_607 0 -9.4393616475216811e-05
GC_10_608 b_10 NI_10 NS_608 0 1.1046320975462246e-04
GC_10_609 b_10 NI_10 NS_609 0 -5.7677931676008635e-06
GC_10_610 b_10 NI_10 NS_610 0 -1.3496240508362586e-05
GC_10_611 b_10 NI_10 NS_611 0 -1.0649463455315817e-05
GC_10_612 b_10 NI_10 NS_612 0 4.9051958911769567e-06
GC_10_613 b_10 NI_10 NS_613 0 2.0406233550466351e-05
GC_10_614 b_10 NI_10 NS_614 0 -4.0948282796942854e-05
GC_10_615 b_10 NI_10 NS_615 0 -4.0245317950035121e-05
GC_10_616 b_10 NI_10 NS_616 0 5.5913555002548786e-05
GC_10_617 b_10 NI_10 NS_617 0 -1.5626950639028778e-02
GC_10_618 b_10 NI_10 NS_618 0 -1.3168205663802925e-03
GC_10_619 b_10 NI_10 NS_619 0 -8.5784258680989879e-04
GC_10_620 b_10 NI_10 NS_620 0 -1.0120647466529502e-03
GC_10_621 b_10 NI_10 NS_621 0 -1.1834877486462598e-03
GC_10_622 b_10 NI_10 NS_622 0 1.3679579038814666e-03
GC_10_623 b_10 NI_10 NS_623 0 8.5002053946324019e-04
GC_10_624 b_10 NI_10 NS_624 0 -7.8518755500926881e-04
GC_10_625 b_10 NI_10 NS_625 0 -3.1542009806875917e-03
GC_10_626 b_10 NI_10 NS_626 0 -8.6413502752787901e-03
GC_10_627 b_10 NI_10 NS_627 0 1.4334396982429955e-04
GC_10_628 b_10 NI_10 NS_628 0 2.9248266007608764e-04
GC_10_629 b_10 NI_10 NS_629 0 1.9539880341973878e-03
GC_10_630 b_10 NI_10 NS_630 0 -2.3240803318472589e-03
GC_10_631 b_10 NI_10 NS_631 0 7.3986093395509995e-04
GC_10_632 b_10 NI_10 NS_632 0 1.7269883996400665e-04
GC_10_633 b_10 NI_10 NS_633 0 9.6201656983447019e-04
GC_10_634 b_10 NI_10 NS_634 0 -1.9843545197016218e-03
GC_10_635 b_10 NI_10 NS_635 0 1.2224896091768836e-03
GC_10_636 b_10 NI_10 NS_636 0 -2.2764590193292853e-03
GC_10_637 b_10 NI_10 NS_637 0 4.0022670476810828e-05
GC_10_638 b_10 NI_10 NS_638 0 8.3464048115018035e-06
GC_10_639 b_10 NI_10 NS_639 0 7.4400237579959486e-03
GC_10_640 b_10 NI_10 NS_640 0 9.9323938492976789e-04
GC_10_641 b_10 NI_10 NS_641 0 -1.2056111177793127e-04
GC_10_642 b_10 NI_10 NS_642 0 4.1547217857106955e-05
GC_10_643 b_10 NI_10 NS_643 0 -1.3571176040859159e-04
GC_10_644 b_10 NI_10 NS_644 0 1.1791348637475406e-04
GC_10_645 b_10 NI_10 NS_645 0 1.8775654067958853e-04
GC_10_646 b_10 NI_10 NS_646 0 -3.8324207868787002e-04
GC_10_647 b_10 NI_10 NS_647 0 3.5053579787665105e-04
GC_10_648 b_10 NI_10 NS_648 0 -1.0949198679199138e-04
GC_10_649 b_10 NI_10 NS_649 0 -7.4695143180210340e-03
GC_10_650 b_10 NI_10 NS_650 0 3.0404032246076061e-03
GC_10_651 b_10 NI_10 NS_651 0 -2.1439477737131220e-04
GC_10_652 b_10 NI_10 NS_652 0 -1.6140356320442937e-04
GC_10_653 b_10 NI_10 NS_653 0 3.8172660632330487e-03
GC_10_654 b_10 NI_10 NS_654 0 4.4515141080362497e-04
GC_10_655 b_10 NI_10 NS_655 0 2.3570074059822404e-03
GC_10_656 b_10 NI_10 NS_656 0 -9.3363739374566939e-04
GC_10_657 b_10 NI_10 NS_657 0 7.5365856719772123e-04
GC_10_658 b_10 NI_10 NS_658 0 3.2995784600058580e-04
GC_10_659 b_10 NI_10 NS_659 0 -2.9544887146700304e-06
GC_10_660 b_10 NI_10 NS_660 0 -4.4539309379401860e-06
GC_10_661 b_10 NI_10 NS_661 0 -1.9883426380251326e-05
GC_10_662 b_10 NI_10 NS_662 0 -4.9842393510494614e-06
GC_10_663 b_10 NI_10 NS_663 0 -3.7260881487981782e-05
GC_10_664 b_10 NI_10 NS_664 0 -7.7416402837566478e-05
GC_10_665 b_10 NI_10 NS_665 0 -2.5277579912313427e-05
GC_10_666 b_10 NI_10 NS_666 0 2.2891817037080432e-06
GC_10_667 b_10 NI_10 NS_667 0 -1.4106412470087479e-05
GC_10_668 b_10 NI_10 NS_668 0 -9.2538625356305751e-06
GC_10_669 b_10 NI_10 NS_669 0 2.3860467510717617e-04
GC_10_670 b_10 NI_10 NS_670 0 -1.3050306293977855e-04
GC_10_671 b_10 NI_10 NS_671 0 -3.9506518624467490e-04
GC_10_672 b_10 NI_10 NS_672 0 9.2451053503236224e-05
GD_10_1 b_10 NI_10 NA_1 0 1.7248625842646629e-03
GD_10_2 b_10 NI_10 NA_2 0 3.9415667803272738e-03
GD_10_3 b_10 NI_10 NA_3 0 -3.4648378884776622e-03
GD_10_4 b_10 NI_10 NA_4 0 3.0061871428501670e-03
GD_10_5 b_10 NI_10 NA_5 0 -9.6464049588868524e-05
GD_10_6 b_10 NI_10 NA_6 0 -3.1486186037240280e-03
GD_10_7 b_10 NI_10 NA_7 0 -1.2216992980835723e-02
GD_10_8 b_10 NI_10 NA_8 0 4.9507838723997413e-03
GD_10_9 b_10 NI_10 NA_9 0 4.2603485398235844e-02
GD_10_10 b_10 NI_10 NA_10 0 9.3932487105311144e-02
GD_10_11 b_10 NI_10 NA_11 0 -5.4675147286476870e-02
GD_10_12 b_10 NI_10 NA_12 0 1.1228841767488370e-02
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 3.2345193180285170e-02
GC_11_2 b_11 NI_11 NS_2 0 -2.1059964198148359e-05
GC_11_3 b_11 NI_11 NS_3 0 2.3040074279715846e-04
GC_11_4 b_11 NI_11 NS_4 0 -5.6559446719548379e-04
GC_11_5 b_11 NI_11 NS_5 0 7.6516420633366807e-04
GC_11_6 b_11 NI_11 NS_6 0 3.5584541722955140e-04
GC_11_7 b_11 NI_11 NS_7 0 1.8691430500480586e-03
GC_11_8 b_11 NI_11 NS_8 0 1.9497909510203994e-03
GC_11_9 b_11 NI_11 NS_9 0 -3.8033075040125948e-04
GC_11_10 b_11 NI_11 NS_10 0 4.2106693176432617e-03
GC_11_11 b_11 NI_11 NS_11 0 -2.3257555751392725e-04
GC_11_12 b_11 NI_11 NS_12 0 5.7504164783841127e-04
GC_11_13 b_11 NI_11 NS_13 0 1.0508309566406087e-03
GC_11_14 b_11 NI_11 NS_14 0 5.8664605060333014e-04
GC_11_15 b_11 NI_11 NS_15 0 1.0300021625476042e-03
GC_11_16 b_11 NI_11 NS_16 0 2.8732096166701119e-04
GC_11_17 b_11 NI_11 NS_17 0 3.6921704061746696e-05
GC_11_18 b_11 NI_11 NS_18 0 5.3304317228771393e-03
GC_11_19 b_11 NI_11 NS_19 0 1.0929009073886689e-03
GC_11_20 b_11 NI_11 NS_20 0 1.9270998397391927e-03
GC_11_21 b_11 NI_11 NS_21 0 3.3144581941224442e-04
GC_11_22 b_11 NI_11 NS_22 0 1.5942086079009666e-04
GC_11_23 b_11 NI_11 NS_23 0 -6.7849043611705089e-03
GC_11_24 b_11 NI_11 NS_24 0 8.9135615988905556e-03
GC_11_25 b_11 NI_11 NS_25 0 -1.5271809998164456e-04
GC_11_26 b_11 NI_11 NS_26 0 -2.6374402912166314e-04
GC_11_27 b_11 NI_11 NS_27 0 -7.3644263703297197e-04
GC_11_28 b_11 NI_11 NS_28 0 -9.9349715198886144e-05
GC_11_29 b_11 NI_11 NS_29 0 -3.7092847758007886e-04
GC_11_30 b_11 NI_11 NS_30 0 -1.4108233965292872e-04
GC_11_31 b_11 NI_11 NS_31 0 -1.1156669776780053e-04
GC_11_32 b_11 NI_11 NS_32 0 2.2538329030579353e-05
GC_11_33 b_11 NI_11 NS_33 0 -8.3646600483811596e-03
GC_11_34 b_11 NI_11 NS_34 0 -4.3034895441439085e-03
GC_11_35 b_11 NI_11 NS_35 0 5.9660640416575302e-05
GC_11_36 b_11 NI_11 NS_36 0 -6.2654333391171441e-05
GC_11_37 b_11 NI_11 NS_37 0 -2.5759488961886310e-04
GC_11_38 b_11 NI_11 NS_38 0 1.5037226128020496e-03
GC_11_39 b_11 NI_11 NS_39 0 3.0373757556221345e-03
GC_11_40 b_11 NI_11 NS_40 0 -4.5808894921753190e-03
GC_11_41 b_11 NI_11 NS_41 0 7.2403686094156278e-05
GC_11_42 b_11 NI_11 NS_42 0 3.4665172275288544e-04
GC_11_43 b_11 NI_11 NS_43 0 1.4136709581717287e-06
GC_11_44 b_11 NI_11 NS_44 0 3.8101517481053902e-06
GC_11_45 b_11 NI_11 NS_45 0 -5.1045094275017345e-06
GC_11_46 b_11 NI_11 NS_46 0 -1.9812760349815932e-05
GC_11_47 b_11 NI_11 NS_47 0 -3.0450303987797399e-04
GC_11_48 b_11 NI_11 NS_48 0 2.7827138924363143e-04
GC_11_49 b_11 NI_11 NS_49 0 1.3734273723039436e-06
GC_11_50 b_11 NI_11 NS_50 0 -4.7309306613029397e-05
GC_11_51 b_11 NI_11 NS_51 0 -3.4617224131407658e-05
GC_11_52 b_11 NI_11 NS_52 0 -7.0181506825600493e-06
GC_11_53 b_11 NI_11 NS_53 0 9.6426075408037387e-05
GC_11_54 b_11 NI_11 NS_54 0 -9.7333428518469947e-05
GC_11_55 b_11 NI_11 NS_55 0 -1.8916155324044478e-04
GC_11_56 b_11 NI_11 NS_56 0 9.9144720726420830e-05
GC_11_57 b_11 NI_11 NS_57 0 -6.3518825150341582e-03
GC_11_58 b_11 NI_11 NS_58 0 -1.0081876760138061e-04
GC_11_59 b_11 NI_11 NS_59 0 2.5384877415710673e-04
GC_11_60 b_11 NI_11 NS_60 0 2.9809391808544266e-04
GC_11_61 b_11 NI_11 NS_61 0 -3.5932983007138232e-04
GC_11_62 b_11 NI_11 NS_62 0 3.0721814472942842e-04
GC_11_63 b_11 NI_11 NS_63 0 -1.7649585074817596e-03
GC_11_64 b_11 NI_11 NS_64 0 2.7455024735844246e-04
GC_11_65 b_11 NI_11 NS_65 0 -1.2020526483094316e-03
GC_11_66 b_11 NI_11 NS_66 0 -2.4964273512978023e-03
GC_11_67 b_11 NI_11 NS_67 0 5.9946031205934105e-04
GC_11_68 b_11 NI_11 NS_68 0 -4.4721532436410897e-04
GC_11_69 b_11 NI_11 NS_69 0 7.3554217786909787e-04
GC_11_70 b_11 NI_11 NS_70 0 -1.7145084796331817e-03
GC_11_71 b_11 NI_11 NS_71 0 3.8518369841143290e-04
GC_11_72 b_11 NI_11 NS_72 0 -1.9544643462083709e-04
GC_11_73 b_11 NI_11 NS_73 0 1.4905749938437564e-03
GC_11_74 b_11 NI_11 NS_74 0 1.1008207424838897e-03
GC_11_75 b_11 NI_11 NS_75 0 -5.3474494476066616e-04
GC_11_76 b_11 NI_11 NS_76 0 9.0367037034517616e-04
GC_11_77 b_11 NI_11 NS_77 0 -1.1872172573023154e-04
GC_11_78 b_11 NI_11 NS_78 0 4.4347108448557610e-05
GC_11_79 b_11 NI_11 NS_79 0 -2.5664879608197125e-03
GC_11_80 b_11 NI_11 NS_80 0 -5.0936308983957370e-04
GC_11_81 b_11 NI_11 NS_81 0 3.1108016566765979e-05
GC_11_82 b_11 NI_11 NS_82 0 6.2462264487393715e-04
GC_11_83 b_11 NI_11 NS_83 0 -3.8495822163263214e-04
GC_11_84 b_11 NI_11 NS_84 0 1.3247920809521538e-05
GC_11_85 b_11 NI_11 NS_85 0 -4.1481098937182513e-04
GC_11_86 b_11 NI_11 NS_86 0 -9.6518399696188974e-05
GC_11_87 b_11 NI_11 NS_87 0 -8.4349460368420457e-05
GC_11_88 b_11 NI_11 NS_88 0 -9.2948657357211882e-05
GC_11_89 b_11 NI_11 NS_89 0 2.9607833226164351e-03
GC_11_90 b_11 NI_11 NS_90 0 -4.5932897099370228e-03
GC_11_91 b_11 NI_11 NS_91 0 1.6884833381501517e-05
GC_11_92 b_11 NI_11 NS_92 0 4.3792659461795640e-05
GC_11_93 b_11 NI_11 NS_93 0 -1.0129361422468947e-03
GC_11_94 b_11 NI_11 NS_94 0 -4.1718160094473368e-04
GC_11_95 b_11 NI_11 NS_95 0 7.6169041996058679e-04
GC_11_96 b_11 NI_11 NS_96 0 1.6985234613840182e-03
GC_11_97 b_11 NI_11 NS_97 0 -1.9284682913094851e-04
GC_11_98 b_11 NI_11 NS_98 0 6.9016590704786454e-05
GC_11_99 b_11 NI_11 NS_99 0 -3.5285770419449568e-06
GC_11_100 b_11 NI_11 NS_100 0 -9.4886666779373745e-07
GC_11_101 b_11 NI_11 NS_101 0 1.0819846895320297e-05
GC_11_102 b_11 NI_11 NS_102 0 7.0055322870792493e-06
GC_11_103 b_11 NI_11 NS_103 0 -5.8573627167774694e-05
GC_11_104 b_11 NI_11 NS_104 0 -2.2009852464749977e-04
GC_11_105 b_11 NI_11 NS_105 0 2.3120321964656591e-05
GC_11_106 b_11 NI_11 NS_106 0 1.6594776746832009e-05
GC_11_107 b_11 NI_11 NS_107 0 1.7087941099957868e-05
GC_11_108 b_11 NI_11 NS_108 0 -9.4796204582604856e-06
GC_11_109 b_11 NI_11 NS_109 0 1.6240348733139500e-05
GC_11_110 b_11 NI_11 NS_110 0 4.8356424693473093e-05
GC_11_111 b_11 NI_11 NS_111 0 6.5092655283625131e-06
GC_11_112 b_11 NI_11 NS_112 0 -7.6064802322564976e-05
GC_11_113 b_11 NI_11 NS_113 0 2.6865503605722336e-02
GC_11_114 b_11 NI_11 NS_114 0 -9.1147608018191875e-06
GC_11_115 b_11 NI_11 NS_115 0 7.2304462123805161e-04
GC_11_116 b_11 NI_11 NS_116 0 -6.2661469541225963e-04
GC_11_117 b_11 NI_11 NS_117 0 3.6818239143609002e-04
GC_11_118 b_11 NI_11 NS_118 0 1.0225473640243881e-03
GC_11_119 b_11 NI_11 NS_119 0 8.8921276972480658e-04
GC_11_120 b_11 NI_11 NS_120 0 2.2914004338159396e-03
GC_11_121 b_11 NI_11 NS_121 0 -2.2939181483885205e-03
GC_11_122 b_11 NI_11 NS_122 0 2.2457940546066085e-03
GC_11_123 b_11 NI_11 NS_123 0 -2.2456681868719707e-04
GC_11_124 b_11 NI_11 NS_124 0 1.5650219517132443e-04
GC_11_125 b_11 NI_11 NS_125 0 1.9356349081290131e-03
GC_11_126 b_11 NI_11 NS_126 0 -6.1778877851996787e-04
GC_11_127 b_11 NI_11 NS_127 0 1.3680151610097270e-03
GC_11_128 b_11 NI_11 NS_128 0 4.3539802342575833e-04
GC_11_129 b_11 NI_11 NS_129 0 -5.6560418246892933e-04
GC_11_130 b_11 NI_11 NS_130 0 3.9670545029511280e-03
GC_11_131 b_11 NI_11 NS_131 0 1.5711343398201823e-03
GC_11_132 b_11 NI_11 NS_132 0 1.9963452962701617e-03
GC_11_133 b_11 NI_11 NS_133 0 4.2452545424470048e-04
GC_11_134 b_11 NI_11 NS_134 0 2.6692915130680672e-04
GC_11_135 b_11 NI_11 NS_135 0 -4.6616642530308084e-03
GC_11_136 b_11 NI_11 NS_136 0 8.8629447378403958e-03
GC_11_137 b_11 NI_11 NS_137 0 -3.5175343472615130e-04
GC_11_138 b_11 NI_11 NS_138 0 -5.7005744886929786e-04
GC_11_139 b_11 NI_11 NS_139 0 -9.6580447283152340e-04
GC_11_140 b_11 NI_11 NS_140 0 4.9223777711219364e-05
GC_11_141 b_11 NI_11 NS_141 0 -4.5987323190148360e-04
GC_11_142 b_11 NI_11 NS_142 0 -1.3566619392521131e-04
GC_11_143 b_11 NI_11 NS_143 0 -1.5010314340280236e-04
GC_11_144 b_11 NI_11 NS_144 0 1.6853737736502163e-05
GC_11_145 b_11 NI_11 NS_145 0 -9.1781170042756835e-03
GC_11_146 b_11 NI_11 NS_146 0 -4.4385164887276564e-03
GC_11_147 b_11 NI_11 NS_147 0 4.8783912430576126e-05
GC_11_148 b_11 NI_11 NS_148 0 -6.2366839353467758e-05
GC_11_149 b_11 NI_11 NS_149 0 -1.2650838807128434e-04
GC_11_150 b_11 NI_11 NS_150 0 1.4402378597652774e-03
GC_11_151 b_11 NI_11 NS_151 0 3.7609136743077922e-03
GC_11_152 b_11 NI_11 NS_152 0 -4.1553736394158505e-03
GC_11_153 b_11 NI_11 NS_153 0 8.2575235934372911e-05
GC_11_154 b_11 NI_11 NS_154 0 3.0350562369078861e-04
GC_11_155 b_11 NI_11 NS_155 0 1.0518228281552034e-06
GC_11_156 b_11 NI_11 NS_156 0 3.7403128709395941e-06
GC_11_157 b_11 NI_11 NS_157 0 -2.3233031573989510e-06
GC_11_158 b_11 NI_11 NS_158 0 -1.6481915753646752e-05
GC_11_159 b_11 NI_11 NS_159 0 -2.4524358388591333e-04
GC_11_160 b_11 NI_11 NS_160 0 1.8847931204388758e-04
GC_11_161 b_11 NI_11 NS_161 0 4.3947344507272098e-06
GC_11_162 b_11 NI_11 NS_162 0 -3.5957957946267051e-05
GC_11_163 b_11 NI_11 NS_163 0 -2.5741989974405352e-05
GC_11_164 b_11 NI_11 NS_164 0 -6.6870901752578558e-06
GC_11_165 b_11 NI_11 NS_165 0 6.8713426889818909e-05
GC_11_166 b_11 NI_11 NS_166 0 -6.7102354469094806e-05
GC_11_167 b_11 NI_11 NS_167 0 -1.3336769739720236e-04
GC_11_168 b_11 NI_11 NS_168 0 6.7183059052160565e-05
GC_11_169 b_11 NI_11 NS_169 0 1.5858636601394317e-03
GC_11_170 b_11 NI_11 NS_170 0 -1.3930469552202328e-04
GC_11_171 b_11 NI_11 NS_171 0 1.6660069711446274e-04
GC_11_172 b_11 NI_11 NS_172 0 5.6245497460988118e-04
GC_11_173 b_11 NI_11 NS_173 0 -5.2813873839795296e-04
GC_11_174 b_11 NI_11 NS_174 0 -1.1100270235549543e-05
GC_11_175 b_11 NI_11 NS_175 0 -1.6224592255486905e-03
GC_11_176 b_11 NI_11 NS_176 0 -2.9776274694647280e-04
GC_11_177 b_11 NI_11 NS_177 0 5.9819465835822940e-04
GC_11_178 b_11 NI_11 NS_178 0 -1.9505061449116427e-03
GC_11_179 b_11 NI_11 NS_179 0 -1.5459692253751469e-05
GC_11_180 b_11 NI_11 NS_180 0 -1.9708618841330765e-04
GC_11_181 b_11 NI_11 NS_181 0 1.1849199735915134e-03
GC_11_182 b_11 NI_11 NS_182 0 -1.2359309433806140e-03
GC_11_183 b_11 NI_11 NS_183 0 7.3022842895232275e-04
GC_11_184 b_11 NI_11 NS_184 0 -2.3178773431841704e-04
GC_11_185 b_11 NI_11 NS_185 0 1.8185155508736517e-03
GC_11_186 b_11 NI_11 NS_186 0 1.9867095240926700e-03
GC_11_187 b_11 NI_11 NS_187 0 -5.4998114947577470e-04
GC_11_188 b_11 NI_11 NS_188 0 2.1768067422876553e-03
GC_11_189 b_11 NI_11 NS_189 0 -1.7623390754204683e-04
GC_11_190 b_11 NI_11 NS_190 0 -1.3365964921572132e-05
GC_11_191 b_11 NI_11 NS_191 0 -1.7125346298856106e-03
GC_11_192 b_11 NI_11 NS_192 0 1.3173825088635726e-03
GC_11_193 b_11 NI_11 NS_193 0 -1.3141239330211804e-05
GC_11_194 b_11 NI_11 NS_194 0 2.9410002192200365e-04
GC_11_195 b_11 NI_11 NS_195 0 -5.4947397875088793e-04
GC_11_196 b_11 NI_11 NS_196 0 9.6961764525898788e-05
GC_11_197 b_11 NI_11 NS_197 0 -3.4944923352633000e-04
GC_11_198 b_11 NI_11 NS_198 0 1.8528832096606921e-06
GC_11_199 b_11 NI_11 NS_199 0 -7.7701770086029918e-05
GC_11_200 b_11 NI_11 NS_200 0 -4.2295818295643913e-05
GC_11_201 b_11 NI_11 NS_201 0 -4.8350120676088327e-04
GC_11_202 b_11 NI_11 NS_202 0 -2.6842009504630527e-03
GC_11_203 b_11 NI_11 NS_203 0 1.8486442492203203e-05
GC_11_204 b_11 NI_11 NS_204 0 -6.2174111640890395e-06
GC_11_205 b_11 NI_11 NS_205 0 -6.3530729613622697e-04
GC_11_206 b_11 NI_11 NS_206 0 1.9393675084681029e-04
GC_11_207 b_11 NI_11 NS_207 0 9.7894910789472138e-04
GC_11_208 b_11 NI_11 NS_208 0 -3.1189658229970003e-04
GC_11_209 b_11 NI_11 NS_209 0 -1.0361976580208971e-04
GC_11_210 b_11 NI_11 NS_210 0 5.9585767990030911e-05
GC_11_211 b_11 NI_11 NS_211 0 -1.2427407089020016e-06
GC_11_212 b_11 NI_11 NS_212 0 7.7525633150641506e-07
GC_11_213 b_11 NI_11 NS_213 0 3.9412766755348963e-06
GC_11_214 b_11 NI_11 NS_214 0 -3.1970582338290403e-07
GC_11_215 b_11 NI_11 NS_215 0 -5.0436767265479588e-05
GC_11_216 b_11 NI_11 NS_216 0 -5.8783799963131927e-05
GC_11_217 b_11 NI_11 NS_217 0 1.1300242728696197e-05
GC_11_218 b_11 NI_11 NS_218 0 2.8132194829248678e-07
GC_11_219 b_11 NI_11 NS_219 0 3.1110831360956457e-06
GC_11_220 b_11 NI_11 NS_220 0 -3.6760171352353435e-06
GC_11_221 b_11 NI_11 NS_221 0 1.9556764542869830e-05
GC_11_222 b_11 NI_11 NS_222 0 -1.9747561453384339e-06
GC_11_223 b_11 NI_11 NS_223 0 -2.3715436457477560e-05
GC_11_224 b_11 NI_11 NS_224 0 -1.8413322119407094e-06
GC_11_225 b_11 NI_11 NS_225 0 6.9540425456234803e-04
GC_11_226 b_11 NI_11 NS_226 0 3.7827142030583870e-05
GC_11_227 b_11 NI_11 NS_227 0 1.2320224963636554e-03
GC_11_228 b_11 NI_11 NS_228 0 -1.3867989218286156e-04
GC_11_229 b_11 NI_11 NS_229 0 -1.1142250211357728e-03
GC_11_230 b_11 NI_11 NS_230 0 1.2983303305714015e-03
GC_11_231 b_11 NI_11 NS_231 0 -9.6308678339310303e-04
GC_11_232 b_11 NI_11 NS_232 0 7.1189469755289438e-04
GC_11_233 b_11 NI_11 NS_233 0 -2.7560385552193403e-03
GC_11_234 b_11 NI_11 NS_234 0 -3.0180073072401058e-03
GC_11_235 b_11 NI_11 NS_235 0 7.1991113400794528e-05
GC_11_236 b_11 NI_11 NS_236 0 -3.2740676926052613e-04
GC_11_237 b_11 NI_11 NS_237 0 2.8165679566524268e-03
GC_11_238 b_11 NI_11 NS_238 0 -1.5940867371299146e-03
GC_11_239 b_11 NI_11 NS_239 0 1.2681648474039526e-03
GC_11_240 b_11 NI_11 NS_240 0 5.1741972193928415e-04
GC_11_241 b_11 NI_11 NS_241 0 -1.3086168403006648e-03
GC_11_242 b_11 NI_11 NS_242 0 4.1156243807015237e-05
GC_11_243 b_11 NI_11 NS_243 0 1.6315819060568355e-03
GC_11_244 b_11 NI_11 NS_244 0 2.4417841598142954e-04
GC_11_245 b_11 NI_11 NS_245 0 4.8154138423240250e-04
GC_11_246 b_11 NI_11 NS_246 0 2.3802634626403940e-04
GC_11_247 b_11 NI_11 NS_247 0 2.1978262805051724e-04
GC_11_248 b_11 NI_11 NS_248 0 5.1342982039380381e-03
GC_11_249 b_11 NI_11 NS_249 0 -3.5469528466643726e-04
GC_11_250 b_11 NI_11 NS_250 0 -6.9365270423744907e-04
GC_11_251 b_11 NI_11 NS_251 0 -8.5901182367222333e-04
GC_11_252 b_11 NI_11 NS_252 0 4.5141393768430474e-05
GC_11_253 b_11 NI_11 NS_253 0 -3.3081418827208100e-04
GC_11_254 b_11 NI_11 NS_254 0 -2.7724700131744295e-04
GC_11_255 b_11 NI_11 NS_255 0 -8.3390310497823348e-05
GC_11_256 b_11 NI_11 NS_256 0 1.0532477204677385e-05
GC_11_257 b_11 NI_11 NS_257 0 -3.4380354148358244e-03
GC_11_258 b_11 NI_11 NS_258 0 -4.7631109611810680e-03
GC_11_259 b_11 NI_11 NS_259 0 2.7475111373268843e-05
GC_11_260 b_11 NI_11 NS_260 0 -5.1795565347352376e-05
GC_11_261 b_11 NI_11 NS_261 0 8.5947956263940627e-05
GC_11_262 b_11 NI_11 NS_262 0 7.8708984805061165e-04
GC_11_263 b_11 NI_11 NS_263 0 2.4790519629065639e-03
GC_11_264 b_11 NI_11 NS_264 0 6.8932619862888513e-04
GC_11_265 b_11 NI_11 NS_265 0 6.0240482963995117e-06
GC_11_266 b_11 NI_11 NS_266 0 3.2036882985167644e-04
GC_11_267 b_11 NI_11 NS_267 0 -8.7571341875453961e-07
GC_11_268 b_11 NI_11 NS_268 0 1.3609419016393678e-06
GC_11_269 b_11 NI_11 NS_269 0 3.2215924590707633e-06
GC_11_270 b_11 NI_11 NS_270 0 -3.3715884641204156e-06
GC_11_271 b_11 NI_11 NS_271 0 -1.0089361858069173e-04
GC_11_272 b_11 NI_11 NS_272 0 1.0649943054278605e-05
GC_11_273 b_11 NI_11 NS_273 0 7.1766640123956785e-06
GC_11_274 b_11 NI_11 NS_274 0 -5.2838506003239976e-06
GC_11_275 b_11 NI_11 NS_275 0 -6.8823445024233530e-06
GC_11_276 b_11 NI_11 NS_276 0 -5.4896806309339152e-06
GC_11_277 b_11 NI_11 NS_277 0 2.1866444239383327e-05
GC_11_278 b_11 NI_11 NS_278 0 -6.6659371106121780e-06
GC_11_279 b_11 NI_11 NS_279 0 -3.5631842337882169e-05
GC_11_280 b_11 NI_11 NS_280 0 7.4023037370398982e-07
GC_11_281 b_11 NI_11 NS_281 0 7.8306304410918903e-03
GC_11_282 b_11 NI_11 NS_282 0 -9.1683925924957973e-05
GC_11_283 b_11 NI_11 NS_283 0 -1.7746160872522728e-04
GC_11_284 b_11 NI_11 NS_284 0 7.1868147592506909e-04
GC_11_285 b_11 NI_11 NS_285 0 -3.1687559950480332e-04
GC_11_286 b_11 NI_11 NS_286 0 -6.9173339832637800e-04
GC_11_287 b_11 NI_11 NS_287 0 -5.4972304468654755e-04
GC_11_288 b_11 NI_11 NS_288 0 -7.7045896933881388e-04
GC_11_289 b_11 NI_11 NS_289 0 2.2332214597003031e-03
GC_11_290 b_11 NI_11 NS_290 0 7.1014888290111058e-04
GC_11_291 b_11 NI_11 NS_291 0 -5.9311172811959934e-04
GC_11_292 b_11 NI_11 NS_292 0 3.0662366387486048e-04
GC_11_293 b_11 NI_11 NS_293 0 5.1812684369132518e-04
GC_11_294 b_11 NI_11 NS_294 0 -6.3159516210515296e-04
GC_11_295 b_11 NI_11 NS_295 0 9.9893440500917956e-04
GC_11_296 b_11 NI_11 NS_296 0 -1.8583036461275755e-04
GC_11_297 b_11 NI_11 NS_297 0 8.3923943504014267e-04
GC_11_298 b_11 NI_11 NS_298 0 2.2099106605656953e-03
GC_11_299 b_11 NI_11 NS_299 0 -1.3060481659067865e-03
GC_11_300 b_11 NI_11 NS_300 0 2.6968060310000180e-03
GC_11_301 b_11 NI_11 NS_301 0 -2.7300723073423545e-04
GC_11_302 b_11 NI_11 NS_302 0 -6.8984088293699882e-05
GC_11_303 b_11 NI_11 NS_303 0 -5.1686945232628850e-04
GC_11_304 b_11 NI_11 NS_304 0 1.3705710614142245e-03
GC_11_305 b_11 NI_11 NS_305 0 5.5089905865704633e-05
GC_11_306 b_11 NI_11 NS_306 0 -1.2475501634155019e-06
GC_11_307 b_11 NI_11 NS_307 0 -7.3218037447783061e-04
GC_11_308 b_11 NI_11 NS_308 0 2.4700416215005640e-04
GC_11_309 b_11 NI_11 NS_309 0 -4.8231904909233110e-04
GC_11_310 b_11 NI_11 NS_310 0 6.0035738309812745e-05
GC_11_311 b_11 NI_11 NS_311 0 -1.1685653964262842e-04
GC_11_312 b_11 NI_11 NS_312 0 -4.0207276257279080e-05
GC_11_313 b_11 NI_11 NS_313 0 -4.7116972503407522e-04
GC_11_314 b_11 NI_11 NS_314 0 -2.7219927015019198e-03
GC_11_315 b_11 NI_11 NS_315 0 2.7566797172455769e-05
GC_11_316 b_11 NI_11 NS_316 0 -2.4079029041491425e-05
GC_11_317 b_11 NI_11 NS_317 0 -8.6665643407938468e-04
GC_11_318 b_11 NI_11 NS_318 0 4.0256217825960020e-04
GC_11_319 b_11 NI_11 NS_319 0 1.0381717063458328e-03
GC_11_320 b_11 NI_11 NS_320 0 2.5633695602932311e-04
GC_11_321 b_11 NI_11 NS_321 0 -1.3608131901744625e-04
GC_11_322 b_11 NI_11 NS_322 0 1.3811464717495661e-04
GC_11_323 b_11 NI_11 NS_323 0 -2.2894717286885097e-06
GC_11_324 b_11 NI_11 NS_324 0 2.5428301028410277e-06
GC_11_325 b_11 NI_11 NS_325 0 3.2788243197843150e-07
GC_11_326 b_11 NI_11 NS_326 0 -3.3797397164917950e-06
GC_11_327 b_11 NI_11 NS_327 0 -5.6560745902107001e-05
GC_11_328 b_11 NI_11 NS_328 0 3.6649605506077448e-05
GC_11_329 b_11 NI_11 NS_329 0 5.6224632493838787e-06
GC_11_330 b_11 NI_11 NS_330 0 -9.4040692107483521e-06
GC_11_331 b_11 NI_11 NS_331 0 -7.7875081784237803e-07
GC_11_332 b_11 NI_11 NS_332 0 -6.4072670727319962e-06
GC_11_333 b_11 NI_11 NS_333 0 2.7637026871451865e-05
GC_11_334 b_11 NI_11 NS_334 0 -3.7206385895602300e-05
GC_11_335 b_11 NI_11 NS_335 0 -5.0132657712862404e-05
GC_11_336 b_11 NI_11 NS_336 0 4.6877754414760336e-05
GC_11_337 b_11 NI_11 NS_337 0 -1.7513274191208829e-02
GC_11_338 b_11 NI_11 NS_338 0 6.2692913950595619e-04
GC_11_339 b_11 NI_11 NS_339 0 8.0498192394140057e-04
GC_11_340 b_11 NI_11 NS_340 0 8.1000824932661814e-04
GC_11_341 b_11 NI_11 NS_341 0 -1.6184484045364360e-03
GC_11_342 b_11 NI_11 NS_342 0 -2.4432493191605120e-03
GC_11_343 b_11 NI_11 NS_343 0 1.2162876038709664e-03
GC_11_344 b_11 NI_11 NS_344 0 -3.6566454444035676e-04
GC_11_345 b_11 NI_11 NS_345 0 4.0419266586437103e-03
GC_11_346 b_11 NI_11 NS_346 0 -4.0562196170599975e-03
GC_11_347 b_11 NI_11 NS_347 0 -3.1815896679098930e-04
GC_11_348 b_11 NI_11 NS_348 0 1.6430966133142917e-04
GC_11_349 b_11 NI_11 NS_349 0 2.5152980162469456e-03
GC_11_350 b_11 NI_11 NS_350 0 -1.6564678125138220e-04
GC_11_351 b_11 NI_11 NS_351 0 1.0452547707192862e-03
GC_11_352 b_11 NI_11 NS_352 0 6.4452650446863372e-04
GC_11_353 b_11 NI_11 NS_353 0 1.0876289110984543e-03
GC_11_354 b_11 NI_11 NS_354 0 -1.5186341414479099e-03
GC_11_355 b_11 NI_11 NS_355 0 2.5713168007458266e-03
GC_11_356 b_11 NI_11 NS_356 0 -1.7437366641506565e-04
GC_11_357 b_11 NI_11 NS_357 0 3.5079276319885876e-04
GC_11_358 b_11 NI_11 NS_358 0 1.7554417196071647e-04
GC_11_359 b_11 NI_11 NS_359 0 2.4325350531653259e-03
GC_11_360 b_11 NI_11 NS_360 0 5.7447965226306540e-03
GC_11_361 b_11 NI_11 NS_361 0 -5.9984672812593894e-05
GC_11_362 b_11 NI_11 NS_362 0 -6.7719109870920666e-04
GC_11_363 b_11 NI_11 NS_363 0 -6.0503983355193443e-04
GC_11_364 b_11 NI_11 NS_364 0 1.8785373372765061e-04
GC_11_365 b_11 NI_11 NS_365 0 -1.6670827904274966e-04
GC_11_366 b_11 NI_11 NS_366 0 -1.0491864427585406e-04
GC_11_367 b_11 NI_11 NS_367 0 -6.3607770944017314e-05
GC_11_368 b_11 NI_11 NS_368 0 2.4854902124881154e-05
GC_11_369 b_11 NI_11 NS_369 0 8.3313264990011939e-04
GC_11_370 b_11 NI_11 NS_370 0 1.0473768561826710e-03
GC_11_371 b_11 NI_11 NS_371 0 1.4736836907659083e-05
GC_11_372 b_11 NI_11 NS_372 0 -3.1671095304953730e-05
GC_11_373 b_11 NI_11 NS_373 0 3.7319105064118595e-04
GC_11_374 b_11 NI_11 NS_374 0 4.1477653696155665e-04
GC_11_375 b_11 NI_11 NS_375 0 -2.2355184734348804e-03
GC_11_376 b_11 NI_11 NS_376 0 5.8076485758390395e-04
GC_11_377 b_11 NI_11 NS_377 0 -1.6288533290265307e-04
GC_11_378 b_11 NI_11 NS_378 0 -2.2751855138437453e-04
GC_11_379 b_11 NI_11 NS_379 0 1.3468051966617057e-06
GC_11_380 b_11 NI_11 NS_380 0 -5.0923232845049700e-07
GC_11_381 b_11 NI_11 NS_381 0 7.3044406817629831e-06
GC_11_382 b_11 NI_11 NS_382 0 9.0616786473155021e-06
GC_11_383 b_11 NI_11 NS_383 0 1.3378574547605630e-04
GC_11_384 b_11 NI_11 NS_384 0 -1.5806843204354306e-04
GC_11_385 b_11 NI_11 NS_385 0 5.9660815147102354e-06
GC_11_386 b_11 NI_11 NS_386 0 2.2325765582598134e-05
GC_11_387 b_11 NI_11 NS_387 0 6.0023983387830244e-06
GC_11_388 b_11 NI_11 NS_388 0 6.8479528774852029e-06
GC_11_389 b_11 NI_11 NS_389 0 -3.7525102279808386e-05
GC_11_390 b_11 NI_11 NS_390 0 2.0239371137989279e-05
GC_11_391 b_11 NI_11 NS_391 0 6.7721926180399719e-05
GC_11_392 b_11 NI_11 NS_392 0 -9.5876283358939877e-06
GC_11_393 b_11 NI_11 NS_393 0 2.6509271169455229e-02
GC_11_394 b_11 NI_11 NS_394 0 -2.8560267373152975e-04
GC_11_395 b_11 NI_11 NS_395 0 -4.6672448184521500e-04
GC_11_396 b_11 NI_11 NS_396 0 5.6166547167500400e-04
GC_11_397 b_11 NI_11 NS_397 0 1.0830866259422260e-03
GC_11_398 b_11 NI_11 NS_398 0 2.4769511767037565e-04
GC_11_399 b_11 NI_11 NS_399 0 -1.1485844227287283e-03
GC_11_400 b_11 NI_11 NS_400 0 9.4539014346810854e-04
GC_11_401 b_11 NI_11 NS_401 0 -2.8069487227110022e-03
GC_11_402 b_11 NI_11 NS_402 0 4.5021822344542958e-03
GC_11_403 b_11 NI_11 NS_403 0 -2.3787033187647950e-04
GC_11_404 b_11 NI_11 NS_404 0 1.4291726896374586e-04
GC_11_405 b_11 NI_11 NS_405 0 4.7113619346138924e-05
GC_11_406 b_11 NI_11 NS_406 0 -1.2076189545111157e-03
GC_11_407 b_11 NI_11 NS_407 0 7.7334494509437096e-04
GC_11_408 b_11 NI_11 NS_408 0 1.3893067117185101e-04
GC_11_409 b_11 NI_11 NS_409 0 -4.8497811809248268e-04
GC_11_410 b_11 NI_11 NS_410 0 7.4306481863390176e-04
GC_11_411 b_11 NI_11 NS_411 0 -1.6970850942716899e-03
GC_11_412 b_11 NI_11 NS_412 0 9.7327851358377170e-04
GC_11_413 b_11 NI_11 NS_413 0 -1.2707743894691825e-04
GC_11_414 b_11 NI_11 NS_414 0 -9.1179174914751495e-05
GC_11_415 b_11 NI_11 NS_415 0 3.3113896435844941e-05
GC_11_416 b_11 NI_11 NS_416 0 2.2189855260738010e-03
GC_11_417 b_11 NI_11 NS_417 0 6.4554428098700511e-05
GC_11_418 b_11 NI_11 NS_418 0 -1.8152559370233584e-04
GC_11_419 b_11 NI_11 NS_419 0 -5.0940186686730139e-04
GC_11_420 b_11 NI_11 NS_420 0 1.5196497028015942e-04
GC_11_421 b_11 NI_11 NS_421 0 -3.0484838175643726e-04
GC_11_422 b_11 NI_11 NS_422 0 1.2518113152990419e-04
GC_11_423 b_11 NI_11 NS_423 0 -9.8987499009788182e-05
GC_11_424 b_11 NI_11 NS_424 0 -1.5066502203278203e-05
GC_11_425 b_11 NI_11 NS_425 0 -1.1915552964813110e-03
GC_11_426 b_11 NI_11 NS_426 0 3.3027167186501369e-04
GC_11_427 b_11 NI_11 NS_427 0 3.0081174530195484e-05
GC_11_428 b_11 NI_11 NS_428 0 -2.1064678215518496e-05
GC_11_429 b_11 NI_11 NS_429 0 -5.1575977597446271e-04
GC_11_430 b_11 NI_11 NS_430 0 5.2073917480612649e-04
GC_11_431 b_11 NI_11 NS_431 0 -1.5817023723714615e-03
GC_11_432 b_11 NI_11 NS_432 0 -1.8552751220747216e-03
GC_11_433 b_11 NI_11 NS_433 0 -1.9381343302402024e-04
GC_11_434 b_11 NI_11 NS_434 0 -6.2506513491129758e-05
GC_11_435 b_11 NI_11 NS_435 0 -3.5796024733112598e-09
GC_11_436 b_11 NI_11 NS_436 0 1.2054900528443924e-06
GC_11_437 b_11 NI_11 NS_437 0 -6.1440954896454758e-06
GC_11_438 b_11 NI_11 NS_438 0 -3.8983646880223630e-06
GC_11_439 b_11 NI_11 NS_439 0 6.7383185378773003e-05
GC_11_440 b_11 NI_11 NS_440 0 1.3609504520204667e-04
GC_11_441 b_11 NI_11 NS_441 0 -9.1000076740416145e-06
GC_11_442 b_11 NI_11 NS_442 0 -1.1808584822019504e-05
GC_11_443 b_11 NI_11 NS_443 0 -4.6496437462752675e-06
GC_11_444 b_11 NI_11 NS_444 0 4.1895675167002972e-06
GC_11_445 b_11 NI_11 NS_445 0 8.5648152682289738e-06
GC_11_446 b_11 NI_11 NS_446 0 -4.9521760414323213e-05
GC_11_447 b_11 NI_11 NS_447 0 -3.2055345758410771e-05
GC_11_448 b_11 NI_11 NS_448 0 7.2202900640079697e-05
GC_11_449 b_11 NI_11 NS_449 0 -1.2339460024625611e-02
GC_11_450 b_11 NI_11 NS_450 0 1.5846354246809064e-03
GC_11_451 b_11 NI_11 NS_451 0 3.7051082345271624e-03
GC_11_452 b_11 NI_11 NS_452 0 2.4603662628618411e-03
GC_11_453 b_11 NI_11 NS_453 0 -5.2611608997405494e-03
GC_11_454 b_11 NI_11 NS_454 0 -6.3979683759243112e-03
GC_11_455 b_11 NI_11 NS_455 0 4.0078752075361577e-03
GC_11_456 b_11 NI_11 NS_456 0 2.5416635664440926e-03
GC_11_457 b_11 NI_11 NS_457 0 1.0136069275778746e-02
GC_11_458 b_11 NI_11 NS_458 0 -9.6415195120836371e-03
GC_11_459 b_11 NI_11 NS_459 0 -6.6842177128774037e-04
GC_11_460 b_11 NI_11 NS_460 0 5.3367257004975144e-04
GC_11_461 b_11 NI_11 NS_461 0 8.6833936288765283e-03
GC_11_462 b_11 NI_11 NS_462 0 3.3057946206565109e-03
GC_11_463 b_11 NI_11 NS_463 0 7.8724626817752990e-04
GC_11_464 b_11 NI_11 NS_464 0 2.0745267491034010e-03
GC_11_465 b_11 NI_11 NS_465 0 7.2191421889323468e-03
GC_11_466 b_11 NI_11 NS_466 0 1.6343651060947238e-03
GC_11_467 b_11 NI_11 NS_467 0 2.5992257205269013e-03
GC_11_468 b_11 NI_11 NS_468 0 4.3715633733234982e-03
GC_11_469 b_11 NI_11 NS_469 0 3.5240276956965592e-04
GC_11_470 b_11 NI_11 NS_470 0 1.0351618503227694e-04
GC_11_471 b_11 NI_11 NS_471 0 -4.5456942019832759e-03
GC_11_472 b_11 NI_11 NS_472 0 1.4407891628132982e-02
GC_11_473 b_11 NI_11 NS_473 0 1.0571347388660494e-03
GC_11_474 b_11 NI_11 NS_474 0 -2.4327580233877580e-05
GC_11_475 b_11 NI_11 NS_475 0 -5.9672236130094798e-04
GC_11_476 b_11 NI_11 NS_476 0 9.1789594268708487e-05
GC_11_477 b_11 NI_11 NS_477 0 -1.7944462537760651e-04
GC_11_478 b_11 NI_11 NS_478 0 2.1211104306922550e-04
GC_11_479 b_11 NI_11 NS_479 0 -7.5002204617307823e-05
GC_11_480 b_11 NI_11 NS_480 0 4.3474499455351532e-05
GC_11_481 b_11 NI_11 NS_481 0 -5.9431781270214701e-03
GC_11_482 b_11 NI_11 NS_482 0 -3.3187183759180107e-03
GC_11_483 b_11 NI_11 NS_483 0 8.5373790590630746e-05
GC_11_484 b_11 NI_11 NS_484 0 -6.5301450676996065e-05
GC_11_485 b_11 NI_11 NS_485 0 -3.4575409487866718e-05
GC_11_486 b_11 NI_11 NS_486 0 1.9728702383123658e-03
GC_11_487 b_11 NI_11 NS_487 0 -2.0814144959693505e-04
GC_11_488 b_11 NI_11 NS_488 0 -1.0923361934796713e-03
GC_11_489 b_11 NI_11 NS_489 0 6.7147092839248387e-05
GC_11_490 b_11 NI_11 NS_490 0 2.9052599824365150e-04
GC_11_491 b_11 NI_11 NS_491 0 -1.9245354080613066e-07
GC_11_492 b_11 NI_11 NS_492 0 7.2388099754010575e-07
GC_11_493 b_11 NI_11 NS_493 0 -1.4758363015936394e-06
GC_11_494 b_11 NI_11 NS_494 0 5.0749362455555511e-07
GC_11_495 b_11 NI_11 NS_495 0 3.5454796719583153e-05
GC_11_496 b_11 NI_11 NS_496 0 8.6835399351839349e-05
GC_11_497 b_11 NI_11 NS_497 0 -4.6804733072873849e-06
GC_11_498 b_11 NI_11 NS_498 0 -7.5284268064740225e-07
GC_11_499 b_11 NI_11 NS_499 0 -5.7916195433476308e-06
GC_11_500 b_11 NI_11 NS_500 0 -4.3944524610903541e-06
GC_11_501 b_11 NI_11 NS_501 0 1.7500238311540825e-05
GC_11_502 b_11 NI_11 NS_502 0 -1.6580121941456485e-05
GC_11_503 b_11 NI_11 NS_503 0 -3.6993400938381457e-05
GC_11_504 b_11 NI_11 NS_504 0 1.7379742673040315e-05
GC_11_505 b_11 NI_11 NS_505 0 5.7434285216554901e-02
GC_11_506 b_11 NI_11 NS_506 0 -7.8096423303072578e-04
GC_11_507 b_11 NI_11 NS_507 0 -1.7649582837868968e-03
GC_11_508 b_11 NI_11 NS_508 0 2.3941417913815747e-03
GC_11_509 b_11 NI_11 NS_509 0 2.8812338170612220e-03
GC_11_510 b_11 NI_11 NS_510 0 2.6566787309154440e-04
GC_11_511 b_11 NI_11 NS_511 0 -5.6069433122299750e-03
GC_11_512 b_11 NI_11 NS_512 0 4.9244666721716423e-04
GC_11_513 b_11 NI_11 NS_513 0 -6.3581741134313306e-03
GC_11_514 b_11 NI_11 NS_514 0 1.0169290054741277e-02
GC_11_515 b_11 NI_11 NS_515 0 -7.6138103010932995e-04
GC_11_516 b_11 NI_11 NS_516 0 3.0400926106163979e-05
GC_11_517 b_11 NI_11 NS_517 0 1.9032017236547271e-03
GC_11_518 b_11 NI_11 NS_518 0 -4.4859297146334388e-03
GC_11_519 b_11 NI_11 NS_519 0 1.0553095129953766e-03
GC_11_520 b_11 NI_11 NS_520 0 1.3589755216437624e-03
GC_11_521 b_11 NI_11 NS_521 0 -9.0134658967045960e-06
GC_11_522 b_11 NI_11 NS_522 0 1.1728772907550050e-03
GC_11_523 b_11 NI_11 NS_523 0 -5.8436637079249979e-03
GC_11_524 b_11 NI_11 NS_524 0 9.4976866331990034e-04
GC_11_525 b_11 NI_11 NS_525 0 -1.5340828563587290e-04
GC_11_526 b_11 NI_11 NS_526 0 -8.1534168087337122e-05
GC_11_527 b_11 NI_11 NS_527 0 1.2920501835581156e-03
GC_11_528 b_11 NI_11 NS_528 0 5.2330587846357276e-03
GC_11_529 b_11 NI_11 NS_529 0 -4.9894056287760077e-04
GC_11_530 b_11 NI_11 NS_530 0 -1.8074639022482012e-04
GC_11_531 b_11 NI_11 NS_531 0 -5.0411159345731759e-04
GC_11_532 b_11 NI_11 NS_532 0 7.6264330709591982e-05
GC_11_533 b_11 NI_11 NS_533 0 -4.5612509097742523e-04
GC_11_534 b_11 NI_11 NS_534 0 4.4236381567472089e-04
GC_11_535 b_11 NI_11 NS_535 0 -2.4602366516807085e-04
GC_11_536 b_11 NI_11 NS_536 0 -4.8690735916357919e-05
GC_11_537 b_11 NI_11 NS_537 0 -7.5535675398481494e-03
GC_11_538 b_11 NI_11 NS_538 0 -1.5776459721911500e-03
GC_11_539 b_11 NI_11 NS_539 0 -2.0328255694833080e-05
GC_11_540 b_11 NI_11 NS_540 0 4.2794299386367548e-05
GC_11_541 b_11 NI_11 NS_541 0 -9.0318469652872268e-05
GC_11_542 b_11 NI_11 NS_542 0 6.4024157100624386e-04
GC_11_543 b_11 NI_11 NS_543 0 -1.6179958643963615e-04
GC_11_544 b_11 NI_11 NS_544 0 -2.5374174946470734e-03
GC_11_545 b_11 NI_11 NS_545 0 3.1862102138717149e-04
GC_11_546 b_11 NI_11 NS_546 0 2.1875096644595680e-04
GC_11_547 b_11 NI_11 NS_547 0 -5.0195635069981616e-07
GC_11_548 b_11 NI_11 NS_548 0 1.2291285014505554e-06
GC_11_549 b_11 NI_11 NS_549 0 -2.3042430254087840e-06
GC_11_550 b_11 NI_11 NS_550 0 -4.7508742159571318e-06
GC_11_551 b_11 NI_11 NS_551 0 -9.4393616475078900e-05
GC_11_552 b_11 NI_11 NS_552 0 1.1046320975460251e-04
GC_11_553 b_11 NI_11 NS_553 0 -5.7677931676093864e-06
GC_11_554 b_11 NI_11 NS_554 0 -1.3496240508348845e-05
GC_11_555 b_11 NI_11 NS_555 0 -1.0649463455309622e-05
GC_11_556 b_11 NI_11 NS_556 0 4.9051958911825276e-06
GC_11_557 b_11 NI_11 NS_557 0 2.0406233550438115e-05
GC_11_558 b_11 NI_11 NS_558 0 -4.0948282796928576e-05
GC_11_559 b_11 NI_11 NS_559 0 -4.0245317949986325e-05
GC_11_560 b_11 NI_11 NS_560 0 5.5913555002541536e-05
GC_11_561 b_11 NI_11 NS_561 0 -5.0772961487054340e-02
GC_11_562 b_11 NI_11 NS_562 0 1.5224376253258941e-02
GC_11_563 b_11 NI_11 NS_563 0 4.2187499672109016e-03
GC_11_564 b_11 NI_11 NS_564 0 2.3075883559298301e-03
GC_11_565 b_11 NI_11 NS_565 0 1.2103046144081446e-02
GC_11_566 b_11 NI_11 NS_566 0 7.9888747121904970e-05
GC_11_567 b_11 NI_11 NS_567 0 -3.1889064069330386e-04
GC_11_568 b_11 NI_11 NS_568 0 2.3868906856476129e-03
GC_11_569 b_11 NI_11 NS_569 0 9.6123307655305787e-03
GC_11_570 b_11 NI_11 NS_570 0 8.0077005170669027e-03
GC_11_571 b_11 NI_11 NS_571 0 -1.6241494538064602e-04
GC_11_572 b_11 NI_11 NS_572 0 5.6148884678374064e-04
GC_11_573 b_11 NI_11 NS_573 0 6.1813587309101159e-03
GC_11_574 b_11 NI_11 NS_574 0 -1.3623871077200361e-03
GC_11_575 b_11 NI_11 NS_575 0 5.6249071523234927e-04
GC_11_576 b_11 NI_11 NS_576 0 1.6319666384646116e-03
GC_11_577 b_11 NI_11 NS_577 0 7.2780520235038232e-03
GC_11_578 b_11 NI_11 NS_578 0 2.2078333715034551e-04
GC_11_579 b_11 NI_11 NS_579 0 3.6729869744357409e-03
GC_11_580 b_11 NI_11 NS_580 0 3.9323199306157538e-03
GC_11_581 b_11 NI_11 NS_581 0 2.3087929367515225e-04
GC_11_582 b_11 NI_11 NS_582 0 1.4362727508414073e-04
GC_11_583 b_11 NI_11 NS_583 0 3.3348259629086587e-03
GC_11_584 b_11 NI_11 NS_584 0 6.7019144379874907e-03
GC_11_585 b_11 NI_11 NS_585 0 3.6049044903672348e-04
GC_11_586 b_11 NI_11 NS_586 0 -3.8014454926639253e-05
GC_11_587 b_11 NI_11 NS_587 0 -3.4114014777627085e-04
GC_11_588 b_11 NI_11 NS_588 0 1.7995715191250218e-04
GC_11_589 b_11 NI_11 NS_589 0 5.9332059725329900e-05
GC_11_590 b_11 NI_11 NS_590 0 -6.0391130817080177e-06
GC_11_591 b_11 NI_11 NS_591 0 1.8055665676252228e-05
GC_11_592 b_11 NI_11 NS_592 0 2.8450865731544846e-05
GC_11_593 b_11 NI_11 NS_593 0 -2.0091379497960320e-03
GC_11_594 b_11 NI_11 NS_594 0 6.5446267675931041e-03
GC_11_595 b_11 NI_11 NS_595 0 -1.9022761224583485e-05
GC_11_596 b_11 NI_11 NS_596 0 -3.8837349851228019e-05
GC_11_597 b_11 NI_11 NS_597 0 1.0755593082989912e-03
GC_11_598 b_11 NI_11 NS_598 0 6.2044481612206343e-04
GC_11_599 b_11 NI_11 NS_599 0 -2.3875310230805471e-03
GC_11_600 b_11 NI_11 NS_600 0 9.2281743085889168e-04
GC_11_601 b_11 NI_11 NS_601 0 3.1058008535684710e-04
GC_11_602 b_11 NI_11 NS_602 0 -2.9841937962163509e-04
GC_11_603 b_11 NI_11 NS_603 0 7.5878324720776135e-07
GC_11_604 b_11 NI_11 NS_604 0 -1.0581265382301363e-06
GC_11_605 b_11 NI_11 NS_605 0 1.3558298220649447e-06
GC_11_606 b_11 NI_11 NS_606 0 1.5431288970308875e-05
GC_11_607 b_11 NI_11 NS_607 0 2.8240765922294921e-04
GC_11_608 b_11 NI_11 NS_608 0 -4.8634242050182695e-05
GC_11_609 b_11 NI_11 NS_609 0 -7.9740011292452571e-06
GC_11_610 b_11 NI_11 NS_610 0 2.8259763302418652e-05
GC_11_611 b_11 NI_11 NS_611 0 4.7569974746711494e-06
GC_11_612 b_11 NI_11 NS_612 0 5.7861301016900678e-06
GC_11_613 b_11 NI_11 NS_613 0 -3.6165844994969412e-05
GC_11_614 b_11 NI_11 NS_614 0 1.3284217551213643e-06
GC_11_615 b_11 NI_11 NS_615 0 5.3175011923343299e-05
GC_11_616 b_11 NI_11 NS_616 0 1.8052846051832169e-05
GC_11_617 b_11 NI_11 NS_617 0 -1.3582688543603018e-02
GC_11_618 b_11 NI_11 NS_618 0 1.2052719573683184e-02
GC_11_619 b_11 NI_11 NS_619 0 -2.2105409811907510e-03
GC_11_620 b_11 NI_11 NS_620 0 1.4361170712965466e-03
GC_11_621 b_11 NI_11 NS_621 0 -2.4024962102804463e-03
GC_11_622 b_11 NI_11 NS_622 0 4.3046295243934747e-03
GC_11_623 b_11 NI_11 NS_623 0 -9.6832476723068557e-04
GC_11_624 b_11 NI_11 NS_624 0 -2.9950257363621367e-03
GC_11_625 b_11 NI_11 NS_625 0 -1.1540951782910589e-02
GC_11_626 b_11 NI_11 NS_626 0 -3.3929374347512514e-03
GC_11_627 b_11 NI_11 NS_627 0 4.0235771144579615e-04
GC_11_628 b_11 NI_11 NS_628 0 -2.3373631167318955e-04
GC_11_629 b_11 NI_11 NS_629 0 3.0822927103608525e-03
GC_11_630 b_11 NI_11 NS_630 0 2.4568279926989099e-04
GC_11_631 b_11 NI_11 NS_631 0 9.7006662314307675e-04
GC_11_632 b_11 NI_11 NS_632 0 6.2935537457243281e-04
GC_11_633 b_11 NI_11 NS_633 0 4.2414245204211295e-03
GC_11_634 b_11 NI_11 NS_634 0 -7.3819591364419706e-04
GC_11_635 b_11 NI_11 NS_635 0 -9.9177062919981584e-04
GC_11_636 b_11 NI_11 NS_636 0 5.5664896419994111e-04
GC_11_637 b_11 NI_11 NS_637 0 -1.4686217756825531e-04
GC_11_638 b_11 NI_11 NS_638 0 -4.1170251036942434e-05
GC_11_639 b_11 NI_11 NS_639 0 4.1927311109715409e-03
GC_11_640 b_11 NI_11 NS_640 0 -5.1482646937652714e-04
GC_11_641 b_11 NI_11 NS_641 0 -4.7934897321347031e-04
GC_11_642 b_11 NI_11 NS_642 0 -1.3502170477012920e-04
GC_11_643 b_11 NI_11 NS_643 0 -2.8903556396718056e-04
GC_11_644 b_11 NI_11 NS_644 0 3.3946579639629768e-05
GC_11_645 b_11 NI_11 NS_645 0 -3.0892356186738905e-04
GC_11_646 b_11 NI_11 NS_646 0 1.2919207991281175e-04
GC_11_647 b_11 NI_11 NS_647 0 -1.2520854911123993e-04
GC_11_648 b_11 NI_11 NS_648 0 -7.4553803634481758e-05
GC_11_649 b_11 NI_11 NS_649 0 -1.8094296549237337e-03
GC_11_650 b_11 NI_11 NS_650 0 1.0904116716386862e-04
GC_11_651 b_11 NI_11 NS_651 0 -1.4746037553868653e-05
GC_11_652 b_11 NI_11 NS_652 0 4.6163425205173620e-05
GC_11_653 b_11 NI_11 NS_653 0 -3.2375448057423990e-04
GC_11_654 b_11 NI_11 NS_654 0 -4.5458078684858079e-05
GC_11_655 b_11 NI_11 NS_655 0 1.8163913488087233e-03
GC_11_656 b_11 NI_11 NS_656 0 -1.4661257866595149e-03
GC_11_657 b_11 NI_11 NS_657 0 1.5834016316656834e-04
GC_11_658 b_11 NI_11 NS_658 0 -1.1143955868347852e-04
GC_11_659 b_11 NI_11 NS_659 0 -9.0760877762409660e-07
GC_11_660 b_11 NI_11 NS_660 0 6.9089364221728316e-07
GC_11_661 b_11 NI_11 NS_661 0 -2.6786912533013064e-06
GC_11_662 b_11 NI_11 NS_662 0 -8.4737008856184624e-06
GC_11_663 b_11 NI_11 NS_663 0 -1.4061721522375868e-04
GC_11_664 b_11 NI_11 NS_664 0 1.2145273835873456e-04
GC_11_665 b_11 NI_11 NS_665 0 1.2056782648452022e-06
GC_11_666 b_11 NI_11 NS_666 0 -2.0553622353589295e-05
GC_11_667 b_11 NI_11 NS_667 0 -4.0578785552966013e-06
GC_11_668 b_11 NI_11 NS_668 0 -4.8001861933182968e-06
GC_11_669 b_11 NI_11 NS_669 0 4.8475210125948711e-05
GC_11_670 b_11 NI_11 NS_670 0 -1.5413466340693061e-05
GC_11_671 b_11 NI_11 NS_671 0 -7.4110994691191780e-05
GC_11_672 b_11 NI_11 NS_672 0 5.8610569926976582e-07
GD_11_1 b_11 NI_11 NA_1 0 -4.0811928009381826e-02
GD_11_2 b_11 NI_11 NA_2 0 1.5285228591892604e-02
GD_11_3 b_11 NI_11 NA_3 0 -3.1130932126016350e-02
GD_11_4 b_11 NI_11 NA_4 0 8.5494315936615985e-04
GD_11_5 b_11 NI_11 NA_5 0 1.9851491321331072e-04
GD_11_6 b_11 NI_11 NA_6 0 -1.2049855159266133e-02
GD_11_7 b_11 NI_11 NA_7 0 5.8730314809781244e-03
GD_11_8 b_11 NI_11 NA_8 0 -2.8015666332145639e-02
GD_11_9 b_11 NI_11 NA_9 0 -2.1712256038408526e-02
GD_11_10 b_11 NI_11 NA_10 0 -5.4675147286465671e-02
GD_11_11 b_11 NI_11 NA_11 0 -1.2698775638146620e-01
GD_11_12 b_11 NI_11 NA_12 0 1.1198585681989760e-02
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -7.7620210888908036e-03
GC_12_2 b_12 NI_12 NS_2 0 -9.4331735254411122e-05
GC_12_3 b_12 NI_12 NS_3 0 2.4035115825604120e-04
GC_12_4 b_12 NI_12 NS_4 0 2.9997188130973131e-04
GC_12_5 b_12 NI_12 NS_5 0 -3.6393067352236119e-04
GC_12_6 b_12 NI_12 NS_6 0 2.9345792259039346e-04
GC_12_7 b_12 NI_12 NS_7 0 -1.7710689390550355e-03
GC_12_8 b_12 NI_12 NS_8 0 2.2436576938433586e-04
GC_12_9 b_12 NI_12 NS_9 0 -1.2042529903519995e-03
GC_12_10 b_12 NI_12 NS_10 0 -2.5335848451690408e-03
GC_12_11 b_12 NI_12 NS_11 0 6.1732082219601676e-04
GC_12_12 b_12 NI_12 NS_12 0 -4.9215614304304930e-04
GC_12_13 b_12 NI_12 NS_13 0 7.0860718599519254e-04
GC_12_14 b_12 NI_12 NS_14 0 -1.6586984946247558e-03
GC_12_15 b_12 NI_12 NS_15 0 3.1036444299962731e-04
GC_12_16 b_12 NI_12 NS_16 0 -1.4334112915041509e-04
GC_12_17 b_12 NI_12 NS_17 0 1.2872285744244642e-03
GC_12_18 b_12 NI_12 NS_18 0 9.4271671193662220e-04
GC_12_19 b_12 NI_12 NS_19 0 -4.8374934929042119e-04
GC_12_20 b_12 NI_12 NS_20 0 7.3696491810933649e-04
GC_12_21 b_12 NI_12 NS_21 0 -8.7836481995074269e-05
GC_12_22 b_12 NI_12 NS_22 0 7.6888173462236206e-05
GC_12_23 b_12 NI_12 NS_23 0 -2.7511100083408898e-03
GC_12_24 b_12 NI_12 NS_24 0 -6.7960325354381689e-04
GC_12_25 b_12 NI_12 NS_25 0 -1.7801832521562350e-06
GC_12_26 b_12 NI_12 NS_26 0 5.7095899183566047e-04
GC_12_27 b_12 NI_12 NS_27 0 -3.9126304968056672e-04
GC_12_28 b_12 NI_12 NS_28 0 -7.5098841359395069e-05
GC_12_29 b_12 NI_12 NS_29 0 -3.6757492688338370e-04
GC_12_30 b_12 NI_12 NS_30 0 -1.4754985017801156e-04
GC_12_31 b_12 NI_12 NS_31 0 -6.3669568592464632e-05
GC_12_32 b_12 NI_12 NS_32 0 -9.7178864548363059e-05
GC_12_33 b_12 NI_12 NS_33 0 3.2029717163201861e-03
GC_12_34 b_12 NI_12 NS_34 0 -4.5270884572636439e-03
GC_12_35 b_12 NI_12 NS_35 0 2.0866877919839087e-05
GC_12_36 b_12 NI_12 NS_36 0 4.9503424064614746e-05
GC_12_37 b_12 NI_12 NS_37 0 -9.9415350544241731e-04
GC_12_38 b_12 NI_12 NS_38 0 -4.6610164850692071e-04
GC_12_39 b_12 NI_12 NS_39 0 1.0041225959399780e-03
GC_12_40 b_12 NI_12 NS_40 0 1.6132437760475974e-03
GC_12_41 b_12 NI_12 NS_41 0 -2.5067919362700843e-04
GC_12_42 b_12 NI_12 NS_42 0 1.2755644886259903e-05
GC_12_43 b_12 NI_12 NS_43 0 -1.5638223732613727e-06
GC_12_44 b_12 NI_12 NS_44 0 -1.1825436905827760e-06
GC_12_45 b_12 NI_12 NS_45 0 7.4144411416685196e-06
GC_12_46 b_12 NI_12 NS_46 0 7.1981130207017337e-06
GC_12_47 b_12 NI_12 NS_47 0 -7.1480713803393834e-05
GC_12_48 b_12 NI_12 NS_48 0 -1.6319146682730617e-04
GC_12_49 b_12 NI_12 NS_49 0 1.5574851173462761e-05
GC_12_50 b_12 NI_12 NS_50 0 1.7159357074947135e-05
GC_12_51 b_12 NI_12 NS_51 0 8.4181572052175475e-06
GC_12_52 b_12 NI_12 NS_52 0 -6.4349542198359015e-06
GC_12_53 b_12 NI_12 NS_53 0 5.2095429431654877e-06
GC_12_54 b_12 NI_12 NS_54 0 6.1062621703059984e-05
GC_12_55 b_12 NI_12 NS_55 0 2.0450563760545726e-05
GC_12_56 b_12 NI_12 NS_56 0 -8.8654192363056794e-05
GC_12_57 b_12 NI_12 NS_57 0 6.5332306778115787e-03
GC_12_58 b_12 NI_12 NS_58 0 -4.6004791693850057e-06
GC_12_59 b_12 NI_12 NS_59 0 -2.2451200675510495e-04
GC_12_60 b_12 NI_12 NS_60 0 1.0290603925398588e-05
GC_12_61 b_12 NI_12 NS_61 0 -5.1957644364583647e-06
GC_12_62 b_12 NI_12 NS_62 0 -2.8521714318297447e-04
GC_12_63 b_12 NI_12 NS_63 0 9.2569461080852162e-04
GC_12_64 b_12 NI_12 NS_64 0 -9.7941643978739800e-04
GC_12_65 b_12 NI_12 NS_65 0 1.8408054698003692e-03
GC_12_66 b_12 NI_12 NS_66 0 1.3644773320639696e-03
GC_12_67 b_12 NI_12 NS_67 0 -6.0706432119444001e-04
GC_12_68 b_12 NI_12 NS_68 0 3.6954344488017985e-04
GC_12_69 b_12 NI_12 NS_69 0 -1.6228634437206371e-05
GC_12_70 b_12 NI_12 NS_70 0 1.6181464691972472e-04
GC_12_71 b_12 NI_12 NS_71 0 3.6050867524345268e-04
GC_12_72 b_12 NI_12 NS_72 0 -1.7203513699822986e-04
GC_12_73 b_12 NI_12 NS_73 0 1.5310678048173340e-03
GC_12_74 b_12 NI_12 NS_74 0 1.6236685147749570e-03
GC_12_75 b_12 NI_12 NS_75 0 -4.2217538500454008e-04
GC_12_76 b_12 NI_12 NS_76 0 6.3770821162007157e-06
GC_12_77 b_12 NI_12 NS_77 0 7.1412911020112091e-05
GC_12_78 b_12 NI_12 NS_78 0 8.0109964101388409e-06
GC_12_79 b_12 NI_12 NS_79 0 1.3339226480306484e-03
GC_12_80 b_12 NI_12 NS_80 0 2.3726207126635000e-03
GC_12_81 b_12 NI_12 NS_81 0 -8.7320947498223636e-05
GC_12_82 b_12 NI_12 NS_82 0 1.0173817586033013e-04
GC_12_83 b_12 NI_12 NS_83 0 -2.9829627394241501e-04
GC_12_84 b_12 NI_12 NS_84 0 2.7549361649735113e-04
GC_12_85 b_12 NI_12 NS_85 0 2.6288256347072729e-05
GC_12_86 b_12 NI_12 NS_86 0 -1.7328847209538675e-04
GC_12_87 b_12 NI_12 NS_87 0 1.1221792263805516e-04
GC_12_88 b_12 NI_12 NS_88 0 4.2270672723582549e-05
GC_12_89 b_12 NI_12 NS_89 0 -3.9389346470410343e-03
GC_12_90 b_12 NI_12 NS_90 0 2.5330233660187367e-03
GC_12_91 b_12 NI_12 NS_91 0 -8.1070847226309584e-05
GC_12_92 b_12 NI_12 NS_92 0 2.3559984151666341e-06
GC_12_93 b_12 NI_12 NS_93 0 1.6437105092914051e-03
GC_12_94 b_12 NI_12 NS_94 0 6.6062319480777391e-04
GC_12_95 b_12 NI_12 NS_95 0 -1.3701144339369948e-03
GC_12_96 b_12 NI_12 NS_96 0 -2.7717461229896895e-03
GC_12_97 b_12 NI_12 NS_97 0 -9.2689362392936223e-05
GC_12_98 b_12 NI_12 NS_98 0 3.8985275793168003e-04
GC_12_99 b_12 NI_12 NS_99 0 4.9482637786764230e-06
GC_12_100 b_12 NI_12 NS_100 0 -1.1087045889487686e-06
GC_12_101 b_12 NI_12 NS_101 0 -1.4236523276800744e-05
GC_12_102 b_12 NI_12 NS_102 0 2.4194250673167976e-05
GC_12_103 b_12 NI_12 NS_103 0 2.2701005965862576e-04
GC_12_104 b_12 NI_12 NS_104 0 6.8932487833697385e-05
GC_12_105 b_12 NI_12 NS_105 0 1.8021726190169944e-06
GC_12_106 b_12 NI_12 NS_106 0 3.3011302570015788e-05
GC_12_107 b_12 NI_12 NS_107 0 -1.4465508678414635e-05
GC_12_108 b_12 NI_12 NS_108 0 2.8840373491444537e-05
GC_12_109 b_12 NI_12 NS_109 0 1.3309326230907735e-04
GC_12_110 b_12 NI_12 NS_110 0 -1.2730198132302313e-04
GC_12_111 b_12 NI_12 NS_111 0 -2.3862282960071819e-04
GC_12_112 b_12 NI_12 NS_112 0 1.3943998138669214e-04
GC_12_113 b_12 NI_12 NS_113 0 1.8343209446144047e-03
GC_12_114 b_12 NI_12 NS_114 0 -1.4045422862675989e-04
GC_12_115 b_12 NI_12 NS_115 0 1.7043545740916586e-04
GC_12_116 b_12 NI_12 NS_116 0 5.6335193925879381e-04
GC_12_117 b_12 NI_12 NS_117 0 -5.2540736870445161e-04
GC_12_118 b_12 NI_12 NS_118 0 -8.3983885505418132e-06
GC_12_119 b_12 NI_12 NS_119 0 -1.6439500113466289e-03
GC_12_120 b_12 NI_12 NS_120 0 -2.9679517304435319e-04
GC_12_121 b_12 NI_12 NS_121 0 6.6223652284027126e-04
GC_12_122 b_12 NI_12 NS_122 0 -1.9688513874583907e-03
GC_12_123 b_12 NI_12 NS_123 0 -1.9852777234534010e-04
GC_12_124 b_12 NI_12 NS_124 0 -2.6793605110251754e-04
GC_12_125 b_12 NI_12 NS_125 0 1.2415093807382467e-03
GC_12_126 b_12 NI_12 NS_126 0 -1.2282972748889531e-03
GC_12_127 b_12 NI_12 NS_127 0 7.4733383889148165e-04
GC_12_128 b_12 NI_12 NS_128 0 -2.2160304251825225e-04
GC_12_129 b_12 NI_12 NS_129 0 1.8707857116181297e-03
GC_12_130 b_12 NI_12 NS_130 0 2.0314576518519032e-03
GC_12_131 b_12 NI_12 NS_131 0 -4.3013844366002435e-04
GC_12_132 b_12 NI_12 NS_132 0 2.2303045855767405e-03
GC_12_133 b_12 NI_12 NS_133 0 -1.8781921884161883e-04
GC_12_134 b_12 NI_12 NS_134 0 -1.1098050345309113e-05
GC_12_135 b_12 NI_12 NS_135 0 -1.7978773910389367e-03
GC_12_136 b_12 NI_12 NS_136 0 1.9533684365740508e-03
GC_12_137 b_12 NI_12 NS_137 0 6.4382667788141048e-06
GC_12_138 b_12 NI_12 NS_138 0 2.4502003338103978e-04
GC_12_139 b_12 NI_12 NS_139 0 -6.4434296997731234e-04
GC_12_140 b_12 NI_12 NS_140 0 1.1840981343246712e-04
GC_12_141 b_12 NI_12 NS_141 0 -4.2460554636680888e-04
GC_12_142 b_12 NI_12 NS_142 0 2.4659134874702948e-05
GC_12_143 b_12 NI_12 NS_143 0 -9.2256356567677923e-05
GC_12_144 b_12 NI_12 NS_144 0 -5.5463596042314138e-05
GC_12_145 b_12 NI_12 NS_145 0 -7.9526760555518976e-04
GC_12_146 b_12 NI_12 NS_146 0 -3.2736039530573357e-03
GC_12_147 b_12 NI_12 NS_147 0 2.8720098436919924e-05
GC_12_148 b_12 NI_12 NS_148 0 -7.4296749632867216e-06
GC_12_149 b_12 NI_12 NS_149 0 -7.0063770688764460e-04
GC_12_150 b_12 NI_12 NS_150 0 2.4396799489557358e-04
GC_12_151 b_12 NI_12 NS_151 0 1.2436848992111473e-03
GC_12_152 b_12 NI_12 NS_152 0 -2.9690449212499144e-04
GC_12_153 b_12 NI_12 NS_153 0 -9.2697154098328943e-05
GC_12_154 b_12 NI_12 NS_154 0 1.2856424565501208e-04
GC_12_155 b_12 NI_12 NS_155 0 -1.9757713893937631e-07
GC_12_156 b_12 NI_12 NS_156 0 2.0347467125190327e-07
GC_12_157 b_12 NI_12 NS_157 0 2.7512744182592581e-06
GC_12_158 b_12 NI_12 NS_158 0 3.3178900146236036e-07
GC_12_159 b_12 NI_12 NS_159 0 -6.5912927937445065e-05
GC_12_160 b_12 NI_12 NS_160 0 -2.4386784367653060e-05
GC_12_161 b_12 NI_12 NS_161 0 6.1590259148895468e-06
GC_12_162 b_12 NI_12 NS_162 0 -7.4028698064469236e-07
GC_12_163 b_12 NI_12 NS_163 0 -3.7118713092022863e-06
GC_12_164 b_12 NI_12 NS_164 0 -9.2754915849637076e-07
GC_12_165 b_12 NI_12 NS_165 0 4.8541134545310648e-06
GC_12_166 b_12 NI_12 NS_166 0 -1.0376135443643529e-05
GC_12_167 b_12 NI_12 NS_167 0 -1.4136928671054673e-05
GC_12_168 b_12 NI_12 NS_168 0 1.1979204006438468e-05
GC_12_169 b_12 NI_12 NS_169 0 3.3050164038179626e-03
GC_12_170 b_12 NI_12 NS_170 0 -4.8021178342958023e-05
GC_12_171 b_12 NI_12 NS_171 0 -3.2253134973445719e-04
GC_12_172 b_12 NI_12 NS_172 0 -9.0109417998017669e-05
GC_12_173 b_12 NI_12 NS_173 0 1.7432495012063574e-04
GC_12_174 b_12 NI_12 NS_174 0 -2.5189239076987634e-04
GC_12_175 b_12 NI_12 NS_175 0 1.1631586436919627e-03
GC_12_176 b_12 NI_12 NS_176 0 -5.8183704093168597e-04
GC_12_177 b_12 NI_12 NS_177 0 3.6968073870633118e-04
GC_12_178 b_12 NI_12 NS_178 0 1.8752666597977342e-03
GC_12_179 b_12 NI_12 NS_179 0 -4.4996178209212421e-04
GC_12_180 b_12 NI_12 NS_180 0 9.0295454406147261e-05
GC_12_181 b_12 NI_12 NS_181 0 -4.5856193887273261e-04
GC_12_182 b_12 NI_12 NS_182 0 -4.6462764736863782e-04
GC_12_183 b_12 NI_12 NS_183 0 3.8048480039441855e-04
GC_12_184 b_12 NI_12 NS_184 0 -1.6482054443329899e-04
GC_12_185 b_12 NI_12 NS_185 0 4.1126070893018467e-04
GC_12_186 b_12 NI_12 NS_186 0 1.4706506396174061e-03
GC_12_187 b_12 NI_12 NS_187 0 -6.3405387300786000e-04
GC_12_188 b_12 NI_12 NS_188 0 -6.6990412337130734e-04
GC_12_189 b_12 NI_12 NS_189 0 7.1833917340240080e-05
GC_12_190 b_12 NI_12 NS_190 0 3.2018601183680614e-05
GC_12_191 b_12 NI_12 NS_191 0 1.4017862101919144e-03
GC_12_192 b_12 NI_12 NS_192 0 1.8753689565740192e-04
GC_12_193 b_12 NI_12 NS_193 0 -1.8068547188373793e-04
GC_12_194 b_12 NI_12 NS_194 0 1.6922299123867571e-04
GC_12_195 b_12 NI_12 NS_195 0 -3.1914150012936208e-04
GC_12_196 b_12 NI_12 NS_196 0 2.3487755375658668e-04
GC_12_197 b_12 NI_12 NS_197 0 1.0396678937727660e-05
GC_12_198 b_12 NI_12 NS_198 0 -2.7177462186973107e-04
GC_12_199 b_12 NI_12 NS_199 0 1.1072171978498458e-04
GC_12_200 b_12 NI_12 NS_200 0 1.2352429771210591e-05
GC_12_201 b_12 NI_12 NS_201 0 -1.7674768436040991e-03
GC_12_202 b_12 NI_12 NS_202 0 2.0872659921675370e-03
GC_12_203 b_12 NI_12 NS_203 0 -8.4304222663081005e-05
GC_12_204 b_12 NI_12 NS_204 0 3.0455192690570750e-05
GC_12_205 b_12 NI_12 NS_205 0 1.2855562465062431e-03
GC_12_206 b_12 NI_12 NS_206 0 2.4229830543309145e-04
GC_12_207 b_12 NI_12 NS_207 0 -8.0060001840222728e-04
GC_12_208 b_12 NI_12 NS_208 0 -1.4584233187652797e-03
GC_12_209 b_12 NI_12 NS_209 0 -2.8962714168130014e-04
GC_12_210 b_12 NI_12 NS_210 0 2.9537996650344560e-04
GC_12_211 b_12 NI_12 NS_211 0 2.9394604000579094e-06
GC_12_212 b_12 NI_12 NS_212 0 -5.7075544580261947e-07
GC_12_213 b_12 NI_12 NS_213 0 -9.2653446333024378e-06
GC_12_214 b_12 NI_12 NS_214 0 2.2410213796723229e-05
GC_12_215 b_12 NI_12 NS_215 0 1.1949593111110797e-04
GC_12_216 b_12 NI_12 NS_216 0 -2.3498513873206219e-05
GC_12_217 b_12 NI_12 NS_217 0 1.1983411701721809e-05
GC_12_218 b_12 NI_12 NS_218 0 3.5313486883429270e-05
GC_12_219 b_12 NI_12 NS_219 0 -7.4874820594847156e-06
GC_12_220 b_12 NI_12 NS_220 0 1.7522848921830285e-05
GC_12_221 b_12 NI_12 NS_221 0 1.5235210457751212e-04
GC_12_222 b_12 NI_12 NS_222 0 -7.2559658131738446e-05
GC_12_223 b_12 NI_12 NS_223 0 -2.4512172561037105e-04
GC_12_224 b_12 NI_12 NS_224 0 4.6970785578731683e-05
GC_12_225 b_12 NI_12 NS_225 0 6.3396374328816164e-03
GC_12_226 b_12 NI_12 NS_226 0 -8.1728957910129216e-05
GC_12_227 b_12 NI_12 NS_227 0 -2.0144037165732248e-04
GC_12_228 b_12 NI_12 NS_228 0 7.0102362090007316e-04
GC_12_229 b_12 NI_12 NS_229 0 -3.1311903075123619e-04
GC_12_230 b_12 NI_12 NS_230 0 -6.9060723758361878e-04
GC_12_231 b_12 NI_12 NS_231 0 -5.2943903449684010e-04
GC_12_232 b_12 NI_12 NS_232 0 -8.6696463104411661e-04
GC_12_233 b_12 NI_12 NS_233 0 2.3194356980047164e-03
GC_12_234 b_12 NI_12 NS_234 0 6.6953672877111245e-04
GC_12_235 b_12 NI_12 NS_235 0 -6.5911680172436459e-04
GC_12_236 b_12 NI_12 NS_236 0 1.9484605950108190e-05
GC_12_237 b_12 NI_12 NS_237 0 4.5461546906658983e-04
GC_12_238 b_12 NI_12 NS_238 0 -4.8104261053527343e-04
GC_12_239 b_12 NI_12 NS_239 0 8.5903802954764082e-04
GC_12_240 b_12 NI_12 NS_240 0 -1.1629004717212635e-04
GC_12_241 b_12 NI_12 NS_241 0 6.7811457395275940e-04
GC_12_242 b_12 NI_12 NS_242 0 1.8218282808834375e-03
GC_12_243 b_12 NI_12 NS_243 0 -1.1267491850533726e-03
GC_12_244 b_12 NI_12 NS_244 0 2.5099798084028879e-03
GC_12_245 b_12 NI_12 NS_245 0 -2.0588961261729861e-04
GC_12_246 b_12 NI_12 NS_246 0 -5.3756855947497666e-05
GC_12_247 b_12 NI_12 NS_247 0 -6.4914850498594629e-04
GC_12_248 b_12 NI_12 NS_248 0 1.2846365322550814e-03
GC_12_249 b_12 NI_12 NS_249 0 3.0226115599127335e-05
GC_12_250 b_12 NI_12 NS_250 0 -2.2046284521070860e-05
GC_12_251 b_12 NI_12 NS_251 0 -6.6066231870577728e-04
GC_12_252 b_12 NI_12 NS_252 0 1.0574583008079969e-04
GC_12_253 b_12 NI_12 NS_253 0 -3.8210948574549157e-04
GC_12_254 b_12 NI_12 NS_254 0 4.5381661684489669e-05
GC_12_255 b_12 NI_12 NS_255 0 -1.0256425862846362e-04
GC_12_256 b_12 NI_12 NS_256 0 -3.9347875639297570e-05
GC_12_257 b_12 NI_12 NS_257 0 -5.7161204689873650e-05
GC_12_258 b_12 NI_12 NS_258 0 -2.6254042120030614e-03
GC_12_259 b_12 NI_12 NS_259 0 3.0917671705282903e-05
GC_12_260 b_12 NI_12 NS_260 0 -1.2756421451869834e-05
GC_12_261 b_12 NI_12 NS_261 0 -8.0844593578457209e-04
GC_12_262 b_12 NI_12 NS_262 0 3.6289713315842861e-04
GC_12_263 b_12 NI_12 NS_263 0 6.7660733409714868e-04
GC_12_264 b_12 NI_12 NS_264 0 4.6428108230172385e-04
GC_12_265 b_12 NI_12 NS_265 0 -1.5657969409619922e-04
GC_12_266 b_12 NI_12 NS_266 0 2.6270286674303506e-04
GC_12_267 b_12 NI_12 NS_267 0 -1.1175792809291493e-06
GC_12_268 b_12 NI_12 NS_268 0 4.9603348190470255e-07
GC_12_269 b_12 NI_12 NS_269 0 -6.1675786959972508e-07
GC_12_270 b_12 NI_12 NS_270 0 -5.0943520818267872e-06
GC_12_271 b_12 NI_12 NS_271 0 -1.6473284938108750e-06
GC_12_272 b_12 NI_12 NS_272 0 4.5927091941131259e-05
GC_12_273 b_12 NI_12 NS_273 0 -2.1796196280708479e-06
GC_12_274 b_12 NI_12 NS_274 0 -8.7083990521325944e-06
GC_12_275 b_12 NI_12 NS_275 0 -6.3290605740795360e-06
GC_12_276 b_12 NI_12 NS_276 0 -5.0551545479343289e-06
GC_12_277 b_12 NI_12 NS_277 0 2.2071775737100396e-05
GC_12_278 b_12 NI_12 NS_278 0 -1.1128590064086238e-05
GC_12_279 b_12 NI_12 NS_279 0 -3.8275351949730056e-05
GC_12_280 b_12 NI_12 NS_280 0 5.6072180722480483e-06
GC_12_281 b_12 NI_12 NS_281 0 -2.3410134868427981e-03
GC_12_282 b_12 NI_12 NS_282 0 -1.4592120124549764e-04
GC_12_283 b_12 NI_12 NS_283 0 -2.9574812599211347e-04
GC_12_284 b_12 NI_12 NS_284 0 -2.2219333376224793e-04
GC_12_285 b_12 NI_12 NS_285 0 3.4396351331093458e-04
GC_12_286 b_12 NI_12 NS_286 0 9.8879390522712638e-05
GC_12_287 b_12 NI_12 NS_287 0 6.5727150602828217e-04
GC_12_288 b_12 NI_12 NS_288 0 3.5060643253941650e-04
GC_12_289 b_12 NI_12 NS_289 0 -2.3804550581441406e-03
GC_12_290 b_12 NI_12 NS_290 0 8.6613055194392698e-04
GC_12_291 b_12 NI_12 NS_291 0 4.2805024029062453e-05
GC_12_292 b_12 NI_12 NS_292 0 -1.3746500196035833e-04
GC_12_293 b_12 NI_12 NS_293 0 -4.6578060797320287e-04
GC_12_294 b_12 NI_12 NS_294 0 -1.4216440208704667e-03
GC_12_295 b_12 NI_12 NS_295 0 3.5578243272979694e-04
GC_12_296 b_12 NI_12 NS_296 0 -2.4250780211551137e-04
GC_12_297 b_12 NI_12 NS_297 0 -8.1205697688906337e-04
GC_12_298 b_12 NI_12 NS_298 0 7.9176137443755039e-04
GC_12_299 b_12 NI_12 NS_299 0 -1.0272272853189114e-03
GC_12_300 b_12 NI_12 NS_300 0 -1.2913300692366885e-03
GC_12_301 b_12 NI_12 NS_301 0 1.1282428361609277e-04
GC_12_302 b_12 NI_12 NS_302 0 4.6795616690101154e-05
GC_12_303 b_12 NI_12 NS_303 0 2.1446308426476116e-03
GC_12_304 b_12 NI_12 NS_304 0 -3.3902611692286314e-03
GC_12_305 b_12 NI_12 NS_305 0 -3.1125597857615568e-04
GC_12_306 b_12 NI_12 NS_306 0 3.2872412443036555e-04
GC_12_307 b_12 NI_12 NS_307 0 -2.7674281535003089e-04
GC_12_308 b_12 NI_12 NS_308 0 2.8375751743667021e-04
GC_12_309 b_12 NI_12 NS_309 0 -4.5507978257570927e-05
GC_12_310 b_12 NI_12 NS_310 0 -5.1070189586874325e-04
GC_12_311 b_12 NI_12 NS_311 0 1.9193616919433327e-04
GC_12_312 b_12 NI_12 NS_312 0 -5.1968389223095792e-05
GC_12_313 b_12 NI_12 NS_313 0 5.0559147052410059e-04
GC_12_314 b_12 NI_12 NS_314 0 2.0558406489626022e-03
GC_12_315 b_12 NI_12 NS_315 0 -1.0539427332938129e-04
GC_12_316 b_12 NI_12 NS_316 0 1.0218758455388260e-04
GC_12_317 b_12 NI_12 NS_317 0 1.3877274826665288e-03
GC_12_318 b_12 NI_12 NS_318 0 -5.7087677839141805e-04
GC_12_319 b_12 NI_12 NS_319 0 -8.9845490945059310e-05
GC_12_320 b_12 NI_12 NS_320 0 -8.0107204920748621e-05
GC_12_321 b_12 NI_12 NS_321 0 -4.6426038117257162e-04
GC_12_322 b_12 NI_12 NS_322 0 3.8565921154693226e-04
GC_12_323 b_12 NI_12 NS_323 0 1.1023303886354479e-06
GC_12_324 b_12 NI_12 NS_324 0 -4.6245681066658601e-06
GC_12_325 b_12 NI_12 NS_325 0 -1.5055318432209844e-06
GC_12_326 b_12 NI_12 NS_326 0 3.3036193134449921e-05
GC_12_327 b_12 NI_12 NS_327 0 4.8184089445370427e-05
GC_12_328 b_12 NI_12 NS_328 0 -1.4853572942128418e-04
GC_12_329 b_12 NI_12 NS_329 0 4.1107244786241730e-05
GC_12_330 b_12 NI_12 NS_330 0 4.8683867301205322e-05
GC_12_331 b_12 NI_12 NS_331 0 3.7451952049427309e-06
GC_12_332 b_12 NI_12 NS_332 0 1.9133957983801656e-05
GC_12_333 b_12 NI_12 NS_333 0 2.3198471715608755e-04
GC_12_334 b_12 NI_12 NS_334 0 -1.1083300977561303e-04
GC_12_335 b_12 NI_12 NS_335 0 -3.7076854327113787e-04
GC_12_336 b_12 NI_12 NS_336 0 6.4778805290128169e-05
GC_12_337 b_12 NI_12 NS_337 0 2.6113910399571342e-02
GC_12_338 b_12 NI_12 NS_338 0 -2.8081568320276038e-04
GC_12_339 b_12 NI_12 NS_339 0 -4.7191378253232688e-04
GC_12_340 b_12 NI_12 NS_340 0 5.6101976288285981e-04
GC_12_341 b_12 NI_12 NS_341 0 1.0796920309498769e-03
GC_12_342 b_12 NI_12 NS_342 0 2.3879991425000105e-04
GC_12_343 b_12 NI_12 NS_343 0 -1.1434196351041990e-03
GC_12_344 b_12 NI_12 NS_344 0 9.1466303617449712e-04
GC_12_345 b_12 NI_12 NS_345 0 -2.7851048566762812e-03
GC_12_346 b_12 NI_12 NS_346 0 4.4659259725294415e-03
GC_12_347 b_12 NI_12 NS_347 0 -3.7630184465388465e-04
GC_12_348 b_12 NI_12 NS_348 0 1.1957781522028629e-04
GC_12_349 b_12 NI_12 NS_349 0 5.7688607417157514e-05
GC_12_350 b_12 NI_12 NS_350 0 -1.2281864553701203e-03
GC_12_351 b_12 NI_12 NS_351 0 7.6765881944247021e-04
GC_12_352 b_12 NI_12 NS_352 0 1.3467173557903881e-04
GC_12_353 b_12 NI_12 NS_353 0 -4.5904687874334400e-04
GC_12_354 b_12 NI_12 NS_354 0 6.9709949778275085e-04
GC_12_355 b_12 NI_12 NS_355 0 -1.6687602019112256e-03
GC_12_356 b_12 NI_12 NS_356 0 9.5919841623460080e-04
GC_12_357 b_12 NI_12 NS_357 0 -1.2970759022220012e-04
GC_12_358 b_12 NI_12 NS_358 0 -8.9930709460961253e-05
GC_12_359 b_12 NI_12 NS_359 0 1.3907437472093553e-04
GC_12_360 b_12 NI_12 NS_360 0 2.1918276102564499e-03
GC_12_361 b_12 NI_12 NS_361 0 5.7125449278595826e-05
GC_12_362 b_12 NI_12 NS_362 0 -1.8310638396023477e-04
GC_12_363 b_12 NI_12 NS_363 0 -5.0642899256671920e-04
GC_12_364 b_12 NI_12 NS_364 0 1.5579893702003062e-04
GC_12_365 b_12 NI_12 NS_365 0 -3.0540480418357689e-04
GC_12_366 b_12 NI_12 NS_366 0 1.2386945641440893e-04
GC_12_367 b_12 NI_12 NS_367 0 -9.8125158265745954e-05
GC_12_368 b_12 NI_12 NS_368 0 -1.7925822106646517e-05
GC_12_369 b_12 NI_12 NS_369 0 -1.0666344494844732e-03
GC_12_370 b_12 NI_12 NS_370 0 4.9152476372611048e-04
GC_12_371 b_12 NI_12 NS_371 0 2.7611644512684139e-05
GC_12_372 b_12 NI_12 NS_372 0 -1.8833014962175021e-05
GC_12_373 b_12 NI_12 NS_373 0 -5.0002447538388434e-04
GC_12_374 b_12 NI_12 NS_374 0 4.8131757480424905e-04
GC_12_375 b_12 NI_12 NS_375 0 -1.7105298186990304e-03
GC_12_376 b_12 NI_12 NS_376 0 -1.7722953190666968e-03
GC_12_377 b_12 NI_12 NS_377 0 -1.9516320925251786e-04
GC_12_378 b_12 NI_12 NS_378 0 -6.8472775576534627e-05
GC_12_379 b_12 NI_12 NS_379 0 -8.5581324187006678e-08
GC_12_380 b_12 NI_12 NS_380 0 1.0152563601777610e-06
GC_12_381 b_12 NI_12 NS_381 0 -6.1146546546886989e-06
GC_12_382 b_12 NI_12 NS_382 0 -3.2297373997486933e-06
GC_12_383 b_12 NI_12 NS_383 0 7.4821653403593527e-05
GC_12_384 b_12 NI_12 NS_384 0 1.2540044745899934e-04
GC_12_385 b_12 NI_12 NS_385 0 -8.7626478164911465e-06
GC_12_386 b_12 NI_12 NS_386 0 -1.0173665950323069e-05
GC_12_387 b_12 NI_12 NS_387 0 -3.7344315344784580e-06
GC_12_388 b_12 NI_12 NS_388 0 3.8930408997559795e-06
GC_12_389 b_12 NI_12 NS_389 0 8.0137038747712679e-06
GC_12_390 b_12 NI_12 NS_390 0 -4.3991496038616188e-05
GC_12_391 b_12 NI_12 NS_391 0 -2.9717983490814752e-05
GC_12_392 b_12 NI_12 NS_392 0 6.4752625915311774e-05
GC_12_393 b_12 NI_12 NS_393 0 -9.1923781034077365e-03
GC_12_394 b_12 NI_12 NS_394 0 -3.8938211451338545e-04
GC_12_395 b_12 NI_12 NS_395 0 -2.0088073306983559e-04
GC_12_396 b_12 NI_12 NS_396 0 -2.5626596970541703e-04
GC_12_397 b_12 NI_12 NS_397 0 -4.5221635030294932e-04
GC_12_398 b_12 NI_12 NS_398 0 4.5388850062820567e-04
GC_12_399 b_12 NI_12 NS_399 0 -2.6344463725562700e-04
GC_12_400 b_12 NI_12 NS_400 0 -2.7046631190481840e-04
GC_12_401 b_12 NI_12 NS_401 0 -8.1399467284000871e-04
GC_12_402 b_12 NI_12 NS_402 0 -3.4082571711303959e-03
GC_12_403 b_12 NI_12 NS_403 0 1.6788045223509388e-04
GC_12_404 b_12 NI_12 NS_404 0 1.7526250150235706e-04
GC_12_405 b_12 NI_12 NS_405 0 3.2045654769386048e-04
GC_12_406 b_12 NI_12 NS_406 0 -5.4830393196586395e-04
GC_12_407 b_12 NI_12 NS_407 0 3.3513751138643477e-04
GC_12_408 b_12 NI_12 NS_408 0 -1.7527674756684619e-04
GC_12_409 b_12 NI_12 NS_409 0 -7.2668002061199990e-04
GC_12_410 b_12 NI_12 NS_410 0 -3.5729647473599618e-04
GC_12_411 b_12 NI_12 NS_411 0 -5.4064369337236456e-04
GC_12_412 b_12 NI_12 NS_412 0 -1.6464202148023625e-03
GC_12_413 b_12 NI_12 NS_413 0 3.9572703324257571e-05
GC_12_414 b_12 NI_12 NS_414 0 3.0058013461995800e-05
GC_12_415 b_12 NI_12 NS_415 0 3.8188818093276814e-03
GC_12_416 b_12 NI_12 NS_416 0 -2.4089955777601055e-03
GC_12_417 b_12 NI_12 NS_417 0 -3.0411111979542437e-04
GC_12_418 b_12 NI_12 NS_418 0 1.0299526214415029e-04
GC_12_419 b_12 NI_12 NS_419 0 -1.2627382383437172e-04
GC_12_420 b_12 NI_12 NS_420 0 1.9055209170995498e-04
GC_12_421 b_12 NI_12 NS_421 0 6.8673979440233424e-05
GC_12_422 b_12 NI_12 NS_422 0 -3.5983483095613822e-04
GC_12_423 b_12 NI_12 NS_423 0 1.5424281531755418e-04
GC_12_424 b_12 NI_12 NS_424 0 -3.1182372873420929e-05
GC_12_425 b_12 NI_12 NS_425 0 1.2365757055083563e-03
GC_12_426 b_12 NI_12 NS_426 0 2.0564199013068689e-03
GC_12_427 b_12 NI_12 NS_427 0 -1.0111765128611800e-04
GC_12_428 b_12 NI_12 NS_428 0 4.2923810168964748e-05
GC_12_429 b_12 NI_12 NS_429 0 1.1568680958851129e-03
GC_12_430 b_12 NI_12 NS_430 0 -5.7811228241716722e-04
GC_12_431 b_12 NI_12 NS_431 0 -5.1286801855619037e-05
GC_12_432 b_12 NI_12 NS_432 0 9.0047981688101328e-04
GC_12_433 b_12 NI_12 NS_433 0 -3.6517973885811893e-04
GC_12_434 b_12 NI_12 NS_434 0 -2.3174511402456903e-05
GC_12_435 b_12 NI_12 NS_435 0 1.3099471393441295e-06
GC_12_436 b_12 NI_12 NS_436 0 -2.6250987448429678e-06
GC_12_437 b_12 NI_12 NS_437 0 -5.4500961228866926e-07
GC_12_438 b_12 NI_12 NS_438 0 1.4278614618036190e-05
GC_12_439 b_12 NI_12 NS_439 0 -8.7080612547065100e-05
GC_12_440 b_12 NI_12 NS_440 0 -1.9499223684507147e-04
GC_12_441 b_12 NI_12 NS_441 0 2.4925786637115916e-05
GC_12_442 b_12 NI_12 NS_442 0 3.0063957453144769e-05
GC_12_443 b_12 NI_12 NS_443 0 3.6416934071095278e-06
GC_12_444 b_12 NI_12 NS_444 0 6.3643839087626126e-06
GC_12_445 b_12 NI_12 NS_445 0 1.4328613965143170e-04
GC_12_446 b_12 NI_12 NS_446 0 -3.4079664260207047e-06
GC_12_447 b_12 NI_12 NS_447 0 -2.0326020729252318e-04
GC_12_448 b_12 NI_12 NS_448 0 -4.8355957809481393e-05
GC_12_449 b_12 NI_12 NS_449 0 5.6746496340048330e-02
GC_12_450 b_12 NI_12 NS_450 0 -7.8728806715628425e-04
GC_12_451 b_12 NI_12 NS_451 0 -1.8256131036095411e-03
GC_12_452 b_12 NI_12 NS_452 0 2.2759316103578148e-03
GC_12_453 b_12 NI_12 NS_453 0 2.8300063910072755e-03
GC_12_454 b_12 NI_12 NS_454 0 2.3731408861845689e-04
GC_12_455 b_12 NI_12 NS_455 0 -5.2608056493074736e-03
GC_12_456 b_12 NI_12 NS_456 0 4.7288411081785790e-04
GC_12_457 b_12 NI_12 NS_457 0 -6.0836554097271362e-03
GC_12_458 b_12 NI_12 NS_458 0 1.0464821360320422e-02
GC_12_459 b_12 NI_12 NS_459 0 -6.3081003831635008e-04
GC_12_460 b_12 NI_12 NS_460 0 -8.4396225365583545e-05
GC_12_461 b_12 NI_12 NS_461 0 1.5620587675219432e-03
GC_12_462 b_12 NI_12 NS_462 0 -4.1083484927379749e-03
GC_12_463 b_12 NI_12 NS_463 0 8.2241960170839493e-04
GC_12_464 b_12 NI_12 NS_464 0 1.2136134837889430e-03
GC_12_465 b_12 NI_12 NS_465 0 -1.2742833565039727e-04
GC_12_466 b_12 NI_12 NS_466 0 8.2893525537653453e-04
GC_12_467 b_12 NI_12 NS_467 0 -5.5432921628299978e-03
GC_12_468 b_12 NI_12 NS_468 0 8.0374405703506808e-04
GC_12_469 b_12 NI_12 NS_469 0 -1.1589360712543446e-04
GC_12_470 b_12 NI_12 NS_470 0 -6.4086897278804232e-05
GC_12_471 b_12 NI_12 NS_471 0 7.6761035014766624e-04
GC_12_472 b_12 NI_12 NS_472 0 4.8048080279917537e-03
GC_12_473 b_12 NI_12 NS_473 0 -3.9895006230969752e-04
GC_12_474 b_12 NI_12 NS_474 0 -1.3836698107617382e-04
GC_12_475 b_12 NI_12 NS_475 0 -4.2774098817740597e-04
GC_12_476 b_12 NI_12 NS_476 0 1.5423701391382360e-05
GC_12_477 b_12 NI_12 NS_477 0 -3.9811863573497555e-04
GC_12_478 b_12 NI_12 NS_478 0 3.3411242004342443e-04
GC_12_479 b_12 NI_12 NS_479 0 -1.9656248381834883e-04
GC_12_480 b_12 NI_12 NS_480 0 -4.3232910920391602e-05
GC_12_481 b_12 NI_12 NS_481 0 -6.1049046588566554e-03
GC_12_482 b_12 NI_12 NS_482 0 -1.0187971846521118e-03
GC_12_483 b_12 NI_12 NS_483 0 -3.9046165131515663e-06
GC_12_484 b_12 NI_12 NS_484 0 2.6099896198596828e-05
GC_12_485 b_12 NI_12 NS_485 0 -2.1995136571282430e-04
GC_12_486 b_12 NI_12 NS_486 0 6.0948943844526344e-04
GC_12_487 b_12 NI_12 NS_487 0 -1.1170299443500501e-03
GC_12_488 b_12 NI_12 NS_488 0 -2.2107386660650571e-03
GC_12_489 b_12 NI_12 NS_489 0 5.7628822108007800e-05
GC_12_490 b_12 NI_12 NS_490 0 1.9491593307861664e-04
GC_12_491 b_12 NI_12 NS_491 0 2.2139502980513901e-06
GC_12_492 b_12 NI_12 NS_492 0 -3.0163817874183924e-07
GC_12_493 b_12 NI_12 NS_493 0 -1.6298160766401427e-06
GC_12_494 b_12 NI_12 NS_494 0 -6.1592170161524771e-06
GC_12_495 b_12 NI_12 NS_495 0 -5.4196328522395994e-05
GC_12_496 b_12 NI_12 NS_496 0 3.8239461186475318e-05
GC_12_497 b_12 NI_12 NS_497 0 3.9962968133833772e-07
GC_12_498 b_12 NI_12 NS_498 0 -8.7100510486682304e-06
GC_12_499 b_12 NI_12 NS_499 0 -9.5715923896351318e-07
GC_12_500 b_12 NI_12 NS_500 0 1.1465102965198915e-06
GC_12_501 b_12 NI_12 NS_501 0 6.2297045956352930e-06
GC_12_502 b_12 NI_12 NS_502 0 1.3998296307910532e-05
GC_12_503 b_12 NI_12 NS_503 0 -1.1852031611562295e-06
GC_12_504 b_12 NI_12 NS_504 0 -2.5956778429955234e-05
GC_12_505 b_12 NI_12 NS_505 0 -1.5626950639046160e-02
GC_12_506 b_12 NI_12 NS_506 0 -1.3168205663801260e-03
GC_12_507 b_12 NI_12 NS_507 0 -8.5784258681008635e-04
GC_12_508 b_12 NI_12 NS_508 0 -1.0120647466529513e-03
GC_12_509 b_12 NI_12 NS_509 0 -1.1834877486464276e-03
GC_12_510 b_12 NI_12 NS_510 0 1.3679579038812189e-03
GC_12_511 b_12 NI_12 NS_511 0 8.5002053946312787e-04
GC_12_512 b_12 NI_12 NS_512 0 -7.8518755501043921e-04
GC_12_513 b_12 NI_12 NS_513 0 -3.1542009806871632e-03
GC_12_514 b_12 NI_12 NS_514 0 -8.6413502752804832e-03
GC_12_515 b_12 NI_12 NS_515 0 1.4334396982543137e-04
GC_12_516 b_12 NI_12 NS_516 0 2.9248266007716019e-04
GC_12_517 b_12 NI_12 NS_517 0 1.9539880341976875e-03
GC_12_518 b_12 NI_12 NS_518 0 -2.3240803318479758e-03
GC_12_519 b_12 NI_12 NS_519 0 7.3986093395498850e-04
GC_12_520 b_12 NI_12 NS_520 0 1.7269883996394607e-04
GC_12_521 b_12 NI_12 NS_521 0 9.6201656983432469e-04
GC_12_522 b_12 NI_12 NS_522 0 -1.9843545197027624e-03
GC_12_523 b_12 NI_12 NS_523 0 1.2224896091769246e-03
GC_12_524 b_12 NI_12 NS_524 0 -2.2764590193300850e-03
GC_12_525 b_12 NI_12 NS_525 0 4.0022670476839342e-05
GC_12_526 b_12 NI_12 NS_526 0 8.3464048115653818e-06
GC_12_527 b_12 NI_12 NS_527 0 7.4400237579965185e-03
GC_12_528 b_12 NI_12 NS_528 0 9.9323938492610567e-04
GC_12_529 b_12 NI_12 NS_529 0 -1.2056111177803640e-04
GC_12_530 b_12 NI_12 NS_530 0 4.1547217857400611e-05
GC_12_531 b_12 NI_12 NS_531 0 -1.3571176040844856e-04
GC_12_532 b_12 NI_12 NS_532 0 1.1791348637467000e-04
GC_12_533 b_12 NI_12 NS_533 0 1.8775654067955811e-04
GC_12_534 b_12 NI_12 NS_534 0 -3.8324207868804425e-04
GC_12_535 b_12 NI_12 NS_535 0 3.5053579787666927e-04
GC_12_536 b_12 NI_12 NS_536 0 -1.0949198679205739e-04
GC_12_537 b_12 NI_12 NS_537 0 -7.4695143180155861e-03
GC_12_538 b_12 NI_12 NS_538 0 3.0404032246071347e-03
GC_12_539 b_12 NI_12 NS_539 0 -2.1439477737132123e-04
GC_12_540 b_12 NI_12 NS_540 0 -1.6140356320436272e-04
GC_12_541 b_12 NI_12 NS_541 0 3.8172660632325374e-03
GC_12_542 b_12 NI_12 NS_542 0 4.4515141080264588e-04
GC_12_543 b_12 NI_12 NS_543 0 2.3570074059827101e-03
GC_12_544 b_12 NI_12 NS_544 0 -9.3363739374300952e-04
GC_12_545 b_12 NI_12 NS_545 0 7.5365856719753052e-04
GC_12_546 b_12 NI_12 NS_546 0 3.2995784600048833e-04
GC_12_547 b_12 NI_12 NS_547 0 -2.9544887146721733e-06
GC_12_548 b_12 NI_12 NS_548 0 -4.4539309379425543e-06
GC_12_549 b_12 NI_12 NS_549 0 -1.9883426380242581e-05
GC_12_550 b_12 NI_12 NS_550 0 -4.9842393510479545e-06
GC_12_551 b_12 NI_12 NS_551 0 -3.7260881488049233e-05
GC_12_552 b_12 NI_12 NS_552 0 -7.7416402837702641e-05
GC_12_553 b_12 NI_12 NS_553 0 -2.5277579912296113e-05
GC_12_554 b_12 NI_12 NS_554 0 2.2891817037125896e-06
GC_12_555 b_12 NI_12 NS_555 0 -1.4106412470080935e-05
GC_12_556 b_12 NI_12 NS_556 0 -9.2538625356390421e-06
GC_12_557 b_12 NI_12 NS_557 0 2.3860467510719593e-04
GC_12_558 b_12 NI_12 NS_558 0 -1.3050306293974933e-04
GC_12_559 b_12 NI_12 NS_559 0 -3.9506518624469013e-04
GC_12_560 b_12 NI_12 NS_560 0 9.2451053503181824e-05
GC_12_561 b_12 NI_12 NS_561 0 -1.3582688543638883e-02
GC_12_562 b_12 NI_12 NS_562 0 1.2052719573684938e-02
GC_12_563 b_12 NI_12 NS_563 0 -2.2105409811910915e-03
GC_12_564 b_12 NI_12 NS_564 0 1.4361170712950777e-03
GC_12_565 b_12 NI_12 NS_565 0 -2.4024962102791856e-03
GC_12_566 b_12 NI_12 NS_566 0 4.3046295243924816e-03
GC_12_567 b_12 NI_12 NS_567 0 -9.6832476722736140e-04
GC_12_568 b_12 NI_12 NS_568 0 -2.9950257363639409e-03
GC_12_569 b_12 NI_12 NS_569 0 -1.1540951782906600e-02
GC_12_570 b_12 NI_12 NS_570 0 -3.3929374347532472e-03
GC_12_571 b_12 NI_12 NS_571 0 4.0235771144307773e-04
GC_12_572 b_12 NI_12 NS_572 0 -2.3373631166888678e-04
GC_12_573 b_12 NI_12 NS_573 0 3.0822927103627499e-03
GC_12_574 b_12 NI_12 NS_574 0 2.4568279926876190e-04
GC_12_575 b_12 NI_12 NS_575 0 9.7006662314289211e-04
GC_12_576 b_12 NI_12 NS_576 0 6.2935537457196454e-04
GC_12_577 b_12 NI_12 NS_577 0 4.2414245204239701e-03
GC_12_578 b_12 NI_12 NS_578 0 -7.3819591364714153e-04
GC_12_579 b_12 NI_12 NS_579 0 -9.9177062919734971e-04
GC_12_580 b_12 NI_12 NS_580 0 5.5664896419894267e-04
GC_12_581 b_12 NI_12 NS_581 0 -1.4686217756839989e-04
GC_12_582 b_12 NI_12 NS_582 0 -4.1170251036843250e-05
GC_12_583 b_12 NI_12 NS_583 0 4.1927311109807150e-03
GC_12_584 b_12 NI_12 NS_584 0 -5.1482646937867874e-04
GC_12_585 b_12 NI_12 NS_585 0 -4.7934897321423109e-04
GC_12_586 b_12 NI_12 NS_586 0 -1.3502170477016796e-04
GC_12_587 b_12 NI_12 NS_587 0 -2.8903556396687406e-04
GC_12_588 b_12 NI_12 NS_588 0 3.3946579639865352e-05
GC_12_589 b_12 NI_12 NS_589 0 -3.0892356186701598e-04
GC_12_590 b_12 NI_12 NS_590 0 1.2919207991262335e-04
GC_12_591 b_12 NI_12 NS_591 0 -1.2520854911108128e-04
GC_12_592 b_12 NI_12 NS_592 0 -7.4553803634474535e-05
GC_12_593 b_12 NI_12 NS_593 0 -1.8094296549172680e-03
GC_12_594 b_12 NI_12 NS_594 0 1.0904116717278156e-04
GC_12_595 b_12 NI_12 NS_595 0 -1.4746037553992392e-05
GC_12_596 b_12 NI_12 NS_596 0 4.6163425205179346e-05
GC_12_597 b_12 NI_12 NS_597 0 -3.2375448057281932e-04
GC_12_598 b_12 NI_12 NS_598 0 -4.5458078686335487e-05
GC_12_599 b_12 NI_12 NS_599 0 1.8163913488044576e-03
GC_12_600 b_12 NI_12 NS_600 0 -1.4661257866545932e-03
GC_12_601 b_12 NI_12 NS_601 0 1.5834016316654357e-04
GC_12_602 b_12 NI_12 NS_602 0 -1.1143955868378034e-04
GC_12_603 b_12 NI_12 NS_603 0 -9.0760877762468836e-07
GC_12_604 b_12 NI_12 NS_604 0 6.9089364221468414e-07
GC_12_605 b_12 NI_12 NS_605 0 -2.6786912532858383e-06
GC_12_606 b_12 NI_12 NS_606 0 -8.4737008856013032e-06
GC_12_607 b_12 NI_12 NS_607 0 -1.4061721522363554e-04
GC_12_608 b_12 NI_12 NS_608 0 1.2145273835835458e-04
GC_12_609 b_12 NI_12 NS_609 0 1.2056782648677182e-06
GC_12_610 b_12 NI_12 NS_610 0 -2.0553622353550911e-05
GC_12_611 b_12 NI_12 NS_611 0 -4.0578785552736805e-06
GC_12_612 b_12 NI_12 NS_612 0 -4.8001861933311666e-06
GC_12_613 b_12 NI_12 NS_613 0 4.8475210125941887e-05
GC_12_614 b_12 NI_12 NS_614 0 -1.5413466340581151e-05
GC_12_615 b_12 NI_12 NS_615 0 -7.4110994691130061e-05
GC_12_616 b_12 NI_12 NS_616 0 5.8610569910796813e-07
GC_12_617 b_12 NI_12 NS_617 0 -8.9312602649792419e-02
GC_12_618 b_12 NI_12 NS_618 0 8.0946383714470601e-03
GC_12_619 b_12 NI_12 NS_619 0 -1.4967636815768918e-04
GC_12_620 b_12 NI_12 NS_620 0 -1.2210924605534090e-03
GC_12_621 b_12 NI_12 NS_621 0 -1.1860367299786410e-03
GC_12_622 b_12 NI_12 NS_622 0 -1.4005686707455583e-03
GC_12_623 b_12 NI_12 NS_623 0 1.6344971057812476e-03
GC_12_624 b_12 NI_12 NS_624 0 2.7039939064248766e-03
GC_12_625 b_12 NI_12 NS_625 0 8.8363914349123898e-03
GC_12_626 b_12 NI_12 NS_626 0 7.7367744929187433e-05
GC_12_627 b_12 NI_12 NS_627 0 7.6828317656542475e-04
GC_12_628 b_12 NI_12 NS_628 0 -7.8080936695229812e-04
GC_12_629 b_12 NI_12 NS_629 0 -9.4907127295546022e-04
GC_12_630 b_12 NI_12 NS_630 0 -2.4481084833010845e-03
GC_12_631 b_12 NI_12 NS_631 0 5.1822551954714628e-04
GC_12_632 b_12 NI_12 NS_632 0 1.7648183813237129e-04
GC_12_633 b_12 NI_12 NS_633 0 1.5009070460137903e-04
GC_12_634 b_12 NI_12 NS_634 0 -1.4178789522131254e-03
GC_12_635 b_12 NI_12 NS_635 0 1.0242871092240593e-03
GC_12_636 b_12 NI_12 NS_636 0 -1.7078757582893388e-03
GC_12_637 b_12 NI_12 NS_637 0 3.8553486523568416e-05
GC_12_638 b_12 NI_12 NS_638 0 -1.4749522111260886e-05
GC_12_639 b_12 NI_12 NS_639 0 3.1746039831607410e-03
GC_12_640 b_12 NI_12 NS_640 0 1.5034801824281041e-03
GC_12_641 b_12 NI_12 NS_641 0 -1.8573984037385840e-05
GC_12_642 b_12 NI_12 NS_642 0 -3.1667327253650130e-05
GC_12_643 b_12 NI_12 NS_643 0 -1.6545586532468661e-04
GC_12_644 b_12 NI_12 NS_644 0 1.0461491194118492e-04
GC_12_645 b_12 NI_12 NS_645 0 1.5063087976755038e-04
GC_12_646 b_12 NI_12 NS_646 0 -1.9442900614526816e-04
GC_12_647 b_12 NI_12 NS_647 0 2.1123050391258860e-04
GC_12_648 b_12 NI_12 NS_648 0 -1.1886647935414002e-05
GC_12_649 b_12 NI_12 NS_649 0 -5.5720565005182576e-03
GC_12_650 b_12 NI_12 NS_650 0 1.8275178204841638e-03
GC_12_651 b_12 NI_12 NS_651 0 -1.2238521374009951e-04
GC_12_652 b_12 NI_12 NS_652 0 -1.1075603994419851e-04
GC_12_653 b_12 NI_12 NS_653 0 2.4179521737174086e-03
GC_12_654 b_12 NI_12 NS_654 0 6.6594364224253964e-04
GC_12_655 b_12 NI_12 NS_655 0 1.8060961614659820e-03
GC_12_656 b_12 NI_12 NS_656 0 -8.6493763770677332e-04
GC_12_657 b_12 NI_12 NS_657 0 4.8305259841672474e-04
GC_12_658 b_12 NI_12 NS_658 0 8.5870506285684047e-05
GC_12_659 b_12 NI_12 NS_659 0 -3.1165917544987164e-07
GC_12_660 b_12 NI_12 NS_660 0 -1.5529148363557479e-06
GC_12_661 b_12 NI_12 NS_661 0 -8.6307810906398913e-06
GC_12_662 b_12 NI_12 NS_662 0 8.6215540052152303e-07
GC_12_663 b_12 NI_12 NS_663 0 -1.8932914327643906e-05
GC_12_664 b_12 NI_12 NS_664 0 -1.1653093317863102e-04
GC_12_665 b_12 NI_12 NS_665 0 -1.2187541833100157e-05
GC_12_666 b_12 NI_12 NS_666 0 6.5368884734210508e-06
GC_12_667 b_12 NI_12 NS_667 0 -9.1202394846432207e-06
GC_12_668 b_12 NI_12 NS_668 0 6.4713251647361220e-06
GC_12_669 b_12 NI_12 NS_669 0 1.1177832148706337e-04
GC_12_670 b_12 NI_12 NS_670 0 -5.0656196300422251e-05
GC_12_671 b_12 NI_12 NS_671 0 -1.7997576078059824e-04
GC_12_672 b_12 NI_12 NS_672 0 3.8915745221929917e-05
GD_12_1 b_12 NI_12 NA_1 0 1.7846885875163806e-02
GD_12_2 b_12 NI_12 NA_2 0 -1.2519126254091678e-02
GD_12_3 b_12 NI_12 NA_3 0 1.3438244043457396e-03
GD_12_4 b_12 NI_12 NA_4 0 -5.4585833604317915e-03
GD_12_5 b_12 NI_12 NA_5 0 -9.3557202206591937e-03
GD_12_6 b_12 NI_12 NA_6 0 5.0915336871086049e-03
GD_12_7 b_12 NI_12 NA_7 0 -2.7059768597434423e-02
GD_12_8 b_12 NI_12 NA_8 0 8.8545031458948324e-03
GD_12_9 b_12 NI_12 NA_9 0 -5.3530411270550728e-02
GD_12_10 b_12 NI_12 NA_10 0 1.1228841767502927e-02
GD_12_11 b_12 NI_12 NA_11 0 1.1198585682005172e-02
GD_12_12 b_12 NI_12 NA_12 0 1.2792535672851610e-01
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 4.1362120035729779e+00
GS_1_1 0 NS_1 NA_1 0 1.3803457954163372e+00
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 2.7078253238558993e+01
GS_2_1 0 NS_2 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 3/4
CS_3 NS_3 0 9.9999999999999998e-13
CS_4 NS_4 0 9.9999999999999998e-13
RS_3 NS_3 0 5.6873212206500213e+01
RS_4 NS_4 0 5.6873212206500220e+01
GL_3 0 NS_3 NS_4 0 4.7960934964359665e-02
GL_4 0 NS_4 NS_3 0 -4.7960934964359665e-02
GS_3_1 0 NS_3 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 5.5832282069998371e+01
RS_6 NS_6 0 5.5832282069998378e+01
GL_5 0 NS_5 NS_6 0 6.1612202840267971e-02
GL_6 0 NS_6 NS_5 0 -6.1612202840267971e-02
GS_5_1 0 NS_5 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 3.4747519722663924e+01
RS_8 NS_8 0 3.4747519722663924e+01
GL_7 0 NS_7 NS_8 0 8.1784427745819094e-02
GL_8 0 NS_8 NS_7 0 -8.1784427745819094e-02
GS_7_1 0 NS_7 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 3.1454928782186034e+01
RS_10 NS_10 0 3.1454928782186034e+01
GL_9 0 NS_9 NS_10 0 1.1192538378623762e-01
GL_10 0 NS_10 NS_9 0 -1.1192538378623762e-01
GS_9_1 0 NS_9 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 2.2209312435826621e+02
RS_12 NS_12 0 2.2209312435826621e+02
GL_11 0 NS_11 NS_12 0 2.9133579865504960e-01
GL_12 0 NS_12 NS_11 0 -2.9133579865504960e-01
GS_11_1 0 NS_11 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 4.4403718965615290e+01
RS_14 NS_14 0 4.4403718965615283e+01
GL_13 0 NS_13 NS_14 0 1.3869030610195973e-01
GL_14 0 NS_14 NS_13 0 -1.3869030610195973e-01
GS_13_1 0 NS_13 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 9.2436417727653946e+01
RS_16 NS_16 0 9.2436417727653946e+01
GL_15 0 NS_15 NS_16 0 1.6009535907039132e-01
GL_16 0 NS_16 NS_15 0 -1.6009535907039132e-01
GS_15_1 0 NS_15 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 5.2247674424140278e+01
RS_18 NS_18 0 5.2247674424140278e+01
GL_17 0 NS_17 NS_18 0 1.7061294296414609e-01
GL_18 0 NS_18 NS_17 0 -1.7061294296414609e-01
GS_17_1 0 NS_17 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 6.3351631924882277e+01
RS_20 NS_20 0 6.3351631924882277e+01
GL_19 0 NS_19 NS_20 0 1.8578563768540060e-01
GL_20 0 NS_20 NS_19 0 -1.8578563768540060e-01
GS_19_1 0 NS_19 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 2.2461363612924958e+02
RS_22 NS_22 0 2.2461363612924956e+02
GL_21 0 NS_21 NS_22 0 2.0090890151880786e-01
GL_22 0 NS_22 NS_21 0 -2.0090890151880786e-01
GS_21_1 0 NS_21 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 6.2323563035856608e+01
RS_24 NS_24 0 6.2323563035856608e+01
GL_23 0 NS_23 NS_24 0 2.0741858581422049e-01
GL_24 0 NS_24 NS_23 0 -2.0741858581422049e-01
GS_23_1 0 NS_23 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 1.5742148578820314e+02
RS_26 NS_26 0 1.5742148578820311e+02
GL_25 0 NS_25 NS_26 0 2.0543767879537947e-01
GL_26 0 NS_26 NS_25 0 -2.0543767879537947e-01
GS_25_1 0 NS_25 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 2.0165146427356075e+02
RS_28 NS_28 0 2.0165146427356075e+02
GL_27 0 NS_27 NS_28 0 2.1530071526798281e-01
GL_28 0 NS_28 NS_27 0 -2.1530071526798281e-01
GS_27_1 0 NS_27 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 2.5655383475382814e+02
RS_30 NS_30 0 2.5655383475382814e+02
GL_29 0 NS_29 NS_30 0 2.2143554872154964e-01
GL_30 0 NS_30 NS_29 0 -2.2143554872154964e-01
GS_29_1 0 NS_29 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 3.7527533273924564e+02
RS_32 NS_32 0 3.7527533273924570e+02
GL_31 0 NS_31 NS_32 0 2.2416553875794559e-01
GL_32 0 NS_32 NS_31 0 -2.2416553875794559e-01
GS_31_1 0 NS_31 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 8.7633211379679196e+01
RS_34 NS_34 0 8.7633211379679196e+01
GL_33 0 NS_33 NS_34 0 2.3541329178654702e-01
GL_34 0 NS_34 NS_33 0 -2.3541329178654702e-01
GS_33_1 0 NS_33 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 4.0937268842404592e+02
RS_36 NS_36 0 4.0937268842404586e+02
GL_35 0 NS_35 NS_36 0 2.2933880932778705e-01
GL_36 0 NS_36 NS_35 0 -2.2933880932778705e-01
GS_35_1 0 NS_35 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 1.8046101089657725e+02
RS_38 NS_38 0 1.8046101089657725e+02
GL_37 0 NS_37 NS_38 0 2.3011433813523779e-01
GL_38 0 NS_38 NS_37 0 -2.3011433813523779e-01
GS_37_1 0 NS_37 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 9.7664924917686449e+01
RS_40 NS_40 0 9.7664924917686449e+01
GL_39 0 NS_39 NS_40 0 2.4746563775454208e-01
GL_40 0 NS_40 NS_39 0 -2.4746563775454208e-01
GS_39_1 0 NS_39 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 2.6057215108102395e+02
RS_42 NS_42 0 2.6057215108102395e+02
GL_41 0 NS_41 NS_42 0 2.3565487776505958e-01
GL_42 0 NS_42 NS_41 0 -2.3565487776505958e-01
GS_41_1 0 NS_41 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 1.4688638444267465e+03
RS_44 NS_44 0 1.4688638444267465e+03
GL_43 0 NS_43 NS_44 0 2.3814510332638331e-01
GL_44 0 NS_44 NS_43 0 -2.3814510332638331e-01
GS_43_1 0 NS_43 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 1.5351229021400181e+03
RS_46 NS_46 0 1.5351229021400181e+03
GL_45 0 NS_45 NS_46 0 2.5027181856001052e-01
GL_46 0 NS_46 NS_45 0 -2.5027181856001052e-01
GS_45_1 0 NS_45 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 4.3650646405920685e+02
RS_48 NS_48 0 4.3650646405920685e+02
GL_47 0 NS_47 NS_48 0 2.4893599896984003e-01
GL_48 0 NS_48 NS_47 0 -2.4893599896984003e-01
GS_47_1 0 NS_47 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 1.1441811687773074e+03
RS_50 NS_50 0 1.1441811687773072e+03
GL_49 0 NS_49 NS_50 0 2.4916499611033449e-01
GL_50 0 NS_50 NS_49 0 -2.4916499611033449e-01
GS_49_1 0 NS_49 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 7.5335118532932768e+02
RS_52 NS_52 0 7.5335118532932768e+02
GL_51 0 NS_51 NS_52 0 2.4298312011423853e-01
GL_52 0 NS_52 NS_51 0 -2.4298312011423853e-01
GS_51_1 0 NS_51 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 1.1346596293114915e+03
RS_54 NS_54 0 1.1346596293114915e+03
GL_53 0 NS_53 NS_54 0 2.4551048269503753e-01
GL_54 0 NS_54 NS_53 0 -2.4551048269503753e-01
GS_53_1 0 NS_53 NA_1 0 1.3803457954163372e+00
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 9.3517666338196523e+02
RS_56 NS_56 0 9.3517666338196523e+02
GL_55 0 NS_55 NS_56 0 2.4538280909205379e-01
GL_56 0 NS_56 NS_55 0 -2.4538280909205379e-01
GS_55_1 0 NS_55 NA_1 0 1.3803457954163372e+00
*
* Real pole n. 57
CS_57 NS_57 0 9.9999999999999998e-13
RS_57 NS_57 0 4.1362120035729779e+00
GS_57_2 0 NS_57 NA_2 0 1.3803457954163372e+00
*
* Real pole n. 58
CS_58 NS_58 0 9.9999999999999998e-13
RS_58 NS_58 0 2.7078253238558993e+01
GS_58_2 0 NS_58 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 5.6873212206500213e+01
RS_60 NS_60 0 5.6873212206500220e+01
GL_59 0 NS_59 NS_60 0 4.7960934964359665e-02
GL_60 0 NS_60 NS_59 0 -4.7960934964359665e-02
GS_59_2 0 NS_59 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 5.5832282069998371e+01
RS_62 NS_62 0 5.5832282069998378e+01
GL_61 0 NS_61 NS_62 0 6.1612202840267971e-02
GL_62 0 NS_62 NS_61 0 -6.1612202840267971e-02
GS_61_2 0 NS_61 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 3.4747519722663924e+01
RS_64 NS_64 0 3.4747519722663924e+01
GL_63 0 NS_63 NS_64 0 8.1784427745819094e-02
GL_64 0 NS_64 NS_63 0 -8.1784427745819094e-02
GS_63_2 0 NS_63 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 3.1454928782186034e+01
RS_66 NS_66 0 3.1454928782186034e+01
GL_65 0 NS_65 NS_66 0 1.1192538378623762e-01
GL_66 0 NS_66 NS_65 0 -1.1192538378623762e-01
GS_65_2 0 NS_65 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 2.2209312435826621e+02
RS_68 NS_68 0 2.2209312435826621e+02
GL_67 0 NS_67 NS_68 0 2.9133579865504960e-01
GL_68 0 NS_68 NS_67 0 -2.9133579865504960e-01
GS_67_2 0 NS_67 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 4.4403718965615290e+01
RS_70 NS_70 0 4.4403718965615283e+01
GL_69 0 NS_69 NS_70 0 1.3869030610195973e-01
GL_70 0 NS_70 NS_69 0 -1.3869030610195973e-01
GS_69_2 0 NS_69 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 9.2436417727653946e+01
RS_72 NS_72 0 9.2436417727653946e+01
GL_71 0 NS_71 NS_72 0 1.6009535907039132e-01
GL_72 0 NS_72 NS_71 0 -1.6009535907039132e-01
GS_71_2 0 NS_71 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 5.2247674424140278e+01
RS_74 NS_74 0 5.2247674424140278e+01
GL_73 0 NS_73 NS_74 0 1.7061294296414609e-01
GL_74 0 NS_74 NS_73 0 -1.7061294296414609e-01
GS_73_2 0 NS_73 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 6.3351631924882277e+01
RS_76 NS_76 0 6.3351631924882277e+01
GL_75 0 NS_75 NS_76 0 1.8578563768540060e-01
GL_76 0 NS_76 NS_75 0 -1.8578563768540060e-01
GS_75_2 0 NS_75 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 2.2461363612924958e+02
RS_78 NS_78 0 2.2461363612924956e+02
GL_77 0 NS_77 NS_78 0 2.0090890151880786e-01
GL_78 0 NS_78 NS_77 0 -2.0090890151880786e-01
GS_77_2 0 NS_77 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 6.2323563035856608e+01
RS_80 NS_80 0 6.2323563035856608e+01
GL_79 0 NS_79 NS_80 0 2.0741858581422049e-01
GL_80 0 NS_80 NS_79 0 -2.0741858581422049e-01
GS_79_2 0 NS_79 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 1.5742148578820314e+02
RS_82 NS_82 0 1.5742148578820311e+02
GL_81 0 NS_81 NS_82 0 2.0543767879537947e-01
GL_82 0 NS_82 NS_81 0 -2.0543767879537947e-01
GS_81_2 0 NS_81 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 2.0165146427356075e+02
RS_84 NS_84 0 2.0165146427356075e+02
GL_83 0 NS_83 NS_84 0 2.1530071526798281e-01
GL_84 0 NS_84 NS_83 0 -2.1530071526798281e-01
GS_83_2 0 NS_83 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 2.5655383475382814e+02
RS_86 NS_86 0 2.5655383475382814e+02
GL_85 0 NS_85 NS_86 0 2.2143554872154964e-01
GL_86 0 NS_86 NS_85 0 -2.2143554872154964e-01
GS_85_2 0 NS_85 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 3.7527533273924564e+02
RS_88 NS_88 0 3.7527533273924570e+02
GL_87 0 NS_87 NS_88 0 2.2416553875794559e-01
GL_88 0 NS_88 NS_87 0 -2.2416553875794559e-01
GS_87_2 0 NS_87 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 8.7633211379679196e+01
RS_90 NS_90 0 8.7633211379679196e+01
GL_89 0 NS_89 NS_90 0 2.3541329178654702e-01
GL_90 0 NS_90 NS_89 0 -2.3541329178654702e-01
GS_89_2 0 NS_89 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 4.0937268842404592e+02
RS_92 NS_92 0 4.0937268842404586e+02
GL_91 0 NS_91 NS_92 0 2.2933880932778705e-01
GL_92 0 NS_92 NS_91 0 -2.2933880932778705e-01
GS_91_2 0 NS_91 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 1.8046101089657725e+02
RS_94 NS_94 0 1.8046101089657725e+02
GL_93 0 NS_93 NS_94 0 2.3011433813523779e-01
GL_94 0 NS_94 NS_93 0 -2.3011433813523779e-01
GS_93_2 0 NS_93 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 9.7664924917686449e+01
RS_96 NS_96 0 9.7664924917686449e+01
GL_95 0 NS_95 NS_96 0 2.4746563775454208e-01
GL_96 0 NS_96 NS_95 0 -2.4746563775454208e-01
GS_95_2 0 NS_95 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 2.6057215108102395e+02
RS_98 NS_98 0 2.6057215108102395e+02
GL_97 0 NS_97 NS_98 0 2.3565487776505958e-01
GL_98 0 NS_98 NS_97 0 -2.3565487776505958e-01
GS_97_2 0 NS_97 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 1.4688638444267465e+03
RS_100 NS_100 0 1.4688638444267465e+03
GL_99 0 NS_99 NS_100 0 2.3814510332638331e-01
GL_100 0 NS_100 NS_99 0 -2.3814510332638331e-01
GS_99_2 0 NS_99 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 1.5351229021400181e+03
RS_102 NS_102 0 1.5351229021400181e+03
GL_101 0 NS_101 NS_102 0 2.5027181856001052e-01
GL_102 0 NS_102 NS_101 0 -2.5027181856001052e-01
GS_101_2 0 NS_101 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 4.3650646405920685e+02
RS_104 NS_104 0 4.3650646405920685e+02
GL_103 0 NS_103 NS_104 0 2.4893599896984003e-01
GL_104 0 NS_104 NS_103 0 -2.4893599896984003e-01
GS_103_2 0 NS_103 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 1.1441811687773074e+03
RS_106 NS_106 0 1.1441811687773072e+03
GL_105 0 NS_105 NS_106 0 2.4916499611033449e-01
GL_106 0 NS_106 NS_105 0 -2.4916499611033449e-01
GS_105_2 0 NS_105 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 7.5335118532932768e+02
RS_108 NS_108 0 7.5335118532932768e+02
GL_107 0 NS_107 NS_108 0 2.4298312011423853e-01
GL_108 0 NS_108 NS_107 0 -2.4298312011423853e-01
GS_107_2 0 NS_107 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 1.1346596293114915e+03
RS_110 NS_110 0 1.1346596293114915e+03
GL_109 0 NS_109 NS_110 0 2.4551048269503753e-01
GL_110 0 NS_110 NS_109 0 -2.4551048269503753e-01
GS_109_2 0 NS_109 NA_2 0 1.3803457954163372e+00
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 9.3517666338196523e+02
RS_112 NS_112 0 9.3517666338196523e+02
GL_111 0 NS_111 NS_112 0 2.4538280909205379e-01
GL_112 0 NS_112 NS_111 0 -2.4538280909205379e-01
GS_111_2 0 NS_111 NA_2 0 1.3803457954163372e+00
*
* Real pole n. 113
CS_113 NS_113 0 9.9999999999999998e-13
RS_113 NS_113 0 4.1362120035729779e+00
GS_113_3 0 NS_113 NA_3 0 1.3803457954163372e+00
*
* Real pole n. 114
CS_114 NS_114 0 9.9999999999999998e-13
RS_114 NS_114 0 2.7078253238558993e+01
GS_114_3 0 NS_114 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 5.6873212206500213e+01
RS_116 NS_116 0 5.6873212206500220e+01
GL_115 0 NS_115 NS_116 0 4.7960934964359665e-02
GL_116 0 NS_116 NS_115 0 -4.7960934964359665e-02
GS_115_3 0 NS_115 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 5.5832282069998371e+01
RS_118 NS_118 0 5.5832282069998378e+01
GL_117 0 NS_117 NS_118 0 6.1612202840267971e-02
GL_118 0 NS_118 NS_117 0 -6.1612202840267971e-02
GS_117_3 0 NS_117 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 3.4747519722663924e+01
RS_120 NS_120 0 3.4747519722663924e+01
GL_119 0 NS_119 NS_120 0 8.1784427745819094e-02
GL_120 0 NS_120 NS_119 0 -8.1784427745819094e-02
GS_119_3 0 NS_119 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 3.1454928782186034e+01
RS_122 NS_122 0 3.1454928782186034e+01
GL_121 0 NS_121 NS_122 0 1.1192538378623762e-01
GL_122 0 NS_122 NS_121 0 -1.1192538378623762e-01
GS_121_3 0 NS_121 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 2.2209312435826621e+02
RS_124 NS_124 0 2.2209312435826621e+02
GL_123 0 NS_123 NS_124 0 2.9133579865504960e-01
GL_124 0 NS_124 NS_123 0 -2.9133579865504960e-01
GS_123_3 0 NS_123 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 4.4403718965615290e+01
RS_126 NS_126 0 4.4403718965615283e+01
GL_125 0 NS_125 NS_126 0 1.3869030610195973e-01
GL_126 0 NS_126 NS_125 0 -1.3869030610195973e-01
GS_125_3 0 NS_125 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 9.2436417727653946e+01
RS_128 NS_128 0 9.2436417727653946e+01
GL_127 0 NS_127 NS_128 0 1.6009535907039132e-01
GL_128 0 NS_128 NS_127 0 -1.6009535907039132e-01
GS_127_3 0 NS_127 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 5.2247674424140278e+01
RS_130 NS_130 0 5.2247674424140278e+01
GL_129 0 NS_129 NS_130 0 1.7061294296414609e-01
GL_130 0 NS_130 NS_129 0 -1.7061294296414609e-01
GS_129_3 0 NS_129 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 6.3351631924882277e+01
RS_132 NS_132 0 6.3351631924882277e+01
GL_131 0 NS_131 NS_132 0 1.8578563768540060e-01
GL_132 0 NS_132 NS_131 0 -1.8578563768540060e-01
GS_131_3 0 NS_131 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 133/134
CS_133 NS_133 0 9.9999999999999998e-13
CS_134 NS_134 0 9.9999999999999998e-13
RS_133 NS_133 0 2.2461363612924958e+02
RS_134 NS_134 0 2.2461363612924956e+02
GL_133 0 NS_133 NS_134 0 2.0090890151880786e-01
GL_134 0 NS_134 NS_133 0 -2.0090890151880786e-01
GS_133_3 0 NS_133 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 6.2323563035856608e+01
RS_136 NS_136 0 6.2323563035856608e+01
GL_135 0 NS_135 NS_136 0 2.0741858581422049e-01
GL_136 0 NS_136 NS_135 0 -2.0741858581422049e-01
GS_135_3 0 NS_135 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 1.5742148578820314e+02
RS_138 NS_138 0 1.5742148578820311e+02
GL_137 0 NS_137 NS_138 0 2.0543767879537947e-01
GL_138 0 NS_138 NS_137 0 -2.0543767879537947e-01
GS_137_3 0 NS_137 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 2.0165146427356075e+02
RS_140 NS_140 0 2.0165146427356075e+02
GL_139 0 NS_139 NS_140 0 2.1530071526798281e-01
GL_140 0 NS_140 NS_139 0 -2.1530071526798281e-01
GS_139_3 0 NS_139 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 2.5655383475382814e+02
RS_142 NS_142 0 2.5655383475382814e+02
GL_141 0 NS_141 NS_142 0 2.2143554872154964e-01
GL_142 0 NS_142 NS_141 0 -2.2143554872154964e-01
GS_141_3 0 NS_141 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 3.7527533273924564e+02
RS_144 NS_144 0 3.7527533273924570e+02
GL_143 0 NS_143 NS_144 0 2.2416553875794559e-01
GL_144 0 NS_144 NS_143 0 -2.2416553875794559e-01
GS_143_3 0 NS_143 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 8.7633211379679196e+01
RS_146 NS_146 0 8.7633211379679196e+01
GL_145 0 NS_145 NS_146 0 2.3541329178654702e-01
GL_146 0 NS_146 NS_145 0 -2.3541329178654702e-01
GS_145_3 0 NS_145 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 4.0937268842404592e+02
RS_148 NS_148 0 4.0937268842404586e+02
GL_147 0 NS_147 NS_148 0 2.2933880932778705e-01
GL_148 0 NS_148 NS_147 0 -2.2933880932778705e-01
GS_147_3 0 NS_147 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 1.8046101089657725e+02
RS_150 NS_150 0 1.8046101089657725e+02
GL_149 0 NS_149 NS_150 0 2.3011433813523779e-01
GL_150 0 NS_150 NS_149 0 -2.3011433813523779e-01
GS_149_3 0 NS_149 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 9.7664924917686449e+01
RS_152 NS_152 0 9.7664924917686449e+01
GL_151 0 NS_151 NS_152 0 2.4746563775454208e-01
GL_152 0 NS_152 NS_151 0 -2.4746563775454208e-01
GS_151_3 0 NS_151 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 2.6057215108102395e+02
RS_154 NS_154 0 2.6057215108102395e+02
GL_153 0 NS_153 NS_154 0 2.3565487776505958e-01
GL_154 0 NS_154 NS_153 0 -2.3565487776505958e-01
GS_153_3 0 NS_153 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 1.4688638444267465e+03
RS_156 NS_156 0 1.4688638444267465e+03
GL_155 0 NS_155 NS_156 0 2.3814510332638331e-01
GL_156 0 NS_156 NS_155 0 -2.3814510332638331e-01
GS_155_3 0 NS_155 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 1.5351229021400181e+03
RS_158 NS_158 0 1.5351229021400181e+03
GL_157 0 NS_157 NS_158 0 2.5027181856001052e-01
GL_158 0 NS_158 NS_157 0 -2.5027181856001052e-01
GS_157_3 0 NS_157 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 4.3650646405920685e+02
RS_160 NS_160 0 4.3650646405920685e+02
GL_159 0 NS_159 NS_160 0 2.4893599896984003e-01
GL_160 0 NS_160 NS_159 0 -2.4893599896984003e-01
GS_159_3 0 NS_159 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 1.1441811687773074e+03
RS_162 NS_162 0 1.1441811687773072e+03
GL_161 0 NS_161 NS_162 0 2.4916499611033449e-01
GL_162 0 NS_162 NS_161 0 -2.4916499611033449e-01
GS_161_3 0 NS_161 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 163/164
CS_163 NS_163 0 9.9999999999999998e-13
CS_164 NS_164 0 9.9999999999999998e-13
RS_163 NS_163 0 7.5335118532932768e+02
RS_164 NS_164 0 7.5335118532932768e+02
GL_163 0 NS_163 NS_164 0 2.4298312011423853e-01
GL_164 0 NS_164 NS_163 0 -2.4298312011423853e-01
GS_163_3 0 NS_163 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 1.1346596293114915e+03
RS_166 NS_166 0 1.1346596293114915e+03
GL_165 0 NS_165 NS_166 0 2.4551048269503753e-01
GL_166 0 NS_166 NS_165 0 -2.4551048269503753e-01
GS_165_3 0 NS_165 NA_3 0 1.3803457954163372e+00
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 9.3517666338196523e+02
RS_168 NS_168 0 9.3517666338196523e+02
GL_167 0 NS_167 NS_168 0 2.4538280909205379e-01
GL_168 0 NS_168 NS_167 0 -2.4538280909205379e-01
GS_167_3 0 NS_167 NA_3 0 1.3803457954163372e+00
*
* Real pole n. 169
CS_169 NS_169 0 9.9999999999999998e-13
RS_169 NS_169 0 4.1362120035729779e+00
GS_169_4 0 NS_169 NA_4 0 1.3803457954163372e+00
*
* Real pole n. 170
CS_170 NS_170 0 9.9999999999999998e-13
RS_170 NS_170 0 2.7078253238558993e+01
GS_170_4 0 NS_170 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 5.6873212206500213e+01
RS_172 NS_172 0 5.6873212206500220e+01
GL_171 0 NS_171 NS_172 0 4.7960934964359665e-02
GL_172 0 NS_172 NS_171 0 -4.7960934964359665e-02
GS_171_4 0 NS_171 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 5.5832282069998371e+01
RS_174 NS_174 0 5.5832282069998378e+01
GL_173 0 NS_173 NS_174 0 6.1612202840267971e-02
GL_174 0 NS_174 NS_173 0 -6.1612202840267971e-02
GS_173_4 0 NS_173 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 3.4747519722663924e+01
RS_176 NS_176 0 3.4747519722663924e+01
GL_175 0 NS_175 NS_176 0 8.1784427745819094e-02
GL_176 0 NS_176 NS_175 0 -8.1784427745819094e-02
GS_175_4 0 NS_175 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 3.1454928782186034e+01
RS_178 NS_178 0 3.1454928782186034e+01
GL_177 0 NS_177 NS_178 0 1.1192538378623762e-01
GL_178 0 NS_178 NS_177 0 -1.1192538378623762e-01
GS_177_4 0 NS_177 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 2.2209312435826621e+02
RS_180 NS_180 0 2.2209312435826621e+02
GL_179 0 NS_179 NS_180 0 2.9133579865504960e-01
GL_180 0 NS_180 NS_179 0 -2.9133579865504960e-01
GS_179_4 0 NS_179 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 181/182
CS_181 NS_181 0 9.9999999999999998e-13
CS_182 NS_182 0 9.9999999999999998e-13
RS_181 NS_181 0 4.4403718965615290e+01
RS_182 NS_182 0 4.4403718965615283e+01
GL_181 0 NS_181 NS_182 0 1.3869030610195973e-01
GL_182 0 NS_182 NS_181 0 -1.3869030610195973e-01
GS_181_4 0 NS_181 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 183/184
CS_183 NS_183 0 9.9999999999999998e-13
CS_184 NS_184 0 9.9999999999999998e-13
RS_183 NS_183 0 9.2436417727653946e+01
RS_184 NS_184 0 9.2436417727653946e+01
GL_183 0 NS_183 NS_184 0 1.6009535907039132e-01
GL_184 0 NS_184 NS_183 0 -1.6009535907039132e-01
GS_183_4 0 NS_183 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 5.2247674424140278e+01
RS_186 NS_186 0 5.2247674424140278e+01
GL_185 0 NS_185 NS_186 0 1.7061294296414609e-01
GL_186 0 NS_186 NS_185 0 -1.7061294296414609e-01
GS_185_4 0 NS_185 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 6.3351631924882277e+01
RS_188 NS_188 0 6.3351631924882277e+01
GL_187 0 NS_187 NS_188 0 1.8578563768540060e-01
GL_188 0 NS_188 NS_187 0 -1.8578563768540060e-01
GS_187_4 0 NS_187 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 2.2461363612924958e+02
RS_190 NS_190 0 2.2461363612924956e+02
GL_189 0 NS_189 NS_190 0 2.0090890151880786e-01
GL_190 0 NS_190 NS_189 0 -2.0090890151880786e-01
GS_189_4 0 NS_189 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 6.2323563035856608e+01
RS_192 NS_192 0 6.2323563035856608e+01
GL_191 0 NS_191 NS_192 0 2.0741858581422049e-01
GL_192 0 NS_192 NS_191 0 -2.0741858581422049e-01
GS_191_4 0 NS_191 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 1.5742148578820314e+02
RS_194 NS_194 0 1.5742148578820311e+02
GL_193 0 NS_193 NS_194 0 2.0543767879537947e-01
GL_194 0 NS_194 NS_193 0 -2.0543767879537947e-01
GS_193_4 0 NS_193 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 2.0165146427356075e+02
RS_196 NS_196 0 2.0165146427356075e+02
GL_195 0 NS_195 NS_196 0 2.1530071526798281e-01
GL_196 0 NS_196 NS_195 0 -2.1530071526798281e-01
GS_195_4 0 NS_195 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 2.5655383475382814e+02
RS_198 NS_198 0 2.5655383475382814e+02
GL_197 0 NS_197 NS_198 0 2.2143554872154964e-01
GL_198 0 NS_198 NS_197 0 -2.2143554872154964e-01
GS_197_4 0 NS_197 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 3.7527533273924564e+02
RS_200 NS_200 0 3.7527533273924570e+02
GL_199 0 NS_199 NS_200 0 2.2416553875794559e-01
GL_200 0 NS_200 NS_199 0 -2.2416553875794559e-01
GS_199_4 0 NS_199 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 201/202
CS_201 NS_201 0 9.9999999999999998e-13
CS_202 NS_202 0 9.9999999999999998e-13
RS_201 NS_201 0 8.7633211379679196e+01
RS_202 NS_202 0 8.7633211379679196e+01
GL_201 0 NS_201 NS_202 0 2.3541329178654702e-01
GL_202 0 NS_202 NS_201 0 -2.3541329178654702e-01
GS_201_4 0 NS_201 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 203/204
CS_203 NS_203 0 9.9999999999999998e-13
CS_204 NS_204 0 9.9999999999999998e-13
RS_203 NS_203 0 4.0937268842404592e+02
RS_204 NS_204 0 4.0937268842404586e+02
GL_203 0 NS_203 NS_204 0 2.2933880932778705e-01
GL_204 0 NS_204 NS_203 0 -2.2933880932778705e-01
GS_203_4 0 NS_203 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 1.8046101089657725e+02
RS_206 NS_206 0 1.8046101089657725e+02
GL_205 0 NS_205 NS_206 0 2.3011433813523779e-01
GL_206 0 NS_206 NS_205 0 -2.3011433813523779e-01
GS_205_4 0 NS_205 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 9.7664924917686449e+01
RS_208 NS_208 0 9.7664924917686449e+01
GL_207 0 NS_207 NS_208 0 2.4746563775454208e-01
GL_208 0 NS_208 NS_207 0 -2.4746563775454208e-01
GS_207_4 0 NS_207 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 2.6057215108102395e+02
RS_210 NS_210 0 2.6057215108102395e+02
GL_209 0 NS_209 NS_210 0 2.3565487776505958e-01
GL_210 0 NS_210 NS_209 0 -2.3565487776505958e-01
GS_209_4 0 NS_209 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 1.4688638444267465e+03
RS_212 NS_212 0 1.4688638444267465e+03
GL_211 0 NS_211 NS_212 0 2.3814510332638331e-01
GL_212 0 NS_212 NS_211 0 -2.3814510332638331e-01
GS_211_4 0 NS_211 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 1.5351229021400181e+03
RS_214 NS_214 0 1.5351229021400181e+03
GL_213 0 NS_213 NS_214 0 2.5027181856001052e-01
GL_214 0 NS_214 NS_213 0 -2.5027181856001052e-01
GS_213_4 0 NS_213 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 4.3650646405920685e+02
RS_216 NS_216 0 4.3650646405920685e+02
GL_215 0 NS_215 NS_216 0 2.4893599896984003e-01
GL_216 0 NS_216 NS_215 0 -2.4893599896984003e-01
GS_215_4 0 NS_215 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 1.1441811687773074e+03
RS_218 NS_218 0 1.1441811687773072e+03
GL_217 0 NS_217 NS_218 0 2.4916499611033449e-01
GL_218 0 NS_218 NS_217 0 -2.4916499611033449e-01
GS_217_4 0 NS_217 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 7.5335118532932768e+02
RS_220 NS_220 0 7.5335118532932768e+02
GL_219 0 NS_219 NS_220 0 2.4298312011423853e-01
GL_220 0 NS_220 NS_219 0 -2.4298312011423853e-01
GS_219_4 0 NS_219 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 221/222
CS_221 NS_221 0 9.9999999999999998e-13
CS_222 NS_222 0 9.9999999999999998e-13
RS_221 NS_221 0 1.1346596293114915e+03
RS_222 NS_222 0 1.1346596293114915e+03
GL_221 0 NS_221 NS_222 0 2.4551048269503753e-01
GL_222 0 NS_222 NS_221 0 -2.4551048269503753e-01
GS_221_4 0 NS_221 NA_4 0 1.3803457954163372e+00
*
* Complex pair n. 223/224
CS_223 NS_223 0 9.9999999999999998e-13
CS_224 NS_224 0 9.9999999999999998e-13
RS_223 NS_223 0 9.3517666338196523e+02
RS_224 NS_224 0 9.3517666338196523e+02
GL_223 0 NS_223 NS_224 0 2.4538280909205379e-01
GL_224 0 NS_224 NS_223 0 -2.4538280909205379e-01
GS_223_4 0 NS_223 NA_4 0 1.3803457954163372e+00
*
* Real pole n. 225
CS_225 NS_225 0 9.9999999999999998e-13
RS_225 NS_225 0 4.1362120035729779e+00
GS_225_5 0 NS_225 NA_5 0 1.3803457954163372e+00
*
* Real pole n. 226
CS_226 NS_226 0 9.9999999999999998e-13
RS_226 NS_226 0 2.7078253238558993e+01
GS_226_5 0 NS_226 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 5.6873212206500213e+01
RS_228 NS_228 0 5.6873212206500220e+01
GL_227 0 NS_227 NS_228 0 4.7960934964359665e-02
GL_228 0 NS_228 NS_227 0 -4.7960934964359665e-02
GS_227_5 0 NS_227 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 229/230
CS_229 NS_229 0 9.9999999999999998e-13
CS_230 NS_230 0 9.9999999999999998e-13
RS_229 NS_229 0 5.5832282069998371e+01
RS_230 NS_230 0 5.5832282069998378e+01
GL_229 0 NS_229 NS_230 0 6.1612202840267971e-02
GL_230 0 NS_230 NS_229 0 -6.1612202840267971e-02
GS_229_5 0 NS_229 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 3.4747519722663924e+01
RS_232 NS_232 0 3.4747519722663924e+01
GL_231 0 NS_231 NS_232 0 8.1784427745819094e-02
GL_232 0 NS_232 NS_231 0 -8.1784427745819094e-02
GS_231_5 0 NS_231 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 3.1454928782186034e+01
RS_234 NS_234 0 3.1454928782186034e+01
GL_233 0 NS_233 NS_234 0 1.1192538378623762e-01
GL_234 0 NS_234 NS_233 0 -1.1192538378623762e-01
GS_233_5 0 NS_233 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 2.2209312435826621e+02
RS_236 NS_236 0 2.2209312435826621e+02
GL_235 0 NS_235 NS_236 0 2.9133579865504960e-01
GL_236 0 NS_236 NS_235 0 -2.9133579865504960e-01
GS_235_5 0 NS_235 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 4.4403718965615290e+01
RS_238 NS_238 0 4.4403718965615283e+01
GL_237 0 NS_237 NS_238 0 1.3869030610195973e-01
GL_238 0 NS_238 NS_237 0 -1.3869030610195973e-01
GS_237_5 0 NS_237 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 9.2436417727653946e+01
RS_240 NS_240 0 9.2436417727653946e+01
GL_239 0 NS_239 NS_240 0 1.6009535907039132e-01
GL_240 0 NS_240 NS_239 0 -1.6009535907039132e-01
GS_239_5 0 NS_239 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 241/242
CS_241 NS_241 0 9.9999999999999998e-13
CS_242 NS_242 0 9.9999999999999998e-13
RS_241 NS_241 0 5.2247674424140278e+01
RS_242 NS_242 0 5.2247674424140278e+01
GL_241 0 NS_241 NS_242 0 1.7061294296414609e-01
GL_242 0 NS_242 NS_241 0 -1.7061294296414609e-01
GS_241_5 0 NS_241 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 243/244
CS_243 NS_243 0 9.9999999999999998e-13
CS_244 NS_244 0 9.9999999999999998e-13
RS_243 NS_243 0 6.3351631924882277e+01
RS_244 NS_244 0 6.3351631924882277e+01
GL_243 0 NS_243 NS_244 0 1.8578563768540060e-01
GL_244 0 NS_244 NS_243 0 -1.8578563768540060e-01
GS_243_5 0 NS_243 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 245/246
CS_245 NS_245 0 9.9999999999999998e-13
CS_246 NS_246 0 9.9999999999999998e-13
RS_245 NS_245 0 2.2461363612924958e+02
RS_246 NS_246 0 2.2461363612924956e+02
GL_245 0 NS_245 NS_246 0 2.0090890151880786e-01
GL_246 0 NS_246 NS_245 0 -2.0090890151880786e-01
GS_245_5 0 NS_245 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 247/248
CS_247 NS_247 0 9.9999999999999998e-13
CS_248 NS_248 0 9.9999999999999998e-13
RS_247 NS_247 0 6.2323563035856608e+01
RS_248 NS_248 0 6.2323563035856608e+01
GL_247 0 NS_247 NS_248 0 2.0741858581422049e-01
GL_248 0 NS_248 NS_247 0 -2.0741858581422049e-01
GS_247_5 0 NS_247 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 249/250
CS_249 NS_249 0 9.9999999999999998e-13
CS_250 NS_250 0 9.9999999999999998e-13
RS_249 NS_249 0 1.5742148578820314e+02
RS_250 NS_250 0 1.5742148578820311e+02
GL_249 0 NS_249 NS_250 0 2.0543767879537947e-01
GL_250 0 NS_250 NS_249 0 -2.0543767879537947e-01
GS_249_5 0 NS_249 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 251/252
CS_251 NS_251 0 9.9999999999999998e-13
CS_252 NS_252 0 9.9999999999999998e-13
RS_251 NS_251 0 2.0165146427356075e+02
RS_252 NS_252 0 2.0165146427356075e+02
GL_251 0 NS_251 NS_252 0 2.1530071526798281e-01
GL_252 0 NS_252 NS_251 0 -2.1530071526798281e-01
GS_251_5 0 NS_251 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 253/254
CS_253 NS_253 0 9.9999999999999998e-13
CS_254 NS_254 0 9.9999999999999998e-13
RS_253 NS_253 0 2.5655383475382814e+02
RS_254 NS_254 0 2.5655383475382814e+02
GL_253 0 NS_253 NS_254 0 2.2143554872154964e-01
GL_254 0 NS_254 NS_253 0 -2.2143554872154964e-01
GS_253_5 0 NS_253 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 255/256
CS_255 NS_255 0 9.9999999999999998e-13
CS_256 NS_256 0 9.9999999999999998e-13
RS_255 NS_255 0 3.7527533273924564e+02
RS_256 NS_256 0 3.7527533273924570e+02
GL_255 0 NS_255 NS_256 0 2.2416553875794559e-01
GL_256 0 NS_256 NS_255 0 -2.2416553875794559e-01
GS_255_5 0 NS_255 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 257/258
CS_257 NS_257 0 9.9999999999999998e-13
CS_258 NS_258 0 9.9999999999999998e-13
RS_257 NS_257 0 8.7633211379679196e+01
RS_258 NS_258 0 8.7633211379679196e+01
GL_257 0 NS_257 NS_258 0 2.3541329178654702e-01
GL_258 0 NS_258 NS_257 0 -2.3541329178654702e-01
GS_257_5 0 NS_257 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 259/260
CS_259 NS_259 0 9.9999999999999998e-13
CS_260 NS_260 0 9.9999999999999998e-13
RS_259 NS_259 0 4.0937268842404592e+02
RS_260 NS_260 0 4.0937268842404586e+02
GL_259 0 NS_259 NS_260 0 2.2933880932778705e-01
GL_260 0 NS_260 NS_259 0 -2.2933880932778705e-01
GS_259_5 0 NS_259 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 261/262
CS_261 NS_261 0 9.9999999999999998e-13
CS_262 NS_262 0 9.9999999999999998e-13
RS_261 NS_261 0 1.8046101089657725e+02
RS_262 NS_262 0 1.8046101089657725e+02
GL_261 0 NS_261 NS_262 0 2.3011433813523779e-01
GL_262 0 NS_262 NS_261 0 -2.3011433813523779e-01
GS_261_5 0 NS_261 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 263/264
CS_263 NS_263 0 9.9999999999999998e-13
CS_264 NS_264 0 9.9999999999999998e-13
RS_263 NS_263 0 9.7664924917686449e+01
RS_264 NS_264 0 9.7664924917686449e+01
GL_263 0 NS_263 NS_264 0 2.4746563775454208e-01
GL_264 0 NS_264 NS_263 0 -2.4746563775454208e-01
GS_263_5 0 NS_263 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 265/266
CS_265 NS_265 0 9.9999999999999998e-13
CS_266 NS_266 0 9.9999999999999998e-13
RS_265 NS_265 0 2.6057215108102395e+02
RS_266 NS_266 0 2.6057215108102395e+02
GL_265 0 NS_265 NS_266 0 2.3565487776505958e-01
GL_266 0 NS_266 NS_265 0 -2.3565487776505958e-01
GS_265_5 0 NS_265 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 267/268
CS_267 NS_267 0 9.9999999999999998e-13
CS_268 NS_268 0 9.9999999999999998e-13
RS_267 NS_267 0 1.4688638444267465e+03
RS_268 NS_268 0 1.4688638444267465e+03
GL_267 0 NS_267 NS_268 0 2.3814510332638331e-01
GL_268 0 NS_268 NS_267 0 -2.3814510332638331e-01
GS_267_5 0 NS_267 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 269/270
CS_269 NS_269 0 9.9999999999999998e-13
CS_270 NS_270 0 9.9999999999999998e-13
RS_269 NS_269 0 1.5351229021400181e+03
RS_270 NS_270 0 1.5351229021400181e+03
GL_269 0 NS_269 NS_270 0 2.5027181856001052e-01
GL_270 0 NS_270 NS_269 0 -2.5027181856001052e-01
GS_269_5 0 NS_269 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 271/272
CS_271 NS_271 0 9.9999999999999998e-13
CS_272 NS_272 0 9.9999999999999998e-13
RS_271 NS_271 0 4.3650646405920685e+02
RS_272 NS_272 0 4.3650646405920685e+02
GL_271 0 NS_271 NS_272 0 2.4893599896984003e-01
GL_272 0 NS_272 NS_271 0 -2.4893599896984003e-01
GS_271_5 0 NS_271 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 273/274
CS_273 NS_273 0 9.9999999999999998e-13
CS_274 NS_274 0 9.9999999999999998e-13
RS_273 NS_273 0 1.1441811687773074e+03
RS_274 NS_274 0 1.1441811687773072e+03
GL_273 0 NS_273 NS_274 0 2.4916499611033449e-01
GL_274 0 NS_274 NS_273 0 -2.4916499611033449e-01
GS_273_5 0 NS_273 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 275/276
CS_275 NS_275 0 9.9999999999999998e-13
CS_276 NS_276 0 9.9999999999999998e-13
RS_275 NS_275 0 7.5335118532932768e+02
RS_276 NS_276 0 7.5335118532932768e+02
GL_275 0 NS_275 NS_276 0 2.4298312011423853e-01
GL_276 0 NS_276 NS_275 0 -2.4298312011423853e-01
GS_275_5 0 NS_275 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 277/278
CS_277 NS_277 0 9.9999999999999998e-13
CS_278 NS_278 0 9.9999999999999998e-13
RS_277 NS_277 0 1.1346596293114915e+03
RS_278 NS_278 0 1.1346596293114915e+03
GL_277 0 NS_277 NS_278 0 2.4551048269503753e-01
GL_278 0 NS_278 NS_277 0 -2.4551048269503753e-01
GS_277_5 0 NS_277 NA_5 0 1.3803457954163372e+00
*
* Complex pair n. 279/280
CS_279 NS_279 0 9.9999999999999998e-13
CS_280 NS_280 0 9.9999999999999998e-13
RS_279 NS_279 0 9.3517666338196523e+02
RS_280 NS_280 0 9.3517666338196523e+02
GL_279 0 NS_279 NS_280 0 2.4538280909205379e-01
GL_280 0 NS_280 NS_279 0 -2.4538280909205379e-01
GS_279_5 0 NS_279 NA_5 0 1.3803457954163372e+00
*
* Real pole n. 281
CS_281 NS_281 0 9.9999999999999998e-13
RS_281 NS_281 0 4.1362120035729779e+00
GS_281_6 0 NS_281 NA_6 0 1.3803457954163372e+00
*
* Real pole n. 282
CS_282 NS_282 0 9.9999999999999998e-13
RS_282 NS_282 0 2.7078253238558993e+01
GS_282_6 0 NS_282 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 283/284
CS_283 NS_283 0 9.9999999999999998e-13
CS_284 NS_284 0 9.9999999999999998e-13
RS_283 NS_283 0 5.6873212206500213e+01
RS_284 NS_284 0 5.6873212206500220e+01
GL_283 0 NS_283 NS_284 0 4.7960934964359665e-02
GL_284 0 NS_284 NS_283 0 -4.7960934964359665e-02
GS_283_6 0 NS_283 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 285/286
CS_285 NS_285 0 9.9999999999999998e-13
CS_286 NS_286 0 9.9999999999999998e-13
RS_285 NS_285 0 5.5832282069998371e+01
RS_286 NS_286 0 5.5832282069998378e+01
GL_285 0 NS_285 NS_286 0 6.1612202840267971e-02
GL_286 0 NS_286 NS_285 0 -6.1612202840267971e-02
GS_285_6 0 NS_285 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 287/288
CS_287 NS_287 0 9.9999999999999998e-13
CS_288 NS_288 0 9.9999999999999998e-13
RS_287 NS_287 0 3.4747519722663924e+01
RS_288 NS_288 0 3.4747519722663924e+01
GL_287 0 NS_287 NS_288 0 8.1784427745819094e-02
GL_288 0 NS_288 NS_287 0 -8.1784427745819094e-02
GS_287_6 0 NS_287 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 289/290
CS_289 NS_289 0 9.9999999999999998e-13
CS_290 NS_290 0 9.9999999999999998e-13
RS_289 NS_289 0 3.1454928782186034e+01
RS_290 NS_290 0 3.1454928782186034e+01
GL_289 0 NS_289 NS_290 0 1.1192538378623762e-01
GL_290 0 NS_290 NS_289 0 -1.1192538378623762e-01
GS_289_6 0 NS_289 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 291/292
CS_291 NS_291 0 9.9999999999999998e-13
CS_292 NS_292 0 9.9999999999999998e-13
RS_291 NS_291 0 2.2209312435826621e+02
RS_292 NS_292 0 2.2209312435826621e+02
GL_291 0 NS_291 NS_292 0 2.9133579865504960e-01
GL_292 0 NS_292 NS_291 0 -2.9133579865504960e-01
GS_291_6 0 NS_291 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 293/294
CS_293 NS_293 0 9.9999999999999998e-13
CS_294 NS_294 0 9.9999999999999998e-13
RS_293 NS_293 0 4.4403718965615290e+01
RS_294 NS_294 0 4.4403718965615283e+01
GL_293 0 NS_293 NS_294 0 1.3869030610195973e-01
GL_294 0 NS_294 NS_293 0 -1.3869030610195973e-01
GS_293_6 0 NS_293 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 295/296
CS_295 NS_295 0 9.9999999999999998e-13
CS_296 NS_296 0 9.9999999999999998e-13
RS_295 NS_295 0 9.2436417727653946e+01
RS_296 NS_296 0 9.2436417727653946e+01
GL_295 0 NS_295 NS_296 0 1.6009535907039132e-01
GL_296 0 NS_296 NS_295 0 -1.6009535907039132e-01
GS_295_6 0 NS_295 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 297/298
CS_297 NS_297 0 9.9999999999999998e-13
CS_298 NS_298 0 9.9999999999999998e-13
RS_297 NS_297 0 5.2247674424140278e+01
RS_298 NS_298 0 5.2247674424140278e+01
GL_297 0 NS_297 NS_298 0 1.7061294296414609e-01
GL_298 0 NS_298 NS_297 0 -1.7061294296414609e-01
GS_297_6 0 NS_297 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 299/300
CS_299 NS_299 0 9.9999999999999998e-13
CS_300 NS_300 0 9.9999999999999998e-13
RS_299 NS_299 0 6.3351631924882277e+01
RS_300 NS_300 0 6.3351631924882277e+01
GL_299 0 NS_299 NS_300 0 1.8578563768540060e-01
GL_300 0 NS_300 NS_299 0 -1.8578563768540060e-01
GS_299_6 0 NS_299 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 301/302
CS_301 NS_301 0 9.9999999999999998e-13
CS_302 NS_302 0 9.9999999999999998e-13
RS_301 NS_301 0 2.2461363612924958e+02
RS_302 NS_302 0 2.2461363612924956e+02
GL_301 0 NS_301 NS_302 0 2.0090890151880786e-01
GL_302 0 NS_302 NS_301 0 -2.0090890151880786e-01
GS_301_6 0 NS_301 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 303/304
CS_303 NS_303 0 9.9999999999999998e-13
CS_304 NS_304 0 9.9999999999999998e-13
RS_303 NS_303 0 6.2323563035856608e+01
RS_304 NS_304 0 6.2323563035856608e+01
GL_303 0 NS_303 NS_304 0 2.0741858581422049e-01
GL_304 0 NS_304 NS_303 0 -2.0741858581422049e-01
GS_303_6 0 NS_303 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 305/306
CS_305 NS_305 0 9.9999999999999998e-13
CS_306 NS_306 0 9.9999999999999998e-13
RS_305 NS_305 0 1.5742148578820314e+02
RS_306 NS_306 0 1.5742148578820311e+02
GL_305 0 NS_305 NS_306 0 2.0543767879537947e-01
GL_306 0 NS_306 NS_305 0 -2.0543767879537947e-01
GS_305_6 0 NS_305 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 307/308
CS_307 NS_307 0 9.9999999999999998e-13
CS_308 NS_308 0 9.9999999999999998e-13
RS_307 NS_307 0 2.0165146427356075e+02
RS_308 NS_308 0 2.0165146427356075e+02
GL_307 0 NS_307 NS_308 0 2.1530071526798281e-01
GL_308 0 NS_308 NS_307 0 -2.1530071526798281e-01
GS_307_6 0 NS_307 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 309/310
CS_309 NS_309 0 9.9999999999999998e-13
CS_310 NS_310 0 9.9999999999999998e-13
RS_309 NS_309 0 2.5655383475382814e+02
RS_310 NS_310 0 2.5655383475382814e+02
GL_309 0 NS_309 NS_310 0 2.2143554872154964e-01
GL_310 0 NS_310 NS_309 0 -2.2143554872154964e-01
GS_309_6 0 NS_309 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 311/312
CS_311 NS_311 0 9.9999999999999998e-13
CS_312 NS_312 0 9.9999999999999998e-13
RS_311 NS_311 0 3.7527533273924564e+02
RS_312 NS_312 0 3.7527533273924570e+02
GL_311 0 NS_311 NS_312 0 2.2416553875794559e-01
GL_312 0 NS_312 NS_311 0 -2.2416553875794559e-01
GS_311_6 0 NS_311 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 313/314
CS_313 NS_313 0 9.9999999999999998e-13
CS_314 NS_314 0 9.9999999999999998e-13
RS_313 NS_313 0 8.7633211379679196e+01
RS_314 NS_314 0 8.7633211379679196e+01
GL_313 0 NS_313 NS_314 0 2.3541329178654702e-01
GL_314 0 NS_314 NS_313 0 -2.3541329178654702e-01
GS_313_6 0 NS_313 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 315/316
CS_315 NS_315 0 9.9999999999999998e-13
CS_316 NS_316 0 9.9999999999999998e-13
RS_315 NS_315 0 4.0937268842404592e+02
RS_316 NS_316 0 4.0937268842404586e+02
GL_315 0 NS_315 NS_316 0 2.2933880932778705e-01
GL_316 0 NS_316 NS_315 0 -2.2933880932778705e-01
GS_315_6 0 NS_315 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 317/318
CS_317 NS_317 0 9.9999999999999998e-13
CS_318 NS_318 0 9.9999999999999998e-13
RS_317 NS_317 0 1.8046101089657725e+02
RS_318 NS_318 0 1.8046101089657725e+02
GL_317 0 NS_317 NS_318 0 2.3011433813523779e-01
GL_318 0 NS_318 NS_317 0 -2.3011433813523779e-01
GS_317_6 0 NS_317 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 319/320
CS_319 NS_319 0 9.9999999999999998e-13
CS_320 NS_320 0 9.9999999999999998e-13
RS_319 NS_319 0 9.7664924917686449e+01
RS_320 NS_320 0 9.7664924917686449e+01
GL_319 0 NS_319 NS_320 0 2.4746563775454208e-01
GL_320 0 NS_320 NS_319 0 -2.4746563775454208e-01
GS_319_6 0 NS_319 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 321/322
CS_321 NS_321 0 9.9999999999999998e-13
CS_322 NS_322 0 9.9999999999999998e-13
RS_321 NS_321 0 2.6057215108102395e+02
RS_322 NS_322 0 2.6057215108102395e+02
GL_321 0 NS_321 NS_322 0 2.3565487776505958e-01
GL_322 0 NS_322 NS_321 0 -2.3565487776505958e-01
GS_321_6 0 NS_321 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 323/324
CS_323 NS_323 0 9.9999999999999998e-13
CS_324 NS_324 0 9.9999999999999998e-13
RS_323 NS_323 0 1.4688638444267465e+03
RS_324 NS_324 0 1.4688638444267465e+03
GL_323 0 NS_323 NS_324 0 2.3814510332638331e-01
GL_324 0 NS_324 NS_323 0 -2.3814510332638331e-01
GS_323_6 0 NS_323 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 325/326
CS_325 NS_325 0 9.9999999999999998e-13
CS_326 NS_326 0 9.9999999999999998e-13
RS_325 NS_325 0 1.5351229021400181e+03
RS_326 NS_326 0 1.5351229021400181e+03
GL_325 0 NS_325 NS_326 0 2.5027181856001052e-01
GL_326 0 NS_326 NS_325 0 -2.5027181856001052e-01
GS_325_6 0 NS_325 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 327/328
CS_327 NS_327 0 9.9999999999999998e-13
CS_328 NS_328 0 9.9999999999999998e-13
RS_327 NS_327 0 4.3650646405920685e+02
RS_328 NS_328 0 4.3650646405920685e+02
GL_327 0 NS_327 NS_328 0 2.4893599896984003e-01
GL_328 0 NS_328 NS_327 0 -2.4893599896984003e-01
GS_327_6 0 NS_327 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 329/330
CS_329 NS_329 0 9.9999999999999998e-13
CS_330 NS_330 0 9.9999999999999998e-13
RS_329 NS_329 0 1.1441811687773074e+03
RS_330 NS_330 0 1.1441811687773072e+03
GL_329 0 NS_329 NS_330 0 2.4916499611033449e-01
GL_330 0 NS_330 NS_329 0 -2.4916499611033449e-01
GS_329_6 0 NS_329 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 331/332
CS_331 NS_331 0 9.9999999999999998e-13
CS_332 NS_332 0 9.9999999999999998e-13
RS_331 NS_331 0 7.5335118532932768e+02
RS_332 NS_332 0 7.5335118532932768e+02
GL_331 0 NS_331 NS_332 0 2.4298312011423853e-01
GL_332 0 NS_332 NS_331 0 -2.4298312011423853e-01
GS_331_6 0 NS_331 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 333/334
CS_333 NS_333 0 9.9999999999999998e-13
CS_334 NS_334 0 9.9999999999999998e-13
RS_333 NS_333 0 1.1346596293114915e+03
RS_334 NS_334 0 1.1346596293114915e+03
GL_333 0 NS_333 NS_334 0 2.4551048269503753e-01
GL_334 0 NS_334 NS_333 0 -2.4551048269503753e-01
GS_333_6 0 NS_333 NA_6 0 1.3803457954163372e+00
*
* Complex pair n. 335/336
CS_335 NS_335 0 9.9999999999999998e-13
CS_336 NS_336 0 9.9999999999999998e-13
RS_335 NS_335 0 9.3517666338196523e+02
RS_336 NS_336 0 9.3517666338196523e+02
GL_335 0 NS_335 NS_336 0 2.4538280909205379e-01
GL_336 0 NS_336 NS_335 0 -2.4538280909205379e-01
GS_335_6 0 NS_335 NA_6 0 1.3803457954163372e+00
*
* Real pole n. 337
CS_337 NS_337 0 9.9999999999999998e-13
RS_337 NS_337 0 4.1362120035729779e+00
GS_337_7 0 NS_337 NA_7 0 1.3803457954163372e+00
*
* Real pole n. 338
CS_338 NS_338 0 9.9999999999999998e-13
RS_338 NS_338 0 2.7078253238558993e+01
GS_338_7 0 NS_338 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 339/340
CS_339 NS_339 0 9.9999999999999998e-13
CS_340 NS_340 0 9.9999999999999998e-13
RS_339 NS_339 0 5.6873212206500213e+01
RS_340 NS_340 0 5.6873212206500220e+01
GL_339 0 NS_339 NS_340 0 4.7960934964359665e-02
GL_340 0 NS_340 NS_339 0 -4.7960934964359665e-02
GS_339_7 0 NS_339 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 341/342
CS_341 NS_341 0 9.9999999999999998e-13
CS_342 NS_342 0 9.9999999999999998e-13
RS_341 NS_341 0 5.5832282069998371e+01
RS_342 NS_342 0 5.5832282069998378e+01
GL_341 0 NS_341 NS_342 0 6.1612202840267971e-02
GL_342 0 NS_342 NS_341 0 -6.1612202840267971e-02
GS_341_7 0 NS_341 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 343/344
CS_343 NS_343 0 9.9999999999999998e-13
CS_344 NS_344 0 9.9999999999999998e-13
RS_343 NS_343 0 3.4747519722663924e+01
RS_344 NS_344 0 3.4747519722663924e+01
GL_343 0 NS_343 NS_344 0 8.1784427745819094e-02
GL_344 0 NS_344 NS_343 0 -8.1784427745819094e-02
GS_343_7 0 NS_343 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 345/346
CS_345 NS_345 0 9.9999999999999998e-13
CS_346 NS_346 0 9.9999999999999998e-13
RS_345 NS_345 0 3.1454928782186034e+01
RS_346 NS_346 0 3.1454928782186034e+01
GL_345 0 NS_345 NS_346 0 1.1192538378623762e-01
GL_346 0 NS_346 NS_345 0 -1.1192538378623762e-01
GS_345_7 0 NS_345 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 347/348
CS_347 NS_347 0 9.9999999999999998e-13
CS_348 NS_348 0 9.9999999999999998e-13
RS_347 NS_347 0 2.2209312435826621e+02
RS_348 NS_348 0 2.2209312435826621e+02
GL_347 0 NS_347 NS_348 0 2.9133579865504960e-01
GL_348 0 NS_348 NS_347 0 -2.9133579865504960e-01
GS_347_7 0 NS_347 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 349/350
CS_349 NS_349 0 9.9999999999999998e-13
CS_350 NS_350 0 9.9999999999999998e-13
RS_349 NS_349 0 4.4403718965615290e+01
RS_350 NS_350 0 4.4403718965615283e+01
GL_349 0 NS_349 NS_350 0 1.3869030610195973e-01
GL_350 0 NS_350 NS_349 0 -1.3869030610195973e-01
GS_349_7 0 NS_349 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 351/352
CS_351 NS_351 0 9.9999999999999998e-13
CS_352 NS_352 0 9.9999999999999998e-13
RS_351 NS_351 0 9.2436417727653946e+01
RS_352 NS_352 0 9.2436417727653946e+01
GL_351 0 NS_351 NS_352 0 1.6009535907039132e-01
GL_352 0 NS_352 NS_351 0 -1.6009535907039132e-01
GS_351_7 0 NS_351 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 353/354
CS_353 NS_353 0 9.9999999999999998e-13
CS_354 NS_354 0 9.9999999999999998e-13
RS_353 NS_353 0 5.2247674424140278e+01
RS_354 NS_354 0 5.2247674424140278e+01
GL_353 0 NS_353 NS_354 0 1.7061294296414609e-01
GL_354 0 NS_354 NS_353 0 -1.7061294296414609e-01
GS_353_7 0 NS_353 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 355/356
CS_355 NS_355 0 9.9999999999999998e-13
CS_356 NS_356 0 9.9999999999999998e-13
RS_355 NS_355 0 6.3351631924882277e+01
RS_356 NS_356 0 6.3351631924882277e+01
GL_355 0 NS_355 NS_356 0 1.8578563768540060e-01
GL_356 0 NS_356 NS_355 0 -1.8578563768540060e-01
GS_355_7 0 NS_355 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 357/358
CS_357 NS_357 0 9.9999999999999998e-13
CS_358 NS_358 0 9.9999999999999998e-13
RS_357 NS_357 0 2.2461363612924958e+02
RS_358 NS_358 0 2.2461363612924956e+02
GL_357 0 NS_357 NS_358 0 2.0090890151880786e-01
GL_358 0 NS_358 NS_357 0 -2.0090890151880786e-01
GS_357_7 0 NS_357 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 359/360
CS_359 NS_359 0 9.9999999999999998e-13
CS_360 NS_360 0 9.9999999999999998e-13
RS_359 NS_359 0 6.2323563035856608e+01
RS_360 NS_360 0 6.2323563035856608e+01
GL_359 0 NS_359 NS_360 0 2.0741858581422049e-01
GL_360 0 NS_360 NS_359 0 -2.0741858581422049e-01
GS_359_7 0 NS_359 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 361/362
CS_361 NS_361 0 9.9999999999999998e-13
CS_362 NS_362 0 9.9999999999999998e-13
RS_361 NS_361 0 1.5742148578820314e+02
RS_362 NS_362 0 1.5742148578820311e+02
GL_361 0 NS_361 NS_362 0 2.0543767879537947e-01
GL_362 0 NS_362 NS_361 0 -2.0543767879537947e-01
GS_361_7 0 NS_361 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 363/364
CS_363 NS_363 0 9.9999999999999998e-13
CS_364 NS_364 0 9.9999999999999998e-13
RS_363 NS_363 0 2.0165146427356075e+02
RS_364 NS_364 0 2.0165146427356075e+02
GL_363 0 NS_363 NS_364 0 2.1530071526798281e-01
GL_364 0 NS_364 NS_363 0 -2.1530071526798281e-01
GS_363_7 0 NS_363 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 365/366
CS_365 NS_365 0 9.9999999999999998e-13
CS_366 NS_366 0 9.9999999999999998e-13
RS_365 NS_365 0 2.5655383475382814e+02
RS_366 NS_366 0 2.5655383475382814e+02
GL_365 0 NS_365 NS_366 0 2.2143554872154964e-01
GL_366 0 NS_366 NS_365 0 -2.2143554872154964e-01
GS_365_7 0 NS_365 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 367/368
CS_367 NS_367 0 9.9999999999999998e-13
CS_368 NS_368 0 9.9999999999999998e-13
RS_367 NS_367 0 3.7527533273924564e+02
RS_368 NS_368 0 3.7527533273924570e+02
GL_367 0 NS_367 NS_368 0 2.2416553875794559e-01
GL_368 0 NS_368 NS_367 0 -2.2416553875794559e-01
GS_367_7 0 NS_367 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 369/370
CS_369 NS_369 0 9.9999999999999998e-13
CS_370 NS_370 0 9.9999999999999998e-13
RS_369 NS_369 0 8.7633211379679196e+01
RS_370 NS_370 0 8.7633211379679196e+01
GL_369 0 NS_369 NS_370 0 2.3541329178654702e-01
GL_370 0 NS_370 NS_369 0 -2.3541329178654702e-01
GS_369_7 0 NS_369 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 371/372
CS_371 NS_371 0 9.9999999999999998e-13
CS_372 NS_372 0 9.9999999999999998e-13
RS_371 NS_371 0 4.0937268842404592e+02
RS_372 NS_372 0 4.0937268842404586e+02
GL_371 0 NS_371 NS_372 0 2.2933880932778705e-01
GL_372 0 NS_372 NS_371 0 -2.2933880932778705e-01
GS_371_7 0 NS_371 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 373/374
CS_373 NS_373 0 9.9999999999999998e-13
CS_374 NS_374 0 9.9999999999999998e-13
RS_373 NS_373 0 1.8046101089657725e+02
RS_374 NS_374 0 1.8046101089657725e+02
GL_373 0 NS_373 NS_374 0 2.3011433813523779e-01
GL_374 0 NS_374 NS_373 0 -2.3011433813523779e-01
GS_373_7 0 NS_373 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 375/376
CS_375 NS_375 0 9.9999999999999998e-13
CS_376 NS_376 0 9.9999999999999998e-13
RS_375 NS_375 0 9.7664924917686449e+01
RS_376 NS_376 0 9.7664924917686449e+01
GL_375 0 NS_375 NS_376 0 2.4746563775454208e-01
GL_376 0 NS_376 NS_375 0 -2.4746563775454208e-01
GS_375_7 0 NS_375 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 377/378
CS_377 NS_377 0 9.9999999999999998e-13
CS_378 NS_378 0 9.9999999999999998e-13
RS_377 NS_377 0 2.6057215108102395e+02
RS_378 NS_378 0 2.6057215108102395e+02
GL_377 0 NS_377 NS_378 0 2.3565487776505958e-01
GL_378 0 NS_378 NS_377 0 -2.3565487776505958e-01
GS_377_7 0 NS_377 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 379/380
CS_379 NS_379 0 9.9999999999999998e-13
CS_380 NS_380 0 9.9999999999999998e-13
RS_379 NS_379 0 1.4688638444267465e+03
RS_380 NS_380 0 1.4688638444267465e+03
GL_379 0 NS_379 NS_380 0 2.3814510332638331e-01
GL_380 0 NS_380 NS_379 0 -2.3814510332638331e-01
GS_379_7 0 NS_379 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 381/382
CS_381 NS_381 0 9.9999999999999998e-13
CS_382 NS_382 0 9.9999999999999998e-13
RS_381 NS_381 0 1.5351229021400181e+03
RS_382 NS_382 0 1.5351229021400181e+03
GL_381 0 NS_381 NS_382 0 2.5027181856001052e-01
GL_382 0 NS_382 NS_381 0 -2.5027181856001052e-01
GS_381_7 0 NS_381 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 383/384
CS_383 NS_383 0 9.9999999999999998e-13
CS_384 NS_384 0 9.9999999999999998e-13
RS_383 NS_383 0 4.3650646405920685e+02
RS_384 NS_384 0 4.3650646405920685e+02
GL_383 0 NS_383 NS_384 0 2.4893599896984003e-01
GL_384 0 NS_384 NS_383 0 -2.4893599896984003e-01
GS_383_7 0 NS_383 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 385/386
CS_385 NS_385 0 9.9999999999999998e-13
CS_386 NS_386 0 9.9999999999999998e-13
RS_385 NS_385 0 1.1441811687773074e+03
RS_386 NS_386 0 1.1441811687773072e+03
GL_385 0 NS_385 NS_386 0 2.4916499611033449e-01
GL_386 0 NS_386 NS_385 0 -2.4916499611033449e-01
GS_385_7 0 NS_385 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 387/388
CS_387 NS_387 0 9.9999999999999998e-13
CS_388 NS_388 0 9.9999999999999998e-13
RS_387 NS_387 0 7.5335118532932768e+02
RS_388 NS_388 0 7.5335118532932768e+02
GL_387 0 NS_387 NS_388 0 2.4298312011423853e-01
GL_388 0 NS_388 NS_387 0 -2.4298312011423853e-01
GS_387_7 0 NS_387 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 389/390
CS_389 NS_389 0 9.9999999999999998e-13
CS_390 NS_390 0 9.9999999999999998e-13
RS_389 NS_389 0 1.1346596293114915e+03
RS_390 NS_390 0 1.1346596293114915e+03
GL_389 0 NS_389 NS_390 0 2.4551048269503753e-01
GL_390 0 NS_390 NS_389 0 -2.4551048269503753e-01
GS_389_7 0 NS_389 NA_7 0 1.3803457954163372e+00
*
* Complex pair n. 391/392
CS_391 NS_391 0 9.9999999999999998e-13
CS_392 NS_392 0 9.9999999999999998e-13
RS_391 NS_391 0 9.3517666338196523e+02
RS_392 NS_392 0 9.3517666338196523e+02
GL_391 0 NS_391 NS_392 0 2.4538280909205379e-01
GL_392 0 NS_392 NS_391 0 -2.4538280909205379e-01
GS_391_7 0 NS_391 NA_7 0 1.3803457954163372e+00
*
* Real pole n. 393
CS_393 NS_393 0 9.9999999999999998e-13
RS_393 NS_393 0 4.1362120035729779e+00
GS_393_8 0 NS_393 NA_8 0 1.3803457954163372e+00
*
* Real pole n. 394
CS_394 NS_394 0 9.9999999999999998e-13
RS_394 NS_394 0 2.7078253238558993e+01
GS_394_8 0 NS_394 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 395/396
CS_395 NS_395 0 9.9999999999999998e-13
CS_396 NS_396 0 9.9999999999999998e-13
RS_395 NS_395 0 5.6873212206500213e+01
RS_396 NS_396 0 5.6873212206500220e+01
GL_395 0 NS_395 NS_396 0 4.7960934964359665e-02
GL_396 0 NS_396 NS_395 0 -4.7960934964359665e-02
GS_395_8 0 NS_395 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 397/398
CS_397 NS_397 0 9.9999999999999998e-13
CS_398 NS_398 0 9.9999999999999998e-13
RS_397 NS_397 0 5.5832282069998371e+01
RS_398 NS_398 0 5.5832282069998378e+01
GL_397 0 NS_397 NS_398 0 6.1612202840267971e-02
GL_398 0 NS_398 NS_397 0 -6.1612202840267971e-02
GS_397_8 0 NS_397 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 399/400
CS_399 NS_399 0 9.9999999999999998e-13
CS_400 NS_400 0 9.9999999999999998e-13
RS_399 NS_399 0 3.4747519722663924e+01
RS_400 NS_400 0 3.4747519722663924e+01
GL_399 0 NS_399 NS_400 0 8.1784427745819094e-02
GL_400 0 NS_400 NS_399 0 -8.1784427745819094e-02
GS_399_8 0 NS_399 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 401/402
CS_401 NS_401 0 9.9999999999999998e-13
CS_402 NS_402 0 9.9999999999999998e-13
RS_401 NS_401 0 3.1454928782186034e+01
RS_402 NS_402 0 3.1454928782186034e+01
GL_401 0 NS_401 NS_402 0 1.1192538378623762e-01
GL_402 0 NS_402 NS_401 0 -1.1192538378623762e-01
GS_401_8 0 NS_401 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 403/404
CS_403 NS_403 0 9.9999999999999998e-13
CS_404 NS_404 0 9.9999999999999998e-13
RS_403 NS_403 0 2.2209312435826621e+02
RS_404 NS_404 0 2.2209312435826621e+02
GL_403 0 NS_403 NS_404 0 2.9133579865504960e-01
GL_404 0 NS_404 NS_403 0 -2.9133579865504960e-01
GS_403_8 0 NS_403 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 405/406
CS_405 NS_405 0 9.9999999999999998e-13
CS_406 NS_406 0 9.9999999999999998e-13
RS_405 NS_405 0 4.4403718965615290e+01
RS_406 NS_406 0 4.4403718965615283e+01
GL_405 0 NS_405 NS_406 0 1.3869030610195973e-01
GL_406 0 NS_406 NS_405 0 -1.3869030610195973e-01
GS_405_8 0 NS_405 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 407/408
CS_407 NS_407 0 9.9999999999999998e-13
CS_408 NS_408 0 9.9999999999999998e-13
RS_407 NS_407 0 9.2436417727653946e+01
RS_408 NS_408 0 9.2436417727653946e+01
GL_407 0 NS_407 NS_408 0 1.6009535907039132e-01
GL_408 0 NS_408 NS_407 0 -1.6009535907039132e-01
GS_407_8 0 NS_407 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 409/410
CS_409 NS_409 0 9.9999999999999998e-13
CS_410 NS_410 0 9.9999999999999998e-13
RS_409 NS_409 0 5.2247674424140278e+01
RS_410 NS_410 0 5.2247674424140278e+01
GL_409 0 NS_409 NS_410 0 1.7061294296414609e-01
GL_410 0 NS_410 NS_409 0 -1.7061294296414609e-01
GS_409_8 0 NS_409 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 411/412
CS_411 NS_411 0 9.9999999999999998e-13
CS_412 NS_412 0 9.9999999999999998e-13
RS_411 NS_411 0 6.3351631924882277e+01
RS_412 NS_412 0 6.3351631924882277e+01
GL_411 0 NS_411 NS_412 0 1.8578563768540060e-01
GL_412 0 NS_412 NS_411 0 -1.8578563768540060e-01
GS_411_8 0 NS_411 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 413/414
CS_413 NS_413 0 9.9999999999999998e-13
CS_414 NS_414 0 9.9999999999999998e-13
RS_413 NS_413 0 2.2461363612924958e+02
RS_414 NS_414 0 2.2461363612924956e+02
GL_413 0 NS_413 NS_414 0 2.0090890151880786e-01
GL_414 0 NS_414 NS_413 0 -2.0090890151880786e-01
GS_413_8 0 NS_413 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 415/416
CS_415 NS_415 0 9.9999999999999998e-13
CS_416 NS_416 0 9.9999999999999998e-13
RS_415 NS_415 0 6.2323563035856608e+01
RS_416 NS_416 0 6.2323563035856608e+01
GL_415 0 NS_415 NS_416 0 2.0741858581422049e-01
GL_416 0 NS_416 NS_415 0 -2.0741858581422049e-01
GS_415_8 0 NS_415 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 417/418
CS_417 NS_417 0 9.9999999999999998e-13
CS_418 NS_418 0 9.9999999999999998e-13
RS_417 NS_417 0 1.5742148578820314e+02
RS_418 NS_418 0 1.5742148578820311e+02
GL_417 0 NS_417 NS_418 0 2.0543767879537947e-01
GL_418 0 NS_418 NS_417 0 -2.0543767879537947e-01
GS_417_8 0 NS_417 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 419/420
CS_419 NS_419 0 9.9999999999999998e-13
CS_420 NS_420 0 9.9999999999999998e-13
RS_419 NS_419 0 2.0165146427356075e+02
RS_420 NS_420 0 2.0165146427356075e+02
GL_419 0 NS_419 NS_420 0 2.1530071526798281e-01
GL_420 0 NS_420 NS_419 0 -2.1530071526798281e-01
GS_419_8 0 NS_419 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 421/422
CS_421 NS_421 0 9.9999999999999998e-13
CS_422 NS_422 0 9.9999999999999998e-13
RS_421 NS_421 0 2.5655383475382814e+02
RS_422 NS_422 0 2.5655383475382814e+02
GL_421 0 NS_421 NS_422 0 2.2143554872154964e-01
GL_422 0 NS_422 NS_421 0 -2.2143554872154964e-01
GS_421_8 0 NS_421 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 423/424
CS_423 NS_423 0 9.9999999999999998e-13
CS_424 NS_424 0 9.9999999999999998e-13
RS_423 NS_423 0 3.7527533273924564e+02
RS_424 NS_424 0 3.7527533273924570e+02
GL_423 0 NS_423 NS_424 0 2.2416553875794559e-01
GL_424 0 NS_424 NS_423 0 -2.2416553875794559e-01
GS_423_8 0 NS_423 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 425/426
CS_425 NS_425 0 9.9999999999999998e-13
CS_426 NS_426 0 9.9999999999999998e-13
RS_425 NS_425 0 8.7633211379679196e+01
RS_426 NS_426 0 8.7633211379679196e+01
GL_425 0 NS_425 NS_426 0 2.3541329178654702e-01
GL_426 0 NS_426 NS_425 0 -2.3541329178654702e-01
GS_425_8 0 NS_425 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 427/428
CS_427 NS_427 0 9.9999999999999998e-13
CS_428 NS_428 0 9.9999999999999998e-13
RS_427 NS_427 0 4.0937268842404592e+02
RS_428 NS_428 0 4.0937268842404586e+02
GL_427 0 NS_427 NS_428 0 2.2933880932778705e-01
GL_428 0 NS_428 NS_427 0 -2.2933880932778705e-01
GS_427_8 0 NS_427 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 429/430
CS_429 NS_429 0 9.9999999999999998e-13
CS_430 NS_430 0 9.9999999999999998e-13
RS_429 NS_429 0 1.8046101089657725e+02
RS_430 NS_430 0 1.8046101089657725e+02
GL_429 0 NS_429 NS_430 0 2.3011433813523779e-01
GL_430 0 NS_430 NS_429 0 -2.3011433813523779e-01
GS_429_8 0 NS_429 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 431/432
CS_431 NS_431 0 9.9999999999999998e-13
CS_432 NS_432 0 9.9999999999999998e-13
RS_431 NS_431 0 9.7664924917686449e+01
RS_432 NS_432 0 9.7664924917686449e+01
GL_431 0 NS_431 NS_432 0 2.4746563775454208e-01
GL_432 0 NS_432 NS_431 0 -2.4746563775454208e-01
GS_431_8 0 NS_431 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 433/434
CS_433 NS_433 0 9.9999999999999998e-13
CS_434 NS_434 0 9.9999999999999998e-13
RS_433 NS_433 0 2.6057215108102395e+02
RS_434 NS_434 0 2.6057215108102395e+02
GL_433 0 NS_433 NS_434 0 2.3565487776505958e-01
GL_434 0 NS_434 NS_433 0 -2.3565487776505958e-01
GS_433_8 0 NS_433 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 435/436
CS_435 NS_435 0 9.9999999999999998e-13
CS_436 NS_436 0 9.9999999999999998e-13
RS_435 NS_435 0 1.4688638444267465e+03
RS_436 NS_436 0 1.4688638444267465e+03
GL_435 0 NS_435 NS_436 0 2.3814510332638331e-01
GL_436 0 NS_436 NS_435 0 -2.3814510332638331e-01
GS_435_8 0 NS_435 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 437/438
CS_437 NS_437 0 9.9999999999999998e-13
CS_438 NS_438 0 9.9999999999999998e-13
RS_437 NS_437 0 1.5351229021400181e+03
RS_438 NS_438 0 1.5351229021400181e+03
GL_437 0 NS_437 NS_438 0 2.5027181856001052e-01
GL_438 0 NS_438 NS_437 0 -2.5027181856001052e-01
GS_437_8 0 NS_437 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 439/440
CS_439 NS_439 0 9.9999999999999998e-13
CS_440 NS_440 0 9.9999999999999998e-13
RS_439 NS_439 0 4.3650646405920685e+02
RS_440 NS_440 0 4.3650646405920685e+02
GL_439 0 NS_439 NS_440 0 2.4893599896984003e-01
GL_440 0 NS_440 NS_439 0 -2.4893599896984003e-01
GS_439_8 0 NS_439 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 441/442
CS_441 NS_441 0 9.9999999999999998e-13
CS_442 NS_442 0 9.9999999999999998e-13
RS_441 NS_441 0 1.1441811687773074e+03
RS_442 NS_442 0 1.1441811687773072e+03
GL_441 0 NS_441 NS_442 0 2.4916499611033449e-01
GL_442 0 NS_442 NS_441 0 -2.4916499611033449e-01
GS_441_8 0 NS_441 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 443/444
CS_443 NS_443 0 9.9999999999999998e-13
CS_444 NS_444 0 9.9999999999999998e-13
RS_443 NS_443 0 7.5335118532932768e+02
RS_444 NS_444 0 7.5335118532932768e+02
GL_443 0 NS_443 NS_444 0 2.4298312011423853e-01
GL_444 0 NS_444 NS_443 0 -2.4298312011423853e-01
GS_443_8 0 NS_443 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 445/446
CS_445 NS_445 0 9.9999999999999998e-13
CS_446 NS_446 0 9.9999999999999998e-13
RS_445 NS_445 0 1.1346596293114915e+03
RS_446 NS_446 0 1.1346596293114915e+03
GL_445 0 NS_445 NS_446 0 2.4551048269503753e-01
GL_446 0 NS_446 NS_445 0 -2.4551048269503753e-01
GS_445_8 0 NS_445 NA_8 0 1.3803457954163372e+00
*
* Complex pair n. 447/448
CS_447 NS_447 0 9.9999999999999998e-13
CS_448 NS_448 0 9.9999999999999998e-13
RS_447 NS_447 0 9.3517666338196523e+02
RS_448 NS_448 0 9.3517666338196523e+02
GL_447 0 NS_447 NS_448 0 2.4538280909205379e-01
GL_448 0 NS_448 NS_447 0 -2.4538280909205379e-01
GS_447_8 0 NS_447 NA_8 0 1.3803457954163372e+00
*
* Real pole n. 449
CS_449 NS_449 0 9.9999999999999998e-13
RS_449 NS_449 0 4.1362120035729779e+00
GS_449_9 0 NS_449 NA_9 0 1.3803457954163372e+00
*
* Real pole n. 450
CS_450 NS_450 0 9.9999999999999998e-13
RS_450 NS_450 0 2.7078253238558993e+01
GS_450_9 0 NS_450 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 451/452
CS_451 NS_451 0 9.9999999999999998e-13
CS_452 NS_452 0 9.9999999999999998e-13
RS_451 NS_451 0 5.6873212206500213e+01
RS_452 NS_452 0 5.6873212206500220e+01
GL_451 0 NS_451 NS_452 0 4.7960934964359665e-02
GL_452 0 NS_452 NS_451 0 -4.7960934964359665e-02
GS_451_9 0 NS_451 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 453/454
CS_453 NS_453 0 9.9999999999999998e-13
CS_454 NS_454 0 9.9999999999999998e-13
RS_453 NS_453 0 5.5832282069998371e+01
RS_454 NS_454 0 5.5832282069998378e+01
GL_453 0 NS_453 NS_454 0 6.1612202840267971e-02
GL_454 0 NS_454 NS_453 0 -6.1612202840267971e-02
GS_453_9 0 NS_453 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 455/456
CS_455 NS_455 0 9.9999999999999998e-13
CS_456 NS_456 0 9.9999999999999998e-13
RS_455 NS_455 0 3.4747519722663924e+01
RS_456 NS_456 0 3.4747519722663924e+01
GL_455 0 NS_455 NS_456 0 8.1784427745819094e-02
GL_456 0 NS_456 NS_455 0 -8.1784427745819094e-02
GS_455_9 0 NS_455 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 457/458
CS_457 NS_457 0 9.9999999999999998e-13
CS_458 NS_458 0 9.9999999999999998e-13
RS_457 NS_457 0 3.1454928782186034e+01
RS_458 NS_458 0 3.1454928782186034e+01
GL_457 0 NS_457 NS_458 0 1.1192538378623762e-01
GL_458 0 NS_458 NS_457 0 -1.1192538378623762e-01
GS_457_9 0 NS_457 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 459/460
CS_459 NS_459 0 9.9999999999999998e-13
CS_460 NS_460 0 9.9999999999999998e-13
RS_459 NS_459 0 2.2209312435826621e+02
RS_460 NS_460 0 2.2209312435826621e+02
GL_459 0 NS_459 NS_460 0 2.9133579865504960e-01
GL_460 0 NS_460 NS_459 0 -2.9133579865504960e-01
GS_459_9 0 NS_459 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 461/462
CS_461 NS_461 0 9.9999999999999998e-13
CS_462 NS_462 0 9.9999999999999998e-13
RS_461 NS_461 0 4.4403718965615290e+01
RS_462 NS_462 0 4.4403718965615283e+01
GL_461 0 NS_461 NS_462 0 1.3869030610195973e-01
GL_462 0 NS_462 NS_461 0 -1.3869030610195973e-01
GS_461_9 0 NS_461 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 463/464
CS_463 NS_463 0 9.9999999999999998e-13
CS_464 NS_464 0 9.9999999999999998e-13
RS_463 NS_463 0 9.2436417727653946e+01
RS_464 NS_464 0 9.2436417727653946e+01
GL_463 0 NS_463 NS_464 0 1.6009535907039132e-01
GL_464 0 NS_464 NS_463 0 -1.6009535907039132e-01
GS_463_9 0 NS_463 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 465/466
CS_465 NS_465 0 9.9999999999999998e-13
CS_466 NS_466 0 9.9999999999999998e-13
RS_465 NS_465 0 5.2247674424140278e+01
RS_466 NS_466 0 5.2247674424140278e+01
GL_465 0 NS_465 NS_466 0 1.7061294296414609e-01
GL_466 0 NS_466 NS_465 0 -1.7061294296414609e-01
GS_465_9 0 NS_465 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 467/468
CS_467 NS_467 0 9.9999999999999998e-13
CS_468 NS_468 0 9.9999999999999998e-13
RS_467 NS_467 0 6.3351631924882277e+01
RS_468 NS_468 0 6.3351631924882277e+01
GL_467 0 NS_467 NS_468 0 1.8578563768540060e-01
GL_468 0 NS_468 NS_467 0 -1.8578563768540060e-01
GS_467_9 0 NS_467 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 469/470
CS_469 NS_469 0 9.9999999999999998e-13
CS_470 NS_470 0 9.9999999999999998e-13
RS_469 NS_469 0 2.2461363612924958e+02
RS_470 NS_470 0 2.2461363612924956e+02
GL_469 0 NS_469 NS_470 0 2.0090890151880786e-01
GL_470 0 NS_470 NS_469 0 -2.0090890151880786e-01
GS_469_9 0 NS_469 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 471/472
CS_471 NS_471 0 9.9999999999999998e-13
CS_472 NS_472 0 9.9999999999999998e-13
RS_471 NS_471 0 6.2323563035856608e+01
RS_472 NS_472 0 6.2323563035856608e+01
GL_471 0 NS_471 NS_472 0 2.0741858581422049e-01
GL_472 0 NS_472 NS_471 0 -2.0741858581422049e-01
GS_471_9 0 NS_471 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 473/474
CS_473 NS_473 0 9.9999999999999998e-13
CS_474 NS_474 0 9.9999999999999998e-13
RS_473 NS_473 0 1.5742148578820314e+02
RS_474 NS_474 0 1.5742148578820311e+02
GL_473 0 NS_473 NS_474 0 2.0543767879537947e-01
GL_474 0 NS_474 NS_473 0 -2.0543767879537947e-01
GS_473_9 0 NS_473 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 475/476
CS_475 NS_475 0 9.9999999999999998e-13
CS_476 NS_476 0 9.9999999999999998e-13
RS_475 NS_475 0 2.0165146427356075e+02
RS_476 NS_476 0 2.0165146427356075e+02
GL_475 0 NS_475 NS_476 0 2.1530071526798281e-01
GL_476 0 NS_476 NS_475 0 -2.1530071526798281e-01
GS_475_9 0 NS_475 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 477/478
CS_477 NS_477 0 9.9999999999999998e-13
CS_478 NS_478 0 9.9999999999999998e-13
RS_477 NS_477 0 2.5655383475382814e+02
RS_478 NS_478 0 2.5655383475382814e+02
GL_477 0 NS_477 NS_478 0 2.2143554872154964e-01
GL_478 0 NS_478 NS_477 0 -2.2143554872154964e-01
GS_477_9 0 NS_477 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 479/480
CS_479 NS_479 0 9.9999999999999998e-13
CS_480 NS_480 0 9.9999999999999998e-13
RS_479 NS_479 0 3.7527533273924564e+02
RS_480 NS_480 0 3.7527533273924570e+02
GL_479 0 NS_479 NS_480 0 2.2416553875794559e-01
GL_480 0 NS_480 NS_479 0 -2.2416553875794559e-01
GS_479_9 0 NS_479 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 481/482
CS_481 NS_481 0 9.9999999999999998e-13
CS_482 NS_482 0 9.9999999999999998e-13
RS_481 NS_481 0 8.7633211379679196e+01
RS_482 NS_482 0 8.7633211379679196e+01
GL_481 0 NS_481 NS_482 0 2.3541329178654702e-01
GL_482 0 NS_482 NS_481 0 -2.3541329178654702e-01
GS_481_9 0 NS_481 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 483/484
CS_483 NS_483 0 9.9999999999999998e-13
CS_484 NS_484 0 9.9999999999999998e-13
RS_483 NS_483 0 4.0937268842404592e+02
RS_484 NS_484 0 4.0937268842404586e+02
GL_483 0 NS_483 NS_484 0 2.2933880932778705e-01
GL_484 0 NS_484 NS_483 0 -2.2933880932778705e-01
GS_483_9 0 NS_483 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 485/486
CS_485 NS_485 0 9.9999999999999998e-13
CS_486 NS_486 0 9.9999999999999998e-13
RS_485 NS_485 0 1.8046101089657725e+02
RS_486 NS_486 0 1.8046101089657725e+02
GL_485 0 NS_485 NS_486 0 2.3011433813523779e-01
GL_486 0 NS_486 NS_485 0 -2.3011433813523779e-01
GS_485_9 0 NS_485 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 487/488
CS_487 NS_487 0 9.9999999999999998e-13
CS_488 NS_488 0 9.9999999999999998e-13
RS_487 NS_487 0 9.7664924917686449e+01
RS_488 NS_488 0 9.7664924917686449e+01
GL_487 0 NS_487 NS_488 0 2.4746563775454208e-01
GL_488 0 NS_488 NS_487 0 -2.4746563775454208e-01
GS_487_9 0 NS_487 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 489/490
CS_489 NS_489 0 9.9999999999999998e-13
CS_490 NS_490 0 9.9999999999999998e-13
RS_489 NS_489 0 2.6057215108102395e+02
RS_490 NS_490 0 2.6057215108102395e+02
GL_489 0 NS_489 NS_490 0 2.3565487776505958e-01
GL_490 0 NS_490 NS_489 0 -2.3565487776505958e-01
GS_489_9 0 NS_489 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 491/492
CS_491 NS_491 0 9.9999999999999998e-13
CS_492 NS_492 0 9.9999999999999998e-13
RS_491 NS_491 0 1.4688638444267465e+03
RS_492 NS_492 0 1.4688638444267465e+03
GL_491 0 NS_491 NS_492 0 2.3814510332638331e-01
GL_492 0 NS_492 NS_491 0 -2.3814510332638331e-01
GS_491_9 0 NS_491 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 493/494
CS_493 NS_493 0 9.9999999999999998e-13
CS_494 NS_494 0 9.9999999999999998e-13
RS_493 NS_493 0 1.5351229021400181e+03
RS_494 NS_494 0 1.5351229021400181e+03
GL_493 0 NS_493 NS_494 0 2.5027181856001052e-01
GL_494 0 NS_494 NS_493 0 -2.5027181856001052e-01
GS_493_9 0 NS_493 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 495/496
CS_495 NS_495 0 9.9999999999999998e-13
CS_496 NS_496 0 9.9999999999999998e-13
RS_495 NS_495 0 4.3650646405920685e+02
RS_496 NS_496 0 4.3650646405920685e+02
GL_495 0 NS_495 NS_496 0 2.4893599896984003e-01
GL_496 0 NS_496 NS_495 0 -2.4893599896984003e-01
GS_495_9 0 NS_495 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 497/498
CS_497 NS_497 0 9.9999999999999998e-13
CS_498 NS_498 0 9.9999999999999998e-13
RS_497 NS_497 0 1.1441811687773074e+03
RS_498 NS_498 0 1.1441811687773072e+03
GL_497 0 NS_497 NS_498 0 2.4916499611033449e-01
GL_498 0 NS_498 NS_497 0 -2.4916499611033449e-01
GS_497_9 0 NS_497 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 499/500
CS_499 NS_499 0 9.9999999999999998e-13
CS_500 NS_500 0 9.9999999999999998e-13
RS_499 NS_499 0 7.5335118532932768e+02
RS_500 NS_500 0 7.5335118532932768e+02
GL_499 0 NS_499 NS_500 0 2.4298312011423853e-01
GL_500 0 NS_500 NS_499 0 -2.4298312011423853e-01
GS_499_9 0 NS_499 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 501/502
CS_501 NS_501 0 9.9999999999999998e-13
CS_502 NS_502 0 9.9999999999999998e-13
RS_501 NS_501 0 1.1346596293114915e+03
RS_502 NS_502 0 1.1346596293114915e+03
GL_501 0 NS_501 NS_502 0 2.4551048269503753e-01
GL_502 0 NS_502 NS_501 0 -2.4551048269503753e-01
GS_501_9 0 NS_501 NA_9 0 1.3803457954163372e+00
*
* Complex pair n. 503/504
CS_503 NS_503 0 9.9999999999999998e-13
CS_504 NS_504 0 9.9999999999999998e-13
RS_503 NS_503 0 9.3517666338196523e+02
RS_504 NS_504 0 9.3517666338196523e+02
GL_503 0 NS_503 NS_504 0 2.4538280909205379e-01
GL_504 0 NS_504 NS_503 0 -2.4538280909205379e-01
GS_503_9 0 NS_503 NA_9 0 1.3803457954163372e+00
*
* Real pole n. 505
CS_505 NS_505 0 9.9999999999999998e-13
RS_505 NS_505 0 4.1362120035729779e+00
GS_505_10 0 NS_505 NA_10 0 1.3803457954163372e+00
*
* Real pole n. 506
CS_506 NS_506 0 9.9999999999999998e-13
RS_506 NS_506 0 2.7078253238558993e+01
GS_506_10 0 NS_506 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 507/508
CS_507 NS_507 0 9.9999999999999998e-13
CS_508 NS_508 0 9.9999999999999998e-13
RS_507 NS_507 0 5.6873212206500213e+01
RS_508 NS_508 0 5.6873212206500220e+01
GL_507 0 NS_507 NS_508 0 4.7960934964359665e-02
GL_508 0 NS_508 NS_507 0 -4.7960934964359665e-02
GS_507_10 0 NS_507 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 509/510
CS_509 NS_509 0 9.9999999999999998e-13
CS_510 NS_510 0 9.9999999999999998e-13
RS_509 NS_509 0 5.5832282069998371e+01
RS_510 NS_510 0 5.5832282069998378e+01
GL_509 0 NS_509 NS_510 0 6.1612202840267971e-02
GL_510 0 NS_510 NS_509 0 -6.1612202840267971e-02
GS_509_10 0 NS_509 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 511/512
CS_511 NS_511 0 9.9999999999999998e-13
CS_512 NS_512 0 9.9999999999999998e-13
RS_511 NS_511 0 3.4747519722663924e+01
RS_512 NS_512 0 3.4747519722663924e+01
GL_511 0 NS_511 NS_512 0 8.1784427745819094e-02
GL_512 0 NS_512 NS_511 0 -8.1784427745819094e-02
GS_511_10 0 NS_511 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 513/514
CS_513 NS_513 0 9.9999999999999998e-13
CS_514 NS_514 0 9.9999999999999998e-13
RS_513 NS_513 0 3.1454928782186034e+01
RS_514 NS_514 0 3.1454928782186034e+01
GL_513 0 NS_513 NS_514 0 1.1192538378623762e-01
GL_514 0 NS_514 NS_513 0 -1.1192538378623762e-01
GS_513_10 0 NS_513 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 515/516
CS_515 NS_515 0 9.9999999999999998e-13
CS_516 NS_516 0 9.9999999999999998e-13
RS_515 NS_515 0 2.2209312435826621e+02
RS_516 NS_516 0 2.2209312435826621e+02
GL_515 0 NS_515 NS_516 0 2.9133579865504960e-01
GL_516 0 NS_516 NS_515 0 -2.9133579865504960e-01
GS_515_10 0 NS_515 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 517/518
CS_517 NS_517 0 9.9999999999999998e-13
CS_518 NS_518 0 9.9999999999999998e-13
RS_517 NS_517 0 4.4403718965615290e+01
RS_518 NS_518 0 4.4403718965615283e+01
GL_517 0 NS_517 NS_518 0 1.3869030610195973e-01
GL_518 0 NS_518 NS_517 0 -1.3869030610195973e-01
GS_517_10 0 NS_517 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 519/520
CS_519 NS_519 0 9.9999999999999998e-13
CS_520 NS_520 0 9.9999999999999998e-13
RS_519 NS_519 0 9.2436417727653946e+01
RS_520 NS_520 0 9.2436417727653946e+01
GL_519 0 NS_519 NS_520 0 1.6009535907039132e-01
GL_520 0 NS_520 NS_519 0 -1.6009535907039132e-01
GS_519_10 0 NS_519 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 521/522
CS_521 NS_521 0 9.9999999999999998e-13
CS_522 NS_522 0 9.9999999999999998e-13
RS_521 NS_521 0 5.2247674424140278e+01
RS_522 NS_522 0 5.2247674424140278e+01
GL_521 0 NS_521 NS_522 0 1.7061294296414609e-01
GL_522 0 NS_522 NS_521 0 -1.7061294296414609e-01
GS_521_10 0 NS_521 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 523/524
CS_523 NS_523 0 9.9999999999999998e-13
CS_524 NS_524 0 9.9999999999999998e-13
RS_523 NS_523 0 6.3351631924882277e+01
RS_524 NS_524 0 6.3351631924882277e+01
GL_523 0 NS_523 NS_524 0 1.8578563768540060e-01
GL_524 0 NS_524 NS_523 0 -1.8578563768540060e-01
GS_523_10 0 NS_523 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 525/526
CS_525 NS_525 0 9.9999999999999998e-13
CS_526 NS_526 0 9.9999999999999998e-13
RS_525 NS_525 0 2.2461363612924958e+02
RS_526 NS_526 0 2.2461363612924956e+02
GL_525 0 NS_525 NS_526 0 2.0090890151880786e-01
GL_526 0 NS_526 NS_525 0 -2.0090890151880786e-01
GS_525_10 0 NS_525 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 527/528
CS_527 NS_527 0 9.9999999999999998e-13
CS_528 NS_528 0 9.9999999999999998e-13
RS_527 NS_527 0 6.2323563035856608e+01
RS_528 NS_528 0 6.2323563035856608e+01
GL_527 0 NS_527 NS_528 0 2.0741858581422049e-01
GL_528 0 NS_528 NS_527 0 -2.0741858581422049e-01
GS_527_10 0 NS_527 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 529/530
CS_529 NS_529 0 9.9999999999999998e-13
CS_530 NS_530 0 9.9999999999999998e-13
RS_529 NS_529 0 1.5742148578820314e+02
RS_530 NS_530 0 1.5742148578820311e+02
GL_529 0 NS_529 NS_530 0 2.0543767879537947e-01
GL_530 0 NS_530 NS_529 0 -2.0543767879537947e-01
GS_529_10 0 NS_529 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 531/532
CS_531 NS_531 0 9.9999999999999998e-13
CS_532 NS_532 0 9.9999999999999998e-13
RS_531 NS_531 0 2.0165146427356075e+02
RS_532 NS_532 0 2.0165146427356075e+02
GL_531 0 NS_531 NS_532 0 2.1530071526798281e-01
GL_532 0 NS_532 NS_531 0 -2.1530071526798281e-01
GS_531_10 0 NS_531 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 533/534
CS_533 NS_533 0 9.9999999999999998e-13
CS_534 NS_534 0 9.9999999999999998e-13
RS_533 NS_533 0 2.5655383475382814e+02
RS_534 NS_534 0 2.5655383475382814e+02
GL_533 0 NS_533 NS_534 0 2.2143554872154964e-01
GL_534 0 NS_534 NS_533 0 -2.2143554872154964e-01
GS_533_10 0 NS_533 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 535/536
CS_535 NS_535 0 9.9999999999999998e-13
CS_536 NS_536 0 9.9999999999999998e-13
RS_535 NS_535 0 3.7527533273924564e+02
RS_536 NS_536 0 3.7527533273924570e+02
GL_535 0 NS_535 NS_536 0 2.2416553875794559e-01
GL_536 0 NS_536 NS_535 0 -2.2416553875794559e-01
GS_535_10 0 NS_535 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 537/538
CS_537 NS_537 0 9.9999999999999998e-13
CS_538 NS_538 0 9.9999999999999998e-13
RS_537 NS_537 0 8.7633211379679196e+01
RS_538 NS_538 0 8.7633211379679196e+01
GL_537 0 NS_537 NS_538 0 2.3541329178654702e-01
GL_538 0 NS_538 NS_537 0 -2.3541329178654702e-01
GS_537_10 0 NS_537 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 539/540
CS_539 NS_539 0 9.9999999999999998e-13
CS_540 NS_540 0 9.9999999999999998e-13
RS_539 NS_539 0 4.0937268842404592e+02
RS_540 NS_540 0 4.0937268842404586e+02
GL_539 0 NS_539 NS_540 0 2.2933880932778705e-01
GL_540 0 NS_540 NS_539 0 -2.2933880932778705e-01
GS_539_10 0 NS_539 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 541/542
CS_541 NS_541 0 9.9999999999999998e-13
CS_542 NS_542 0 9.9999999999999998e-13
RS_541 NS_541 0 1.8046101089657725e+02
RS_542 NS_542 0 1.8046101089657725e+02
GL_541 0 NS_541 NS_542 0 2.3011433813523779e-01
GL_542 0 NS_542 NS_541 0 -2.3011433813523779e-01
GS_541_10 0 NS_541 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 543/544
CS_543 NS_543 0 9.9999999999999998e-13
CS_544 NS_544 0 9.9999999999999998e-13
RS_543 NS_543 0 9.7664924917686449e+01
RS_544 NS_544 0 9.7664924917686449e+01
GL_543 0 NS_543 NS_544 0 2.4746563775454208e-01
GL_544 0 NS_544 NS_543 0 -2.4746563775454208e-01
GS_543_10 0 NS_543 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 545/546
CS_545 NS_545 0 9.9999999999999998e-13
CS_546 NS_546 0 9.9999999999999998e-13
RS_545 NS_545 0 2.6057215108102395e+02
RS_546 NS_546 0 2.6057215108102395e+02
GL_545 0 NS_545 NS_546 0 2.3565487776505958e-01
GL_546 0 NS_546 NS_545 0 -2.3565487776505958e-01
GS_545_10 0 NS_545 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 547/548
CS_547 NS_547 0 9.9999999999999998e-13
CS_548 NS_548 0 9.9999999999999998e-13
RS_547 NS_547 0 1.4688638444267465e+03
RS_548 NS_548 0 1.4688638444267465e+03
GL_547 0 NS_547 NS_548 0 2.3814510332638331e-01
GL_548 0 NS_548 NS_547 0 -2.3814510332638331e-01
GS_547_10 0 NS_547 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 549/550
CS_549 NS_549 0 9.9999999999999998e-13
CS_550 NS_550 0 9.9999999999999998e-13
RS_549 NS_549 0 1.5351229021400181e+03
RS_550 NS_550 0 1.5351229021400181e+03
GL_549 0 NS_549 NS_550 0 2.5027181856001052e-01
GL_550 0 NS_550 NS_549 0 -2.5027181856001052e-01
GS_549_10 0 NS_549 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 551/552
CS_551 NS_551 0 9.9999999999999998e-13
CS_552 NS_552 0 9.9999999999999998e-13
RS_551 NS_551 0 4.3650646405920685e+02
RS_552 NS_552 0 4.3650646405920685e+02
GL_551 0 NS_551 NS_552 0 2.4893599896984003e-01
GL_552 0 NS_552 NS_551 0 -2.4893599896984003e-01
GS_551_10 0 NS_551 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 553/554
CS_553 NS_553 0 9.9999999999999998e-13
CS_554 NS_554 0 9.9999999999999998e-13
RS_553 NS_553 0 1.1441811687773074e+03
RS_554 NS_554 0 1.1441811687773072e+03
GL_553 0 NS_553 NS_554 0 2.4916499611033449e-01
GL_554 0 NS_554 NS_553 0 -2.4916499611033449e-01
GS_553_10 0 NS_553 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 555/556
CS_555 NS_555 0 9.9999999999999998e-13
CS_556 NS_556 0 9.9999999999999998e-13
RS_555 NS_555 0 7.5335118532932768e+02
RS_556 NS_556 0 7.5335118532932768e+02
GL_555 0 NS_555 NS_556 0 2.4298312011423853e-01
GL_556 0 NS_556 NS_555 0 -2.4298312011423853e-01
GS_555_10 0 NS_555 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 557/558
CS_557 NS_557 0 9.9999999999999998e-13
CS_558 NS_558 0 9.9999999999999998e-13
RS_557 NS_557 0 1.1346596293114915e+03
RS_558 NS_558 0 1.1346596293114915e+03
GL_557 0 NS_557 NS_558 0 2.4551048269503753e-01
GL_558 0 NS_558 NS_557 0 -2.4551048269503753e-01
GS_557_10 0 NS_557 NA_10 0 1.3803457954163372e+00
*
* Complex pair n. 559/560
CS_559 NS_559 0 9.9999999999999998e-13
CS_560 NS_560 0 9.9999999999999998e-13
RS_559 NS_559 0 9.3517666338196523e+02
RS_560 NS_560 0 9.3517666338196523e+02
GL_559 0 NS_559 NS_560 0 2.4538280909205379e-01
GL_560 0 NS_560 NS_559 0 -2.4538280909205379e-01
GS_559_10 0 NS_559 NA_10 0 1.3803457954163372e+00
*
* Real pole n. 561
CS_561 NS_561 0 9.9999999999999998e-13
RS_561 NS_561 0 4.1362120035729779e+00
GS_561_11 0 NS_561 NA_11 0 1.3803457954163372e+00
*
* Real pole n. 562
CS_562 NS_562 0 9.9999999999999998e-13
RS_562 NS_562 0 2.7078253238558993e+01
GS_562_11 0 NS_562 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 563/564
CS_563 NS_563 0 9.9999999999999998e-13
CS_564 NS_564 0 9.9999999999999998e-13
RS_563 NS_563 0 5.6873212206500213e+01
RS_564 NS_564 0 5.6873212206500220e+01
GL_563 0 NS_563 NS_564 0 4.7960934964359665e-02
GL_564 0 NS_564 NS_563 0 -4.7960934964359665e-02
GS_563_11 0 NS_563 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 565/566
CS_565 NS_565 0 9.9999999999999998e-13
CS_566 NS_566 0 9.9999999999999998e-13
RS_565 NS_565 0 5.5832282069998371e+01
RS_566 NS_566 0 5.5832282069998378e+01
GL_565 0 NS_565 NS_566 0 6.1612202840267971e-02
GL_566 0 NS_566 NS_565 0 -6.1612202840267971e-02
GS_565_11 0 NS_565 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 567/568
CS_567 NS_567 0 9.9999999999999998e-13
CS_568 NS_568 0 9.9999999999999998e-13
RS_567 NS_567 0 3.4747519722663924e+01
RS_568 NS_568 0 3.4747519722663924e+01
GL_567 0 NS_567 NS_568 0 8.1784427745819094e-02
GL_568 0 NS_568 NS_567 0 -8.1784427745819094e-02
GS_567_11 0 NS_567 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 569/570
CS_569 NS_569 0 9.9999999999999998e-13
CS_570 NS_570 0 9.9999999999999998e-13
RS_569 NS_569 0 3.1454928782186034e+01
RS_570 NS_570 0 3.1454928782186034e+01
GL_569 0 NS_569 NS_570 0 1.1192538378623762e-01
GL_570 0 NS_570 NS_569 0 -1.1192538378623762e-01
GS_569_11 0 NS_569 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 571/572
CS_571 NS_571 0 9.9999999999999998e-13
CS_572 NS_572 0 9.9999999999999998e-13
RS_571 NS_571 0 2.2209312435826621e+02
RS_572 NS_572 0 2.2209312435826621e+02
GL_571 0 NS_571 NS_572 0 2.9133579865504960e-01
GL_572 0 NS_572 NS_571 0 -2.9133579865504960e-01
GS_571_11 0 NS_571 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 573/574
CS_573 NS_573 0 9.9999999999999998e-13
CS_574 NS_574 0 9.9999999999999998e-13
RS_573 NS_573 0 4.4403718965615290e+01
RS_574 NS_574 0 4.4403718965615283e+01
GL_573 0 NS_573 NS_574 0 1.3869030610195973e-01
GL_574 0 NS_574 NS_573 0 -1.3869030610195973e-01
GS_573_11 0 NS_573 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 575/576
CS_575 NS_575 0 9.9999999999999998e-13
CS_576 NS_576 0 9.9999999999999998e-13
RS_575 NS_575 0 9.2436417727653946e+01
RS_576 NS_576 0 9.2436417727653946e+01
GL_575 0 NS_575 NS_576 0 1.6009535907039132e-01
GL_576 0 NS_576 NS_575 0 -1.6009535907039132e-01
GS_575_11 0 NS_575 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 577/578
CS_577 NS_577 0 9.9999999999999998e-13
CS_578 NS_578 0 9.9999999999999998e-13
RS_577 NS_577 0 5.2247674424140278e+01
RS_578 NS_578 0 5.2247674424140278e+01
GL_577 0 NS_577 NS_578 0 1.7061294296414609e-01
GL_578 0 NS_578 NS_577 0 -1.7061294296414609e-01
GS_577_11 0 NS_577 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 579/580
CS_579 NS_579 0 9.9999999999999998e-13
CS_580 NS_580 0 9.9999999999999998e-13
RS_579 NS_579 0 6.3351631924882277e+01
RS_580 NS_580 0 6.3351631924882277e+01
GL_579 0 NS_579 NS_580 0 1.8578563768540060e-01
GL_580 0 NS_580 NS_579 0 -1.8578563768540060e-01
GS_579_11 0 NS_579 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 581/582
CS_581 NS_581 0 9.9999999999999998e-13
CS_582 NS_582 0 9.9999999999999998e-13
RS_581 NS_581 0 2.2461363612924958e+02
RS_582 NS_582 0 2.2461363612924956e+02
GL_581 0 NS_581 NS_582 0 2.0090890151880786e-01
GL_582 0 NS_582 NS_581 0 -2.0090890151880786e-01
GS_581_11 0 NS_581 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 583/584
CS_583 NS_583 0 9.9999999999999998e-13
CS_584 NS_584 0 9.9999999999999998e-13
RS_583 NS_583 0 6.2323563035856608e+01
RS_584 NS_584 0 6.2323563035856608e+01
GL_583 0 NS_583 NS_584 0 2.0741858581422049e-01
GL_584 0 NS_584 NS_583 0 -2.0741858581422049e-01
GS_583_11 0 NS_583 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 585/586
CS_585 NS_585 0 9.9999999999999998e-13
CS_586 NS_586 0 9.9999999999999998e-13
RS_585 NS_585 0 1.5742148578820314e+02
RS_586 NS_586 0 1.5742148578820311e+02
GL_585 0 NS_585 NS_586 0 2.0543767879537947e-01
GL_586 0 NS_586 NS_585 0 -2.0543767879537947e-01
GS_585_11 0 NS_585 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 587/588
CS_587 NS_587 0 9.9999999999999998e-13
CS_588 NS_588 0 9.9999999999999998e-13
RS_587 NS_587 0 2.0165146427356075e+02
RS_588 NS_588 0 2.0165146427356075e+02
GL_587 0 NS_587 NS_588 0 2.1530071526798281e-01
GL_588 0 NS_588 NS_587 0 -2.1530071526798281e-01
GS_587_11 0 NS_587 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 589/590
CS_589 NS_589 0 9.9999999999999998e-13
CS_590 NS_590 0 9.9999999999999998e-13
RS_589 NS_589 0 2.5655383475382814e+02
RS_590 NS_590 0 2.5655383475382814e+02
GL_589 0 NS_589 NS_590 0 2.2143554872154964e-01
GL_590 0 NS_590 NS_589 0 -2.2143554872154964e-01
GS_589_11 0 NS_589 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 591/592
CS_591 NS_591 0 9.9999999999999998e-13
CS_592 NS_592 0 9.9999999999999998e-13
RS_591 NS_591 0 3.7527533273924564e+02
RS_592 NS_592 0 3.7527533273924570e+02
GL_591 0 NS_591 NS_592 0 2.2416553875794559e-01
GL_592 0 NS_592 NS_591 0 -2.2416553875794559e-01
GS_591_11 0 NS_591 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 593/594
CS_593 NS_593 0 9.9999999999999998e-13
CS_594 NS_594 0 9.9999999999999998e-13
RS_593 NS_593 0 8.7633211379679196e+01
RS_594 NS_594 0 8.7633211379679196e+01
GL_593 0 NS_593 NS_594 0 2.3541329178654702e-01
GL_594 0 NS_594 NS_593 0 -2.3541329178654702e-01
GS_593_11 0 NS_593 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 595/596
CS_595 NS_595 0 9.9999999999999998e-13
CS_596 NS_596 0 9.9999999999999998e-13
RS_595 NS_595 0 4.0937268842404592e+02
RS_596 NS_596 0 4.0937268842404586e+02
GL_595 0 NS_595 NS_596 0 2.2933880932778705e-01
GL_596 0 NS_596 NS_595 0 -2.2933880932778705e-01
GS_595_11 0 NS_595 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 597/598
CS_597 NS_597 0 9.9999999999999998e-13
CS_598 NS_598 0 9.9999999999999998e-13
RS_597 NS_597 0 1.8046101089657725e+02
RS_598 NS_598 0 1.8046101089657725e+02
GL_597 0 NS_597 NS_598 0 2.3011433813523779e-01
GL_598 0 NS_598 NS_597 0 -2.3011433813523779e-01
GS_597_11 0 NS_597 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 599/600
CS_599 NS_599 0 9.9999999999999998e-13
CS_600 NS_600 0 9.9999999999999998e-13
RS_599 NS_599 0 9.7664924917686449e+01
RS_600 NS_600 0 9.7664924917686449e+01
GL_599 0 NS_599 NS_600 0 2.4746563775454208e-01
GL_600 0 NS_600 NS_599 0 -2.4746563775454208e-01
GS_599_11 0 NS_599 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 601/602
CS_601 NS_601 0 9.9999999999999998e-13
CS_602 NS_602 0 9.9999999999999998e-13
RS_601 NS_601 0 2.6057215108102395e+02
RS_602 NS_602 0 2.6057215108102395e+02
GL_601 0 NS_601 NS_602 0 2.3565487776505958e-01
GL_602 0 NS_602 NS_601 0 -2.3565487776505958e-01
GS_601_11 0 NS_601 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 603/604
CS_603 NS_603 0 9.9999999999999998e-13
CS_604 NS_604 0 9.9999999999999998e-13
RS_603 NS_603 0 1.4688638444267465e+03
RS_604 NS_604 0 1.4688638444267465e+03
GL_603 0 NS_603 NS_604 0 2.3814510332638331e-01
GL_604 0 NS_604 NS_603 0 -2.3814510332638331e-01
GS_603_11 0 NS_603 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 605/606
CS_605 NS_605 0 9.9999999999999998e-13
CS_606 NS_606 0 9.9999999999999998e-13
RS_605 NS_605 0 1.5351229021400181e+03
RS_606 NS_606 0 1.5351229021400181e+03
GL_605 0 NS_605 NS_606 0 2.5027181856001052e-01
GL_606 0 NS_606 NS_605 0 -2.5027181856001052e-01
GS_605_11 0 NS_605 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 607/608
CS_607 NS_607 0 9.9999999999999998e-13
CS_608 NS_608 0 9.9999999999999998e-13
RS_607 NS_607 0 4.3650646405920685e+02
RS_608 NS_608 0 4.3650646405920685e+02
GL_607 0 NS_607 NS_608 0 2.4893599896984003e-01
GL_608 0 NS_608 NS_607 0 -2.4893599896984003e-01
GS_607_11 0 NS_607 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 609/610
CS_609 NS_609 0 9.9999999999999998e-13
CS_610 NS_610 0 9.9999999999999998e-13
RS_609 NS_609 0 1.1441811687773074e+03
RS_610 NS_610 0 1.1441811687773072e+03
GL_609 0 NS_609 NS_610 0 2.4916499611033449e-01
GL_610 0 NS_610 NS_609 0 -2.4916499611033449e-01
GS_609_11 0 NS_609 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 611/612
CS_611 NS_611 0 9.9999999999999998e-13
CS_612 NS_612 0 9.9999999999999998e-13
RS_611 NS_611 0 7.5335118532932768e+02
RS_612 NS_612 0 7.5335118532932768e+02
GL_611 0 NS_611 NS_612 0 2.4298312011423853e-01
GL_612 0 NS_612 NS_611 0 -2.4298312011423853e-01
GS_611_11 0 NS_611 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 613/614
CS_613 NS_613 0 9.9999999999999998e-13
CS_614 NS_614 0 9.9999999999999998e-13
RS_613 NS_613 0 1.1346596293114915e+03
RS_614 NS_614 0 1.1346596293114915e+03
GL_613 0 NS_613 NS_614 0 2.4551048269503753e-01
GL_614 0 NS_614 NS_613 0 -2.4551048269503753e-01
GS_613_11 0 NS_613 NA_11 0 1.3803457954163372e+00
*
* Complex pair n. 615/616
CS_615 NS_615 0 9.9999999999999998e-13
CS_616 NS_616 0 9.9999999999999998e-13
RS_615 NS_615 0 9.3517666338196523e+02
RS_616 NS_616 0 9.3517666338196523e+02
GL_615 0 NS_615 NS_616 0 2.4538280909205379e-01
GL_616 0 NS_616 NS_615 0 -2.4538280909205379e-01
GS_615_11 0 NS_615 NA_11 0 1.3803457954163372e+00
*
* Real pole n. 617
CS_617 NS_617 0 9.9999999999999998e-13
RS_617 NS_617 0 4.1362120035729779e+00
GS_617_12 0 NS_617 NA_12 0 1.3803457954163372e+00
*
* Real pole n. 618
CS_618 NS_618 0 9.9999999999999998e-13
RS_618 NS_618 0 2.7078253238558993e+01
GS_618_12 0 NS_618 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 619/620
CS_619 NS_619 0 9.9999999999999998e-13
CS_620 NS_620 0 9.9999999999999998e-13
RS_619 NS_619 0 5.6873212206500213e+01
RS_620 NS_620 0 5.6873212206500220e+01
GL_619 0 NS_619 NS_620 0 4.7960934964359665e-02
GL_620 0 NS_620 NS_619 0 -4.7960934964359665e-02
GS_619_12 0 NS_619 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 621/622
CS_621 NS_621 0 9.9999999999999998e-13
CS_622 NS_622 0 9.9999999999999998e-13
RS_621 NS_621 0 5.5832282069998371e+01
RS_622 NS_622 0 5.5832282069998378e+01
GL_621 0 NS_621 NS_622 0 6.1612202840267971e-02
GL_622 0 NS_622 NS_621 0 -6.1612202840267971e-02
GS_621_12 0 NS_621 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 623/624
CS_623 NS_623 0 9.9999999999999998e-13
CS_624 NS_624 0 9.9999999999999998e-13
RS_623 NS_623 0 3.4747519722663924e+01
RS_624 NS_624 0 3.4747519722663924e+01
GL_623 0 NS_623 NS_624 0 8.1784427745819094e-02
GL_624 0 NS_624 NS_623 0 -8.1784427745819094e-02
GS_623_12 0 NS_623 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 625/626
CS_625 NS_625 0 9.9999999999999998e-13
CS_626 NS_626 0 9.9999999999999998e-13
RS_625 NS_625 0 3.1454928782186034e+01
RS_626 NS_626 0 3.1454928782186034e+01
GL_625 0 NS_625 NS_626 0 1.1192538378623762e-01
GL_626 0 NS_626 NS_625 0 -1.1192538378623762e-01
GS_625_12 0 NS_625 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 627/628
CS_627 NS_627 0 9.9999999999999998e-13
CS_628 NS_628 0 9.9999999999999998e-13
RS_627 NS_627 0 2.2209312435826621e+02
RS_628 NS_628 0 2.2209312435826621e+02
GL_627 0 NS_627 NS_628 0 2.9133579865504960e-01
GL_628 0 NS_628 NS_627 0 -2.9133579865504960e-01
GS_627_12 0 NS_627 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 629/630
CS_629 NS_629 0 9.9999999999999998e-13
CS_630 NS_630 0 9.9999999999999998e-13
RS_629 NS_629 0 4.4403718965615290e+01
RS_630 NS_630 0 4.4403718965615283e+01
GL_629 0 NS_629 NS_630 0 1.3869030610195973e-01
GL_630 0 NS_630 NS_629 0 -1.3869030610195973e-01
GS_629_12 0 NS_629 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 631/632
CS_631 NS_631 0 9.9999999999999998e-13
CS_632 NS_632 0 9.9999999999999998e-13
RS_631 NS_631 0 9.2436417727653946e+01
RS_632 NS_632 0 9.2436417727653946e+01
GL_631 0 NS_631 NS_632 0 1.6009535907039132e-01
GL_632 0 NS_632 NS_631 0 -1.6009535907039132e-01
GS_631_12 0 NS_631 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 633/634
CS_633 NS_633 0 9.9999999999999998e-13
CS_634 NS_634 0 9.9999999999999998e-13
RS_633 NS_633 0 5.2247674424140278e+01
RS_634 NS_634 0 5.2247674424140278e+01
GL_633 0 NS_633 NS_634 0 1.7061294296414609e-01
GL_634 0 NS_634 NS_633 0 -1.7061294296414609e-01
GS_633_12 0 NS_633 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 635/636
CS_635 NS_635 0 9.9999999999999998e-13
CS_636 NS_636 0 9.9999999999999998e-13
RS_635 NS_635 0 6.3351631924882277e+01
RS_636 NS_636 0 6.3351631924882277e+01
GL_635 0 NS_635 NS_636 0 1.8578563768540060e-01
GL_636 0 NS_636 NS_635 0 -1.8578563768540060e-01
GS_635_12 0 NS_635 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 637/638
CS_637 NS_637 0 9.9999999999999998e-13
CS_638 NS_638 0 9.9999999999999998e-13
RS_637 NS_637 0 2.2461363612924958e+02
RS_638 NS_638 0 2.2461363612924956e+02
GL_637 0 NS_637 NS_638 0 2.0090890151880786e-01
GL_638 0 NS_638 NS_637 0 -2.0090890151880786e-01
GS_637_12 0 NS_637 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 639/640
CS_639 NS_639 0 9.9999999999999998e-13
CS_640 NS_640 0 9.9999999999999998e-13
RS_639 NS_639 0 6.2323563035856608e+01
RS_640 NS_640 0 6.2323563035856608e+01
GL_639 0 NS_639 NS_640 0 2.0741858581422049e-01
GL_640 0 NS_640 NS_639 0 -2.0741858581422049e-01
GS_639_12 0 NS_639 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 641/642
CS_641 NS_641 0 9.9999999999999998e-13
CS_642 NS_642 0 9.9999999999999998e-13
RS_641 NS_641 0 1.5742148578820314e+02
RS_642 NS_642 0 1.5742148578820311e+02
GL_641 0 NS_641 NS_642 0 2.0543767879537947e-01
GL_642 0 NS_642 NS_641 0 -2.0543767879537947e-01
GS_641_12 0 NS_641 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 643/644
CS_643 NS_643 0 9.9999999999999998e-13
CS_644 NS_644 0 9.9999999999999998e-13
RS_643 NS_643 0 2.0165146427356075e+02
RS_644 NS_644 0 2.0165146427356075e+02
GL_643 0 NS_643 NS_644 0 2.1530071526798281e-01
GL_644 0 NS_644 NS_643 0 -2.1530071526798281e-01
GS_643_12 0 NS_643 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 645/646
CS_645 NS_645 0 9.9999999999999998e-13
CS_646 NS_646 0 9.9999999999999998e-13
RS_645 NS_645 0 2.5655383475382814e+02
RS_646 NS_646 0 2.5655383475382814e+02
GL_645 0 NS_645 NS_646 0 2.2143554872154964e-01
GL_646 0 NS_646 NS_645 0 -2.2143554872154964e-01
GS_645_12 0 NS_645 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 647/648
CS_647 NS_647 0 9.9999999999999998e-13
CS_648 NS_648 0 9.9999999999999998e-13
RS_647 NS_647 0 3.7527533273924564e+02
RS_648 NS_648 0 3.7527533273924570e+02
GL_647 0 NS_647 NS_648 0 2.2416553875794559e-01
GL_648 0 NS_648 NS_647 0 -2.2416553875794559e-01
GS_647_12 0 NS_647 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 649/650
CS_649 NS_649 0 9.9999999999999998e-13
CS_650 NS_650 0 9.9999999999999998e-13
RS_649 NS_649 0 8.7633211379679196e+01
RS_650 NS_650 0 8.7633211379679196e+01
GL_649 0 NS_649 NS_650 0 2.3541329178654702e-01
GL_650 0 NS_650 NS_649 0 -2.3541329178654702e-01
GS_649_12 0 NS_649 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 651/652
CS_651 NS_651 0 9.9999999999999998e-13
CS_652 NS_652 0 9.9999999999999998e-13
RS_651 NS_651 0 4.0937268842404592e+02
RS_652 NS_652 0 4.0937268842404586e+02
GL_651 0 NS_651 NS_652 0 2.2933880932778705e-01
GL_652 0 NS_652 NS_651 0 -2.2933880932778705e-01
GS_651_12 0 NS_651 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 653/654
CS_653 NS_653 0 9.9999999999999998e-13
CS_654 NS_654 0 9.9999999999999998e-13
RS_653 NS_653 0 1.8046101089657725e+02
RS_654 NS_654 0 1.8046101089657725e+02
GL_653 0 NS_653 NS_654 0 2.3011433813523779e-01
GL_654 0 NS_654 NS_653 0 -2.3011433813523779e-01
GS_653_12 0 NS_653 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 655/656
CS_655 NS_655 0 9.9999999999999998e-13
CS_656 NS_656 0 9.9999999999999998e-13
RS_655 NS_655 0 9.7664924917686449e+01
RS_656 NS_656 0 9.7664924917686449e+01
GL_655 0 NS_655 NS_656 0 2.4746563775454208e-01
GL_656 0 NS_656 NS_655 0 -2.4746563775454208e-01
GS_655_12 0 NS_655 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 657/658
CS_657 NS_657 0 9.9999999999999998e-13
CS_658 NS_658 0 9.9999999999999998e-13
RS_657 NS_657 0 2.6057215108102395e+02
RS_658 NS_658 0 2.6057215108102395e+02
GL_657 0 NS_657 NS_658 0 2.3565487776505958e-01
GL_658 0 NS_658 NS_657 0 -2.3565487776505958e-01
GS_657_12 0 NS_657 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 659/660
CS_659 NS_659 0 9.9999999999999998e-13
CS_660 NS_660 0 9.9999999999999998e-13
RS_659 NS_659 0 1.4688638444267465e+03
RS_660 NS_660 0 1.4688638444267465e+03
GL_659 0 NS_659 NS_660 0 2.3814510332638331e-01
GL_660 0 NS_660 NS_659 0 -2.3814510332638331e-01
GS_659_12 0 NS_659 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 661/662
CS_661 NS_661 0 9.9999999999999998e-13
CS_662 NS_662 0 9.9999999999999998e-13
RS_661 NS_661 0 1.5351229021400181e+03
RS_662 NS_662 0 1.5351229021400181e+03
GL_661 0 NS_661 NS_662 0 2.5027181856001052e-01
GL_662 0 NS_662 NS_661 0 -2.5027181856001052e-01
GS_661_12 0 NS_661 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 663/664
CS_663 NS_663 0 9.9999999999999998e-13
CS_664 NS_664 0 9.9999999999999998e-13
RS_663 NS_663 0 4.3650646405920685e+02
RS_664 NS_664 0 4.3650646405920685e+02
GL_663 0 NS_663 NS_664 0 2.4893599896984003e-01
GL_664 0 NS_664 NS_663 0 -2.4893599896984003e-01
GS_663_12 0 NS_663 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 665/666
CS_665 NS_665 0 9.9999999999999998e-13
CS_666 NS_666 0 9.9999999999999998e-13
RS_665 NS_665 0 1.1441811687773074e+03
RS_666 NS_666 0 1.1441811687773072e+03
GL_665 0 NS_665 NS_666 0 2.4916499611033449e-01
GL_666 0 NS_666 NS_665 0 -2.4916499611033449e-01
GS_665_12 0 NS_665 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 667/668
CS_667 NS_667 0 9.9999999999999998e-13
CS_668 NS_668 0 9.9999999999999998e-13
RS_667 NS_667 0 7.5335118532932768e+02
RS_668 NS_668 0 7.5335118532932768e+02
GL_667 0 NS_667 NS_668 0 2.4298312011423853e-01
GL_668 0 NS_668 NS_667 0 -2.4298312011423853e-01
GS_667_12 0 NS_667 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 669/670
CS_669 NS_669 0 9.9999999999999998e-13
CS_670 NS_670 0 9.9999999999999998e-13
RS_669 NS_669 0 1.1346596293114915e+03
RS_670 NS_670 0 1.1346596293114915e+03
GL_669 0 NS_669 NS_670 0 2.4551048269503753e-01
GL_670 0 NS_670 NS_669 0 -2.4551048269503753e-01
GS_669_12 0 NS_669 NA_12 0 1.3803457954163372e+00
*
* Complex pair n. 671/672
CS_671 NS_671 0 9.9999999999999998e-13
CS_672 NS_672 0 9.9999999999999998e-13
RS_671 NS_671 0 9.3517666338196523e+02
RS_672 NS_672 0 9.3517666338196523e+02
GL_671 0 NS_671 NS_672 0 2.4538280909205379e-01
GL_672 0 NS_672 NS_671 0 -2.4538280909205379e-01
GS_671_12 0 NS_671 NA_12 0 1.3803457954163372e+00
*
******************************


.ends
*******************
* End of subcircuit
*******************
