**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 5.0000e+10 Hz
** Order: [2 2 12] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_5_C4escape_1mm_lowloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 2.3570668663388930e-01
GC_1_2 b_1 NI_1 NS_2 0 -8.4010544545778465e-04
GC_1_3 b_1 NI_1 NS_3 0 2.7374984727719345e-05
GC_1_4 b_1 NI_1 NS_4 0 -3.2161878972044406e-06
GC_1_5 b_1 NI_1 NS_5 0 -3.6342079653281378e-11
GC_1_6 b_1 NI_1 NS_6 0 -2.0793641311401382e-07
GC_1_7 b_1 NI_1 NS_7 0 -2.8744441872469061e-02
GC_1_8 b_1 NI_1 NS_8 0 1.2390377328845991e-02
GC_1_9 b_1 NI_1 NS_9 0 -1.4922286225268777e-02
GC_1_10 b_1 NI_1 NS_10 0 6.1041338156985876e-02
GC_1_11 b_1 NI_1 NS_11 0 -1.4475757340506115e-01
GC_1_12 b_1 NI_1 NS_12 0 7.1004783037250290e-03
GC_1_13 b_1 NI_1 NS_13 0 -1.6611346106465083e-01
GC_1_14 b_1 NI_1 NS_14 0 7.7902861713077798e-04
GC_1_15 b_1 NI_1 NS_15 0 -1.0081659731066468e-05
GC_1_16 b_1 NI_1 NS_16 0 4.4063523266782311e-06
GC_1_17 b_1 NI_1 NS_17 0 5.2198179209087209e-09
GC_1_18 b_1 NI_1 NS_18 0 1.7216700246894972e-07
GC_1_19 b_1 NI_1 NS_19 0 -5.0680331321099704e-02
GC_1_20 b_1 NI_1 NS_20 0 -5.0185253865991208e-02
GC_1_21 b_1 NI_1 NS_21 0 -1.8088788753475835e-02
GC_1_22 b_1 NI_1 NS_22 0 -7.4854183411212721e-02
GC_1_23 b_1 NI_1 NS_23 0 1.2153117050980806e-01
GC_1_24 b_1 NI_1 NS_24 0 -5.5012505951577565e-03
GC_1_25 b_1 NI_1 NS_25 0 4.5236596312690024e-02
GC_1_26 b_1 NI_1 NS_26 0 -2.1070046701493784e-04
GC_1_27 b_1 NI_1 NS_27 0 9.0931533075683065e-08
GC_1_28 b_1 NI_1 NS_28 0 -5.9499118600443202e-07
GC_1_29 b_1 NI_1 NS_29 0 -9.2850173516625123e-10
GC_1_30 b_1 NI_1 NS_30 0 -3.1475501608521995e-08
GC_1_31 b_1 NI_1 NS_31 0 -2.4219574873819351e-02
GC_1_32 b_1 NI_1 NS_32 0 -1.3397402435310471e-02
GC_1_33 b_1 NI_1 NS_33 0 1.4226423965900658e-02
GC_1_34 b_1 NI_1 NS_34 0 1.4703248392188239e-02
GC_1_35 b_1 NI_1 NS_35 0 -4.2182686774170808e-02
GC_1_36 b_1 NI_1 NS_36 0 5.9539176072512159e-03
GC_1_37 b_1 NI_1 NS_37 0 7.5494009814382410e-03
GC_1_38 b_1 NI_1 NS_38 0 -2.7274248920791646e-05
GC_1_39 b_1 NI_1 NS_39 0 4.2560345478428432e-06
GC_1_40 b_1 NI_1 NS_40 0 2.4799676438072629e-07
GC_1_41 b_1 NI_1 NS_41 0 7.3564845517219324e-10
GC_1_42 b_1 NI_1 NS_42 0 2.6666789328783997e-08
GC_1_43 b_1 NI_1 NS_43 0 -1.0895505433459920e-03
GC_1_44 b_1 NI_1 NS_44 0 -2.2178362519627956e-03
GC_1_45 b_1 NI_1 NS_45 0 -8.3883402209483583e-04
GC_1_46 b_1 NI_1 NS_46 0 3.4881190119098668e-03
GC_1_47 b_1 NI_1 NS_47 0 -5.7609883454454959e-03
GC_1_48 b_1 NI_1 NS_48 0 -2.7574507399449276e-03
GC_1_49 b_1 NI_1 NS_49 0 1.9940450669753878e-03
GC_1_50 b_1 NI_1 NS_50 0 -1.9462391435495011e-05
GC_1_51 b_1 NI_1 NS_51 0 -1.0455009281010323e-07
GC_1_52 b_1 NI_1 NS_52 0 -6.8160731890698158e-08
GC_1_53 b_1 NI_1 NS_53 0 9.1715214433407238e-11
GC_1_54 b_1 NI_1 NS_54 0 -2.0392073028864459e-09
GC_1_55 b_1 NI_1 NS_55 0 -1.4091128216253124e-03
GC_1_56 b_1 NI_1 NS_56 0 -2.4181058681136997e-03
GC_1_57 b_1 NI_1 NS_57 0 -4.2763972822347941e-04
GC_1_58 b_1 NI_1 NS_58 0 9.4093353859239629e-04
GC_1_59 b_1 NI_1 NS_59 0 -1.9912210582245940e-03
GC_1_60 b_1 NI_1 NS_60 0 1.7387157438808005e-03
GC_1_61 b_1 NI_1 NS_61 0 1.1232215200473128e-02
GC_1_62 b_1 NI_1 NS_62 0 -3.6178680468245924e-05
GC_1_63 b_1 NI_1 NS_63 0 3.6314268619149565e-06
GC_1_64 b_1 NI_1 NS_64 0 4.0783744767332475e-08
GC_1_65 b_1 NI_1 NS_65 0 -1.2220708203606243e-10
GC_1_66 b_1 NI_1 NS_66 0 2.9772099887489882e-09
GC_1_67 b_1 NI_1 NS_67 0 -2.2240758283006180e-03
GC_1_68 b_1 NI_1 NS_68 0 -4.2734794317932792e-03
GC_1_69 b_1 NI_1 NS_69 0 -2.3598799437846039e-03
GC_1_70 b_1 NI_1 NS_70 0 1.1521787502172056e-02
GC_1_71 b_1 NI_1 NS_71 0 -5.8123245305420155e-03
GC_1_72 b_1 NI_1 NS_72 0 -4.7340954847290041e-03
GC_1_73 b_1 NI_1 NS_73 0 5.0793347024182508e-03
GC_1_74 b_1 NI_1 NS_74 0 -1.8527002064135352e-05
GC_1_75 b_1 NI_1 NS_75 0 7.3020106218857066e-07
GC_1_76 b_1 NI_1 NS_76 0 -1.2333468738861062e-08
GC_1_77 b_1 NI_1 NS_77 0 1.3409497951777571e-10
GC_1_78 b_1 NI_1 NS_78 0 9.6871385307572226e-10
GC_1_79 b_1 NI_1 NS_79 0 9.0804996991243766e-04
GC_1_80 b_1 NI_1 NS_80 0 -1.9384015433813687e-03
GC_1_81 b_1 NI_1 NS_81 0 -4.6724832406139167e-03
GC_1_82 b_1 NI_1 NS_82 0 3.6650264593364934e-04
GC_1_83 b_1 NI_1 NS_83 0 -2.4149410524096121e-03
GC_1_84 b_1 NI_1 NS_84 0 3.0592314905037170e-03
GC_1_85 b_1 NI_1 NS_85 0 4.2229117175287762e-03
GC_1_86 b_1 NI_1 NS_86 0 -1.0991487995477852e-05
GC_1_87 b_1 NI_1 NS_87 0 9.2608130318116273e-07
GC_1_88 b_1 NI_1 NS_88 0 -2.5038099377662873e-09
GC_1_89 b_1 NI_1 NS_89 0 -1.4961375483256356e-10
GC_1_90 b_1 NI_1 NS_90 0 -4.2561761425112620e-10
GC_1_91 b_1 NI_1 NS_91 0 -3.5777259588668360e-04
GC_1_92 b_1 NI_1 NS_92 0 -1.3121073042401041e-03
GC_1_93 b_1 NI_1 NS_93 0 -1.0810765362368384e-03
GC_1_94 b_1 NI_1 NS_94 0 2.8527419811876483e-03
GC_1_95 b_1 NI_1 NS_95 0 -2.6788953815839074e-03
GC_1_96 b_1 NI_1 NS_96 0 -1.6454226974031260e-03
GC_1_97 b_1 NI_1 NS_97 0 -2.1459727371715077e-04
GC_1_98 b_1 NI_1 NS_98 0 -2.2224597112709023e-06
GC_1_99 b_1 NI_1 NS_99 0 4.5685942728962303e-08
GC_1_100 b_1 NI_1 NS_100 0 -1.0948939631836215e-10
GC_1_101 b_1 NI_1 NS_101 0 6.0712633900744335e-11
GC_1_102 b_1 NI_1 NS_102 0 4.8266786419268324e-11
GC_1_103 b_1 NI_1 NS_103 0 4.0681431252768290e-04
GC_1_104 b_1 NI_1 NS_104 0 -3.9665454064615916e-04
GC_1_105 b_1 NI_1 NS_105 0 -9.8081005320829837e-04
GC_1_106 b_1 NI_1 NS_106 0 -2.1225315491809788e-04
GC_1_107 b_1 NI_1 NS_107 0 4.2995262367454863e-04
GC_1_108 b_1 NI_1 NS_108 0 7.9393648435952370e-04
GC_1_109 b_1 NI_1 NS_109 0 4.8857469954766337e-04
GC_1_110 b_1 NI_1 NS_110 0 -2.9269411706606577e-06
GC_1_111 b_1 NI_1 NS_111 0 2.7250880793919761e-07
GC_1_112 b_1 NI_1 NS_112 0 -2.9640707871932108e-09
GC_1_113 b_1 NI_1 NS_113 0 -6.3831790750589672e-11
GC_1_114 b_1 NI_1 NS_114 0 4.9128944011563055e-11
GC_1_115 b_1 NI_1 NS_115 0 5.1373569525717754e-04
GC_1_116 b_1 NI_1 NS_116 0 -1.4982876484090241e-04
GC_1_117 b_1 NI_1 NS_117 0 -1.7726119573908977e-04
GC_1_118 b_1 NI_1 NS_118 0 -1.0127027008045551e-03
GC_1_119 b_1 NI_1 NS_119 0 -1.2278958845585734e-03
GC_1_120 b_1 NI_1 NS_120 0 -1.1792200207786840e-03
GC_1_121 b_1 NI_1 NS_121 0 -2.1577210029994276e-03
GC_1_122 b_1 NI_1 NS_122 0 3.0993750460521559e-06
GC_1_123 b_1 NI_1 NS_123 0 -1.6353131701991469e-07
GC_1_124 b_1 NI_1 NS_124 0 2.6448825414085440e-09
GC_1_125 b_1 NI_1 NS_125 0 2.6359893768848937e-11
GC_1_126 b_1 NI_1 NS_126 0 1.1477633726101760e-11
GC_1_127 b_1 NI_1 NS_127 0 2.0971550901842731e-04
GC_1_128 b_1 NI_1 NS_128 0 -2.8336000025675490e-06
GC_1_129 b_1 NI_1 NS_129 0 1.7091525342660067e-04
GC_1_130 b_1 NI_1 NS_130 0 -3.1346924350710140e-04
GC_1_131 b_1 NI_1 NS_131 0 1.5860769723682450e-03
GC_1_132 b_1 NI_1 NS_132 0 2.6011044260328305e-04
GC_1_133 b_1 NI_1 NS_133 0 4.2805970620410320e-05
GC_1_134 b_1 NI_1 NS_134 0 -7.1924074158393002e-07
GC_1_135 b_1 NI_1 NS_135 0 7.4135880506759587e-08
GC_1_136 b_1 NI_1 NS_136 0 -2.2966872381477048e-09
GC_1_137 b_1 NI_1 NS_137 0 -2.5681030698796296e-11
GC_1_138 b_1 NI_1 NS_138 0 -3.8702609047179875e-11
GC_1_139 b_1 NI_1 NS_139 0 2.8894597880845289e-04
GC_1_140 b_1 NI_1 NS_140 0 -5.4017262361909358e-06
GC_1_141 b_1 NI_1 NS_141 0 -2.3718108638547864e-05
GC_1_142 b_1 NI_1 NS_142 0 -6.8477759459401662e-04
GC_1_143 b_1 NI_1 NS_143 0 -5.2270867254624101e-04
GC_1_144 b_1 NI_1 NS_144 0 -5.5975475294921338e-04
GD_1_1 b_1 NI_1 NA_1 0 -4.9038961964207199e-02
GD_1_2 b_1 NI_1 NA_2 0 1.3127130336541257e-01
GD_1_3 b_1 NI_1 NA_3 0 5.1203296378591313e-02
GD_1_4 b_1 NI_1 NA_4 0 8.1621036869574773e-05
GD_1_5 b_1 NI_1 NA_5 0 6.1769019055698390e-03
GD_1_6 b_1 NI_1 NA_6 0 -3.4042808120793376e-04
GD_1_7 b_1 NI_1 NA_7 0 1.8866867543062143e-03
GD_1_8 b_1 NI_1 NA_8 0 1.3928245167370127e-06
GD_1_9 b_1 NI_1 NA_9 0 4.3455189490313736e-04
GD_1_10 b_1 NI_1 NA_10 0 3.6756584344559032e-04
GD_1_11 b_1 NI_1 NA_11 0 1.7347950858974674e-04
GD_1_12 b_1 NI_1 NA_12 0 1.9112395209383893e-04
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 -1.6608623964194033e-01
GC_2_2 b_2 NI_2 NS_2 0 7.7890708372751918e-04
GC_2_3 b_2 NI_2 NS_3 0 -1.0072864343609636e-05
GC_2_4 b_2 NI_2 NS_4 0 4.4062190384374240e-06
GC_2_5 b_2 NI_2 NS_5 0 5.2191421142557424e-09
GC_2_6 b_2 NI_2 NS_6 0 1.7217944742127099e-07
GC_2_7 b_2 NI_2 NS_7 0 -5.0685203973367468e-02
GC_2_8 b_2 NI_2 NS_8 0 -5.0184467201051852e-02
GC_2_9 b_2 NI_2 NS_9 0 -1.8090295009315097e-02
GC_2_10 b_2 NI_2 NS_10 0 -7.4849279883038258e-02
GC_2_11 b_2 NI_2 NS_11 0 1.2151243066283066e-01
GC_2_12 b_2 NI_2 NS_12 0 -5.5027614042469156e-03
GC_2_13 b_2 NI_2 NS_13 0 2.3570668663388908e-01
GC_2_14 b_2 NI_2 NS_14 0 -8.4010544545778400e-04
GC_2_15 b_2 NI_2 NS_15 0 2.7374984727719318e-05
GC_2_16 b_2 NI_2 NS_16 0 -3.2161878972044406e-06
GC_2_17 b_2 NI_2 NS_17 0 -3.6342079653280195e-11
GC_2_18 b_2 NI_2 NS_18 0 -2.0793641311401382e-07
GC_2_19 b_2 NI_2 NS_19 0 -2.8744441872469041e-02
GC_2_20 b_2 NI_2 NS_20 0 1.2390377328846000e-02
GC_2_21 b_2 NI_2 NS_21 0 -1.4922286225268745e-02
GC_2_22 b_2 NI_2 NS_22 0 6.1041338156985848e-02
GC_2_23 b_2 NI_2 NS_23 0 -1.4475757340506104e-01
GC_2_24 b_2 NI_2 NS_24 0 7.1004783037250316e-03
GC_2_25 b_2 NI_2 NS_25 0 7.5502213177796361e-03
GC_2_26 b_2 NI_2 NS_26 0 -2.7274646182327268e-05
GC_2_27 b_2 NI_2 NS_27 0 4.2562733409240906e-06
GC_2_28 b_2 NI_2 NS_28 0 2.4799800012840749e-07
GC_2_29 b_2 NI_2 NS_29 0 7.3566439729811976e-10
GC_2_30 b_2 NI_2 NS_30 0 2.6666996797230032e-08
GC_2_31 b_2 NI_2 NS_31 0 -1.0908140553623344e-03
GC_2_32 b_2 NI_2 NS_32 0 -2.2177922953377084e-03
GC_2_33 b_2 NI_2 NS_33 0 -8.3820605107892232e-04
GC_2_34 b_2 NI_2 NS_34 0 3.4882218294716091e-03
GC_2_35 b_2 NI_2 NS_35 0 -5.7618594233832055e-03
GC_2_36 b_2 NI_2 NS_36 0 -2.7577440833783814e-03
GC_2_37 b_2 NI_2 NS_37 0 4.5219151572628152e-02
GC_2_38 b_2 NI_2 NS_38 0 -2.1057586660610023e-04
GC_2_39 b_2 NI_2 NS_39 0 7.7884043058683377e-08
GC_2_40 b_2 NI_2 NS_40 0 -5.9496941217256012e-07
GC_2_41 b_2 NI_2 NS_41 0 -9.2824700639792962e-10
GC_2_42 b_2 NI_2 NS_42 0 -3.1476537919672348e-08
GC_2_43 b_2 NI_2 NS_43 0 -2.4219196566716228e-02
GC_2_44 b_2 NI_2 NS_44 0 -1.3397006587585499e-02
GC_2_45 b_2 NI_2 NS_45 0 1.4228525743463867e-02
GC_2_46 b_2 NI_2 NS_46 0 1.4700417927940624e-02
GC_2_47 b_2 NI_2 NS_47 0 -4.2169601446526081e-02
GC_2_48 b_2 NI_2 NS_48 0 5.9572256931884580e-03
GC_2_49 b_2 NI_2 NS_49 0 1.1240410865458966e-02
GC_2_50 b_2 NI_2 NS_50 0 -3.6204409215825214e-05
GC_2_51 b_2 NI_2 NS_51 0 3.6329437451189333e-06
GC_2_52 b_2 NI_2 NS_52 0 4.0773193251769918e-08
GC_2_53 b_2 NI_2 NS_53 0 -1.2221732377706014e-10
GC_2_54 b_2 NI_2 NS_54 0 2.9776677409534936e-09
GC_2_55 b_2 NI_2 NS_55 0 -2.2253617755250152e-03
GC_2_56 b_2 NI_2 NS_56 0 -4.2733161579852205e-03
GC_2_57 b_2 NI_2 NS_57 0 -2.3606294851509172e-03
GC_2_58 b_2 NI_2 NS_58 0 1.1523556896708810e-02
GC_2_59 b_2 NI_2 NS_59 0 -5.8176620945913950e-03
GC_2_60 b_2 NI_2 NS_60 0 -4.7341058509362205e-03
GC_2_61 b_2 NI_2 NS_61 0 1.8898177479772140e-03
GC_2_62 b_2 NI_2 NS_62 0 -1.9085620350725712e-05
GC_2_63 b_2 NI_2 NS_63 0 -1.3316160116580309e-07
GC_2_64 b_2 NI_2 NS_64 0 -6.8073536308518638e-08
GC_2_65 b_2 NI_2 NS_65 0 9.2131101705471007e-11
GC_2_66 b_2 NI_2 NS_66 0 -2.0425137780993355e-09
GC_2_67 b_2 NI_2 NS_67 0 -1.3991083666175478e-03
GC_2_68 b_2 NI_2 NS_68 0 -2.4217865717782762e-03
GC_2_69 b_2 NI_2 NS_69 0 -4.1843602527255348e-04
GC_2_70 b_2 NI_2 NS_70 0 9.1462938177173394e-04
GC_2_71 b_2 NI_2 NS_71 0 -1.9249489511344302e-03
GC_2_72 b_2 NI_2 NS_72 0 1.7404125697702830e-03
GC_2_73 b_2 NI_2 NS_73 0 4.2309798861081627e-03
GC_2_74 b_2 NI_2 NS_74 0 -1.1007814111019868e-05
GC_2_75 b_2 NI_2 NS_75 0 9.2772587899198388e-07
GC_2_76 b_2 NI_2 NS_76 0 -2.5046969741600412e-09
GC_2_77 b_2 NI_2 NS_77 0 -1.4960896144930879e-10
GC_2_78 b_2 NI_2 NS_78 0 -4.2477304474345856e-10
GC_2_79 b_2 NI_2 NS_79 0 -3.6268377919282239e-04
GC_2_80 b_2 NI_2 NS_80 0 -1.3120923075894571e-03
GC_2_81 b_2 NI_2 NS_81 0 -1.0797800003135988e-03
GC_2_82 b_2 NI_2 NS_82 0 2.8544950052259706e-03
GC_2_83 b_2 NI_2 NS_83 0 -2.6850997141922594e-03
GC_2_84 b_2 NI_2 NS_84 0 -1.6462129944013646e-03
GC_2_85 b_2 NI_2 NS_85 0 5.0774235533640995e-03
GC_2_86 b_2 NI_2 NS_86 0 -1.8520284736360316e-05
GC_2_87 b_2 NI_2 NS_87 0 7.2948407184465606e-07
GC_2_88 b_2 NI_2 NS_88 0 -1.2332554169245561e-08
GC_2_89 b_2 NI_2 NS_89 0 1.3410380654892966e-10
GC_2_90 b_2 NI_2 NS_90 0 9.6867128364204112e-10
GC_2_91 b_2 NI_2 NS_91 0 9.0821366128556748e-04
GC_2_92 b_2 NI_2 NS_92 0 -1.9384486570403845e-03
GC_2_93 b_2 NI_2 NS_93 0 -4.6722913951591548e-03
GC_2_94 b_2 NI_2 NS_94 0 3.6602325269617425e-04
GC_2_95 b_2 NI_2 NS_95 0 -2.4137135025500732e-03
GC_2_96 b_2 NI_2 NS_96 0 3.0592687143752646e-03
GC_2_97 b_2 NI_2 NS_97 0 4.8886184048031018e-04
GC_2_98 b_2 NI_2 NS_98 0 -2.9276272509574688e-06
GC_2_99 b_2 NI_2 NS_99 0 2.7255353955707310e-07
GC_2_100 b_2 NI_2 NS_100 0 -2.9640988286863260e-09
GC_2_101 b_2 NI_2 NS_101 0 -6.3831889412397356e-11
GC_2_102 b_2 NI_2 NS_102 0 4.9149286004319241e-11
GC_2_103 b_2 NI_2 NS_103 0 5.1365524859266546e-04
GC_2_104 b_2 NI_2 NS_104 0 -1.4980104250861699e-04
GC_2_105 b_2 NI_2 NS_105 0 -1.7724777100441218e-04
GC_2_106 b_2 NI_2 NS_106 0 -1.0126566845846420e-03
GC_2_107 b_2 NI_2 NS_107 0 -1.2280970289211173e-03
GC_2_108 b_2 NI_2 NS_108 0 -1.1792311158617167e-03
GC_2_109 b_2 NI_2 NS_109 0 -2.1052848236954145e-04
GC_2_110 b_2 NI_2 NS_110 0 -2.2379586722491984e-06
GC_2_111 b_2 NI_2 NS_111 0 4.5991303339166450e-08
GC_2_112 b_2 NI_2 NS_112 0 -1.2154974888510499e-10
GC_2_113 b_2 NI_2 NS_113 0 6.0706441484927148e-11
GC_2_114 b_2 NI_2 NS_114 0 4.8867575781271705e-11
GC_2_115 b_2 NI_2 NS_115 0 4.0508612046811289e-04
GC_2_116 b_2 NI_2 NS_116 0 -3.9700991042814122e-04
GC_2_117 b_2 NI_2 NS_117 0 -9.8073459376479388e-04
GC_2_118 b_2 NI_2 NS_118 0 -2.0966682644267879e-04
GC_2_119 b_2 NI_2 NS_119 0 4.2797076888303944e-04
GC_2_120 b_2 NI_2 NS_120 0 7.9429805014927756e-04
GC_2_121 b_2 NI_2 NS_121 0 4.8622050608137950e-05
GC_2_122 b_2 NI_2 NS_122 0 -7.3649343052453844e-07
GC_2_123 b_2 NI_2 NS_123 0 7.5254857401842110e-08
GC_2_124 b_2 NI_2 NS_124 0 -2.3063069853452410e-09
GC_2_125 b_2 NI_2 NS_125 0 -2.5694409591291924e-11
GC_2_126 b_2 NI_2 NS_126 0 -3.8290943258831747e-11
GC_2_127 b_2 NI_2 NS_127 0 2.8807983957665966e-04
GC_2_128 b_2 NI_2 NS_128 0 -5.9053451549561750e-06
GC_2_129 b_2 NI_2 NS_129 0 -2.4850639691884564e-05
GC_2_130 b_2 NI_2 NS_130 0 -6.8327333054448618e-04
GC_2_131 b_2 NI_2 NS_131 0 -5.2640450789824447e-04
GC_2_132 b_2 NI_2 NS_132 0 -5.5958812640004069e-04
GC_2_133 b_2 NI_2 NS_133 0 -2.1577211853650081e-03
GC_2_134 b_2 NI_2 NS_134 0 3.0993760920596358e-06
GC_2_135 b_2 NI_2 NS_135 0 -1.6353137276362475e-07
GC_2_136 b_2 NI_2 NS_136 0 2.6448827222114630e-09
GC_2_137 b_2 NI_2 NS_137 0 2.6359893148453891e-11
GC_2_138 b_2 NI_2 NS_138 0 1.1477656455424175e-11
GC_2_139 b_2 NI_2 NS_139 0 2.0971551819487229e-04
GC_2_140 b_2 NI_2 NS_140 0 -2.8336009838994721e-06
GC_2_141 b_2 NI_2 NS_141 0 1.7091529086114084e-04
GC_2_142 b_2 NI_2 NS_142 0 -3.1346926906069303e-04
GC_2_143 b_2 NI_2 NS_143 0 1.5860771058445022e-03
GC_2_144 b_2 NI_2 NS_144 0 2.6011047108747559e-04
GD_2_1 b_2 NI_2 NA_1 0 1.3127070861022236e-01
GD_2_2 b_2 NI_2 NA_2 0 -4.9038961964207199e-02
GD_2_3 b_2 NI_2 NA_3 0 8.3026773874449671e-05
GD_2_4 b_2 NI_2 NA_4 0 5.1203280119930090e-02
GD_2_5 b_2 NI_2 NA_5 0 -3.4091753277603725e-04
GD_2_6 b_2 NI_2 NA_6 0 6.1934623387746371e-03
GD_2_7 b_2 NI_2 NA_7 0 5.6840734381250982e-06
GD_2_8 b_2 NI_2 NA_8 0 1.8869350544172465e-03
GD_2_9 b_2 NI_2 NA_9 0 3.6757421084058258e-04
GD_2_10 b_2 NI_2 NA_10 0 4.3422080676758023e-04
GD_2_11 b_2 NI_2 NA_11 0 1.9132631673239979e-04
GD_2_12 b_2 NI_2 NA_12 0 1.7347945530799661e-04
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 4.5219151572654930e-02
GC_3_2 b_3 NI_3 NS_2 0 -2.1057586660623931e-04
GC_3_3 b_3 NI_3 NS_3 0 7.7884043066978265e-08
GC_3_4 b_3 NI_3 NS_4 0 -5.9496941217264630e-07
GC_3_5 b_3 NI_3 NS_5 0 -9.2824700639807727e-10
GC_3_6 b_3 NI_3 NS_6 0 -3.1476537919670455e-08
GC_3_7 b_3 NI_3 NS_7 0 -2.4219196566718341e-02
GC_3_8 b_3 NI_3 NS_8 0 -1.3397006587586866e-02
GC_3_9 b_3 NI_3 NS_9 0 1.4228525743458934e-02
GC_3_10 b_3 NI_3 NS_10 0 1.4700417927944825e-02
GC_3_11 b_3 NI_3 NS_11 0 -4.2169601446544698e-02
GC_3_12 b_3 NI_3 NS_12 0 5.9572256931867580e-03
GC_3_13 b_3 NI_3 NS_13 0 7.5494009814375601e-03
GC_3_14 b_3 NI_3 NS_14 0 -2.7274248920788072e-05
GC_3_15 b_3 NI_3 NS_15 0 4.2560345478426229e-06
GC_3_16 b_3 NI_3 NS_16 0 2.4799676438072877e-07
GC_3_17 b_3 NI_3 NS_17 0 7.3564845517220037e-10
GC_3_18 b_3 NI_3 NS_18 0 2.6666789328783904e-08
GC_3_19 b_3 NI_3 NS_19 0 -1.0895505433459378e-03
GC_3_20 b_3 NI_3 NS_20 0 -2.2178362519627601e-03
GC_3_21 b_3 NI_3 NS_21 0 -8.3883402209471007e-04
GC_3_22 b_3 NI_3 NS_22 0 3.4881190119097597e-03
GC_3_23 b_3 NI_3 NS_23 0 -5.7609883454450206e-03
GC_3_24 b_3 NI_3 NS_24 0 -2.7574507399448847e-03
GC_3_25 b_3 NI_3 NS_25 0 2.2400105485780514e-01
GC_3_26 b_3 NI_3 NS_26 0 -8.4675553269946227e-04
GC_3_27 b_3 NI_3 NS_27 0 3.0352474013254748e-05
GC_3_28 b_3 NI_3 NS_28 0 -3.3545498139811098e-06
GC_3_29 b_3 NI_3 NS_29 0 -7.7377662634893383e-10
GC_3_30 b_3 NI_3 NS_30 0 -2.0977090495226983e-07
GC_3_31 b_3 NI_3 NS_31 0 -2.4709039419403236e-02
GC_3_32 b_3 NI_3 NS_32 0 1.1897477639964151e-02
GC_3_33 b_3 NI_3 NS_33 0 -1.7546761669663572e-02
GC_3_34 b_3 NI_3 NS_34 0 5.6447029253653705e-02
GC_3_35 b_3 NI_3 NS_35 0 -1.3690354412518746e-01
GC_3_36 b_3 NI_3 NS_36 0 5.8883036864623628e-03
GC_3_37 b_3 NI_3 NS_37 0 -1.6867780301683724e-01
GC_3_38 b_3 NI_3 NS_38 0 8.1246322261204341e-04
GC_3_39 b_3 NI_3 NS_39 0 -1.1179390577396567e-05
GC_3_40 b_3 NI_3 NS_40 0 4.5242887577049176e-06
GC_3_41 b_3 NI_3 NS_41 0 5.7758219077500001e-09
GC_3_42 b_3 NI_3 NS_42 0 1.7340084729978262e-07
GC_3_43 b_3 NI_3 NS_43 0 -5.1296415736924512e-02
GC_3_44 b_3 NI_3 NS_44 0 -5.2321760270435176e-02
GC_3_45 b_3 NI_3 NS_45 0 -1.8162016821413079e-02
GC_3_46 b_3 NI_3 NS_46 0 -6.9460381710532496e-02
GC_3_47 b_3 NI_3 NS_47 0 1.2462992102311668e-01
GC_3_48 b_3 NI_3 NS_48 0 -7.4284013215734843e-03
GC_3_49 b_3 NI_3 NS_49 0 4.1960218127016009e-02
GC_3_50 b_3 NI_3 NS_50 0 -1.7447852091881613e-04
GC_3_51 b_3 NI_3 NS_51 0 5.8276866677410436e-07
GC_3_52 b_3 NI_3 NS_52 0 -5.1406387598215356e-07
GC_3_53 b_3 NI_3 NS_53 0 -7.6687074069403291e-10
GC_3_54 b_3 NI_3 NS_54 0 -3.2399426650528637e-08
GC_3_55 b_3 NI_3 NS_55 0 -1.5013437542708466e-02
GC_3_56 b_3 NI_3 NS_56 0 -9.2415775847938374e-03
GC_3_57 b_3 NI_3 NS_57 0 3.6749590497664759e-03
GC_3_58 b_3 NI_3 NS_58 0 1.1740794560460278e-02
GC_3_59 b_3 NI_3 NS_59 0 -3.3755311019172937e-02
GC_3_60 b_3 NI_3 NS_60 0 6.8939494554820444e-03
GC_3_61 b_3 NI_3 NS_61 0 -3.8427833840465218e-05
GC_3_62 b_3 NI_3 NS_62 0 8.7915602743908825e-07
GC_3_63 b_3 NI_3 NS_63 0 3.4293646431783969e-06
GC_3_64 b_3 NI_3 NS_64 0 2.8834921354275517e-07
GC_3_65 b_3 NI_3 NS_65 0 6.8381255791821818e-10
GC_3_66 b_3 NI_3 NS_66 0 2.9367357115525777e-08
GC_3_67 b_3 NI_3 NS_67 0 1.8799404109772437e-04
GC_3_68 b_3 NI_3 NS_68 0 -2.3622944715187980e-03
GC_3_69 b_3 NI_3 NS_69 0 -7.4633007088286850e-04
GC_3_70 b_3 NI_3 NS_70 0 1.3586658879689961e-03
GC_3_71 b_3 NI_3 NS_71 0 -9.8950220351403241e-04
GC_3_72 b_3 NI_3 NS_72 0 -2.9418881994748842e-03
GC_3_73 b_3 NI_3 NS_73 0 1.2344693231432387e-03
GC_3_74 b_3 NI_3 NS_74 0 -1.9200283107505086e-05
GC_3_75 b_3 NI_3 NS_75 0 -1.6566663336701651e-07
GC_3_76 b_3 NI_3 NS_76 0 -7.2745805088193404e-08
GC_3_77 b_3 NI_3 NS_77 0 8.4510116726162204e-11
GC_3_78 b_3 NI_3 NS_78 0 -2.2770251841955457e-09
GC_3_79 b_3 NI_3 NS_79 0 -1.3091991431276278e-03
GC_3_80 b_3 NI_3 NS_80 0 -2.3678855533673048e-03
GC_3_81 b_3 NI_3 NS_81 0 -3.5156966654086963e-04
GC_3_82 b_3 NI_3 NS_82 0 7.8836348668976730e-04
GC_3_83 b_3 NI_3 NS_83 0 -1.4416385043292594e-03
GC_3_84 b_3 NI_3 NS_84 0 1.7754268146023509e-03
GC_3_85 b_3 NI_3 NS_85 0 1.0864869893323369e-02
GC_3_86 b_3 NI_3 NS_86 0 -3.5600313658916289e-05
GC_3_87 b_3 NI_3 NS_87 0 3.6569520974268640e-06
GC_3_88 b_3 NI_3 NS_88 0 4.5406804423305742e-08
GC_3_89 b_3 NI_3 NS_89 0 -1.1479621821222492e-10
GC_3_90 b_3 NI_3 NS_90 0 3.2124786200041588e-09
GC_3_91 b_3 NI_3 NS_91 0 -1.8532606679503958e-03
GC_3_92 b_3 NI_3 NS_92 0 -4.1629141639127889e-03
GC_3_93 b_3 NI_3 NS_93 0 -2.2907019740573613e-03
GC_3_94 b_3 NI_3 NS_94 0 1.0457048295577830e-02
GC_3_95 b_3 NI_3 NS_95 0 -6.1522854209501952e-03
GC_3_96 b_3 NI_3 NS_96 0 -5.2206586038885394e-03
GC_3_97 b_3 NI_3 NS_97 0 1.3427743835554243e-03
GC_3_98 b_3 NI_3 NS_98 0 -9.1430271645803999e-06
GC_3_99 b_3 NI_3 NS_99 0 2.1359225935005602e-07
GC_3_100 b_3 NI_3 NS_100 0 -1.3119145181212020e-08
GC_3_101 b_3 NI_3 NS_101 0 1.1305781924862017e-10
GC_3_102 b_3 NI_3 NS_102 0 -1.8759296753003879e-10
GC_3_103 b_3 NI_3 NS_103 0 6.6878987263333022e-04
GC_3_104 b_3 NI_3 NS_104 0 -1.1220537732613901e-03
GC_3_105 b_3 NI_3 NS_105 0 -2.6054955647411399e-03
GC_3_106 b_3 NI_3 NS_106 0 3.9275190003531151e-05
GC_3_107 b_3 NI_3 NS_107 0 -1.5513279108814919e-04
GC_3_108 b_3 NI_3 NS_108 0 2.0670225004262087e-03
GC_3_109 b_3 NI_3 NS_109 0 2.3309835117911121e-03
GC_3_110 b_3 NI_3 NS_110 0 -6.0826371747049156e-06
GC_3_111 b_3 NI_3 NS_111 0 6.8137038605141341e-07
GC_3_112 b_3 NI_3 NS_112 0 4.6378329350682919e-09
GC_3_113 b_3 NI_3 NS_113 0 -1.2227884430301900e-10
GC_3_114 b_3 NI_3 NS_114 0 4.8737609485881588e-10
GC_3_115 b_3 NI_3 NS_115 0 8.0147215419040567e-06
GC_3_116 b_3 NI_3 NS_116 0 -8.0132596263998311e-04
GC_3_117 b_3 NI_3 NS_117 0 -6.2479285238258887e-04
GC_3_118 b_3 NI_3 NS_118 0 1.1738291695825636e-03
GC_3_119 b_3 NI_3 NS_119 0 -1.8495675702562588e-03
GC_3_120 b_3 NI_3 NS_120 0 -1.4232095103738447e-03
GC_3_121 b_3 NI_3 NS_121 0 -2.1049773460758388e-04
GC_3_122 b_3 NI_3 NS_122 0 -2.2380207134908103e-06
GC_3_123 b_3 NI_3 NS_123 0 4.5996143605990624e-08
GC_3_124 b_3 NI_3 NS_124 0 -1.2161408969525485e-10
GC_3_125 b_3 NI_3 NS_125 0 6.0706361631602354e-11
GC_3_126 b_3 NI_3 NS_126 0 4.8871300124999698e-11
GC_3_127 b_3 NI_3 NS_127 0 4.0508114612046984e-04
GC_3_128 b_3 NI_3 NS_128 0 -3.9700694111525684e-04
GC_3_129 b_3 NI_3 NS_129 0 -9.8073584786316764e-04
GC_3_130 b_3 NI_3 NS_130 0 -2.0965712540449975e-04
GC_3_131 b_3 NI_3 NS_131 0 4.2795362311702582e-04
GC_3_132 b_3 NI_3 NS_132 0 7.9430098508268931e-04
GC_3_133 b_3 NI_3 NS_133 0 4.8857161828666225e-04
GC_3_134 b_3 NI_3 NS_134 0 -2.9269714395746898e-06
GC_3_135 b_3 NI_3 NS_135 0 2.7250927761157655e-07
GC_3_136 b_3 NI_3 NS_136 0 -2.9640647231678041e-09
GC_3_137 b_3 NI_3 NS_137 0 -6.3831825804353647e-11
GC_3_138 b_3 NI_3 NS_138 0 4.9127728082677267e-11
GC_3_139 b_3 NI_3 NS_139 0 5.1373640083183755e-04
GC_3_140 b_3 NI_3 NS_140 0 -1.4982946193365420e-04
GC_3_141 b_3 NI_3 NS_141 0 -1.7726205497256976e-04
GC_3_142 b_3 NI_3 NS_142 0 -1.0127064845121142e-03
GC_3_143 b_3 NI_3 NS_143 0 -1.2278958749630674e-03
GC_3_144 b_3 NI_3 NS_144 0 -1.1792220317923896e-03
GD_3_1 b_3 NI_3 NA_1 0 5.1203280119930090e-02
GD_3_2 b_3 NI_3 NA_2 0 8.1621036869574773e-05
GD_3_3 b_3 NI_3 NA_3 0 -5.0105576251450769e-02
GD_3_4 b_3 NI_3 NA_4 0 1.3167218838765501e-01
GD_3_5 b_3 NI_3 NA_5 0 3.0480814121245335e-02
GD_3_6 b_3 NI_3 NA_6 0 1.9047963175751633e-03
GD_3_7 b_3 NI_3 NA_7 0 6.1354669900258669e-03
GD_3_8 b_3 NI_3 NA_8 0 -1.0917433071322557e-04
GD_3_9 b_3 NI_3 NA_9 0 1.2057088590888020e-03
GD_3_10 b_3 NI_3 NA_10 0 1.9265549640022528e-04
GD_3_11 b_3 NI_3 NA_11 0 4.3421261987482102e-04
GD_3_12 b_3 NI_3 NA_12 0 3.6757071204543998e-04
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 7.5502213177791348e-03
GC_4_2 b_4 NI_4 NS_2 0 -2.7274646182324710e-05
GC_4_3 b_4 NI_4 NS_3 0 4.2562733409239356e-06
GC_4_4 b_4 NI_4 NS_4 0 2.4799800012840913e-07
GC_4_5 b_4 NI_4 NS_5 0 7.3566439729812504e-10
GC_4_6 b_4 NI_4 NS_6 0 2.6666996797229976e-08
GC_4_7 b_4 NI_4 NS_7 0 -1.0908140553622932e-03
GC_4_8 b_4 NI_4 NS_8 0 -2.2177922953376828e-03
GC_4_9 b_4 NI_4 NS_9 0 -8.3820605107882984e-04
GC_4_10 b_4 NI_4 NS_10 0 3.4882218294715272e-03
GC_4_11 b_4 NI_4 NS_11 0 -5.7618594233828594e-03
GC_4_12 b_4 NI_4 NS_12 0 -2.7577440833783519e-03
GC_4_13 b_4 NI_4 NS_13 0 4.5236596312707010e-02
GC_4_14 b_4 NI_4 NS_14 0 -2.1070046701502807e-04
GC_4_15 b_4 NI_4 NS_15 0 9.0931533081122155e-08
GC_4_16 b_4 NI_4 NS_16 0 -5.9499118600448824e-07
GC_4_17 b_4 NI_4 NS_17 0 -9.2850173516634439e-10
GC_4_18 b_4 NI_4 NS_18 0 -3.1475501608520672e-08
GC_4_19 b_4 NI_4 NS_19 0 -2.4219574873820655e-02
GC_4_20 b_4 NI_4 NS_20 0 -1.3397402435311340e-02
GC_4_21 b_4 NI_4 NS_21 0 1.4226423965897518e-02
GC_4_22 b_4 NI_4 NS_22 0 1.4703248392190851e-02
GC_4_23 b_4 NI_4 NS_23 0 -4.2182686774182666e-02
GC_4_24 b_4 NI_4 NS_24 0 5.9539176072500796e-03
GC_4_25 b_4 NI_4 NS_25 0 -1.6870756753929878e-01
GC_4_26 b_4 NI_4 NS_26 0 8.1259529273994106e-04
GC_4_27 b_4 NI_4 NS_27 0 -1.1189045452148097e-05
GC_4_28 b_4 NI_4 NS_28 0 4.5244375117713460e-06
GC_4_29 b_4 NI_4 NS_29 0 5.7765932853712857e-09
GC_4_30 b_4 NI_4 NS_30 0 1.7338694523172418e-07
GC_4_31 b_4 NI_4 NS_31 0 -5.1291394864950136e-02
GC_4_32 b_4 NI_4 NS_32 0 -5.2322489627015974e-02
GC_4_33 b_4 NI_4 NS_33 0 -1.8160001863470804e-02
GC_4_34 b_4 NI_4 NS_34 0 -6.9465921970294511e-02
GC_4_35 b_4 NI_4 NS_35 0 1.2465020281629673e-01
GC_4_36 b_4 NI_4 NS_36 0 -7.4269932529971109e-03
GC_4_37 b_4 NI_4 NS_37 0 2.2400105485780444e-01
GC_4_38 b_4 NI_4 NS_38 0 -8.4675553269945793e-04
GC_4_39 b_4 NI_4 NS_39 0 3.0352474013254446e-05
GC_4_40 b_4 NI_4 NS_40 0 -3.3545498139811047e-06
GC_4_41 b_4 NI_4 NS_41 0 -7.7377662634891998e-10
GC_4_42 b_4 NI_4 NS_42 0 -2.0977090495227007e-07
GC_4_43 b_4 NI_4 NS_43 0 -2.4709039419403184e-02
GC_4_44 b_4 NI_4 NS_44 0 1.1897477639964189e-02
GC_4_45 b_4 NI_4 NS_45 0 -1.7546761669663437e-02
GC_4_46 b_4 NI_4 NS_46 0 5.6447029253653601e-02
GC_4_47 b_4 NI_4 NS_47 0 -1.3690354412518693e-01
GC_4_48 b_4 NI_4 NS_48 0 5.8883036864624217e-03
GC_4_49 b_4 NI_4 NS_49 0 -4.6313538296786372e-05
GC_4_50 b_4 NI_4 NS_50 0 8.9285863710816954e-07
GC_4_51 b_4 NI_4 NS_51 0 3.4279736785855222e-06
GC_4_52 b_4 NI_4 NS_52 0 2.8834756814752495e-07
GC_4_53 b_4 NI_4 NS_53 0 6.8376263973803614e-10
GC_4_54 b_4 NI_4 NS_54 0 2.9366421298113370e-08
GC_4_55 b_4 NI_4 NS_55 0 1.9289161270081770e-04
GC_4_56 b_4 NI_4 NS_56 0 -2.3626302485197166e-03
GC_4_57 b_4 NI_4 NS_57 0 -7.4794277244121454e-04
GC_4_58 b_4 NI_4 NS_58 0 1.3568457708203292e-03
GC_4_59 b_4 NI_4 NS_59 0 -9.8353568198989534e-04
GC_4_60 b_4 NI_4 NS_60 0 -2.9411785379371549e-03
GC_4_61 b_4 NI_4 NS_61 0 4.1946210944911841e-02
GC_4_62 b_4 NI_4 NS_62 0 -1.7440790712237717e-04
GC_4_63 b_4 NI_4 NS_63 0 5.7870694062224707e-07
GC_4_64 b_4 NI_4 NS_64 0 -5.1402801784243172e-07
GC_4_65 b_4 NI_4 NS_65 0 -7.6679736106973107e-10
GC_4_66 b_4 NI_4 NS_66 0 -3.2399885749940067e-08
GC_4_67 b_4 NI_4 NS_67 0 -1.5011412662759240e-02
GC_4_68 b_4 NI_4 NS_68 0 -9.2416847845086803e-03
GC_4_69 b_4 NI_4 NS_69 0 3.6761996000868867e-03
GC_4_70 b_4 NI_4 NS_70 0 1.1736911457164906e-02
GC_4_71 b_4 NI_4 NS_71 0 -3.3746472994047060e-02
GC_4_72 b_4 NI_4 NS_72 0 6.8943052033932648e-03
GC_4_73 b_4 NI_4 NS_73 0 1.0862657108896334e-02
GC_4_74 b_4 NI_4 NS_74 0 -3.5594961285054492e-05
GC_4_75 b_4 NI_4 NS_75 0 3.6565786357074271e-06
GC_4_76 b_4 NI_4 NS_76 0 4.5410354544762035e-08
GC_4_77 b_4 NI_4 NS_77 0 -1.1479122905349591e-10
GC_4_78 b_4 NI_4 NS_78 0 3.2123773313228768e-09
GC_4_79 b_4 NI_4 NS_79 0 -1.8529868530461294e-03
GC_4_80 b_4 NI_4 NS_80 0 -4.1628218413725616e-03
GC_4_81 b_4 NI_4 NS_81 0 -2.2902858853000333e-03
GC_4_82 b_4 NI_4 NS_82 0 1.0456459067221419e-02
GC_4_83 b_4 NI_4 NS_83 0 -6.1509419875855984e-03
GC_4_84 b_4 NI_4 NS_84 0 -5.2208012896741212e-03
GC_4_85 b_4 NI_4 NS_85 0 1.3272923611955280e-03
GC_4_86 b_4 NI_4 NS_86 0 -1.9513537791416618e-05
GC_4_87 b_4 NI_4 NS_87 0 -1.4173732170615312e-07
GC_4_88 b_4 NI_4 NS_88 0 -7.2811867814749793e-08
GC_4_89 b_4 NI_4 NS_89 0 8.4168105259141097e-11
GC_4_90 b_4 NI_4 NS_90 0 -2.2741008081358438e-09
GC_4_91 b_4 NI_4 NS_91 0 -1.3174943893732075e-03
GC_4_92 b_4 NI_4 NS_92 0 -2.3639656911624480e-03
GC_4_93 b_4 NI_4 NS_93 0 -3.5982957995161580e-04
GC_4_94 b_4 NI_4 NS_94 0 8.1127988160130220e-04
GC_4_95 b_4 NI_4 NS_95 0 -1.5004813369986878e-03
GC_4_96 b_4 NI_4 NS_96 0 1.7745055080583805e-03
GC_4_97 b_4 NI_4 NS_97 0 2.3226481820087870e-03
GC_4_98 b_4 NI_4 NS_98 0 -6.0665490999815356e-06
GC_4_99 b_4 NI_4 NS_99 0 6.7996611247155293e-07
GC_4_100 b_4 NI_4 NS_100 0 4.6420344461670317e-09
GC_4_101 b_4 NI_4 NS_101 0 -1.2227704227296991e-10
GC_4_102 b_4 NI_4 NS_102 0 4.8672326643990640e-10
GC_4_103 b_4 NI_4 NS_103 0 1.1437261314637998e-05
GC_4_104 b_4 NI_4 NS_104 0 -8.0083496624703849e-04
GC_4_105 b_4 NI_4 NS_105 0 -6.2462121898572323e-04
GC_4_106 b_4 NI_4 NS_106 0 1.1716323368556529e-03
GC_4_107 b_4 NI_4 NS_107 0 -1.8438019473260684e-03
GC_4_108 b_4 NI_4 NS_108 0 -1.4230868201696298e-03
GC_4_109 b_4 NI_4 NS_109 0 1.3427748968819525e-03
GC_4_110 b_4 NI_4 NS_110 0 -9.1430283847191564e-06
GC_4_111 b_4 NI_4 NS_111 0 2.1359231110147520e-07
GC_4_112 b_4 NI_4 NS_112 0 -1.3119146083236503e-08
GC_4_113 b_4 NI_4 NS_113 0 1.1305781787425029e-10
GC_4_114 b_4 NI_4 NS_114 0 -1.8759295463952842e-10
GC_4_115 b_4 NI_4 NS_115 0 6.6878979204935149e-04
GC_4_116 b_4 NI_4 NS_116 0 -1.1220537134256515e-03
GC_4_117 b_4 NI_4 NS_117 0 -2.6054955707281017e-03
GC_4_118 b_4 NI_4 NS_118 0 3.9275352642242243e-05
GC_4_119 b_4 NI_4 NS_119 0 -1.5513308558024456e-04
GC_4_120 b_4 NI_4 NS_120 0 2.0670225277402642e-03
GC_4_121 b_4 NI_4 NS_121 0 4.8885680058605001e-04
GC_4_122 b_4 NI_4 NS_122 0 -2.9276499663681166e-06
GC_4_123 b_4 NI_4 NS_123 0 2.7255376274662447e-07
GC_4_124 b_4 NI_4 NS_124 0 -2.9640930480894485e-09
GC_4_125 b_4 NI_4 NS_125 0 -6.3831920742698793e-11
GC_4_126 b_4 NI_4 NS_126 0 4.9148072146145028e-11
GC_4_127 b_4 NI_4 NS_127 0 5.1365613651502013e-04
GC_4_128 b_4 NI_4 NS_128 0 -1.4980161287909922e-04
GC_4_129 b_4 NI_4 NS_129 0 -1.7724826999802724e-04
GC_4_130 b_4 NI_4 NS_130 0 -1.0126608130872046e-03
GC_4_131 b_4 NI_4 NS_131 0 -1.2280956717391244e-03
GC_4_132 b_4 NI_4 NS_132 0 -1.1792330381222972e-03
GC_4_133 b_4 NI_4 NS_133 0 -2.1456487219706749e-04
GC_4_134 b_4 NI_4 NS_134 0 -2.2225270019474541e-06
GC_4_135 b_4 NI_4 NS_135 0 4.5691122514726061e-08
GC_4_136 b_4 NI_4 NS_136 0 -1.0955584598740775e-10
GC_4_137 b_4 NI_4 NS_137 0 6.0712532389070971e-11
GC_4_138 b_4 NI_4 NS_138 0 4.8270500099370263e-11
GC_4_139 b_4 NI_4 NS_139 0 4.0680910269778295e-04
GC_4_140 b_4 NI_4 NS_140 0 -3.9665146070817650e-04
GC_4_141 b_4 NI_4 NS_141 0 -9.8081136861491599e-04
GC_4_142 b_4 NI_4 NS_142 0 -2.1224297956274208e-04
GC_4_143 b_4 NI_4 NS_143 0 4.2993451182912198e-04
GC_4_144 b_4 NI_4 NS_144 0 7.9393952040583812e-04
GD_4_1 b_4 NI_4 NA_1 0 8.3026773874449671e-05
GD_4_2 b_4 NI_4 NA_2 0 5.1203296378591313e-02
GD_4_3 b_4 NI_4 NA_3 0 1.3167311490746747e-01
GD_4_4 b_4 NI_4 NA_4 0 -5.0105576251450769e-02
GD_4_5 b_4 NI_4 NA_5 0 1.9010413155636076e-03
GD_4_6 b_4 NI_4 NA_6 0 3.0482291068286357e-02
GD_4_7 b_4 NI_4 NA_7 0 -1.0908552512925597e-04
GD_4_8 b_4 NI_4 NA_8 0 6.1194615955975414e-03
GD_4_9 b_4 NI_4 NA_9 0 1.8991362176736312e-04
GD_4_10 b_4 NI_4 NA_10 0 1.2057087294470997e-03
GD_4_11 b_4 NI_4 NA_11 0 3.6757908566745939e-04
GD_4_12 b_4 NI_4 NA_12 0 4.3454315334320230e-04
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 1.8898177479834708e-03
GC_5_2 b_5 NI_5 NS_2 0 -1.9085620350758262e-05
GC_5_3 b_5 NI_5 NS_3 0 -1.3316160116385870e-07
GC_5_4 b_5 NI_5 NS_4 0 -6.8073536308539019e-08
GC_5_5 b_5 NI_5 NS_5 0 9.2131101705440776e-11
GC_5_6 b_5 NI_5 NS_6 0 -2.0425137780989141e-09
GC_5_7 b_5 NI_5 NS_7 0 -1.3991083666180435e-03
GC_5_8 b_5 NI_5 NS_8 0 -2.4217865717785949e-03
GC_5_9 b_5 NI_5 NS_9 0 -4.1843602527370539e-04
GC_5_10 b_5 NI_5 NS_10 0 9.1462938177271883e-04
GC_5_11 b_5 NI_5 NS_11 0 -1.9249489511387813e-03
GC_5_12 b_5 NI_5 NS_12 0 1.7404125697698871e-03
GC_5_13 b_5 NI_5 NS_13 0 1.1232215200467516e-02
GC_5_14 b_5 NI_5 NS_14 0 -3.6178680468216508e-05
GC_5_15 b_5 NI_5 NS_15 0 3.6314268619131934e-06
GC_5_16 b_5 NI_5 NS_16 0 4.0783744767350858e-08
GC_5_17 b_5 NI_5 NS_17 0 -1.2220708203603570e-10
GC_5_18 b_5 NI_5 NS_18 0 2.9772099887485928e-09
GC_5_19 b_5 NI_5 NS_19 0 -2.2240758283001778e-03
GC_5_20 b_5 NI_5 NS_20 0 -4.2734794317929922e-03
GC_5_21 b_5 NI_5 NS_21 0 -2.3598799437835691e-03
GC_5_22 b_5 NI_5 NS_22 0 1.1521787502171180e-02
GC_5_23 b_5 NI_5 NS_23 0 -5.8123245305381072e-03
GC_5_24 b_5 NI_5 NS_24 0 -4.7340954847286416e-03
GC_5_25 b_5 NI_5 NS_25 0 4.1946210944949103e-02
GC_5_26 b_5 NI_5 NS_26 0 -1.7440790712257051e-04
GC_5_27 b_5 NI_5 NS_27 0 5.7870694063377720e-07
GC_5_28 b_5 NI_5 NS_28 0 -5.1402801784255221e-07
GC_5_29 b_5 NI_5 NS_29 0 -7.6679736106994076e-10
GC_5_30 b_5 NI_5 NS_30 0 -3.2399885749937480e-08
GC_5_31 b_5 NI_5 NS_31 0 -1.5011412662762189e-02
GC_5_32 b_5 NI_5 NS_32 0 -9.2416847845105832e-03
GC_5_33 b_5 NI_5 NS_33 0 3.6761996000800228e-03
GC_5_34 b_5 NI_5 NS_34 0 1.1736911457170769e-02
GC_5_35 b_5 NI_5 NS_35 0 -3.3746472994072969e-02
GC_5_36 b_5 NI_5 NS_36 0 6.8943052033909125e-03
GC_5_37 b_5 NI_5 NS_37 0 -3.8427833841871469e-05
GC_5_38 b_5 NI_5 NS_38 0 8.7915602744649090e-07
GC_5_39 b_5 NI_5 NS_39 0 3.4293646431779433e-06
GC_5_40 b_5 NI_5 NS_40 0 2.8834921354276036e-07
GC_5_41 b_5 NI_5 NS_41 0 6.8381255791823193e-10
GC_5_42 b_5 NI_5 NS_42 0 2.9367357115525621e-08
GC_5_43 b_5 NI_5 NS_43 0 1.8799404109783605e-04
GC_5_44 b_5 NI_5 NS_44 0 -2.3622944715187269e-03
GC_5_45 b_5 NI_5 NS_45 0 -7.4633007088261024e-04
GC_5_46 b_5 NI_5 NS_46 0 1.3586658879687745e-03
GC_5_47 b_5 NI_5 NS_47 0 -9.8950220351305446e-04
GC_5_48 b_5 NI_5 NS_48 0 -2.9418881994747949e-03
GC_5_49 b_5 NI_5 NS_49 0 2.2000009389390668e-01
GC_5_50 b_5 NI_5 NS_50 0 -8.4117219569839602e-04
GC_5_51 b_5 NI_5 NS_51 0 3.0177538065481025e-05
GC_5_52 b_5 NI_5 NS_52 0 -3.3623526249797337e-06
GC_5_53 b_5 NI_5 NS_53 0 -8.0226494635996835e-10
GC_5_54 b_5 NI_5 NS_54 0 -2.1007102462669761e-07
GC_5_55 b_5 NI_5 NS_55 0 -2.4188099030426638e-02
GC_5_56 b_5 NI_5 NS_56 0 1.1786350780877933e-02
GC_5_57 b_5 NI_5 NS_57 0 -1.7257681342090533e-02
GC_5_58 b_5 NI_5 NS_58 0 5.5409688512598421e-02
GC_5_59 b_5 NI_5 NS_59 0 -1.3437382346476356e-01
GC_5_60 b_5 NI_5 NS_60 0 5.8053021877571753e-03
GC_5_61 b_5 NI_5 NS_61 0 -1.7636412290295697e-01
GC_5_62 b_5 NI_5 NS_62 0 8.6547518201292458e-04
GC_5_63 b_5 NI_5 NS_63 0 -1.5390117042153797e-05
GC_5_64 b_5 NI_5 NS_64 0 4.6154846005047276e-06
GC_5_65 b_5 NI_5 NS_65 0 6.2868134723974044e-09
GC_5_66 b_5 NI_5 NS_66 0 1.6582384401838644e-07
GC_5_67 b_5 NI_5 NS_67 0 -5.0273987508574786e-02
GC_5_68 b_5 NI_5 NS_68 0 -5.1965674064694080e-02
GC_5_69 b_5 NI_5 NS_69 0 -1.6950175224523075e-02
GC_5_70 b_5 NI_5 NS_70 0 -7.2073581381944640e-02
GC_5_71 b_5 NI_5 NS_71 0 1.2915680926872447e-01
GC_5_72 b_5 NI_5 NS_72 0 -7.4441654867010215e-03
GC_5_73 b_5 NI_5 NS_73 0 4.8536552541238967e-02
GC_5_74 b_5 NI_5 NS_74 0 -2.2743854750332100e-04
GC_5_75 b_5 NI_5 NS_75 0 8.3302383914318666e-07
GC_5_76 b_5 NI_5 NS_76 0 -6.3071450988624545e-07
GC_5_77 b_5 NI_5 NS_77 0 -9.7210182641320204e-10
GC_5_78 b_5 NI_5 NS_78 0 -3.2569423280656212e-08
GC_5_79 b_5 NI_5 NS_79 0 -2.3416311478099080e-02
GC_5_80 b_5 NI_5 NS_80 0 -1.3900300372963768e-02
GC_5_81 b_5 NI_5 NS_81 0 1.1403223908453214e-02
GC_5_82 b_5 NI_5 NS_82 0 1.4942438470155767e-02
GC_5_83 b_5 NI_5 NS_83 0 -4.3469993171037571e-02
GC_5_84 b_5 NI_5 NS_84 0 7.5391534381776945e-03
GC_5_85 b_5 NI_5 NS_85 0 5.4819587052257349e-03
GC_5_86 b_5 NI_5 NS_86 0 -1.7137352684306397e-05
GC_5_87 b_5 NI_5 NS_87 0 3.9073369516379621e-06
GC_5_88 b_5 NI_5 NS_88 0 2.8019717805331460e-07
GC_5_89 b_5 NI_5 NS_89 0 7.9554769583068835e-10
GC_5_90 b_5 NI_5 NS_90 0 2.7616182962561345e-08
GC_5_91 b_5 NI_5 NS_91 0 -3.6662534007919780e-04
GC_5_92 b_5 NI_5 NS_92 0 -2.0511587923623537e-03
GC_5_93 b_5 NI_5 NS_93 0 -7.3145786443027251e-04
GC_5_94 b_5 NI_5 NS_94 0 1.4824773703910621e-03
GC_5_95 b_5 NI_5 NS_95 0 -5.1593039959526099e-03
GC_5_96 b_5 NI_5 NS_96 0 -3.0581719914394736e-03
GC_5_97 b_5 NI_5 NS_97 0 1.3273205919093396e-03
GC_5_98 b_5 NI_5 NS_98 0 -1.9513663171605448e-05
GC_5_99 b_5 NI_5 NS_99 0 -1.4172560971485596e-07
GC_5_100 b_5 NI_5 NS_100 0 -7.2812366939657940e-08
GC_5_101 b_5 NI_5 NS_101 0 8.4153281785307944e-11
GC_5_102 b_5 NI_5 NS_102 0 -2.2739453061637985e-09
GC_5_103 b_5 NI_5 NS_103 0 -1.3174988886496698e-03
GC_5_104 b_5 NI_5 NS_104 0 -2.3639640757188484e-03
GC_5_105 b_5 NI_5 NS_105 0 -3.5983148418215440e-04
GC_5_106 b_5 NI_5 NS_106 0 8.1128675830275884e-04
GC_5_107 b_5 NI_5 NS_107 0 -1.5004987608067076e-03
GC_5_108 b_5 NI_5 NS_108 0 1.7745062024234601e-03
GC_5_109 b_5 NI_5 NS_109 0 1.0864943270449887e-02
GC_5_110 b_5 NI_5 NS_110 0 -3.5600529508431843e-05
GC_5_111 b_5 NI_5 NS_111 0 3.6569563861731139e-06
GC_5_112 b_5 NI_5 NS_112 0 4.5407222612022546e-08
GC_5_113 b_5 NI_5 NS_113 0 -1.1478141557247145e-10
GC_5_114 b_5 NI_5 NS_114 0 3.2123229186354735e-09
GC_5_115 b_5 NI_5 NS_115 0 -1.8532685974524058e-03
GC_5_116 b_5 NI_5 NS_116 0 -4.1629108672277242e-03
GC_5_117 b_5 NI_5 NS_117 0 -2.2907093992697073e-03
GC_5_118 b_5 NI_5 NS_118 0 1.0457063710973519e-02
GC_5_119 b_5 NI_5 NS_119 0 -6.1523321214198203e-03
GC_5_120 b_5 NI_5 NS_120 0 -5.2206578141558149e-03
GC_5_121 b_5 NI_5 NS_121 0 5.0776152495564083e-03
GC_5_122 b_5 NI_5 NS_122 0 -1.8520847161729861e-05
GC_5_123 b_5 NI_5 NS_123 0 7.2952520166529483e-07
GC_5_124 b_5 NI_5 NS_124 0 -1.2333156060169070e-08
GC_5_125 b_5 NI_5 NS_125 0 1.3410093802497754e-10
GC_5_126 b_5 NI_5 NS_126 0 9.6871019294210781e-10
GC_5_127 b_5 NI_5 NS_127 0 9.0818992255816311e-04
GC_5_128 b_5 NI_5 NS_128 0 -1.9384358581755799e-03
GC_5_129 b_5 NI_5 NS_129 0 -4.6723063311410185e-03
GC_5_130 b_5 NI_5 NS_130 0 3.6607765509906221e-04
GC_5_131 b_5 NI_5 NS_131 0 -2.4138258019113503e-03
GC_5_132 b_5 NI_5 NS_132 0 3.0592774774284275e-03
GC_5_133 b_5 NI_5 NS_133 0 4.2228725450485626e-03
GC_5_134 b_5 NI_5 NS_134 0 -1.0991489590242371e-05
GC_5_135 b_5 NI_5 NS_135 0 9.2608169996248885e-07
GC_5_136 b_5 NI_5 NS_136 0 -2.5038170766799749e-09
GC_5_137 b_5 NI_5 NS_137 0 -1.4961183510655973e-10
GC_5_138 b_5 NI_5 NS_138 0 -4.2562873433720577e-10
GC_5_139 b_5 NI_5 NS_139 0 -3.5777178697689050e-04
GC_5_140 b_5 NI_5 NS_140 0 -1.3121060881780616e-03
GC_5_141 b_5 NI_5 NS_141 0 -1.0810728105758868e-03
GC_5_142 b_5 NI_5 NS_142 0 2.8527296137076316e-03
GC_5_143 b_5 NI_5 NS_143 0 -2.6788727572075442e-03
GC_5_144 b_5 NI_5 NS_144 0 -1.6454282606839260e-03
GD_5_1 b_5 NI_5 NA_1 0 6.1934623387746371e-03
GD_5_2 b_5 NI_5 NA_2 0 -3.4042808120793376e-04
GD_5_3 b_5 NI_5 NA_3 0 3.0482291068286357e-02
GD_5_4 b_5 NI_5 NA_4 0 1.9047963175751633e-03
GD_5_5 b_5 NI_5 NA_5 0 -4.9495926725586142e-02
GD_5_6 b_5 NI_5 NA_6 0 1.3241931555769479e-01
GD_5_7 b_5 NI_5 NA_7 0 5.0627972643333595e-02
GD_5_8 b_5 NI_5 NA_8 0 6.8938798190542390e-04
GD_5_9 b_5 NI_5 NA_9 0 6.1194575195962549e-03
GD_5_10 b_5 NI_5 NA_10 0 -1.0918537265261697e-04
GD_5_11 b_5 NI_5 NA_11 0 1.8868877227967388e-03
GD_5_12 b_5 NI_5 NA_12 0 1.4129039939162737e-06
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 1.1240410865452905e-02
GC_6_2 b_6 NI_6 NS_2 0 -3.6204409215794484e-05
GC_6_3 b_6 NI_6 NS_3 0 3.6329437451171258e-06
GC_6_4 b_6 NI_6 NS_4 0 4.0773193251788765e-08
GC_6_5 b_6 NI_6 NS_5 0 -1.2221732377703168e-10
GC_6_6 b_6 NI_6 NS_6 0 2.9776677409531403e-09
GC_6_7 b_6 NI_6 NS_7 0 -2.2253617755245234e-03
GC_6_8 b_6 NI_6 NS_8 0 -4.2733161579849117e-03
GC_6_9 b_6 NI_6 NS_9 0 -2.3606294851498013e-03
GC_6_10 b_6 NI_6 NS_10 0 1.1523556896707839e-02
GC_6_11 b_6 NI_6 NS_11 0 -5.8176620945871943e-03
GC_6_12 b_6 NI_6 NS_12 0 -4.7341058509358588e-03
GC_6_13 b_6 NI_6 NS_13 0 1.9940450669817871e-03
GC_6_14 b_6 NI_6 NS_14 0 -1.9462391435527825e-05
GC_6_15 b_6 NI_6 NS_15 0 -1.0455009280815954e-07
GC_6_16 b_6 NI_6 NS_16 0 -6.8160731890718514e-08
GC_6_17 b_6 NI_6 NS_17 0 9.1715214433376542e-11
GC_6_18 b_6 NI_6 NS_18 0 -2.0392073028860489e-09
GC_6_19 b_6 NI_6 NS_19 0 -1.4091128216258267e-03
GC_6_20 b_6 NI_6 NS_20 0 -2.4181058681140258e-03
GC_6_21 b_6 NI_6 NS_21 0 -4.2763972822465685e-04
GC_6_22 b_6 NI_6 NS_22 0 9.4093353859341750e-04
GC_6_23 b_6 NI_6 NS_23 0 -1.9912210582290341e-03
GC_6_24 b_6 NI_6 NS_24 0 1.7387157438804096e-03
GC_6_25 b_6 NI_6 NS_25 0 -4.6313538298730665e-05
GC_6_26 b_6 NI_6 NS_26 0 8.9285863711813880e-07
GC_6_27 b_6 NI_6 NS_27 0 3.4279736785849204e-06
GC_6_28 b_6 NI_6 NS_28 0 2.8834756814753173e-07
GC_6_29 b_6 NI_6 NS_29 0 6.8376263973805537e-10
GC_6_30 b_6 NI_6 NS_30 0 2.9366421298113178e-08
GC_6_31 b_6 NI_6 NS_31 0 1.9289161270097629e-04
GC_6_32 b_6 NI_6 NS_32 0 -2.3626302485196182e-03
GC_6_33 b_6 NI_6 NS_33 0 -7.4794277244085783e-04
GC_6_34 b_6 NI_6 NS_34 0 1.3568457708200152e-03
GC_6_35 b_6 NI_6 NS_35 0 -9.8353568198854854e-04
GC_6_36 b_6 NI_6 NS_36 0 -2.9411785379370383e-03
GC_6_37 b_6 NI_6 NS_37 0 4.1960218127047831e-02
GC_6_38 b_6 NI_6 NS_38 0 -1.7447852091897321e-04
GC_6_39 b_6 NI_6 NS_39 0 5.8276866678319663e-07
GC_6_40 b_6 NI_6 NS_40 0 -5.1406387598224864e-07
GC_6_41 b_6 NI_6 NS_41 0 -7.6687074069421365e-10
GC_6_42 b_6 NI_6 NS_42 0 -3.2399426650526983e-08
GC_6_43 b_6 NI_6 NS_43 0 -1.5013437542711115e-02
GC_6_44 b_6 NI_6 NS_44 0 -9.2415775847954594e-03
GC_6_45 b_6 NI_6 NS_45 0 3.6749590497606255e-03
GC_6_46 b_6 NI_6 NS_46 0 1.1740794560465525e-02
GC_6_47 b_6 NI_6 NS_47 0 -3.3755311019194899e-02
GC_6_48 b_6 NI_6 NS_48 0 6.8939494554802775e-03
GC_6_49 b_6 NI_6 NS_49 0 -1.7636209667358269e-01
GC_6_50 b_6 NI_6 NS_50 0 8.6546748574712392e-04
GC_6_51 b_6 NI_6 NS_51 0 -1.5389453476708602e-05
GC_6_52 b_6 NI_6 NS_52 0 4.6154719441345791e-06
GC_6_53 b_6 NI_6 NS_53 0 6.2867337300986555e-09
GC_6_54 b_6 NI_6 NS_54 0 1.6582502673964577e-07
GC_6_55 b_6 NI_6 NS_55 0 -5.0274107512396200e-02
GC_6_56 b_6 NI_6 NS_56 0 -5.1965750863517970e-02
GC_6_57 b_6 NI_6 NS_57 0 -1.6950620652552578e-02
GC_6_58 b_6 NI_6 NS_58 0 -7.2073025574349942e-02
GC_6_59 b_6 NI_6 NS_59 0 1.2915561439930526e-01
GC_6_60 b_6 NI_6 NS_60 0 -7.4440371012940085e-03
GC_6_61 b_6 NI_6 NS_61 0 2.2000009389389838e-01
GC_6_62 b_6 NI_6 NS_62 0 -8.4117219569817235e-04
GC_6_63 b_6 NI_6 NS_63 0 3.0177538065455302e-05
GC_6_64 b_6 NI_6 NS_64 0 -3.3623526249792250e-06
GC_6_65 b_6 NI_6 NS_65 0 -8.0226494634976870e-10
GC_6_66 b_6 NI_6 NS_66 0 -2.1007102462674936e-07
GC_6_67 b_6 NI_6 NS_67 0 -2.4188099030426152e-02
GC_6_68 b_6 NI_6 NS_68 0 1.1786350780876647e-02
GC_6_69 b_6 NI_6 NS_69 0 -1.7257681342091276e-02
GC_6_70 b_6 NI_6 NS_70 0 5.5409688512597477e-02
GC_6_71 b_6 NI_6 NS_71 0 -1.3437382346475743e-01
GC_6_72 b_6 NI_6 NS_72 0 5.8053021877602137e-03
GC_6_73 b_6 NI_6 NS_73 0 5.4843824144410729e-03
GC_6_74 b_6 NI_6 NS_74 0 -1.7139696260601074e-05
GC_6_75 b_6 NI_6 NS_75 0 3.9079478424632787e-06
GC_6_76 b_6 NI_6 NS_76 0 2.8019695410546820e-07
GC_6_77 b_6 NI_6 NS_77 0 7.9557076700303995e-10
GC_6_78 b_6 NI_6 NS_78 0 2.7616671162318015e-08
GC_6_79 b_6 NI_6 NS_79 0 -3.6911708103831063e-04
GC_6_80 b_6 NI_6 NS_80 0 -2.0512083117273637e-03
GC_6_81 b_6 NI_6 NS_81 0 -7.3054742329536936e-04
GC_6_82 b_6 NI_6 NS_82 0 1.4830214422838844e-03
GC_6_83 b_6 NI_6 NS_83 0 -5.1614094384650373e-03
GC_6_84 b_6 NI_6 NS_84 0 -3.0585858755697200e-03
GC_6_85 b_6 NI_6 NS_85 0 4.8536551962246002e-02
GC_6_86 b_6 NI_6 NS_86 0 -2.2743853783404314e-04
GC_6_87 b_6 NI_6 NS_87 0 8.3302345961160922e-07
GC_6_88 b_6 NI_6 NS_88 0 -6.3071451646566461e-07
GC_6_89 b_6 NI_6 NS_89 0 -9.7210183423082645e-10
GC_6_90 b_6 NI_6 NS_90 0 -3.2569422867599954e-08
GC_6_91 b_6 NI_6 NS_91 0 -2.3416311619223407e-02
GC_6_92 b_6 NI_6 NS_92 0 -1.3900300261699803e-02
GC_6_93 b_6 NI_6 NS_93 0 1.1403224112185866e-02
GC_6_94 b_6 NI_6 NS_94 0 1.4942438711044382e-02
GC_6_95 b_6 NI_6 NS_95 0 -4.3469992548393510e-02
GC_6_96 b_6 NI_6 NS_96 0 7.5391537497767206e-03
GC_6_97 b_6 NI_6 NS_97 0 1.0862693856980195e-02
GC_6_98 b_6 NI_6 NS_98 0 -3.5594952491940069e-05
GC_6_99 b_6 NI_6 NS_99 0 3.6565670975767611e-06
GC_6_100 b_6 NI_6 NS_100 0 4.5410903815680037e-08
GC_6_101 b_6 NI_6 NS_101 0 -1.1477636020363388e-10
GC_6_102 b_6 NI_6 NS_102 0 3.2122170325728598e-09
GC_6_103 b_6 NI_6 NS_103 0 -1.8529917409112549e-03
GC_6_104 b_6 NI_6 NS_104 0 -4.1628193438068119e-03
GC_6_105 b_6 NI_6 NS_105 0 -2.2902894265693658e-03
GC_6_106 b_6 NI_6 NS_106 0 1.0456468031387152e-02
GC_6_107 b_6 NI_6 NS_107 0 -6.1509639060060269e-03
GC_6_108 b_6 NI_6 NS_108 0 -5.2207980239416312e-03
GC_6_109 b_6 NI_6 NS_109 0 1.2344750425225665e-03
GC_6_110 b_6 NI_6 NS_110 0 -1.9200359762749084e-05
GC_6_111 b_6 NI_6 NS_111 0 -1.6565620384704142e-07
GC_6_112 b_6 NI_6 NS_112 0 -7.2746318345653761e-08
GC_6_113 b_6 NI_6 NS_113 0 8.4495288985347639e-11
GC_6_114 b_6 NI_6 NS_114 0 -2.2768686473884669e-09
GC_6_115 b_6 NI_6 NS_115 0 -1.3092006272324250e-03
GC_6_116 b_6 NI_6 NS_116 0 -2.3678852794048457e-03
GC_6_117 b_6 NI_6 NS_117 0 -3.5157008440983502e-04
GC_6_118 b_6 NI_6 NS_118 0 7.8836385719273155e-04
GC_6_119 b_6 NI_6 NS_119 0 -1.4416426295163160e-03
GC_6_120 b_6 NI_6 NS_120 0 1.7754263218758349e-03
GC_6_121 b_6 NI_6 NS_121 0 4.2309469671519620e-03
GC_6_122 b_6 NI_6 NS_122 0 -1.1007839912098661e-05
GC_6_123 b_6 NI_6 NS_123 0 9.2772769406622697e-07
GC_6_124 b_6 NI_6 NS_124 0 -2.5047091134672579e-09
GC_6_125 b_6 NI_6 NS_125 0 -1.4960708293035260e-10
GC_6_126 b_6 NI_6 NS_126 0 -4.2478288251201136e-10
GC_6_127 b_6 NI_6 NS_127 0 -3.6268360075236179e-04
GC_6_128 b_6 NI_6 NS_128 0 -1.3120905163259207e-03
GC_6_129 b_6 NI_6 NS_129 0 -1.0797766428347136e-03
GC_6_130 b_6 NI_6 NS_130 0 2.8544842384299121e-03
GC_6_131 b_6 NI_6 NS_131 0 -2.6850808468543981e-03
GC_6_132 b_6 NI_6 NS_132 0 -1.6462183999218494e-03
GC_6_133 b_6 NI_6 NS_133 0 5.0795379504729758e-03
GC_6_134 b_6 NI_6 NS_134 0 -1.8527609238793777e-05
GC_6_135 b_6 NI_6 NS_135 0 7.3024486498347187e-07
GC_6_136 b_6 NI_6 NS_136 0 -1.2334102731167366e-08
GC_6_137 b_6 NI_6 NS_137 0 1.3409208913866477e-10
GC_6_138 b_6 NI_6 NS_138 0 9.6875331338746038e-10
GC_6_139 b_6 NI_6 NS_139 0 9.0802500331060301e-04
GC_6_140 b_6 NI_6 NS_140 0 -1.9383887053155738e-03
GC_6_141 b_6 NI_6 NS_141 0 -4.6724996511191032e-03
GC_6_142 b_6 NI_6 NS_142 0 3.6655965392259871e-04
GC_6_143 b_6 NI_6 NS_143 0 -2.4150607677583904e-03
GC_6_144 b_6 NI_6 NS_144 0 3.0592401847397799e-03
GD_6_1 b_6 NI_6 NA_1 0 -3.4091753277603725e-04
GD_6_2 b_6 NI_6 NA_2 0 6.1769019055698390e-03
GD_6_3 b_6 NI_6 NA_3 0 1.9010413155636076e-03
GD_6_4 b_6 NI_6 NA_4 0 3.0480814121245335e-02
GD_6_5 b_6 NI_6 NA_5 0 1.3241906596251396e-01
GD_6_6 b_6 NI_6 NA_6 0 -4.9495926725583152e-02
GD_6_7 b_6 NI_6 NA_7 0 6.9207054480047332e-04
GD_6_8 b_6 NI_6 NA_8 0 5.0627972593922363e-02
GD_6_9 b_6 NI_6 NA_9 0 -1.0909158462998901e-04
GD_6_10 b_6 NI_6 NA_10 0 6.1354681668953012e-03
GD_6_11 b_6 NI_6 NA_11 0 5.7024688927638791e-06
GD_6_12 b_6 NI_6 NA_12 0 1.8866381493710604e-03
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 5.0774235420953349e-03
GC_7_2 b_7 NI_7 NS_2 0 -1.8520284682846519e-05
GC_7_3 b_7 NI_7 NS_3 0 7.2948406855790119e-07
GC_7_4 b_7 NI_7 NS_4 0 -1.2332554139063901e-08
GC_7_5 b_7 NI_7 NS_5 0 1.3410380658016804e-10
GC_7_6 b_7 NI_7 NS_6 0 9.6867128240810044e-10
GC_7_7 b_7 NI_7 NS_7 0 9.0821366229434410e-04
GC_7_8 b_7 NI_7 NS_8 0 -1.9384486570375560e-03
GC_7_9 b_7 NI_7 NS_9 0 -4.6722913936610658e-03
GC_7_10 b_7 NI_7 NS_10 0 3.6602325052776573e-04
GC_7_11 b_7 NI_7 NS_11 0 -2.4137134950620196e-03
GC_7_12 b_7 NI_7 NS_12 0 3.0592687147877810e-03
GC_7_13 b_7 NI_7 NS_13 0 4.2229117175261194e-03
GC_7_14 b_7 NI_7 NS_14 0 -1.0991487995464384e-05
GC_7_15 b_7 NI_7 NS_15 0 9.2608130318037170e-07
GC_7_16 b_7 NI_7 NS_16 0 -2.5038099377580639e-09
GC_7_17 b_7 NI_7 NS_17 0 -1.4961375483255348e-10
GC_7_18 b_7 NI_7 NS_18 0 -4.2561761425126976e-10
GC_7_19 b_7 NI_7 NS_19 0 -3.5777259588646790e-04
GC_7_20 b_7 NI_7 NS_20 0 -1.3121073042399688e-03
GC_7_21 b_7 NI_7 NS_21 0 -1.0810765362363494e-03
GC_7_22 b_7 NI_7 NS_22 0 2.8527419811872194e-03
GC_7_23 b_7 NI_7 NS_23 0 -2.6788953815820664e-03
GC_7_24 b_7 NI_7 NS_24 0 -1.6454226974029680e-03
GC_7_25 b_7 NI_7 NS_25 0 1.3272923548825065e-03
GC_7_26 b_7 NI_7 NS_26 0 -1.9513537742268748e-05
GC_7_27 b_7 NI_7 NS_27 0 -1.4173732668011283e-07
GC_7_28 b_7 NI_7 NS_28 0 -7.2811867607184634e-08
GC_7_29 b_7 NI_7 NS_29 0 8.4168119310904388e-11
GC_7_30 b_7 NI_7 NS_30 0 -2.2741008491701402e-09
GC_7_31 b_7 NI_7 NS_31 0 -1.3174943888856563e-03
GC_7_32 b_7 NI_7 NS_32 0 -2.3639656912217586e-03
GC_7_33 b_7 NI_7 NS_33 0 -3.5982957920942162e-04
GC_7_34 b_7 NI_7 NS_34 0 8.1127988056163341e-04
GC_7_35 b_7 NI_7 NS_35 0 -1.5004813326640215e-03
GC_7_36 b_7 NI_7 NS_36 0 1.7745055086073058e-03
GC_7_37 b_7 NI_7 NS_37 0 1.0864869893314776e-02
GC_7_38 b_7 NI_7 NS_38 0 -3.5600313658873544e-05
GC_7_39 b_7 NI_7 NS_39 0 3.6569520974243818e-06
GC_7_40 b_7 NI_7 NS_40 0 4.5406804423331716e-08
GC_7_41 b_7 NI_7 NS_41 0 -1.1479621821218453e-10
GC_7_42 b_7 NI_7 NS_42 0 3.2124786200037212e-09
GC_7_43 b_7 NI_7 NS_43 0 -1.8532606679496841e-03
GC_7_44 b_7 NI_7 NS_44 0 -4.1629141639123518e-03
GC_7_45 b_7 NI_7 NS_45 0 -2.2907019740557805e-03
GC_7_46 b_7 NI_7 NS_46 0 1.0457048295576421e-02
GC_7_47 b_7 NI_7 NS_47 0 -6.1522854209442581e-03
GC_7_48 b_7 NI_7 NS_48 0 -5.2206586038880546e-03
GC_7_49 b_7 NI_7 NS_49 0 4.8536551962305566e-02
GC_7_50 b_7 NI_7 NS_50 0 -2.2743853783433872e-04
GC_7_51 b_7 NI_7 NS_51 0 8.3302345962877668e-07
GC_7_52 b_7 NI_7 NS_52 0 -6.3071451646584354e-07
GC_7_53 b_7 NI_7 NS_53 0 -9.7210183423116105e-10
GC_7_54 b_7 NI_7 NS_54 0 -3.2569422867596731e-08
GC_7_55 b_7 NI_7 NS_55 0 -2.3416311619228334e-02
GC_7_56 b_7 NI_7 NS_56 0 -1.3900300261702841e-02
GC_7_57 b_7 NI_7 NS_57 0 1.1403224112174912e-02
GC_7_58 b_7 NI_7 NS_58 0 1.4942438711054155e-02
GC_7_59 b_7 NI_7 NS_59 0 -4.3469992548434665e-02
GC_7_60 b_7 NI_7 NS_60 0 7.5391537497733647e-03
GC_7_61 b_7 NI_7 NS_61 0 5.4819587047321584e-03
GC_7_62 b_7 NI_7 NS_62 0 -1.7137352682025479e-05
GC_7_63 b_7 NI_7 NS_63 0 3.9073369514989877e-06
GC_7_64 b_7 NI_7 NS_64 0 2.8019717805478743e-07
GC_7_65 b_7 NI_7 NS_65 0 7.9554769583424916e-10
GC_7_66 b_7 NI_7 NS_66 0 2.7616182962482806e-08
GC_7_67 b_7 NI_7 NS_67 0 -3.6662534003352654e-04
GC_7_68 b_7 NI_7 NS_68 0 -2.0511587923489494e-03
GC_7_69 b_7 NI_7 NS_69 0 -7.3145786435236705e-04
GC_7_70 b_7 NI_7 NS_70 0 1.4824773702964960e-03
GC_7_71 b_7 NI_7 NS_71 0 -5.1593039956222579e-03
GC_7_72 b_7 NI_7 NS_72 0 -3.0581719914217855e-03
GC_7_73 b_7 NI_7 NS_73 0 2.2000012094882873e-01
GC_7_74 b_7 NI_7 NS_74 0 -8.4117228611806387e-04
GC_7_75 b_7 NI_7 NS_75 0 3.0177543234324138e-05
GC_7_76 b_7 NI_7 NS_76 0 -3.3623526868368786e-06
GC_7_77 b_7 NI_7 NS_77 0 -8.0226512044408508e-10
GC_7_78 b_7 NI_7 NS_78 0 -2.1007102099711095e-07
GC_7_79 b_7 NI_7 NS_79 0 -2.4188102219297271e-02
GC_7_80 b_7 NI_7 NS_80 0 1.1786351174973177e-02
GC_7_81 b_7 NI_7 NS_81 0 -1.7257684471469113e-02
GC_7_82 b_7 NI_7 NS_82 0 5.5409695305402212e-02
GC_7_83 b_7 NI_7 NS_83 0 -1.3437384032485303e-01
GC_7_84 b_7 NI_7 NS_84 0 5.8053026351617566e-03
GC_7_85 b_7 NI_7 NS_85 0 -1.7636408134268197e-01
GC_7_86 b_7 NI_7 NS_86 0 8.6547493395085857e-04
GC_7_87 b_7 NI_7 NS_87 0 -1.5390096193926349e-05
GC_7_88 b_7 NI_7 NS_88 0 4.6154841806943552e-06
GC_7_89 b_7 NI_7 NS_89 0 6.2868109382599931e-09
GC_7_90 b_7 NI_7 NS_90 0 1.6582388483023826e-07
GC_7_91 b_7 NI_7 NS_91 0 -5.0273992194559504e-02
GC_7_92 b_7 NI_7 NS_92 0 -5.1965672154779270e-02
GC_7_93 b_7 NI_7 NS_93 0 -1.6950178423066124e-02
GC_7_94 b_7 NI_7 NS_94 0 -7.2073572147318174e-02
GC_7_95 b_7 NI_7 NS_95 0 1.2915678239637368e-01
GC_7_96 b_7 NI_7 NS_96 0 -7.4441671225573504e-03
GC_7_97 b_7 NI_7 NS_97 0 4.1946350052475614e-02
GC_7_98 b_7 NI_7 NS_98 0 -1.7440834779712671e-04
GC_7_99 b_7 NI_7 NS_99 0 5.7873283473280193e-07
GC_7_100 b_7 NI_7 NS_100 0 -5.1402838048937752e-07
GC_7_101 b_7 NI_7 NS_101 0 -7.6680262802050697e-10
GC_7_102 b_7 NI_7 NS_102 0 -3.2399854190571301e-08
GC_7_103 b_7 NI_7 NS_103 0 -1.5011431217309442e-02
GC_7_104 b_7 NI_7 NS_104 0 -9.2416782120910528e-03
GC_7_105 b_7 NI_7 NS_105 0 3.6761889300958375e-03
GC_7_106 b_7 NI_7 NS_106 0 1.1736949771054314e-02
GC_7_107 b_7 NI_7 NS_107 0 -3.3746557294655845e-02
GC_7_108 b_7 NI_7 NS_108 0 6.8943091498476182e-03
GC_7_109 b_7 NI_7 NS_109 0 -3.8369878990799497e-05
GC_7_110 b_7 NI_7 NS_110 0 8.7899445061528892e-07
GC_7_111 b_7 NI_7 NS_111 0 3.4293754233098523e-06
GC_7_112 b_7 NI_7 NS_112 0 2.8834905730743922e-07
GC_7_113 b_7 NI_7 NS_113 0 6.8381509573633570e-10
GC_7_114 b_7 NI_7 NS_114 0 2.9367357449012790e-08
GC_7_115 b_7 NI_7 NS_115 0 1.8798474525441274e-04
GC_7_116 b_7 NI_7 NS_116 0 -2.3622896214915610e-03
GC_7_117 b_7 NI_7 NS_117 0 -7.4633196007450875e-04
GC_7_118 b_7 NI_7 NS_118 0 1.3586848279842204e-03
GC_7_119 b_7 NI_7 NS_119 0 -9.8953529302121725e-04
GC_7_120 b_7 NI_7 NS_120 0 -2.9418847595874585e-03
GC_7_121 b_7 NI_7 NS_121 0 1.8902852114441341e-03
GC_7_122 b_7 NI_7 NS_122 0 -1.9088488299260968e-05
GC_7_123 b_7 NI_7 NS_123 0 -1.3292016220294169e-07
GC_7_124 b_7 NI_7 NS_124 0 -6.8074241105348643e-08
GC_7_125 b_7 NI_7 NS_125 0 9.2132931544714500e-11
GC_7_126 b_7 NI_7 NS_126 0 -2.0426275497231071e-09
GC_7_127 b_7 NI_7 NS_127 0 -1.3991584083405404e-03
GC_7_128 b_7 NI_7 NS_128 0 -2.4217634439046070e-03
GC_7_129 b_7 NI_7 NS_129 0 -4.1847029932917516e-04
GC_7_130 b_7 NI_7 NS_130 0 9.1473296049794661e-04
GC_7_131 b_7 NI_7 NS_131 0 -1.9252501810574070e-03
GC_7_132 b_7 NI_7 NS_132 0 1.7403948149612471e-03
GC_7_133 b_7 NI_7 NS_133 0 1.1232822465062492e-02
GC_7_134 b_7 NI_7 NS_134 0 -3.6181922855782127e-05
GC_7_135 b_7 NI_7 NS_135 0 3.6316863346934909e-06
GC_7_136 b_7 NI_7 NS_136 0 4.0782959677011086e-08
GC_7_137 b_7 NI_7 NS_137 0 -1.2220518439263678e-10
GC_7_138 b_7 NI_7 NS_138 0 2.9770982973319697e-09
GC_7_139 b_7 NI_7 NS_139 0 -2.2241447075952419e-03
GC_7_140 b_7 NI_7 NS_140 0 -4.2734433260865267e-03
GC_7_141 b_7 NI_7 NS_141 0 -2.3599194525801797e-03
GC_7_142 b_7 NI_7 NS_142 0 1.1521932537318921e-02
GC_7_143 b_7 NI_7 NS_143 0 -5.8127072235763435e-03
GC_7_144 b_7 NI_7 NS_144 0 -4.7341063236883254e-03
GD_7_1 b_7 NI_7 NA_1 0 1.8869350555708140e-03
GD_7_2 b_7 NI_7 NA_2 0 1.3928245167370127e-06
GD_7_3 b_7 NI_7 NA_3 0 6.1194615963220417e-03
GD_7_4 b_7 NI_7 NA_4 0 -1.0917433071322557e-04
GD_7_5 b_7 NI_7 NA_5 0 5.0627972593922363e-02
GD_7_6 b_7 NI_7 NA_6 0 6.8938798193227200e-04
GD_7_7 b_7 NI_7 NA_7 0 -4.9495930321987937e-02
GD_7_8 b_7 NI_7 NA_8 0 1.3241930911043559e-01
GD_7_9 b_7 NI_7 NA_9 0 3.0482265331857241e-02
GD_7_10 b_7 NI_7 NA_10 0 1.9047819960769322e-03
GD_7_11 b_7 NI_7 NA_11 0 6.1933763447625089e-03
GD_7_12 b_7 NI_7 NA_12 0 -3.4055192441957705e-04
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 4.2309798798352491e-03
GC_8_2 b_8 NI_8 NS_2 0 -1.1007814058955084e-05
GC_8_3 b_8 NI_8 NS_3 0 9.2772587358764930e-07
GC_8_4 b_8 NI_8 NS_4 0 -2.5046967603839722e-09
GC_8_5 b_8 NI_8 NS_5 0 -1.4960896131719678e-10
GC_8_6 b_8 NI_8 NS_6 0 -4.2477306506130037e-10
GC_8_7 b_8 NI_8 NS_7 0 -3.6268377873436880e-04
GC_8_8 b_8 NI_8 NS_8 0 -1.3120923076184042e-03
GC_8_9 b_8 NI_8 NS_9 0 -1.0797799995486627e-03
GC_8_10 b_8 NI_8 NS_10 0 2.8544950042564362e-03
GC_8_11 b_8 NI_8 NS_11 0 -2.6850997098346900e-03
GC_8_12 b_8 NI_8 NS_12 0 -1.6462129937818203e-03
GC_8_13 b_8 NI_8 NS_13 0 5.0793347063051233e-03
GC_8_14 b_8 NI_8 NS_14 0 -1.8527002080211008e-05
GC_8_15 b_8 NI_8 NS_15 0 7.3020106124476568e-07
GC_8_16 b_8 NI_8 NS_16 0 -1.2333468557248498e-08
GC_8_17 b_8 NI_8 NS_17 0 1.3409497978786207e-10
GC_8_18 b_8 NI_8 NS_18 0 9.6871384450632902e-10
GC_8_19 b_8 NI_8 NS_19 0 9.0804996959010912e-04
GC_8_20 b_8 NI_8 NS_20 0 -1.9384015433245114e-03
GC_8_21 b_8 NI_8 NS_21 0 -4.6724832410655779e-03
GC_8_22 b_8 NI_8 NS_22 0 3.6650264663568049e-04
GC_8_23 b_8 NI_8 NS_23 0 -2.4149410550241292e-03
GC_8_24 b_8 NI_8 NS_24 0 3.0592314903017822e-03
GC_8_25 b_8 NI_8 NS_25 0 1.0862657108892712e-02
GC_8_26 b_8 NI_8 NS_26 0 -3.5594961285035186e-05
GC_8_27 b_8 NI_8 NS_27 0 3.6565786357062598e-06
GC_8_28 b_8 NI_8 NS_28 0 4.5410354544774218e-08
GC_8_29 b_8 NI_8 NS_29 0 -1.1479122905347837e-10
GC_8_30 b_8 NI_8 NS_30 0 3.2123773313226009e-09
GC_8_31 b_8 NI_8 NS_31 0 -1.8529868530458499e-03
GC_8_32 b_8 NI_8 NS_32 0 -4.1628218413723760e-03
GC_8_33 b_8 NI_8 NS_33 0 -2.2902858852993650e-03
GC_8_34 b_8 NI_8 NS_34 0 1.0456459067220864e-02
GC_8_35 b_8 NI_8 NS_35 0 -6.1509419875830675e-03
GC_8_36 b_8 NI_8 NS_36 0 -5.2208012896738784e-03
GC_8_37 b_8 NI_8 NS_37 0 1.2344693291192273e-03
GC_8_38 b_8 NI_8 NS_38 0 -1.9200283190478177e-05
GC_8_39 b_8 NI_8 NS_39 0 -1.6566662509038994e-07
GC_8_40 b_8 NI_8 NS_40 0 -7.2745804917330447e-08
GC_8_41 b_8 NI_8 NS_41 0 8.4510117988408283e-11
GC_8_42 b_8 NI_8 NS_42 0 -2.2770252483671977e-09
GC_8_43 b_8 NI_8 NS_43 0 -1.3091991432067867e-03
GC_8_44 b_8 NI_8 NS_44 0 -2.3678855538198647e-03
GC_8_45 b_8 NI_8 NS_45 0 -3.5156966773381196e-04
GC_8_46 b_8 NI_8 NS_46 0 7.8836348673197269e-04
GC_8_47 b_8 NI_8 NS_47 0 -1.4416385091777849e-03
GC_8_48 b_8 NI_8 NS_48 0 1.7754268130705563e-03
GC_8_49 b_8 NI_8 NS_49 0 5.4843824144467142e-03
GC_8_50 b_8 NI_8 NS_50 0 -1.7139696260626732e-05
GC_8_51 b_8 NI_8 NS_51 0 3.9079478424647975e-06
GC_8_52 b_8 NI_8 NS_52 0 2.8019695410545401e-07
GC_8_53 b_8 NI_8 NS_53 0 7.9557076700317540e-10
GC_8_54 b_8 NI_8 NS_54 0 2.7616671162318326e-08
GC_8_55 b_8 NI_8 NS_55 0 -3.6911708103883241e-04
GC_8_56 b_8 NI_8 NS_56 0 -2.0512083117275315e-03
GC_8_57 b_8 NI_8 NS_57 0 -7.3054742329627640e-04
GC_8_58 b_8 NI_8 NS_58 0 1.4830214422849593e-03
GC_8_59 b_8 NI_8 NS_59 0 -5.1614094384688182e-03
GC_8_60 b_8 NI_8 NS_60 0 -3.0585858755699203e-03
GC_8_61 b_8 NI_8 NS_61 0 4.8536552541218497e-02
GC_8_62 b_8 NI_8 NS_62 0 -2.2743854750322125e-04
GC_8_63 b_8 NI_8 NS_63 0 8.3302383913746824e-07
GC_8_64 b_8 NI_8 NS_64 0 -6.3071450988618584e-07
GC_8_65 b_8 NI_8 NS_65 0 -9.7210182641308706e-10
GC_8_66 b_8 NI_8 NS_66 0 -3.2569423280657185e-08
GC_8_67 b_8 NI_8 NS_67 0 -2.3416311478097359e-02
GC_8_68 b_8 NI_8 NS_68 0 -1.3900300372962726e-02
GC_8_69 b_8 NI_8 NS_69 0 1.1403223908456977e-02
GC_8_70 b_8 NI_8 NS_70 0 1.4942438470152352e-02
GC_8_71 b_8 NI_8 NS_71 0 -4.3469993171023451e-02
GC_8_72 b_8 NI_8 NS_72 0 7.5391534381787908e-03
GC_8_73 b_8 NI_8 NS_73 0 -1.7636204531709326e-01
GC_8_74 b_8 NI_8 NS_74 0 8.6546710599174465e-04
GC_8_75 b_8 NI_8 NS_75 0 -1.5389421994267642e-05
GC_8_76 b_8 NI_8 NS_76 0 4.6154713342139433e-06
GC_8_77 b_8 NI_8 NS_77 0 6.2867302578610220e-09
GC_8_78 b_8 NI_8 NS_78 0 1.6582508491266824e-07
GC_8_79 b_8 NI_8 NS_79 0 -5.0274110916476558e-02
GC_8_80 b_8 NI_8 NS_80 0 -5.1965752474653480e-02
GC_8_81 b_8 NI_8 NS_81 0 -1.6950628911070922e-02
GC_8_82 b_8 NI_8 NS_82 0 -7.2073018679154568e-02
GC_8_83 b_8 NI_8 NS_83 0 1.2915557785434265e-01
GC_8_84 b_8 NI_8 NS_84 0 -7.4440424295501000e-03
GC_8_85 b_8 NI_8 NS_85 0 2.2000012097140700e-01
GC_8_86 b_8 NI_8 NS_86 0 -8.4117228609275339e-04
GC_8_87 b_8 NI_8 NS_87 0 3.0177543230751136e-05
GC_8_88 b_8 NI_8 NS_88 0 -3.3623526874322140e-06
GC_8_89 b_8 NI_8 NS_89 0 -8.0226512191254791e-10
GC_8_90 b_8 NI_8 NS_90 0 -2.1007102096480771e-07
GC_8_91 b_8 NI_8 NS_91 0 -2.4188102222222240e-02
GC_8_92 b_8 NI_8 NS_92 0 1.1786351176150314e-02
GC_8_93 b_8 NI_8 NS_93 0 -1.7257684473435723e-02
GC_8_94 b_8 NI_8 NS_94 0 5.5409695312003418e-02
GC_8_95 b_8 NI_8 NS_95 0 -1.3437384033800689e-01
GC_8_96 b_8 NI_8 NS_96 0 5.8053026372330814e-03
GC_8_97 b_8 NI_8 NS_97 0 -4.6256029091385129e-05
GC_8_98 b_8 NI_8 NS_98 0 8.9271627124154266e-07
GC_8_99 b_8 NI_8 NS_99 0 3.4279827431127183e-06
GC_8_100 b_8 NI_8 NS_100 0 2.8834742544733974e-07
GC_8_101 b_8 NI_8 NS_101 0 6.8376516474789621e-10
GC_8_102 b_8 NI_8 NS_102 0 2.9366421721859141e-08
GC_8_103 b_8 NI_8 NS_103 0 1.9288203279010084e-04
GC_8_104 b_8 NI_8 NS_104 0 -2.3626255197072769e-03
GC_8_105 b_8 NI_8 NS_105 0 -7.4794460845667909e-04
GC_8_106 b_8 NI_8 NS_106 0 1.3568651552256822e-03
GC_8_107 b_8 NI_8 NS_107 0 -9.8356816670829624e-04
GC_8_108 b_8 NI_8 NS_108 0 -2.9411746040699741e-03
GC_8_109 b_8 NI_8 NS_109 0 4.1960295689752368e-02
GC_8_110 b_8 NI_8 NS_110 0 -1.7447883246396453e-04
GC_8_111 b_8 NI_8 NS_111 0 5.8278955020046512e-07
GC_8_112 b_8 NI_8 NS_112 0 -5.1406421246803046e-07
GC_8_113 b_8 NI_8 NS_113 0 -7.6687603356963428e-10
GC_8_114 b_8 NI_8 NS_114 0 -3.2399395551951267e-08
GC_8_115 b_8 NI_8 NS_115 0 -1.5013447283019224e-02
GC_8_116 b_8 NI_8 NS_116 0 -9.2415751361634990e-03
GC_8_117 b_8 NI_8 NS_117 0 3.6749520987320004e-03
GC_8_118 b_8 NI_8 NS_118 0 1.1740814065974681e-02
GC_8_119 b_8 NI_8 NS_119 0 -3.3755359599609694e-02
GC_8_120 b_8 NI_8 NS_120 0 6.8939495835625992e-03
GC_8_121 b_8 NI_8 NS_121 0 1.1241001810520410e-02
GC_8_122 b_8 NI_8 NS_122 0 -3.6207626975927611e-05
GC_8_123 b_8 NI_8 NS_123 0 3.6332029796775134e-06
GC_8_124 b_8 NI_8 NS_124 0 4.0772385705428225e-08
GC_8_125 b_8 NI_8 NS_125 0 -1.2221549402619504e-10
GC_8_126 b_8 NI_8 NS_126 0 2.9775577025116685e-09
GC_8_127 b_8 NI_8 NS_127 0 -2.2254286062979457e-03
GC_8_128 b_8 NI_8 NS_128 0 -4.2732797415505654e-03
GC_8_129 b_8 NI_8 NS_129 0 -2.3606664513181877e-03
GC_8_130 b_8 NI_8 NS_130 0 1.1523697443942335e-02
GC_8_131 b_8 NI_8 NS_131 0 -5.8180349138055743e-03
GC_8_132 b_8 NI_8 NS_132 0 -4.7341176873562808e-03
GC_8_133 b_8 NI_8 NS_133 0 1.9945303200888812e-03
GC_8_134 b_8 NI_8 NS_134 0 -1.9465309958756369e-05
GC_8_135 b_8 NI_8 NS_135 0 -1.0430733282720278e-07
GC_8_136 b_8 NI_8 NS_136 0 -6.8161397846871874e-08
GC_8_137 b_8 NI_8 NS_137 0 9.1717140375285405e-11
GC_8_138 b_8 NI_8 NS_138 0 -2.0393257383904818e-09
GC_8_139 b_8 NI_8 NS_139 0 -1.4091648215697401e-03
GC_8_140 b_8 NI_8 NS_140 0 -2.4180821574154867e-03
GC_8_141 b_8 NI_8 NS_141 0 -4.2767569372560807e-04
GC_8_142 b_8 NI_8 NS_142 0 9.4104142098488594e-04
GC_8_143 b_8 NI_8 NS_143 0 -1.9915333986704939e-03
GC_8_144 b_8 NI_8 NS_144 0 1.7386982752066768e-03
GD_8_1 b_8 NI_8 NA_1 0 5.6840740902168033e-06
GD_8_2 b_8 NI_8 NA_2 0 1.8866867537985870e-03
GD_8_3 b_8 NI_8 NA_3 0 -1.0908552512925597e-04
GD_8_4 b_8 NI_8 NA_4 0 6.1354669904669246e-03
GD_8_5 b_8 NI_8 NA_5 0 6.9207054480018644e-04
GD_8_6 b_8 NI_8 NA_6 0 5.0627972643333595e-02
GD_8_7 b_8 NI_8 NA_7 0 1.3241906414361970e-01
GD_8_8 b_8 NI_8 NA_8 0 -4.9495930326954700e-02
GD_8_9 b_8 NI_8 NA_9 0 1.9010271344699601e-03
GD_8_10 b_8 NI_8 NA_10 0 3.0480802347834325e-02
GD_8_11 b_8 NI_8 NA_11 0 -3.4103988353148914e-04
GD_8_12 b_8 NI_8 NA_12 0 6.1768124883823626e-03
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 -2.1052848153026935e-04
GC_9_2 b_9 NI_9 NS_2 0 -2.2379586797911221e-06
GC_9_3 b_9 NI_9 NS_3 0 4.5991304048799298e-08
GC_9_4 b_9 NI_9 NS_4 0 -1.2154977113660121e-10
GC_9_5 b_9 NI_9 NS_5 0 6.0706441090385156e-11
GC_9_6 b_9 NI_9 NS_6 0 4.8867581069696708e-11
GC_9_7 b_9 NI_9 NS_7 0 4.0508612041620449e-04
GC_9_8 b_9 NI_9 NS_8 0 -3.9700991043333244e-04
GC_9_9 b_9 NI_9 NS_9 0 -9.8073459387535995e-04
GC_9_10 b_9 NI_9 NS_10 0 -2.0966682633599806e-04
GC_9_11 b_9 NI_9 NS_11 0 4.2797076828173018e-04
GC_9_12 b_9 NI_9 NS_12 0 7.9429805004137028e-04
GC_9_13 b_9 NI_9 NS_13 0 4.8857469948701136e-04
GC_9_14 b_9 NI_9 NS_14 0 -2.9269411704293042e-06
GC_9_15 b_9 NI_9 NS_15 0 2.7250880790060975e-07
GC_9_16 b_9 NI_9 NS_16 0 -2.9640707771797598e-09
GC_9_17 b_9 NI_9 NS_17 0 -6.3831790599590281e-11
GC_9_18 b_9 NI_9 NS_18 0 4.9128941340308061e-11
GC_9_19 b_9 NI_9 NS_19 0 5.1373569526465908e-04
GC_9_20 b_9 NI_9 NS_20 0 -1.4982876484489314e-04
GC_9_21 b_9 NI_9 NS_21 0 -1.7726119573521675e-04
GC_9_22 b_9 NI_9 NS_22 0 -1.0127027008214045e-03
GC_9_23 b_9 NI_9 NS_23 0 -1.2278958845223626e-03
GC_9_24 b_9 NI_9 NS_24 0 -1.1792200207808483e-03
GC_9_25 b_9 NI_9 NS_25 0 1.3427748959051237e-03
GC_9_26 b_9 NI_9 NS_26 0 -9.1430283810851225e-06
GC_9_27 b_9 NI_9 NS_27 0 2.1359231098526490e-07
GC_9_28 b_9 NI_9 NS_28 0 -1.3119146083541649e-08
GC_9_29 b_9 NI_9 NS_29 0 1.1305781787352071e-10
GC_9_30 b_9 NI_9 NS_30 0 -1.8759295460792236e-10
GC_9_31 b_9 NI_9 NS_31 0 6.6878979212585366e-04
GC_9_32 b_9 NI_9 NS_32 0 -1.1220537134049226e-03
GC_9_33 b_9 NI_9 NS_33 0 -2.6054955705728786e-03
GC_9_34 b_9 NI_9 NS_34 0 3.9275352479384479e-05
GC_9_35 b_9 NI_9 NS_35 0 -1.5513308491436407e-04
GC_9_36 b_9 NI_9 NS_36 0 2.0670225277805705e-03
GC_9_37 b_9 NI_9 NS_37 0 2.3309835117901485e-03
GC_9_38 b_9 NI_9 NS_38 0 -6.0826371746999266e-06
GC_9_39 b_9 NI_9 NS_39 0 6.8137038605111631e-07
GC_9_40 b_9 NI_9 NS_40 0 4.6378329350714062e-09
GC_9_41 b_9 NI_9 NS_41 0 -1.2227884430301515e-10
GC_9_42 b_9 NI_9 NS_42 0 4.8737609485875716e-10
GC_9_43 b_9 NI_9 NS_43 0 8.0147215419808589e-06
GC_9_44 b_9 NI_9 NS_44 0 -8.0132596263993400e-04
GC_9_45 b_9 NI_9 NS_45 0 -6.2479285238241161e-04
GC_9_46 b_9 NI_9 NS_46 0 1.1738291695824110e-03
GC_9_47 b_9 NI_9 NS_47 0 -1.8495675702555894e-03
GC_9_48 b_9 NI_9 NS_48 0 -1.4232095103737842e-03
GC_9_49 b_9 NI_9 NS_49 0 1.2344750425246221e-03
GC_9_50 b_9 NI_9 NS_50 0 -1.9200359762760583e-05
GC_9_51 b_9 NI_9 NS_51 0 -1.6565620384632677e-07
GC_9_52 b_9 NI_9 NS_52 0 -7.2746318345661239e-08
GC_9_53 b_9 NI_9 NS_53 0 8.4495288985337364e-11
GC_9_54 b_9 NI_9 NS_54 0 -2.2768686473882705e-09
GC_9_55 b_9 NI_9 NS_55 0 -1.3092006272325746e-03
GC_9_56 b_9 NI_9 NS_56 0 -2.3678852794049516e-03
GC_9_57 b_9 NI_9 NS_57 0 -3.5157008441021471e-04
GC_9_58 b_9 NI_9 NS_58 0 7.8836385719303112e-04
GC_9_59 b_9 NI_9 NS_59 0 -1.4416426295177614e-03
GC_9_60 b_9 NI_9 NS_60 0 1.7754263218756805e-03
GC_9_61 b_9 NI_9 NS_61 0 1.0864943270447619e-02
GC_9_62 b_9 NI_9 NS_62 0 -3.5600529508420270e-05
GC_9_63 b_9 NI_9 NS_63 0 3.6569563861724312e-06
GC_9_64 b_9 NI_9 NS_64 0 4.5407222612029687e-08
GC_9_65 b_9 NI_9 NS_65 0 -1.1478141557246069e-10
GC_9_66 b_9 NI_9 NS_66 0 3.2123229186353370e-09
GC_9_67 b_9 NI_9 NS_67 0 -1.8532685974522222e-03
GC_9_68 b_9 NI_9 NS_68 0 -4.1629108672276089e-03
GC_9_69 b_9 NI_9 NS_69 0 -2.2907093992692901e-03
GC_9_70 b_9 NI_9 NS_70 0 1.0457063710973156e-02
GC_9_71 b_9 NI_9 NS_71 0 -6.1523321214182469e-03
GC_9_72 b_9 NI_9 NS_72 0 -5.2206578141556778e-03
GC_9_73 b_9 NI_9 NS_73 0 4.1960295689779721e-02
GC_9_74 b_9 NI_9 NS_74 0 -1.7447883246410163e-04
GC_9_75 b_9 NI_9 NS_75 0 5.8278955020847742e-07
GC_9_76 b_9 NI_9 NS_76 0 -5.1406421246811442e-07
GC_9_77 b_9 NI_9 NS_77 0 -7.6687603356978907e-10
GC_9_78 b_9 NI_9 NS_78 0 -3.2399395551949698e-08
GC_9_79 b_9 NI_9 NS_79 0 -1.5013447283021465e-02
GC_9_80 b_9 NI_9 NS_80 0 -9.2415751361648920e-03
GC_9_81 b_9 NI_9 NS_81 0 3.6749520987269702e-03
GC_9_82 b_9 NI_9 NS_82 0 1.1740814065979131e-02
GC_9_83 b_9 NI_9 NS_83 0 -3.3755359599628616e-02
GC_9_84 b_9 NI_9 NS_84 0 6.8939495835610180e-03
GC_9_85 b_9 NI_9 NS_85 0 -3.8369878989959667e-05
GC_9_86 b_9 NI_9 NS_86 0 8.7899445061142243e-07
GC_9_87 b_9 NI_9 NS_87 0 3.4293754233100692e-06
GC_9_88 b_9 NI_9 NS_88 0 2.8834905730743678e-07
GC_9_89 b_9 NI_9 NS_89 0 6.8381509573632753e-10
GC_9_90 b_9 NI_9 NS_90 0 2.9367357449012823e-08
GC_9_91 b_9 NI_9 NS_91 0 1.8798474525433731e-04
GC_9_92 b_9 NI_9 NS_92 0 -2.3622896214916030e-03
GC_9_93 b_9 NI_9 NS_93 0 -7.4633196007466217e-04
GC_9_94 b_9 NI_9 NS_94 0 1.3586848279843688e-03
GC_9_95 b_9 NI_9 NS_95 0 -9.8953529302179036e-04
GC_9_96 b_9 NI_9 NS_96 0 -2.9418847595874958e-03
GC_9_97 b_9 NI_9 NS_97 0 2.2400108303505370e-01
GC_9_98 b_9 NI_9 NS_98 0 -8.4675561262135646e-04
GC_9_99 b_9 NI_9 NS_99 0 3.0352476750355526e-05
GC_9_100 b_9 NI_9 NS_100 0 -3.3545496870844934e-06
GC_9_101 b_9 NI_9 NS_101 0 -7.7375340993698707e-10
GC_9_102 b_9 NI_9 NS_102 0 -2.0977095889152244e-07
GC_9_103 b_9 NI_9 NS_103 0 -2.4709043054827007e-02
GC_9_104 b_9 NI_9 NS_104 0 1.1897478167225910e-02
GC_9_105 b_9 NI_9 NS_105 0 -1.7546764642470628e-02
GC_9_106 b_9 NI_9 NS_106 0 5.6447036755187377e-02
GC_9_107 b_9 NI_9 NS_107 0 -1.3690356146642885e-01
GC_9_108 b_9 NI_9 NS_108 0 5.8883044032311217e-03
GC_9_109 b_9 NI_9 NS_109 0 -1.6867773860048016e-01
GC_9_110 b_9 NI_9 NS_110 0 8.1246271128150983e-04
GC_9_111 b_9 NI_9 NS_111 0 -1.1179346634451217e-05
GC_9_112 b_9 NI_9 NS_112 0 4.5242878230459427e-06
GC_9_113 b_9 NI_9 NS_113 0 5.7757966030295800e-09
GC_9_114 b_9 NI_9 NS_114 0 1.7340096968452293e-07
GC_9_115 b_9 NI_9 NS_115 0 -5.1296420120694443e-02
GC_9_116 b_9 NI_9 NS_116 0 -5.2321761979893307e-02
GC_9_117 b_9 NI_9 NS_117 0 -1.8162026636973919e-02
GC_9_118 b_9 NI_9 NS_118 0 -6.9460373104216599e-02
GC_9_119 b_9 NI_9 NS_119 0 1.2462987502525150e-01
GC_9_120 b_9 NI_9 NS_120 0 -7.4284086228288432e-03
GC_9_121 b_9 NI_9 NS_121 0 4.5219216564568135e-02
GC_9_122 b_9 NI_9 NS_122 0 -2.1057606527248267e-04
GC_9_123 b_9 NI_9 NS_123 0 7.7895297476854829e-08
GC_9_124 b_9 NI_9 NS_124 0 -5.9496955626725141e-07
GC_9_125 b_9 NI_9 NS_125 0 -9.2824714312299078e-10
GC_9_126 b_9 NI_9 NS_126 0 -3.1476532821460468e-08
GC_9_127 b_9 NI_9 NS_127 0 -2.4219205289253799e-02
GC_9_128 b_9 NI_9 NS_128 0 -1.3397004326800306e-02
GC_9_129 b_9 NI_9 NS_129 0 1.4228520026941773e-02
GC_9_130 b_9 NI_9 NS_130 0 1.4700435691788399e-02
GC_9_131 b_9 NI_9 NS_131 0 -4.2169641053321869e-02
GC_9_132 b_9 NI_9 NS_132 0 5.9572275103232939e-03
GC_9_133 b_9 NI_9 NS_133 0 7.5494467118858918e-03
GC_9_134 b_9 NI_9 NS_134 0 -2.7274375597351259e-05
GC_9_135 b_9 NI_9 NS_135 0 4.2560422141462619e-06
GC_9_136 b_9 NI_9 NS_136 0 2.4799665090828933e-07
GC_9_137 b_9 NI_9 NS_137 0 7.3564826584918451e-10
GC_9_138 b_9 NI_9 NS_138 0 2.6666795432527012e-08
GC_9_139 b_9 NI_9 NS_139 0 -1.0895574383373784e-03
GC_9_140 b_9 NI_9 NS_140 0 -2.2178332659894906e-03
GC_9_141 b_9 NI_9 NS_141 0 -8.3883646034535030e-04
GC_9_142 b_9 NI_9 NS_142 0 3.4881331257413323e-03
GC_9_143 b_9 NI_9 NS_143 0 -5.7610150436300783e-03
GC_9_144 b_9 NI_9 NS_144 0 -2.7574484406131098e-03
GD_9_1 b_9 NI_9 NA_1 0 4.3422080670183578e-04
GD_9_2 b_9 NI_9 NA_2 0 3.6756584346027334e-04
GD_9_3 b_9 NI_9 NA_3 0 1.2057087295072448e-03
GD_9_4 b_9 NI_9 NA_4 0 1.9265549640022528e-04
GD_9_5 b_9 NI_9 NA_5 0 6.1354681668953012e-03
GD_9_6 b_9 NI_9 NA_6 0 -1.0918537265261697e-04
GD_9_7 b_9 NI_9 NA_7 0 3.0480802347834325e-02
GD_9_8 b_9 NI_9 NA_8 0 1.9047819960769322e-03
GD_9_9 b_9 NI_9 NA_9 0 -5.0105580198010882e-02
GD_9_10 b_9 NI_9 NA_10 0 1.3167218582495305e-01
GD_9_11 b_9 NI_9 NA_11 0 5.1203269514768841e-02
GD_9_12 b_9 NI_9 NA_12 0 8.1611027282107659e-05
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 4.8886184218286343e-04
GC_10_2 b_10 NI_10 NS_2 0 -2.9276272512430129e-06
GC_10_3 b_10 NI_10 NS_3 0 2.7255353944077531e-07
GC_10_4 b_10 NI_10 NS_4 0 -2.9640988258279848e-09
GC_10_5 b_10 NI_10 NS_5 0 -6.3831889409291383e-11
GC_10_6 b_10 NI_10 NS_6 0 4.9149285984524311e-11
GC_10_7 b_10 NI_10 NS_7 0 5.1365524828289523e-04
GC_10_8 b_10 NI_10 NS_8 0 -1.4980104231320662e-04
GC_10_9 b_10 NI_10 NS_9 0 -1.7724777101623619e-04
GC_10_10 b_10 NI_10 NS_10 0 -1.0126566839038730e-03
GC_10_11 b_10 NI_10 NS_11 0 -1.2280970297915297e-03
GC_10_12 b_10 NI_10 NS_12 0 -1.1792311156218068e-03
GC_10_13 b_10 NI_10 NS_13 0 -2.1459728878750735e-04
GC_10_14 b_10 NI_10 NS_14 0 -2.2224595469260280e-06
GC_10_15 b_10 NI_10 NS_15 0 4.5685930043921610e-08
GC_10_16 b_10 NI_10 NS_16 0 -1.0948931468039835e-10
GC_10_17 b_10 NI_10 NS_17 0 6.0712634212579044e-11
GC_10_18 b_10 NI_10 NS_18 0 4.8266785235884902e-11
GC_10_19 b_10 NI_10 NS_19 0 4.0681431310652944e-04
GC_10_20 b_10 NI_10 NS_20 0 -3.9665454009978280e-04
GC_10_21 b_10 NI_10 NS_21 0 -9.8081005079664850e-04
GC_10_22 b_10 NI_10 NS_22 0 -2.1225315595396364e-04
GC_10_23 b_10 NI_10 NS_23 0 4.2995263517617765e-04
GC_10_24 b_10 NI_10 NS_24 0 7.9393648726596062e-04
GC_10_25 b_10 NI_10 NS_25 0 2.3226481820075745e-03
GC_10_26 b_10 NI_10 NS_26 0 -6.0665490999753319e-06
GC_10_27 b_10 NI_10 NS_27 0 6.7996611247118616e-07
GC_10_28 b_10 NI_10 NS_28 0 4.6420344461708773e-09
GC_10_29 b_10 NI_10 NS_29 0 -1.2227704227296513e-10
GC_10_30 b_10 NI_10 NS_30 0 4.8672326643983815e-10
GC_10_31 b_10 NI_10 NS_31 0 1.1437261314735881e-05
GC_10_32 b_10 NI_10 NS_32 0 -8.0083496624697669e-04
GC_10_33 b_10 NI_10 NS_33 0 -6.2462121898550042e-04
GC_10_34 b_10 NI_10 NS_34 0 1.1716323368554588e-03
GC_10_35 b_10 NI_10 NS_35 0 -1.8438019473252273e-03
GC_10_36 b_10 NI_10 NS_36 0 -1.4230868201695558e-03
GC_10_37 b_10 NI_10 NS_37 0 1.3427743835553699e-03
GC_10_38 b_10 NI_10 NS_38 0 -9.1430271645834272e-06
GC_10_39 b_10 NI_10 NS_39 0 2.1359225935050415e-07
GC_10_40 b_10 NI_10 NS_40 0 -1.3119145181220647e-08
GC_10_41 b_10 NI_10 NS_41 0 1.1305781924860101e-10
GC_10_42 b_10 NI_10 NS_42 0 -1.8759296752958280e-10
GC_10_43 b_10 NI_10 NS_43 0 6.6878987263332501e-04
GC_10_44 b_10 NI_10 NS_44 0 -1.1220537732613697e-03
GC_10_45 b_10 NI_10 NS_45 0 -2.6054955647410996e-03
GC_10_46 b_10 NI_10 NS_46 0 3.9275190003536172e-05
GC_10_47 b_10 NI_10 NS_47 0 -1.5513279108810853e-04
GC_10_48 b_10 NI_10 NS_48 0 2.0670225004261814e-03
GC_10_49 b_10 NI_10 NS_49 0 1.0862693856977834e-02
GC_10_50 b_10 NI_10 NS_50 0 -3.5594952491927790e-05
GC_10_51 b_10 NI_10 NS_51 0 3.6565670975760292e-06
GC_10_52 b_10 NI_10 NS_52 0 4.5410903815687680e-08
GC_10_53 b_10 NI_10 NS_53 0 -1.1477636020362258e-10
GC_10_54 b_10 NI_10 NS_54 0 3.2122170325727006e-09
GC_10_55 b_10 NI_10 NS_55 0 -1.8529917409110682e-03
GC_10_56 b_10 NI_10 NS_56 0 -4.1628193438066913e-03
GC_10_57 b_10 NI_10 NS_57 0 -2.2902894265689308e-03
GC_10_58 b_10 NI_10 NS_58 0 1.0456468031386780e-02
GC_10_59 b_10 NI_10 NS_59 0 -6.1509639060043841e-03
GC_10_60 b_10 NI_10 NS_60 0 -5.2207980239414803e-03
GC_10_61 b_10 NI_10 NS_61 0 1.3273205919123274e-03
GC_10_62 b_10 NI_10 NS_62 0 -1.9513663171619962e-05
GC_10_63 b_10 NI_10 NS_63 0 -1.4172560971402439e-07
GC_10_64 b_10 NI_10 NS_64 0 -7.2812366939666702e-08
GC_10_65 b_10 NI_10 NS_65 0 8.4153281785293752e-11
GC_10_66 b_10 NI_10 NS_66 0 -2.2739453061636711e-09
GC_10_67 b_10 NI_10 NS_67 0 -1.3174988886499230e-03
GC_10_68 b_10 NI_10 NS_68 0 -2.3639640757190002e-03
GC_10_69 b_10 NI_10 NS_69 0 -3.5983148418270268e-04
GC_10_70 b_10 NI_10 NS_70 0 8.1128675830325974e-04
GC_10_71 b_10 NI_10 NS_71 0 -1.5004987608087646e-03
GC_10_72 b_10 NI_10 NS_72 0 1.7745062024233018e-03
GC_10_73 b_10 NI_10 NS_73 0 -4.6256029092880881e-05
GC_10_74 b_10 NI_10 NS_74 0 8.9271627124896859e-07
GC_10_75 b_10 NI_10 NS_75 0 3.4279827431122795e-06
GC_10_76 b_10 NI_10 NS_76 0 2.8834742544734472e-07
GC_10_77 b_10 NI_10 NS_77 0 6.8376516474791100e-10
GC_10_78 b_10 NI_10 NS_78 0 2.9366421721859022e-08
GC_10_79 b_10 NI_10 NS_79 0 1.9288203279022671e-04
GC_10_80 b_10 NI_10 NS_80 0 -2.3626255197072015e-03
GC_10_81 b_10 NI_10 NS_81 0 -7.4794460845640533e-04
GC_10_82 b_10 NI_10 NS_82 0 1.3568651552254337e-03
GC_10_83 b_10 NI_10 NS_83 0 -9.8356816670726473e-04
GC_10_84 b_10 NI_10 NS_84 0 -2.9411746040698926e-03
GC_10_85 b_10 NI_10 NS_85 0 4.1946350052461764e-02
GC_10_86 b_10 NI_10 NS_86 0 -1.7440834779706131e-04
GC_10_87 b_10 NI_10 NS_87 0 5.7873283472912718e-07
GC_10_88 b_10 NI_10 NS_88 0 -5.1402838048933909e-07
GC_10_89 b_10 NI_10 NS_89 0 -7.6680262802042776e-10
GC_10_90 b_10 NI_10 NS_90 0 -3.2399854190571804e-08
GC_10_91 b_10 NI_10 NS_91 0 -1.5011431217308240e-02
GC_10_92 b_10 NI_10 NS_92 0 -9.2416782120903485e-03
GC_10_93 b_10 NI_10 NS_93 0 3.6761889300983789e-03
GC_10_94 b_10 NI_10 NS_94 0 1.1736949771051941e-02
GC_10_95 b_10 NI_10 NS_95 0 -3.3746557294646339e-02
GC_10_96 b_10 NI_10 NS_96 0 6.8943091498482947e-03
GC_10_97 b_10 NI_10 NS_97 0 -1.6870749289315806e-01
GC_10_98 b_10 NI_10 NS_98 0 8.1259476657962967e-04
GC_10_99 b_10 NI_10 NS_99 0 -1.1189001963630187e-05
GC_10_100 b_10 NI_10 NS_100 0 4.5244366122383310e-06
GC_10_101 b_10 NI_10 NS_101 0 5.7765682383489782e-09
GC_10_102 b_10 NI_10 NS_102 0 1.7338706376541180e-07
GC_10_103 b_10 NI_10 NS_103 0 -5.1291400589785541e-02
GC_10_104 b_10 NI_10 NS_104 0 -5.2322491294981378e-02
GC_10_105 b_10 NI_10 NS_105 0 -1.8160012978416653e-02
GC_10_106 b_10 NI_10 NS_106 0 -6.9465910528827959e-02
GC_10_107 b_10 NI_10 NS_107 0 1.2465015063600025e-01
GC_10_108 b_10 NI_10 NS_108 0 -7.4269999898423063e-03
GC_10_109 b_10 NI_10 NS_109 0 2.2400108304469904e-01
GC_10_110 b_10 NI_10 NS_110 0 -8.4675561269350003e-04
GC_10_111 b_10 NI_10 NS_111 0 3.0352476755602631e-05
GC_10_112 b_10 NI_10 NS_112 0 -3.3545496871478637e-06
GC_10_113 b_10 NI_10 NS_113 0 -7.7375341011387003e-10
GC_10_114 b_10 NI_10 NS_114 0 -2.0977095888755740e-07
GC_10_115 b_10 NI_10 NS_115 0 -2.4709043055414447e-02
GC_10_116 b_10 NI_10 NS_116 0 1.1897478167111546e-02
GC_10_117 b_10 NI_10 NS_117 0 -1.7546764643830471e-02
GC_10_118 b_10 NI_10 NS_118 0 5.6447036756404799e-02
GC_10_119 b_10 NI_10 NS_119 0 -1.3690356147332902e-01
GC_10_120 b_10 NI_10 NS_120 0 5.8883044021247211e-03
GC_10_121 b_10 NI_10 NS_121 0 7.5502705389227402e-03
GC_10_122 b_10 NI_10 NS_122 0 -2.7274797372547591e-05
GC_10_123 b_10 NI_10 NS_123 0 4.2562823888301434e-06
GC_10_124 b_10 NI_10 NS_124 0 2.4799787114815247e-07
GC_10_125 b_10 NI_10 NS_125 0 7.3566416678482008e-10
GC_10_126 b_10 NI_10 NS_126 0 2.6667003816917148e-08
GC_10_127 b_10 NI_10 NS_127 0 -1.0908210560917611e-03
GC_10_128 b_10 NI_10 NS_128 0 -2.2177893724464812e-03
GC_10_129 b_10 NI_10 NS_129 0 -8.3820905902373731e-04
GC_10_130 b_10 NI_10 NS_130 0 3.4882361911381878e-03
GC_10_131 b_10 NI_10 NS_131 0 -5.7618887277548292e-03
GC_10_132 b_10 NI_10 NS_132 0 -2.7577422718693153e-03
GC_10_133 b_10 NI_10 NS_133 0 4.5236646748357985e-02
GC_10_134 b_10 NI_10 NS_134 0 -2.1070060598431795e-04
GC_10_135 b_10 NI_10 NS_135 0 9.0938068987294190e-08
GC_10_136 b_10 NI_10 NS_136 0 -5.9499129271737305e-07
GC_10_137 b_10 NI_10 NS_137 0 -9.2850190469968645e-10
GC_10_138 b_10 NI_10 NS_138 0 -3.1475498806714499e-08
GC_10_139 b_10 NI_10 NS_139 0 -2.4219581420572737e-02
GC_10_140 b_10 NI_10 NS_140 0 -1.3397401890606718e-02
GC_10_141 b_10 NI_10 NS_141 0 1.4226418210207221e-02
GC_10_142 b_10 NI_10 NS_142 0 1.4703261453936804e-02
GC_10_143 b_10 NI_10 NS_143 0 -4.2182718075536647e-02
GC_10_144 b_10 NI_10 NS_144 0 5.9539188515264569e-03
GD_10_1 b_10 NI_10 NA_1 0 3.6757421026674376e-04
GD_10_2 b_10 NI_10 NA_2 0 4.3455189505917400e-04
GD_10_3 b_10 NI_10 NA_3 0 1.8991362176736312e-04
GD_10_4 b_10 NI_10 NA_4 0 1.2057088590887749e-03
GD_10_5 b_10 NI_10 NA_5 0 -1.0909158462998901e-04
GD_10_6 b_10 NI_10 NA_6 0 6.1194575195962549e-03
GD_10_7 b_10 NI_10 NA_7 0 1.9010271344699601e-03
GD_10_8 b_10 NI_10 NA_8 0 3.0482265331857241e-02
GD_10_9 b_10 NI_10 NA_9 0 1.3167311108266844e-01
GD_10_10 b_10 NI_10 NA_10 0 -5.0105580198682755e-02
GD_10_11 b_10 NI_10 NA_11 0 8.3016615741810017e-05
GD_10_12 b_10 NI_10 NA_12 0 5.1203290464629132e-02
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 -2.1577211839931719e-03
GC_11_2 b_11 NI_11 NS_2 0 3.0993760839374144e-06
GC_11_3 b_11 NI_11 NS_3 0 -1.6353137296808818e-07
GC_11_4 b_11 NI_11 NS_4 0 2.6448827552497201e-09
GC_11_5 b_11 NI_11 NS_5 0 2.6359893505563552e-11
GC_11_6 b_11 NI_11 NS_6 0 1.1477651613103090e-11
GC_11_7 b_11 NI_11 NS_7 0 2.0971551828687907e-04
GC_11_8 b_11 NI_11 NS_8 0 -2.8336012300654078e-06
GC_11_9 b_11 NI_11 NS_9 0 1.7091529040415531e-04
GC_11_10 b_11 NI_11 NS_10 0 -3.1346926928302912e-04
GC_11_11 b_11 NI_11 NS_11 0 1.5860771045782146e-03
GC_11_12 b_11 NI_11 NS_12 0 2.6011047068382137e-04
GC_11_13 b_11 NI_11 NS_13 0 4.2805972161945910e-05
GC_11_14 b_11 NI_11 NS_14 0 -7.1924075308640832e-07
GC_11_15 b_11 NI_11 NS_15 0 7.4135881607495300e-08
GC_11_16 b_11 NI_11 NS_16 0 -2.2966872760649932e-09
GC_11_17 b_11 NI_11 NS_17 0 -2.5681030904620268e-11
GC_11_18 b_11 NI_11 NS_18 0 -3.8702601439812786e-11
GC_11_19 b_11 NI_11 NS_19 0 2.8894597869208281e-04
GC_11_20 b_11 NI_11 NS_20 0 -5.4017262289654102e-06
GC_11_21 b_11 NI_11 NS_21 0 -2.3718108828354571e-05
GC_11_22 b_11 NI_11 NS_22 0 -6.8477759434932379e-04
GC_11_23 b_11 NI_11 NS_23 0 -5.2270867361140199e-04
GC_11_24 b_11 NI_11 NS_24 0 -5.5975475308537399e-04
GC_11_25 b_11 NI_11 NS_25 0 -2.1456487044199684e-04
GC_11_26 b_11 NI_11 NS_26 0 -2.2225270179232197e-06
GC_11_27 b_11 NI_11 NS_27 0 4.5691123600918278e-08
GC_11_28 b_11 NI_11 NS_28 0 -1.0955582683552472e-10
GC_11_29 b_11 NI_11 NS_29 0 6.0712532184624881e-11
GC_11_30 b_11 NI_11 NS_30 0 4.8270504438239686e-11
GC_11_31 b_11 NI_11 NS_31 0 4.0680910259012867e-04
GC_11_32 b_11 NI_11 NS_32 0 -3.9665146071601382e-04
GC_11_33 b_11 NI_11 NS_33 0 -9.8081136884206437e-04
GC_11_34 b_11 NI_11 NS_34 0 -2.1224297933959005e-04
GC_11_35 b_11 NI_11 NS_35 0 4.2993451057162343e-04
GC_11_36 b_11 NI_11 NS_36 0 7.9393952017462106e-04
GC_11_37 b_11 NI_11 NS_37 0 4.8857161821362302e-04
GC_11_38 b_11 NI_11 NS_38 0 -2.9269714399491402e-06
GC_11_39 b_11 NI_11 NS_39 0 2.7250927762800168e-07
GC_11_40 b_11 NI_11 NS_40 0 -2.9640647041570363e-09
GC_11_41 b_11 NI_11 NS_41 0 -6.3831825704813369e-11
GC_11_42 b_11 NI_11 NS_42 0 4.9127724261925249e-11
GC_11_43 b_11 NI_11 NS_43 0 5.1373640084780459e-04
GC_11_44 b_11 NI_11 NS_44 0 -1.4982946194841008e-04
GC_11_45 b_11 NI_11 NS_45 0 -1.7726205497755064e-04
GC_11_46 b_11 NI_11 NS_46 0 -1.0127064845497928e-03
GC_11_47 b_11 NI_11 NS_47 0 -1.2278958749332746e-03
GC_11_48 b_11 NI_11 NS_48 0 -1.1792220318134789e-03
GC_11_49 b_11 NI_11 NS_49 0 5.0795379492554089e-03
GC_11_50 b_11 NI_11 NS_50 0 -1.8527609225408898e-05
GC_11_51 b_11 NI_11 NS_51 0 7.3024486340435618e-07
GC_11_52 b_11 NI_11 NS_52 0 -1.2334102656940115e-08
GC_11_53 b_11 NI_11 NS_53 0 1.3409209295977843e-10
GC_11_54 b_11 NI_11 NS_54 0 9.6875329730628076e-10
GC_11_55 b_11 NI_11 NS_55 0 9.0802500338216859e-04
GC_11_56 b_11 NI_11 NS_56 0 -1.9383887053115443e-03
GC_11_57 b_11 NI_11 NS_57 0 -4.6724996509654865e-03
GC_11_58 b_11 NI_11 NS_58 0 3.6655965377647493e-04
GC_11_59 b_11 NI_11 NS_59 0 -2.4150607668786384e-03
GC_11_60 b_11 NI_11 NS_60 0 3.0592401849205354e-03
GC_11_61 b_11 NI_11 NS_61 0 4.2228725450482235e-03
GC_11_62 b_11 NI_11 NS_62 0 -1.0991489590240789e-05
GC_11_63 b_11 NI_11 NS_63 0 9.2608169996240097e-07
GC_11_64 b_11 NI_11 NS_64 0 -2.5038170766790563e-09
GC_11_65 b_11 NI_11 NS_65 0 -1.4961183510655854e-10
GC_11_66 b_11 NI_11 NS_66 0 -4.2562873433721425e-10
GC_11_67 b_11 NI_11 NS_67 0 -3.5777178697686069e-04
GC_11_68 b_11 NI_11 NS_68 0 -1.3121060881780442e-03
GC_11_69 b_11 NI_11 NS_69 0 -1.0810728105758248e-03
GC_11_70 b_11 NI_11 NS_70 0 2.8527296137075722e-03
GC_11_71 b_11 NI_11 NS_71 0 -2.6788727572073122e-03
GC_11_72 b_11 NI_11 NS_72 0 -1.6454282606839104e-03
GC_11_73 b_11 NI_11 NS_73 0 1.9945303200913436e-03
GC_11_74 b_11 NI_11 NS_74 0 -1.9465309958768163e-05
GC_11_75 b_11 NI_11 NS_75 0 -1.0430733282653326e-07
GC_11_76 b_11 NI_11 NS_76 0 -6.8161397846878914e-08
GC_11_77 b_11 NI_11 NS_77 0 9.1717140375273889e-11
GC_11_78 b_11 NI_11 NS_78 0 -2.0393257383903887e-09
GC_11_79 b_11 NI_11 NS_79 0 -1.4091648215699513e-03
GC_11_80 b_11 NI_11 NS_80 0 -2.4180821574156116e-03
GC_11_81 b_11 NI_11 NS_81 0 -4.2767569372605975e-04
GC_11_82 b_11 NI_11 NS_82 0 9.4104142098530390e-04
GC_11_83 b_11 NI_11 NS_83 0 -1.9915333986721857e-03
GC_11_84 b_11 NI_11 NS_84 0 1.7386982752065515e-03
GC_11_85 b_11 NI_11 NS_85 0 1.1232822465064834e-02
GC_11_86 b_11 NI_11 NS_86 0 -3.6181922855793504e-05
GC_11_87 b_11 NI_11 NS_87 0 3.6316863346941432e-06
GC_11_88 b_11 NI_11 NS_88 0 4.0782959677004270e-08
GC_11_89 b_11 NI_11 NS_89 0 -1.2220518439264754e-10
GC_11_90 b_11 NI_11 NS_90 0 2.9770982973320711e-09
GC_11_91 b_11 NI_11 NS_91 0 -2.2241447075954392e-03
GC_11_92 b_11 NI_11 NS_92 0 -4.2734433260866473e-03
GC_11_93 b_11 NI_11 NS_93 0 -2.3599194525806100e-03
GC_11_94 b_11 NI_11 NS_94 0 1.1521932537319309e-02
GC_11_95 b_11 NI_11 NS_95 0 -5.8127072235779559e-03
GC_11_96 b_11 NI_11 NS_96 0 -4.7341063236884503e-03
GC_11_97 b_11 NI_11 NS_97 0 4.5236646748349221e-02
GC_11_98 b_11 NI_11 NS_98 0 -2.1070060598427369e-04
GC_11_99 b_11 NI_11 NS_99 0 9.0938068984701370e-08
GC_11_100 b_11 NI_11 NS_100 0 -5.9499129271734615e-07
GC_11_101 b_11 NI_11 NS_101 0 -9.2850190469963785e-10
GC_11_102 b_11 NI_11 NS_102 0 -3.1475498806715028e-08
GC_11_103 b_11 NI_11 NS_103 0 -2.4219581420572026e-02
GC_11_104 b_11 NI_11 NS_104 0 -1.3397401890606269e-02
GC_11_105 b_11 NI_11 NS_105 0 1.4226418210208836e-02
GC_11_106 b_11 NI_11 NS_106 0 1.4703261453935388e-02
GC_11_107 b_11 NI_11 NS_107 0 -4.2182718075530576e-02
GC_11_108 b_11 NI_11 NS_108 0 5.9539188515269729e-03
GC_11_109 b_11 NI_11 NS_109 0 7.5494467118860376e-03
GC_11_110 b_11 NI_11 NS_110 0 -2.7274375597352113e-05
GC_11_111 b_11 NI_11 NS_111 0 4.2560422141463169e-06
GC_11_112 b_11 NI_11 NS_112 0 2.4799665090828870e-07
GC_11_113 b_11 NI_11 NS_113 0 7.3564826584918306e-10
GC_11_114 b_11 NI_11 NS_114 0 2.6666795432527045e-08
GC_11_115 b_11 NI_11 NS_115 0 -1.0895574383373884e-03
GC_11_116 b_11 NI_11 NS_116 0 -2.2178332659894980e-03
GC_11_117 b_11 NI_11 NS_117 0 -8.3883646034537719e-04
GC_11_118 b_11 NI_11 NS_118 0 3.4881331257413523e-03
GC_11_119 b_11 NI_11 NS_119 0 -5.7610150436301806e-03
GC_11_120 b_11 NI_11 NS_120 0 -2.7574484406131215e-03
GC_11_121 b_11 NI_11 NS_121 0 2.3570671292937803e-01
GC_11_122 b_11 NI_11 NS_122 0 -8.4010550972380468e-04
GC_11_123 b_11 NI_11 NS_123 0 2.7374986306266388e-05
GC_11_124 b_11 NI_11 NS_124 0 -3.2161877407040324e-06
GC_11_125 b_11 NI_11 NS_125 0 -3.6319368783948096e-11
GC_11_126 b_11 NI_11 NS_126 0 -2.0793646988908162e-07
GC_11_127 b_11 NI_11 NS_127 0 -2.8744445536320443e-02
GC_11_128 b_11 NI_11 NS_128 0 1.2390377859696383e-02
GC_11_129 b_11 NI_11 NS_129 0 -1.4922288901499157e-02
GC_11_130 b_11 NI_11 NS_130 0 6.1041345666854908e-02
GC_11_131 b_11 NI_11 NS_131 0 -1.4475758926399993e-01
GC_11_132 b_11 NI_11 NS_132 0 7.1004793766956571e-03
GC_11_133 b_11 NI_11 NS_133 0 -1.6611341697246579e-01
GC_11_134 b_11 NI_11 NS_134 0 7.7902840579039800e-04
GC_11_135 b_11 NI_11 NS_135 0 -1.0081643537581333e-05
GC_11_136 b_11 NI_11 NS_136 0 4.4063519578991585e-06
GC_11_137 b_11 NI_11 NS_137 0 5.2197958395111431e-09
GC_11_138 b_11 NI_11 NS_138 0 1.7216707023088985e-07
GC_11_139 b_11 NI_11 NS_139 0 -5.0680336461358756e-02
GC_11_140 b_11 NI_11 NS_140 0 -5.0185253008319865e-02
GC_11_141 b_11 NI_11 NS_141 0 -1.8088793263708908e-02
GC_11_142 b_11 NI_11 NS_142 0 -7.4854172974320468e-02
GC_11_143 b_11 NI_11 NS_143 0 1.2153114236378983e-01
GC_11_144 b_11 NI_11 NS_144 0 -5.5012512937953990e-03
GD_11_1 b_11 NI_11 NA_1 0 1.7347945566864654e-04
GD_11_2 b_11 NI_11 NA_2 0 1.9112395193547616e-04
GD_11_3 b_11 NI_11 NA_3 0 4.3454315319714422e-04
GD_11_4 b_11 NI_11 NA_4 0 3.6757071208514774e-04
GD_11_5 b_11 NI_11 NA_5 0 1.8866381494708033e-03
GD_11_6 b_11 NI_11 NA_6 0 1.4129039939162737e-06
GD_11_7 b_11 NI_11 NA_7 0 6.1768124883823626e-03
GD_11_8 b_11 NI_11 NA_8 0 -3.4055192441957705e-04
GD_11_9 b_11 NI_11 NA_9 0 5.1203290464629132e-02
GD_11_10 b_11 NI_11 NA_10 0 8.1611027282107659e-05
GD_11_11 b_11 NI_11 NA_11 0 -4.9038965748759836e-02
GD_11_12 b_11 NI_11 NA_12 0 1.3127129754717567e-01
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 4.8622047272097664e-05
GC_12_2 b_12 NI_12 NS_2 0 -7.3649342468998693e-07
GC_12_3 b_12 NI_12 NS_3 0 7.5254857654443998e-08
GC_12_4 b_12 NI_12 NS_4 0 -2.3063069974402201e-09
GC_12_5 b_12 NI_12 NS_5 0 -2.5694409643499076e-11
GC_12_6 b_12 NI_12 NS_6 0 -3.8290941719243816e-11
GC_12_7 b_12 NI_12 NS_7 0 2.8807983988923488e-04
GC_12_8 b_12 NI_12 NS_8 0 -5.9053451373167138e-06
GC_12_9 b_12 NI_12 NS_9 0 -2.4850639203513637e-05
GC_12_10 b_12 NI_12 NS_10 0 -6.8327333122159700e-04
GC_12_11 b_12 NI_12 NS_11 0 -5.2640450572609128e-04
GC_12_12 b_12 NI_12 NS_12 0 -5.5958812642674632e-04
GC_12_13 b_12 NI_12 NS_13 0 -2.1577210030624358e-03
GC_12_14 b_12 NI_12 NS_14 0 3.0993750469310796e-06
GC_12_15 b_12 NI_12 NS_15 0 -1.6353131712779337e-07
GC_12_16 b_12 NI_12 NS_16 0 2.6448825461724617e-09
GC_12_17 b_12 NI_12 NS_17 0 2.6359893802132872e-11
GC_12_18 b_12 NI_12 NS_18 0 1.1477632502211604e-11
GC_12_19 b_12 NI_12 NS_19 0 2.0971550902044029e-04
GC_12_20 b_12 NI_12 NS_20 0 -2.8335999999038578e-06
GC_12_21 b_12 NI_12 NS_21 0 1.7091525343691352e-04
GC_12_22 b_12 NI_12 NS_22 0 -3.1346924351043477e-04
GC_12_23 b_12 NI_12 NS_23 0 1.5860769724171358e-03
GC_12_24 b_12 NI_12 NS_24 0 2.6011044261725473e-04
GC_12_25 b_12 NI_12 NS_25 0 4.8885680418179675e-04
GC_12_26 b_12 NI_12 NS_26 0 -2.9276499694755417e-06
GC_12_27 b_12 NI_12 NS_27 0 2.7255376258029648e-07
GC_12_28 b_12 NI_12 NS_28 0 -2.9640930729646795e-09
GC_12_29 b_12 NI_12 NS_29 0 -6.3831920924437805e-11
GC_12_30 b_12 NI_12 NS_30 0 4.9148079017427237e-11
GC_12_31 b_12 NI_12 NS_31 0 5.1365613590942827e-04
GC_12_32 b_12 NI_12 NS_32 0 -1.4980161247207419e-04
GC_12_33 b_12 NI_12 NS_33 0 -1.7724827003658600e-04
GC_12_34 b_12 NI_12 NS_34 0 -1.0126608117921297e-03
GC_12_35 b_12 NI_12 NS_35 0 -1.2280956736773435e-03
GC_12_36 b_12 NI_12 NS_36 0 -1.1792330377420192e-03
GC_12_37 b_12 NI_12 NS_37 0 -2.1049773338333068e-04
GC_12_38 b_12 NI_12 NS_38 0 -2.2380207210140922e-06
GC_12_39 b_12 NI_12 NS_39 0 4.5996143851677559e-08
GC_12_40 b_12 NI_12 NS_40 0 -1.2161406282576222e-10
GC_12_41 b_12 NI_12 NS_41 0 6.0706361674066886e-11
GC_12_42 b_12 NI_12 NS_42 0 4.8871298860227436e-11
GC_12_43 b_12 NI_12 NS_43 0 4.0508114602980094e-04
GC_12_44 b_12 NI_12 NS_44 0 -3.9700694111081221e-04
GC_12_45 b_12 NI_12 NS_45 0 -9.8073584801670844e-04
GC_12_46 b_12 NI_12 NS_46 0 -2.0965712521093028e-04
GC_12_47 b_12 NI_12 NS_47 0 4.2795362227107561e-04
GC_12_48 b_12 NI_12 NS_48 0 7.9430098498113610e-04
GC_12_49 b_12 NI_12 NS_49 0 4.2309469671519698e-03
GC_12_50 b_12 NI_12 NS_50 0 -1.1007839912098722e-05
GC_12_51 b_12 NI_12 NS_51 0 9.2772769406623174e-07
GC_12_52 b_12 NI_12 NS_52 0 -2.5047091134673051e-09
GC_12_53 b_12 NI_12 NS_53 0 -1.4960708293035270e-10
GC_12_54 b_12 NI_12 NS_54 0 -4.2478288251200888e-10
GC_12_55 b_12 NI_12 NS_55 0 -3.6268360075236179e-04
GC_12_56 b_12 NI_12 NS_56 0 -1.3120905163259216e-03
GC_12_57 b_12 NI_12 NS_57 0 -1.0797766428347147e-03
GC_12_58 b_12 NI_12 NS_58 0 2.8544842384299121e-03
GC_12_59 b_12 NI_12 NS_59 0 -2.6850808468544029e-03
GC_12_60 b_12 NI_12 NS_60 0 -1.6462183999218507e-03
GC_12_61 b_12 NI_12 NS_61 0 5.0776152607535140e-03
GC_12_62 b_12 NI_12 NS_62 0 -1.8520847216593090e-05
GC_12_63 b_12 NI_12 NS_63 0 7.2952520508934103e-07
GC_12_64 b_12 NI_12 NS_64 0 -1.2333156092250799e-08
GC_12_65 b_12 NI_12 NS_65 0 1.3410093799093430e-10
GC_12_66 b_12 NI_12 NS_66 0 9.6871019425497310e-10
GC_12_67 b_12 NI_12 NS_67 0 9.0818992158010325e-04
GC_12_68 b_12 NI_12 NS_68 0 -1.9384358581965165e-03
GC_12_69 b_12 NI_12 NS_69 0 -4.6723063326488653e-03
GC_12_70 b_12 NI_12 NS_70 0 3.6607765720108893e-04
GC_12_71 b_12 NI_12 NS_71 0 -2.4138258093903899e-03
GC_12_72 b_12 NI_12 NS_72 0 3.0592774769665609e-03
GC_12_73 b_12 NI_12 NS_73 0 1.1241001810519038e-02
GC_12_74 b_12 NI_12 NS_74 0 -3.6207626975921607e-05
GC_12_75 b_12 NI_12 NS_75 0 3.6332029796771953e-06
GC_12_76 b_12 NI_12 NS_76 0 4.0772385705431561e-08
GC_12_77 b_12 NI_12 NS_77 0 -1.2221549402618897e-10
GC_12_78 b_12 NI_12 NS_78 0 2.9775577025116573e-09
GC_12_79 b_12 NI_12 NS_79 0 -2.2254286062978186e-03
GC_12_80 b_12 NI_12 NS_80 0 -4.2732797415504960e-03
GC_12_81 b_12 NI_12 NS_81 0 -2.3606664513179361e-03
GC_12_82 b_12 NI_12 NS_82 0 1.1523697443942086e-02
GC_12_83 b_12 NI_12 NS_83 0 -5.8180349138046428e-03
GC_12_84 b_12 NI_12 NS_84 0 -4.7341176873562279e-03
GC_12_85 b_12 NI_12 NS_85 0 1.8902852114406274e-03
GC_12_86 b_12 NI_12 NS_86 0 -1.9088488299243346e-05
GC_12_87 b_12 NI_12 NS_87 0 -1.3292016220397298e-07
GC_12_88 b_12 NI_12 NS_88 0 -6.8074241105337830e-08
GC_12_89 b_12 NI_12 NS_89 0 9.2132931544731225e-11
GC_12_90 b_12 NI_12 NS_90 0 -2.0426275497232986e-09
GC_12_91 b_12 NI_12 NS_91 0 -1.3991584083402526e-03
GC_12_92 b_12 NI_12 NS_92 0 -2.4217634439044284e-03
GC_12_93 b_12 NI_12 NS_93 0 -4.1847029932853044e-04
GC_12_94 b_12 NI_12 NS_94 0 9.1473296049737632e-04
GC_12_95 b_12 NI_12 NS_95 0 -1.9252501810549810e-03
GC_12_96 b_12 NI_12 NS_96 0 1.7403948149614505e-03
GC_12_97 b_12 NI_12 NS_97 0 7.5502705389232112e-03
GC_12_98 b_12 NI_12 NS_98 0 -2.7274797372550003e-05
GC_12_99 b_12 NI_12 NS_99 0 4.2562823888302908e-06
GC_12_100 b_12 NI_12 NS_100 0 2.4799787114815083e-07
GC_12_101 b_12 NI_12 NS_101 0 7.3566416678481533e-10
GC_12_102 b_12 NI_12 NS_102 0 2.6667003816917208e-08
GC_12_103 b_12 NI_12 NS_103 0 -1.0908210560917992e-03
GC_12_104 b_12 NI_12 NS_104 0 -2.2177893724465050e-03
GC_12_105 b_12 NI_12 NS_105 0 -8.3820905902382416e-04
GC_12_106 b_12 NI_12 NS_106 0 3.4882361911382645e-03
GC_12_107 b_12 NI_12 NS_107 0 -5.7618887277551562e-03
GC_12_108 b_12 NI_12 NS_108 0 -2.7577422718693444e-03
GC_12_109 b_12 NI_12 NS_109 0 4.5219216564554202e-02
GC_12_110 b_12 NI_12 NS_110 0 -2.1057606527240459e-04
GC_12_111 b_12 NI_12 NS_111 0 7.7895297472005539e-08
GC_12_112 b_12 NI_12 NS_112 0 -5.9496955626720143e-07
GC_12_113 b_12 NI_12 NS_113 0 -9.2824714312291551e-10
GC_12_114 b_12 NI_12 NS_114 0 -3.1476532821461844e-08
GC_12_115 b_12 NI_12 NS_115 0 -2.4219205289252789e-02
GC_12_116 b_12 NI_12 NS_116 0 -1.3397004326799588e-02
GC_12_117 b_12 NI_12 NS_117 0 1.4228520026944353e-02
GC_12_118 b_12 NI_12 NS_118 0 1.4700435691786383e-02
GC_12_119 b_12 NI_12 NS_119 0 -4.2169641053312057e-02
GC_12_120 b_12 NI_12 NS_120 0 5.9572275103243512e-03
GC_12_121 b_12 NI_12 NS_121 0 -1.6608617735824427e-01
GC_12_122 b_12 NI_12 NS_122 0 7.7890676686796377e-04
GC_12_123 b_12 NI_12 NS_123 0 -1.0072840362803416e-05
GC_12_124 b_12 NI_12 NS_124 0 4.4062185453954594e-06
GC_12_125 b_12 NI_12 NS_125 0 5.2191194672547786e-09
GC_12_126 b_12 NI_12 NS_126 0 1.7217952677952029e-07
GC_12_127 b_12 NI_12 NS_127 0 -5.0685210612998001e-02
GC_12_128 b_12 NI_12 NS_128 0 -5.0184465999200199e-02
GC_12_129 b_12 NI_12 NS_129 0 -1.8090301563193894e-02
GC_12_130 b_12 NI_12 NS_130 0 -7.4849266062242015e-02
GC_12_131 b_12 NI_12 NS_131 0 1.2151239037284675e-01
GC_12_132 b_12 NI_12 NS_132 0 -5.5027630745757309e-03
GC_12_133 b_12 NI_12 NS_133 0 2.3570671292936693e-01
GC_12_134 b_12 NI_12 NS_134 0 -8.4010550972372575e-04
GC_12_135 b_12 NI_12 NS_135 0 2.7374986306260662e-05
GC_12_136 b_12 NI_12 NS_136 0 -3.2161877407039308e-06
GC_12_137 b_12 NI_12 NS_137 0 -3.6319368781243829e-11
GC_12_138 b_12 NI_12 NS_138 0 -2.0793646988909369e-07
GC_12_139 b_12 NI_12 NS_139 0 -2.8744445536320030e-02
GC_12_140 b_12 NI_12 NS_140 0 1.2390377859696726e-02
GC_12_141 b_12 NI_12 NS_141 0 -1.4922288901497266e-02
GC_12_142 b_12 NI_12 NS_142 0 6.1041345666853937e-02
GC_12_143 b_12 NI_12 NS_143 0 -1.4475758926399171e-01
GC_12_144 b_12 NI_12 NS_144 0 7.1004793766970527e-03
GD_12_1 b_12 NI_12 NA_1 0 1.9132631705418956e-04
GD_12_2 b_12 NI_12 NA_2 0 1.7347950858952109e-04
GD_12_3 b_12 NI_12 NA_3 0 3.6757908454782549e-04
GD_12_4 b_12 NI_12 NA_4 0 4.3421261974659542e-04
GD_12_5 b_12 NI_12 NA_5 0 5.7024688927638791e-06
GD_12_6 b_12 NI_12 NA_6 0 1.8868877216893063e-03
GD_12_7 b_12 NI_12 NA_7 0 -3.4103988353148914e-04
GD_12_8 b_12 NI_12 NA_8 0 6.1933763447625089e-03
GD_12_9 b_12 NI_12 NA_9 0 8.3016615741810017e-05
GD_12_10 b_12 NI_12 NA_10 0 5.1203269514768841e-02
GD_12_11 b_12 NI_12 NA_11 0 1.3127070018746739e-01
GD_12_12 b_12 NI_12 NA_12 0 -4.9038965748758996e-02
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 3.8414975773197675e+00
GS_1_1 0 NS_1 NA_1 0 1.8633417190798034e+00
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 1.1313231168287849e+01
GS_2_1 0 NS_2 NA_1 0 1.8633417190798034e+00
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 2.1781270883655303e+01
GS_3_1 0 NS_3 NA_1 0 1.8633417190798034e+00
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 1.0756159933866989e+02
GS_4_1 0 NS_4 NA_1 0 1.8633417190798034e+00
*
* Real pole n. 5
CS_5 NS_5 0 9.9999999999999998e-13
RS_5 NS_5 0 5.3815059877326075e+03
GS_5_1 0 NS_5 NA_1 0 1.8633417190798034e+00
*
* Real pole n. 6
CS_6 NS_6 0 9.9999999999999998e-13
RS_6 NS_6 0 5.6074140450118989e+02
GS_6_1 0 NS_6 NA_1 0 1.8633417190798034e+00
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 4.2779650153465623e+00
RS_8 NS_8 0 4.2779650153465614e+00
GL_7 0 NS_7 NS_8 0 4.3075440120031583e-01
GL_8 0 NS_8 NS_7 0 -4.3075440120031583e-01
GS_7_1 0 NS_7 NA_1 0 1.8633417190798034e+00
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 3.7856278017814375e+00
RS_10 NS_10 0 3.7856278017814371e+00
GL_9 0 NS_9 NS_10 0 2.4382319655162871e-01
GL_10 0 NS_10 NS_9 0 -2.4382319655162871e-01
GS_9_1 0 NS_9 NA_1 0 1.8633417190798034e+00
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 4.8594901345377242e+00
RS_12 NS_12 0 4.8594901345377242e+00
GL_11 0 NS_11 NS_12 0 4.8770313856068365e-02
GL_12 0 NS_12 NS_11 0 -4.8770313856068365e-02
GS_11_1 0 NS_11 NA_1 0 1.8633417190798034e+00
*
* Real pole n. 13
CS_13 NS_13 0 9.9999999999999998e-13
RS_13 NS_13 0 3.8414975773197675e+00
GS_13_2 0 NS_13 NA_2 0 1.8633417190798034e+00
*
* Real pole n. 14
CS_14 NS_14 0 9.9999999999999998e-13
RS_14 NS_14 0 1.1313231168287849e+01
GS_14_2 0 NS_14 NA_2 0 1.8633417190798034e+00
*
* Real pole n. 15
CS_15 NS_15 0 9.9999999999999998e-13
RS_15 NS_15 0 2.1781270883655303e+01
GS_15_2 0 NS_15 NA_2 0 1.8633417190798034e+00
*
* Real pole n. 16
CS_16 NS_16 0 9.9999999999999998e-13
RS_16 NS_16 0 1.0756159933866989e+02
GS_16_2 0 NS_16 NA_2 0 1.8633417190798034e+00
*
* Real pole n. 17
CS_17 NS_17 0 9.9999999999999998e-13
RS_17 NS_17 0 5.3815059877326075e+03
GS_17_2 0 NS_17 NA_2 0 1.8633417190798034e+00
*
* Real pole n. 18
CS_18 NS_18 0 9.9999999999999998e-13
RS_18 NS_18 0 5.6074140450118989e+02
GS_18_2 0 NS_18 NA_2 0 1.8633417190798034e+00
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 4.2779650153465623e+00
RS_20 NS_20 0 4.2779650153465614e+00
GL_19 0 NS_19 NS_20 0 4.3075440120031583e-01
GL_20 0 NS_20 NS_19 0 -4.3075440120031583e-01
GS_19_2 0 NS_19 NA_2 0 1.8633417190798034e+00
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 3.7856278017814375e+00
RS_22 NS_22 0 3.7856278017814371e+00
GL_21 0 NS_21 NS_22 0 2.4382319655162871e-01
GL_22 0 NS_22 NS_21 0 -2.4382319655162871e-01
GS_21_2 0 NS_21 NA_2 0 1.8633417190798034e+00
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 4.8594901345377242e+00
RS_24 NS_24 0 4.8594901345377242e+00
GL_23 0 NS_23 NS_24 0 4.8770313856068365e-02
GL_24 0 NS_24 NS_23 0 -4.8770313856068365e-02
GS_23_2 0 NS_23 NA_2 0 1.8633417190798034e+00
*
* Real pole n. 25
CS_25 NS_25 0 9.9999999999999998e-13
RS_25 NS_25 0 3.8414975773197675e+00
GS_25_3 0 NS_25 NA_3 0 1.8633417190798034e+00
*
* Real pole n. 26
CS_26 NS_26 0 9.9999999999999998e-13
RS_26 NS_26 0 1.1313231168287849e+01
GS_26_3 0 NS_26 NA_3 0 1.8633417190798034e+00
*
* Real pole n. 27
CS_27 NS_27 0 9.9999999999999998e-13
RS_27 NS_27 0 2.1781270883655303e+01
GS_27_3 0 NS_27 NA_3 0 1.8633417190798034e+00
*
* Real pole n. 28
CS_28 NS_28 0 9.9999999999999998e-13
RS_28 NS_28 0 1.0756159933866989e+02
GS_28_3 0 NS_28 NA_3 0 1.8633417190798034e+00
*
* Real pole n. 29
CS_29 NS_29 0 9.9999999999999998e-13
RS_29 NS_29 0 5.3815059877326075e+03
GS_29_3 0 NS_29 NA_3 0 1.8633417190798034e+00
*
* Real pole n. 30
CS_30 NS_30 0 9.9999999999999998e-13
RS_30 NS_30 0 5.6074140450118989e+02
GS_30_3 0 NS_30 NA_3 0 1.8633417190798034e+00
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 4.2779650153465623e+00
RS_32 NS_32 0 4.2779650153465614e+00
GL_31 0 NS_31 NS_32 0 4.3075440120031583e-01
GL_32 0 NS_32 NS_31 0 -4.3075440120031583e-01
GS_31_3 0 NS_31 NA_3 0 1.8633417190798034e+00
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 3.7856278017814375e+00
RS_34 NS_34 0 3.7856278017814371e+00
GL_33 0 NS_33 NS_34 0 2.4382319655162871e-01
GL_34 0 NS_34 NS_33 0 -2.4382319655162871e-01
GS_33_3 0 NS_33 NA_3 0 1.8633417190798034e+00
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 4.8594901345377242e+00
RS_36 NS_36 0 4.8594901345377242e+00
GL_35 0 NS_35 NS_36 0 4.8770313856068365e-02
GL_36 0 NS_36 NS_35 0 -4.8770313856068365e-02
GS_35_3 0 NS_35 NA_3 0 1.8633417190798034e+00
*
* Real pole n. 37
CS_37 NS_37 0 9.9999999999999998e-13
RS_37 NS_37 0 3.8414975773197675e+00
GS_37_4 0 NS_37 NA_4 0 1.8633417190798034e+00
*
* Real pole n. 38
CS_38 NS_38 0 9.9999999999999998e-13
RS_38 NS_38 0 1.1313231168287849e+01
GS_38_4 0 NS_38 NA_4 0 1.8633417190798034e+00
*
* Real pole n. 39
CS_39 NS_39 0 9.9999999999999998e-13
RS_39 NS_39 0 2.1781270883655303e+01
GS_39_4 0 NS_39 NA_4 0 1.8633417190798034e+00
*
* Real pole n. 40
CS_40 NS_40 0 9.9999999999999998e-13
RS_40 NS_40 0 1.0756159933866989e+02
GS_40_4 0 NS_40 NA_4 0 1.8633417190798034e+00
*
* Real pole n. 41
CS_41 NS_41 0 9.9999999999999998e-13
RS_41 NS_41 0 5.3815059877326075e+03
GS_41_4 0 NS_41 NA_4 0 1.8633417190798034e+00
*
* Real pole n. 42
CS_42 NS_42 0 9.9999999999999998e-13
RS_42 NS_42 0 5.6074140450118989e+02
GS_42_4 0 NS_42 NA_4 0 1.8633417190798034e+00
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 4.2779650153465623e+00
RS_44 NS_44 0 4.2779650153465614e+00
GL_43 0 NS_43 NS_44 0 4.3075440120031583e-01
GL_44 0 NS_44 NS_43 0 -4.3075440120031583e-01
GS_43_4 0 NS_43 NA_4 0 1.8633417190798034e+00
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 3.7856278017814375e+00
RS_46 NS_46 0 3.7856278017814371e+00
GL_45 0 NS_45 NS_46 0 2.4382319655162871e-01
GL_46 0 NS_46 NS_45 0 -2.4382319655162871e-01
GS_45_4 0 NS_45 NA_4 0 1.8633417190798034e+00
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 4.8594901345377242e+00
RS_48 NS_48 0 4.8594901345377242e+00
GL_47 0 NS_47 NS_48 0 4.8770313856068365e-02
GL_48 0 NS_48 NS_47 0 -4.8770313856068365e-02
GS_47_4 0 NS_47 NA_4 0 1.8633417190798034e+00
*
* Real pole n. 49
CS_49 NS_49 0 9.9999999999999998e-13
RS_49 NS_49 0 3.8414975773197675e+00
GS_49_5 0 NS_49 NA_5 0 1.8633417190798034e+00
*
* Real pole n. 50
CS_50 NS_50 0 9.9999999999999998e-13
RS_50 NS_50 0 1.1313231168287849e+01
GS_50_5 0 NS_50 NA_5 0 1.8633417190798034e+00
*
* Real pole n. 51
CS_51 NS_51 0 9.9999999999999998e-13
RS_51 NS_51 0 2.1781270883655303e+01
GS_51_5 0 NS_51 NA_5 0 1.8633417190798034e+00
*
* Real pole n. 52
CS_52 NS_52 0 9.9999999999999998e-13
RS_52 NS_52 0 1.0756159933866989e+02
GS_52_5 0 NS_52 NA_5 0 1.8633417190798034e+00
*
* Real pole n. 53
CS_53 NS_53 0 9.9999999999999998e-13
RS_53 NS_53 0 5.3815059877326075e+03
GS_53_5 0 NS_53 NA_5 0 1.8633417190798034e+00
*
* Real pole n. 54
CS_54 NS_54 0 9.9999999999999998e-13
RS_54 NS_54 0 5.6074140450118989e+02
GS_54_5 0 NS_54 NA_5 0 1.8633417190798034e+00
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 4.2779650153465623e+00
RS_56 NS_56 0 4.2779650153465614e+00
GL_55 0 NS_55 NS_56 0 4.3075440120031583e-01
GL_56 0 NS_56 NS_55 0 -4.3075440120031583e-01
GS_55_5 0 NS_55 NA_5 0 1.8633417190798034e+00
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 3.7856278017814375e+00
RS_58 NS_58 0 3.7856278017814371e+00
GL_57 0 NS_57 NS_58 0 2.4382319655162871e-01
GL_58 0 NS_58 NS_57 0 -2.4382319655162871e-01
GS_57_5 0 NS_57 NA_5 0 1.8633417190798034e+00
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 4.8594901345377242e+00
RS_60 NS_60 0 4.8594901345377242e+00
GL_59 0 NS_59 NS_60 0 4.8770313856068365e-02
GL_60 0 NS_60 NS_59 0 -4.8770313856068365e-02
GS_59_5 0 NS_59 NA_5 0 1.8633417190798034e+00
*
* Real pole n. 61
CS_61 NS_61 0 9.9999999999999998e-13
RS_61 NS_61 0 3.8414975773197675e+00
GS_61_6 0 NS_61 NA_6 0 1.8633417190798034e+00
*
* Real pole n. 62
CS_62 NS_62 0 9.9999999999999998e-13
RS_62 NS_62 0 1.1313231168287849e+01
GS_62_6 0 NS_62 NA_6 0 1.8633417190798034e+00
*
* Real pole n. 63
CS_63 NS_63 0 9.9999999999999998e-13
RS_63 NS_63 0 2.1781270883655303e+01
GS_63_6 0 NS_63 NA_6 0 1.8633417190798034e+00
*
* Real pole n. 64
CS_64 NS_64 0 9.9999999999999998e-13
RS_64 NS_64 0 1.0756159933866989e+02
GS_64_6 0 NS_64 NA_6 0 1.8633417190798034e+00
*
* Real pole n. 65
CS_65 NS_65 0 9.9999999999999998e-13
RS_65 NS_65 0 5.3815059877326075e+03
GS_65_6 0 NS_65 NA_6 0 1.8633417190798034e+00
*
* Real pole n. 66
CS_66 NS_66 0 9.9999999999999998e-13
RS_66 NS_66 0 5.6074140450118989e+02
GS_66_6 0 NS_66 NA_6 0 1.8633417190798034e+00
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 4.2779650153465623e+00
RS_68 NS_68 0 4.2779650153465614e+00
GL_67 0 NS_67 NS_68 0 4.3075440120031583e-01
GL_68 0 NS_68 NS_67 0 -4.3075440120031583e-01
GS_67_6 0 NS_67 NA_6 0 1.8633417190798034e+00
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 3.7856278017814375e+00
RS_70 NS_70 0 3.7856278017814371e+00
GL_69 0 NS_69 NS_70 0 2.4382319655162871e-01
GL_70 0 NS_70 NS_69 0 -2.4382319655162871e-01
GS_69_6 0 NS_69 NA_6 0 1.8633417190798034e+00
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 4.8594901345377242e+00
RS_72 NS_72 0 4.8594901345377242e+00
GL_71 0 NS_71 NS_72 0 4.8770313856068365e-02
GL_72 0 NS_72 NS_71 0 -4.8770313856068365e-02
GS_71_6 0 NS_71 NA_6 0 1.8633417190798034e+00
*
* Real pole n. 73
CS_73 NS_73 0 9.9999999999999998e-13
RS_73 NS_73 0 3.8414975773197675e+00
GS_73_7 0 NS_73 NA_7 0 1.8633417190798034e+00
*
* Real pole n. 74
CS_74 NS_74 0 9.9999999999999998e-13
RS_74 NS_74 0 1.1313231168287849e+01
GS_74_7 0 NS_74 NA_7 0 1.8633417190798034e+00
*
* Real pole n. 75
CS_75 NS_75 0 9.9999999999999998e-13
RS_75 NS_75 0 2.1781270883655303e+01
GS_75_7 0 NS_75 NA_7 0 1.8633417190798034e+00
*
* Real pole n. 76
CS_76 NS_76 0 9.9999999999999998e-13
RS_76 NS_76 0 1.0756159933866989e+02
GS_76_7 0 NS_76 NA_7 0 1.8633417190798034e+00
*
* Real pole n. 77
CS_77 NS_77 0 9.9999999999999998e-13
RS_77 NS_77 0 5.3815059877326075e+03
GS_77_7 0 NS_77 NA_7 0 1.8633417190798034e+00
*
* Real pole n. 78
CS_78 NS_78 0 9.9999999999999998e-13
RS_78 NS_78 0 5.6074140450118989e+02
GS_78_7 0 NS_78 NA_7 0 1.8633417190798034e+00
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 4.2779650153465623e+00
RS_80 NS_80 0 4.2779650153465614e+00
GL_79 0 NS_79 NS_80 0 4.3075440120031583e-01
GL_80 0 NS_80 NS_79 0 -4.3075440120031583e-01
GS_79_7 0 NS_79 NA_7 0 1.8633417190798034e+00
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 3.7856278017814375e+00
RS_82 NS_82 0 3.7856278017814371e+00
GL_81 0 NS_81 NS_82 0 2.4382319655162871e-01
GL_82 0 NS_82 NS_81 0 -2.4382319655162871e-01
GS_81_7 0 NS_81 NA_7 0 1.8633417190798034e+00
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 4.8594901345377242e+00
RS_84 NS_84 0 4.8594901345377242e+00
GL_83 0 NS_83 NS_84 0 4.8770313856068365e-02
GL_84 0 NS_84 NS_83 0 -4.8770313856068365e-02
GS_83_7 0 NS_83 NA_7 0 1.8633417190798034e+00
*
* Real pole n. 85
CS_85 NS_85 0 9.9999999999999998e-13
RS_85 NS_85 0 3.8414975773197675e+00
GS_85_8 0 NS_85 NA_8 0 1.8633417190798034e+00
*
* Real pole n. 86
CS_86 NS_86 0 9.9999999999999998e-13
RS_86 NS_86 0 1.1313231168287849e+01
GS_86_8 0 NS_86 NA_8 0 1.8633417190798034e+00
*
* Real pole n. 87
CS_87 NS_87 0 9.9999999999999998e-13
RS_87 NS_87 0 2.1781270883655303e+01
GS_87_8 0 NS_87 NA_8 0 1.8633417190798034e+00
*
* Real pole n. 88
CS_88 NS_88 0 9.9999999999999998e-13
RS_88 NS_88 0 1.0756159933866989e+02
GS_88_8 0 NS_88 NA_8 0 1.8633417190798034e+00
*
* Real pole n. 89
CS_89 NS_89 0 9.9999999999999998e-13
RS_89 NS_89 0 5.3815059877326075e+03
GS_89_8 0 NS_89 NA_8 0 1.8633417190798034e+00
*
* Real pole n. 90
CS_90 NS_90 0 9.9999999999999998e-13
RS_90 NS_90 0 5.6074140450118989e+02
GS_90_8 0 NS_90 NA_8 0 1.8633417190798034e+00
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 4.2779650153465623e+00
RS_92 NS_92 0 4.2779650153465614e+00
GL_91 0 NS_91 NS_92 0 4.3075440120031583e-01
GL_92 0 NS_92 NS_91 0 -4.3075440120031583e-01
GS_91_8 0 NS_91 NA_8 0 1.8633417190798034e+00
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 3.7856278017814375e+00
RS_94 NS_94 0 3.7856278017814371e+00
GL_93 0 NS_93 NS_94 0 2.4382319655162871e-01
GL_94 0 NS_94 NS_93 0 -2.4382319655162871e-01
GS_93_8 0 NS_93 NA_8 0 1.8633417190798034e+00
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 4.8594901345377242e+00
RS_96 NS_96 0 4.8594901345377242e+00
GL_95 0 NS_95 NS_96 0 4.8770313856068365e-02
GL_96 0 NS_96 NS_95 0 -4.8770313856068365e-02
GS_95_8 0 NS_95 NA_8 0 1.8633417190798034e+00
*
* Real pole n. 97
CS_97 NS_97 0 9.9999999999999998e-13
RS_97 NS_97 0 3.8414975773197675e+00
GS_97_9 0 NS_97 NA_9 0 1.8633417190798034e+00
*
* Real pole n. 98
CS_98 NS_98 0 9.9999999999999998e-13
RS_98 NS_98 0 1.1313231168287849e+01
GS_98_9 0 NS_98 NA_9 0 1.8633417190798034e+00
*
* Real pole n. 99
CS_99 NS_99 0 9.9999999999999998e-13
RS_99 NS_99 0 2.1781270883655303e+01
GS_99_9 0 NS_99 NA_9 0 1.8633417190798034e+00
*
* Real pole n. 100
CS_100 NS_100 0 9.9999999999999998e-13
RS_100 NS_100 0 1.0756159933866989e+02
GS_100_9 0 NS_100 NA_9 0 1.8633417190798034e+00
*
* Real pole n. 101
CS_101 NS_101 0 9.9999999999999998e-13
RS_101 NS_101 0 5.3815059877326075e+03
GS_101_9 0 NS_101 NA_9 0 1.8633417190798034e+00
*
* Real pole n. 102
CS_102 NS_102 0 9.9999999999999998e-13
RS_102 NS_102 0 5.6074140450118989e+02
GS_102_9 0 NS_102 NA_9 0 1.8633417190798034e+00
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 4.2779650153465623e+00
RS_104 NS_104 0 4.2779650153465614e+00
GL_103 0 NS_103 NS_104 0 4.3075440120031583e-01
GL_104 0 NS_104 NS_103 0 -4.3075440120031583e-01
GS_103_9 0 NS_103 NA_9 0 1.8633417190798034e+00
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 3.7856278017814375e+00
RS_106 NS_106 0 3.7856278017814371e+00
GL_105 0 NS_105 NS_106 0 2.4382319655162871e-01
GL_106 0 NS_106 NS_105 0 -2.4382319655162871e-01
GS_105_9 0 NS_105 NA_9 0 1.8633417190798034e+00
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 4.8594901345377242e+00
RS_108 NS_108 0 4.8594901345377242e+00
GL_107 0 NS_107 NS_108 0 4.8770313856068365e-02
GL_108 0 NS_108 NS_107 0 -4.8770313856068365e-02
GS_107_9 0 NS_107 NA_9 0 1.8633417190798034e+00
*
* Real pole n. 109
CS_109 NS_109 0 9.9999999999999998e-13
RS_109 NS_109 0 3.8414975773197675e+00
GS_109_10 0 NS_109 NA_10 0 1.8633417190798034e+00
*
* Real pole n. 110
CS_110 NS_110 0 9.9999999999999998e-13
RS_110 NS_110 0 1.1313231168287849e+01
GS_110_10 0 NS_110 NA_10 0 1.8633417190798034e+00
*
* Real pole n. 111
CS_111 NS_111 0 9.9999999999999998e-13
RS_111 NS_111 0 2.1781270883655303e+01
GS_111_10 0 NS_111 NA_10 0 1.8633417190798034e+00
*
* Real pole n. 112
CS_112 NS_112 0 9.9999999999999998e-13
RS_112 NS_112 0 1.0756159933866989e+02
GS_112_10 0 NS_112 NA_10 0 1.8633417190798034e+00
*
* Real pole n. 113
CS_113 NS_113 0 9.9999999999999998e-13
RS_113 NS_113 0 5.3815059877326075e+03
GS_113_10 0 NS_113 NA_10 0 1.8633417190798034e+00
*
* Real pole n. 114
CS_114 NS_114 0 9.9999999999999998e-13
RS_114 NS_114 0 5.6074140450118989e+02
GS_114_10 0 NS_114 NA_10 0 1.8633417190798034e+00
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 4.2779650153465623e+00
RS_116 NS_116 0 4.2779650153465614e+00
GL_115 0 NS_115 NS_116 0 4.3075440120031583e-01
GL_116 0 NS_116 NS_115 0 -4.3075440120031583e-01
GS_115_10 0 NS_115 NA_10 0 1.8633417190798034e+00
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 3.7856278017814375e+00
RS_118 NS_118 0 3.7856278017814371e+00
GL_117 0 NS_117 NS_118 0 2.4382319655162871e-01
GL_118 0 NS_118 NS_117 0 -2.4382319655162871e-01
GS_117_10 0 NS_117 NA_10 0 1.8633417190798034e+00
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 4.8594901345377242e+00
RS_120 NS_120 0 4.8594901345377242e+00
GL_119 0 NS_119 NS_120 0 4.8770313856068365e-02
GL_120 0 NS_120 NS_119 0 -4.8770313856068365e-02
GS_119_10 0 NS_119 NA_10 0 1.8633417190798034e+00
*
* Real pole n. 121
CS_121 NS_121 0 9.9999999999999998e-13
RS_121 NS_121 0 3.8414975773197675e+00
GS_121_11 0 NS_121 NA_11 0 1.8633417190798034e+00
*
* Real pole n. 122
CS_122 NS_122 0 9.9999999999999998e-13
RS_122 NS_122 0 1.1313231168287849e+01
GS_122_11 0 NS_122 NA_11 0 1.8633417190798034e+00
*
* Real pole n. 123
CS_123 NS_123 0 9.9999999999999998e-13
RS_123 NS_123 0 2.1781270883655303e+01
GS_123_11 0 NS_123 NA_11 0 1.8633417190798034e+00
*
* Real pole n. 124
CS_124 NS_124 0 9.9999999999999998e-13
RS_124 NS_124 0 1.0756159933866989e+02
GS_124_11 0 NS_124 NA_11 0 1.8633417190798034e+00
*
* Real pole n. 125
CS_125 NS_125 0 9.9999999999999998e-13
RS_125 NS_125 0 5.3815059877326075e+03
GS_125_11 0 NS_125 NA_11 0 1.8633417190798034e+00
*
* Real pole n. 126
CS_126 NS_126 0 9.9999999999999998e-13
RS_126 NS_126 0 5.6074140450118989e+02
GS_126_11 0 NS_126 NA_11 0 1.8633417190798034e+00
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 4.2779650153465623e+00
RS_128 NS_128 0 4.2779650153465614e+00
GL_127 0 NS_127 NS_128 0 4.3075440120031583e-01
GL_128 0 NS_128 NS_127 0 -4.3075440120031583e-01
GS_127_11 0 NS_127 NA_11 0 1.8633417190798034e+00
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 3.7856278017814375e+00
RS_130 NS_130 0 3.7856278017814371e+00
GL_129 0 NS_129 NS_130 0 2.4382319655162871e-01
GL_130 0 NS_130 NS_129 0 -2.4382319655162871e-01
GS_129_11 0 NS_129 NA_11 0 1.8633417190798034e+00
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 4.8594901345377242e+00
RS_132 NS_132 0 4.8594901345377242e+00
GL_131 0 NS_131 NS_132 0 4.8770313856068365e-02
GL_132 0 NS_132 NS_131 0 -4.8770313856068365e-02
GS_131_11 0 NS_131 NA_11 0 1.8633417190798034e+00
*
* Real pole n. 133
CS_133 NS_133 0 9.9999999999999998e-13
RS_133 NS_133 0 3.8414975773197675e+00
GS_133_12 0 NS_133 NA_12 0 1.8633417190798034e+00
*
* Real pole n. 134
CS_134 NS_134 0 9.9999999999999998e-13
RS_134 NS_134 0 1.1313231168287849e+01
GS_134_12 0 NS_134 NA_12 0 1.8633417190798034e+00
*
* Real pole n. 135
CS_135 NS_135 0 9.9999999999999998e-13
RS_135 NS_135 0 2.1781270883655303e+01
GS_135_12 0 NS_135 NA_12 0 1.8633417190798034e+00
*
* Real pole n. 136
CS_136 NS_136 0 9.9999999999999998e-13
RS_136 NS_136 0 1.0756159933866989e+02
GS_136_12 0 NS_136 NA_12 0 1.8633417190798034e+00
*
* Real pole n. 137
CS_137 NS_137 0 9.9999999999999998e-13
RS_137 NS_137 0 5.3815059877326075e+03
GS_137_12 0 NS_137 NA_12 0 1.8633417190798034e+00
*
* Real pole n. 138
CS_138 NS_138 0 9.9999999999999998e-13
RS_138 NS_138 0 5.6074140450118989e+02
GS_138_12 0 NS_138 NA_12 0 1.8633417190798034e+00
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 4.2779650153465623e+00
RS_140 NS_140 0 4.2779650153465614e+00
GL_139 0 NS_139 NS_140 0 4.3075440120031583e-01
GL_140 0 NS_140 NS_139 0 -4.3075440120031583e-01
GS_139_12 0 NS_139 NA_12 0 1.8633417190798034e+00
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 3.7856278017814375e+00
RS_142 NS_142 0 3.7856278017814371e+00
GL_141 0 NS_141 NS_142 0 2.4382319655162871e-01
GL_142 0 NS_142 NS_141 0 -2.4382319655162871e-01
GS_141_12 0 NS_141 NA_12 0 1.8633417190798034e+00
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 4.8594901345377242e+00
RS_144 NS_144 0 4.8594901345377242e+00
GL_143 0 NS_143 NS_144 0 4.8770313856068365e-02
GL_144 0 NS_144 NS_143 0 -4.8770313856068365e-02
GS_143_12 0 NS_143 NA_12 0 1.8633417190798034e+00
*
******************************


.ends
*******************
* End of subcircuit
*******************
