**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [2 2 10] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** n/a - passivity was not enforced
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_4_C4escape_1mm_highloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 5.2859301621601310e-02
GC_1_2 b_1 NI_1 NS_2 0 -1.3064761545831007e-02
GC_1_3 b_1 NI_1 NS_3 0 5.9279803764012493e-05
GC_1_4 b_1 NI_1 NS_4 0 -1.3381678614826348e-05
GC_1_5 b_1 NI_1 NS_5 0 -8.5088506889302727e-09
GC_1_6 b_1 NI_1 NS_6 0 -1.3098057513172002e-06
GC_1_7 b_1 NI_1 NS_7 0 -1.9013504529624933e-03
GC_1_8 b_1 NI_1 NS_8 0 4.2717664707473306e-03
GC_1_9 b_1 NI_1 NS_9 0 -1.3200522438650462e-02
GC_1_10 b_1 NI_1 NS_10 0 2.3506099807481265e-02
GC_1_11 b_1 NI_1 NS_11 0 -1.7979744716375870e-01
GC_1_12 b_1 NI_1 NS_12 0 5.6387268071270834e-02
GC_1_13 b_1 NI_1 NS_13 0 -2.6203527603905889e-04
GC_1_14 b_1 NI_1 NS_14 0 8.7772980712331344e-05
GC_1_15 b_1 NI_1 NS_15 0 6.1883623643798174e-08
GC_1_16 b_1 NI_1 NS_16 0 6.3236589811054525e-08
GC_1_17 b_1 NI_1 NS_17 0 -3.2557534419983103e-02
GC_1_18 b_1 NI_1 NS_18 0 -6.1488507846060435e-02
GC_1_19 b_1 NI_1 NS_19 0 8.4503795400059825e-02
GC_1_20 b_1 NI_1 NS_20 0 -1.0099190995628843e-01
GC_1_21 b_1 NI_1 NS_21 0 -7.0303330590827115e-03
GC_1_22 b_1 NI_1 NS_22 0 -4.4850017400638060e-03
GC_1_23 b_1 NI_1 NS_23 0 -1.6071362626906194e-05
GC_1_24 b_1 NI_1 NS_24 0 -2.4812561109900059e-06
GC_1_25 b_1 NI_1 NS_25 0 -2.2962509480293271e-09
GC_1_26 b_1 NI_1 NS_26 0 -3.9507715081732348e-07
GC_1_27 b_1 NI_1 NS_27 0 1.7173864573176683e-03
GC_1_28 b_1 NI_1 NS_28 0 -1.3398639507239605e-02
GC_1_29 b_1 NI_1 NS_29 0 5.8796835844652567e-03
GC_1_30 b_1 NI_1 NS_30 0 1.3002224138356774e-02
GC_1_31 b_1 NI_1 NS_31 0 -1.3075307274922842e-03
GC_1_32 b_1 NI_1 NS_32 0 1.1612753497448833e-03
GC_1_33 b_1 NI_1 NS_33 0 -5.2062560447287294e-06
GC_1_34 b_1 NI_1 NS_34 0 -1.3604705060372988e-07
GC_1_35 b_1 NI_1 NS_35 0 1.8849443440605641e-09
GC_1_36 b_1 NI_1 NS_36 0 1.0944625790218953e-07
GC_1_37 b_1 NI_1 NS_37 0 2.1791749868034795e-03
GC_1_38 b_1 NI_1 NS_38 0 -5.3352870929134898e-04
GC_1_39 b_1 NI_1 NS_39 0 -2.6656372835813101e-03
GC_1_40 b_1 NI_1 NS_40 0 -1.2467026618913151e-03
GC_1_41 b_1 NI_1 NS_41 0 -2.7882340457254899e-03
GC_1_42 b_1 NI_1 NS_42 0 -5.7603257060246760e-04
GC_1_43 b_1 NI_1 NS_43 0 -2.2832322525186888e-06
GC_1_44 b_1 NI_1 NS_44 0 5.2509674129389776e-08
GC_1_45 b_1 NI_1 NS_45 0 1.0694927813137638e-10
GC_1_46 b_1 NI_1 NS_46 0 -3.1757470645053139e-08
GC_1_47 b_1 NI_1 NS_47 0 5.7218330748787141e-04
GC_1_48 b_1 NI_1 NS_48 0 -1.1815750180375708e-03
GC_1_49 b_1 NI_1 NS_49 0 2.0454127164122879e-03
GC_1_50 b_1 NI_1 NS_50 0 -7.0599483380387278e-05
GC_1_51 b_1 NI_1 NS_51 0 4.4879461587188715e-04
GC_1_52 b_1 NI_1 NS_52 0 1.7423941774537904e-03
GC_1_53 b_1 NI_1 NS_53 0 2.5851612781879403e-06
GC_1_54 b_1 NI_1 NS_54 0 6.8465792549908691e-08
GC_1_55 b_1 NI_1 NS_55 0 -1.1309071083045831e-10
GC_1_56 b_1 NI_1 NS_56 0 2.8407691385166663e-08
GC_1_57 b_1 NI_1 NS_57 0 3.2315056701227090e-03
GC_1_58 b_1 NI_1 NS_58 0 -2.7458384256641893e-04
GC_1_59 b_1 NI_1 NS_59 0 -5.7928527581335354e-03
GC_1_60 b_1 NI_1 NS_60 0 -1.0206293933180512e-03
GC_1_61 b_1 NI_1 NS_61 0 -1.8083805680269159e-03
GC_1_62 b_1 NI_1 NS_62 0 -4.2589675325296254e-04
GC_1_63 b_1 NI_1 NS_63 0 -1.7713896485539640e-06
GC_1_64 b_1 NI_1 NS_64 0 2.3182273074637414e-07
GC_1_65 b_1 NI_1 NS_65 0 2.3510236112728134e-10
GC_1_66 b_1 NI_1 NS_66 0 -4.8108770705629611e-09
GC_1_67 b_1 NI_1 NS_67 0 3.9570368448633568e-04
GC_1_68 b_1 NI_1 NS_68 0 4.5789574721321875e-04
GC_1_69 b_1 NI_1 NS_69 0 1.7011466517145200e-03
GC_1_70 b_1 NI_1 NS_70 0 -1.8054253450967015e-03
GC_1_71 b_1 NI_1 NS_71 0 1.7726806265213851e-04
GC_1_72 b_1 NI_1 NS_72 0 5.7708080829966266e-04
GC_1_73 b_1 NI_1 NS_73 0 3.8452142880391208e-07
GC_1_74 b_1 NI_1 NS_74 0 5.5176060545675808e-09
GC_1_75 b_1 NI_1 NS_75 0 -2.1149653085821725e-10
GC_1_76 b_1 NI_1 NS_76 0 1.1310143202669461e-09
GC_1_77 b_1 NI_1 NS_77 0 5.7502414607187187e-04
GC_1_78 b_1 NI_1 NS_78 0 7.6086239297994577e-05
GC_1_79 b_1 NI_1 NS_79 0 -1.1522858676960759e-03
GC_1_80 b_1 NI_1 NS_80 0 2.9496670632460673e-04
GC_1_81 b_1 NI_1 NS_81 0 -1.5078854548084765e-04
GC_1_82 b_1 NI_1 NS_82 0 -2.5231272645266737e-04
GC_1_83 b_1 NI_1 NS_83 0 -3.1462006780480187e-07
GC_1_84 b_1 NI_1 NS_84 0 4.4620488362912420e-08
GC_1_85 b_1 NI_1 NS_85 0 1.0763234468196428e-10
GC_1_86 b_1 NI_1 NS_86 0 5.2939954377662918e-11
GC_1_87 b_1 NI_1 NS_87 0 8.6961757586850603e-05
GC_1_88 b_1 NI_1 NS_88 0 1.6484274725236408e-04
GC_1_89 b_1 NI_1 NS_89 0 3.1650314601421183e-04
GC_1_90 b_1 NI_1 NS_90 0 -5.7170825778301215e-04
GC_1_91 b_1 NI_1 NS_91 0 -6.8110663934043062e-05
GC_1_92 b_1 NI_1 NS_92 0 3.4263860861849440e-04
GC_1_93 b_1 NI_1 NS_93 0 -2.0423855983249287e-08
GC_1_94 b_1 NI_1 NS_94 0 1.4259177777872977e-08
GC_1_95 b_1 NI_1 NS_95 0 -1.0175926760562784e-10
GC_1_96 b_1 NI_1 NS_96 0 -9.1086072048921074e-10
GC_1_97 b_1 NI_1 NS_97 0 -5.6814754007499051e-05
GC_1_98 b_1 NI_1 NS_98 0 1.2051224837869429e-04
GC_1_99 b_1 NI_1 NS_99 0 2.1893798623872612e-05
GC_1_100 b_1 NI_1 NS_100 0 5.8520957279704835e-04
GC_1_101 b_1 NI_1 NS_101 0 2.9950568709309313e-04
GC_1_102 b_1 NI_1 NS_102 0 -1.6297487896081727e-04
GC_1_103 b_1 NI_1 NS_103 0 3.2148093910201142e-08
GC_1_104 b_1 NI_1 NS_104 0 -1.0198415394417565e-08
GC_1_105 b_1 NI_1 NS_105 0 3.8755172796953024e-11
GC_1_106 b_1 NI_1 NS_106 0 9.2512210389744349e-10
GC_1_107 b_1 NI_1 NS_107 0 -2.7773871197578423e-06
GC_1_108 b_1 NI_1 NS_108 0 1.7958982134132495e-05
GC_1_109 b_1 NI_1 NS_109 0 -1.1314384074756495e-04
GC_1_110 b_1 NI_1 NS_110 0 -1.0759340696470801e-04
GC_1_111 b_1 NI_1 NS_111 0 -9.7220809498346766e-05
GC_1_112 b_1 NI_1 NS_112 0 1.3616955559621417e-04
GC_1_113 b_1 NI_1 NS_113 0 -8.0289895940418349e-09
GC_1_114 b_1 NI_1 NS_114 0 8.0786405512087354e-09
GC_1_115 b_1 NI_1 NS_115 0 -3.8739547827781783e-11
GC_1_116 b_1 NI_1 NS_116 0 -8.7101973761499855e-10
GC_1_117 b_1 NI_1 NS_117 0 -4.7013291556070843e-05
GC_1_118 b_1 NI_1 NS_118 0 4.5272529151951507e-05
GC_1_119 b_1 NI_1 NS_119 0 8.8826450853963002e-05
GC_1_120 b_1 NI_1 NS_120 0 2.2568047343720499e-04
GD_1_1 b_1 NI_1 NA_1 0 -1.3863812267786419e-02
GD_1_2 b_1 NI_1 NA_2 0 1.9655245108939828e-02
GD_1_3 b_1 NI_1 NA_3 0 3.1099222062001709e-02
GD_1_4 b_1 NI_1 NA_4 0 3.7223665651837500e-04
GD_1_5 b_1 NI_1 NA_5 0 3.8585855893856912e-03
GD_1_6 b_1 NI_1 NA_6 0 2.3520227332051908e-04
GD_1_7 b_1 NI_1 NA_7 0 4.3463287813285756e-04
GD_1_8 b_1 NI_1 NA_8 0 -1.3166542884561320e-04
GD_1_9 b_1 NI_1 NA_9 0 3.9136900122655807e-05
GD_1_10 b_1 NI_1 NA_10 0 -1.6522435545847635e-04
GD_1_11 b_1 NI_1 NA_11 0 -1.5547960944828617e-06
GD_1_12 b_1 NI_1 NA_12 0 -5.5599313327973641e-05
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 -1.7980244990755068e-01
GC_2_2 b_2 NI_2 NS_2 0 5.6388736466444656e-02
GC_2_3 b_2 NI_2 NS_3 0 -2.6204708171640540e-04
GC_2_4 b_2 NI_2 NS_4 0 8.7776591566488985e-05
GC_2_5 b_2 NI_2 NS_5 0 6.1886780823697295e-08
GC_2_6 b_2 NI_2 NS_6 0 6.3073454044695431e-08
GC_2_7 b_2 NI_2 NS_7 0 -3.2559836401256544e-02
GC_2_8 b_2 NI_2 NS_8 0 -6.1491335348565879e-02
GC_2_9 b_2 NI_2 NS_9 0 8.4505078097955946e-02
GC_2_10 b_2 NI_2 NS_10 0 -1.0099134515478536e-01
GC_2_11 b_2 NI_2 NS_11 0 5.2859301621601310e-02
GC_2_12 b_2 NI_2 NS_12 0 -1.3064761545831007e-02
GC_2_13 b_2 NI_2 NS_13 0 5.9279803764012493e-05
GC_2_14 b_2 NI_2 NS_14 0 -1.3381678614826348e-05
GC_2_15 b_2 NI_2 NS_15 0 -8.5088506889302727e-09
GC_2_16 b_2 NI_2 NS_16 0 -1.3098057513172002e-06
GC_2_17 b_2 NI_2 NS_17 0 -1.9013504529624933e-03
GC_2_18 b_2 NI_2 NS_18 0 4.2717664707473306e-03
GC_2_19 b_2 NI_2 NS_19 0 -1.3200522438650462e-02
GC_2_20 b_2 NI_2 NS_20 0 2.3506099807481265e-02
GC_2_21 b_2 NI_2 NS_21 0 -1.3064076650635922e-03
GC_2_22 b_2 NI_2 NS_22 0 1.1609671570068636e-03
GC_2_23 b_2 NI_2 NS_23 0 -5.2046701074105827e-06
GC_2_24 b_2 NI_2 NS_24 0 -1.3622416252452102e-07
GC_2_25 b_2 NI_2 NS_25 0 1.8849506907402238e-09
GC_2_26 b_2 NI_2 NS_26 0 1.0944781804581485e-07
GC_2_27 b_2 NI_2 NS_27 0 2.1789912091479606e-03
GC_2_28 b_2 NI_2 NS_28 0 -5.3354771307407233e-04
GC_2_29 b_2 NI_2 NS_29 0 -2.6661110234395880e-03
GC_2_30 b_2 NI_2 NS_30 0 -1.2464190329196801e-03
GC_2_31 b_2 NI_2 NS_31 0 -7.0548319716035521e-03
GC_2_32 b_2 NI_2 NS_32 0 -4.4830559052310833e-03
GC_2_33 b_2 NI_2 NS_33 0 -1.6084432710801727e-05
GC_2_34 b_2 NI_2 NS_34 0 -2.4819199509575522e-06
GC_2_35 b_2 NI_2 NS_35 0 -2.2944151022451606e-09
GC_2_36 b_2 NI_2 NS_36 0 -3.9506216110263826e-07
GC_2_37 b_2 NI_2 NS_37 0 1.7171964151413931e-03
GC_2_38 b_2 NI_2 NS_38 0 -1.3406034021209086e-02
GC_2_39 b_2 NI_2 NS_39 0 5.8860653819341538e-03
GC_2_40 b_2 NI_2 NS_40 0 1.2986713716173895e-02
GC_2_41 b_2 NI_2 NS_41 0 4.4221077296529839e-04
GC_2_42 b_2 NI_2 NS_42 0 1.7436489372742686e-03
GC_2_43 b_2 NI_2 NS_43 0 2.5868934374718469e-06
GC_2_44 b_2 NI_2 NS_44 0 6.8132163790513363e-08
GC_2_45 b_2 NI_2 NS_45 0 -1.1317491206945763e-10
GC_2_46 b_2 NI_2 NS_46 0 2.8413703378657205e-08
GC_2_47 b_2 NI_2 NS_47 0 3.2308596094018337e-03
GC_2_48 b_2 NI_2 NS_48 0 -2.7670604659806134e-04
GC_2_49 b_2 NI_2 NS_49 0 -5.7911556532728430e-03
GC_2_50 b_2 NI_2 NS_50 0 -1.0224888052617921e-03
GC_2_51 b_2 NI_2 NS_51 0 -2.7969920567862752e-03
GC_2_52 b_2 NI_2 NS_52 0 -5.7452506927769273e-04
GC_2_53 b_2 NI_2 NS_53 0 -2.2977364695200834e-06
GC_2_54 b_2 NI_2 NS_54 0 5.4639600786713524e-08
GC_2_55 b_2 NI_2 NS_55 0 1.0754501521530430e-10
GC_2_56 b_2 NI_2 NS_56 0 -3.1810271387062057e-08
GC_2_57 b_2 NI_2 NS_57 0 5.7236763104545954e-04
GC_2_58 b_2 NI_2 NS_58 0 -1.1831822711651785e-03
GC_2_59 b_2 NI_2 NS_59 0 2.0484023784160615e-03
GC_2_60 b_2 NI_2 NS_60 0 -7.4431985879680877e-05
GC_2_61 b_2 NI_2 NS_61 0 1.7512171572988327e-04
GC_2_62 b_2 NI_2 NS_62 0 5.7758963987158138e-04
GC_2_63 b_2 NI_2 NS_63 0 3.8256035183627728e-07
GC_2_64 b_2 NI_2 NS_64 0 5.8909093128057647e-09
GC_2_65 b_2 NI_2 NS_65 0 -2.1145808913900906e-10
GC_2_66 b_2 NI_2 NS_66 0 1.1273506148340423e-09
GC_2_67 b_2 NI_2 NS_67 0 5.7479252341689562e-04
GC_2_68 b_2 NI_2 NS_68 0 7.5485693406342991e-05
GC_2_69 b_2 NI_2 NS_69 0 -1.1516162709818746e-03
GC_2_70 b_2 NI_2 NS_70 0 2.9456704838688692e-04
GC_2_71 b_2 NI_2 NS_71 0 -1.8103086080908442e-03
GC_2_72 b_2 NI_2 NS_72 0 -4.2554411892932811e-04
GC_2_73 b_2 NI_2 NS_73 0 -1.7770576628909205e-06
GC_2_74 b_2 NI_2 NS_74 0 2.3274736994592285e-07
GC_2_75 b_2 NI_2 NS_75 0 2.3522415508806004e-10
GC_2_76 b_2 NI_2 NS_76 0 -4.8289272699913976e-09
GC_2_77 b_2 NI_2 NS_77 0 3.9578755176589793e-04
GC_2_78 b_2 NI_2 NS_78 0 4.5729849441930533e-04
GC_2_79 b_2 NI_2 NS_79 0 1.7014914530512301e-03
GC_2_80 b_2 NI_2 NS_80 0 -1.8063081690673948e-03
GC_2_81 b_2 NI_2 NS_81 0 -6.8799613938542152e-05
GC_2_82 b_2 NI_2 NS_82 0 3.4277166450000614e-04
GC_2_83 b_2 NI_2 NS_83 0 -2.0714519939758428e-08
GC_2_84 b_2 NI_2 NS_84 0 1.4344062583856994e-08
GC_2_85 b_2 NI_2 NS_85 0 -1.0174748616111340e-10
GC_2_86 b_2 NI_2 NS_86 0 -9.1239918190250832e-10
GC_2_87 b_2 NI_2 NS_87 0 -5.6845011500187794e-05
GC_2_88 b_2 NI_2 NS_88 0 1.2033342580408023e-04
GC_2_89 b_2 NI_2 NS_89 0 2.2093533547946310e-05
GC_2_90 b_2 NI_2 NS_90 0 5.8499452995802725e-04
GC_2_91 b_2 NI_2 NS_91 0 -1.5096395792225386e-04
GC_2_92 b_2 NI_2 NS_92 0 -2.5228975229088128e-04
GC_2_93 b_2 NI_2 NS_93 0 -3.1553261516787772e-07
GC_2_94 b_2 NI_2 NS_94 0 4.4725458220605296e-08
GC_2_95 b_2 NI_2 NS_95 0 1.0764361019824762e-10
GC_2_96 b_2 NI_2 NS_96 0 5.1109993696245445e-11
GC_2_97 b_2 NI_2 NS_97 0 8.6978354446912569e-05
GC_2_98 b_2 NI_2 NS_98 0 1.6471009113755645e-04
GC_2_99 b_2 NI_2 NS_99 0 3.1642735768477100e-04
GC_2_100 b_2 NI_2 NS_100 0 -5.7184015220568447e-04
GC_2_101 b_2 NI_2 NS_101 0 -9.7681611493678598e-05
GC_2_102 b_2 NI_2 NS_102 0 1.3625652411588271e-04
GC_2_103 b_2 NI_2 NS_103 0 -8.2304077755972315e-09
GC_2_104 b_2 NI_2 NS_104 0 8.1286055351795112e-09
GC_2_105 b_2 NI_2 NS_105 0 -3.8731874586279440e-11
GC_2_106 b_2 NI_2 NS_106 0 -8.7182408139556192e-10
GC_2_107 b_2 NI_2 NS_107 0 -4.6992204407757525e-05
GC_2_108 b_2 NI_2 NS_108 0 4.5214859426022167e-05
GC_2_109 b_2 NI_2 NS_109 0 8.8993848083572329e-05
GC_2_110 b_2 NI_2 NS_110 0 2.2551044614933105e-04
GC_2_111 b_2 NI_2 NS_111 0 2.9949897747088552e-04
GC_2_112 b_2 NI_2 NS_112 0 -1.6297325967750130e-04
GC_2_113 b_2 NI_2 NS_113 0 3.2141973059138642e-08
GC_2_114 b_2 NI_2 NS_114 0 -1.0197462899819804e-08
GC_2_115 b_2 NI_2 NS_115 0 3.8755308880426955e-11
GC_2_116 b_2 NI_2 NS_116 0 9.2510731016750194e-10
GC_2_117 b_2 NI_2 NS_117 0 -2.7765464681837651e-06
GC_2_118 b_2 NI_2 NS_118 0 1.7958537920894944e-05
GC_2_119 b_2 NI_2 NS_119 0 -1.1314121306781161e-04
GC_2_120 b_2 NI_2 NS_120 0 -1.0759536368278283e-04
GD_2_1 b_2 NI_2 NA_1 0 1.9658445259010188e-02
GD_2_2 b_2 NI_2 NA_2 0 -1.3863812267786419e-02
GD_2_3 b_2 NI_2 NA_3 0 3.7211526732520192e-04
GD_2_4 b_2 NI_2 NA_4 0 3.1107304579876829e-02
GD_2_5 b_2 NI_2 NA_5 0 2.3853587052750537e-04
GD_2_6 b_2 NI_2 NA_6 0 3.8606050553713798e-03
GD_2_7 b_2 NI_2 NA_7 0 -1.3079564415693494e-04
GD_2_8 b_2 NI_2 NA_8 0 4.3529775617166675e-04
GD_2_9 b_2 NI_2 NA_9 0 -1.6493460942386661e-04
GD_2_10 b_2 NI_2 NA_10 0 3.9293699158599537e-05
GD_2_11 b_2 NI_2 NA_11 0 -5.5459114778578140e-05
GD_2_12 b_2 NI_2 NA_12 0 -1.5538174042610196e-06
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 -7.0548319716035521e-03
GC_3_2 b_3 NI_3 NS_2 0 -4.4830559052310833e-03
GC_3_3 b_3 NI_3 NS_3 0 -1.6084432710801727e-05
GC_3_4 b_3 NI_3 NS_4 0 -2.4819199509575522e-06
GC_3_5 b_3 NI_3 NS_5 0 -2.2944151022451606e-09
GC_3_6 b_3 NI_3 NS_6 0 -3.9506216110263826e-07
GC_3_7 b_3 NI_3 NS_7 0 1.7171964151413931e-03
GC_3_8 b_3 NI_3 NS_8 0 -1.3406034021209086e-02
GC_3_9 b_3 NI_3 NS_9 0 5.8860653819341538e-03
GC_3_10 b_3 NI_3 NS_10 0 1.2986713716173895e-02
GC_3_11 b_3 NI_3 NS_11 0 -1.3075307274922842e-03
GC_3_12 b_3 NI_3 NS_12 0 1.1612753497448833e-03
GC_3_13 b_3 NI_3 NS_13 0 -5.2062560447287294e-06
GC_3_14 b_3 NI_3 NS_14 0 -1.3604705060372988e-07
GC_3_15 b_3 NI_3 NS_15 0 1.8849443440605641e-09
GC_3_16 b_3 NI_3 NS_16 0 1.0944625790218953e-07
GC_3_17 b_3 NI_3 NS_17 0 2.1791749868034795e-03
GC_3_18 b_3 NI_3 NS_18 0 -5.3352870929134898e-04
GC_3_19 b_3 NI_3 NS_19 0 -2.6656372835813101e-03
GC_3_20 b_3 NI_3 NS_20 0 -1.2467026618913151e-03
GC_3_21 b_3 NI_3 NS_21 0 5.3616779120527064e-02
GC_3_22 b_3 NI_3 NS_22 0 -1.2804945067003930e-02
GC_3_23 b_3 NI_3 NS_23 0 6.3940087657096697e-05
GC_3_24 b_3 NI_3 NS_24 0 -1.3871599455596756e-05
GC_3_25 b_3 NI_3 NS_25 0 -1.0851117673452737e-08
GC_3_26 b_3 NI_3 NS_26 0 -1.2971657354454211e-06
GC_3_27 b_3 NI_3 NS_27 0 -1.9507878599407341e-03
GC_3_28 b_3 NI_3 NS_28 0 7.0862888731600430e-03
GC_3_29 b_3 NI_3 NS_29 0 -1.3281287280820304e-02
GC_3_30 b_3 NI_3 NS_30 0 1.9983224645311447e-02
GC_3_31 b_3 NI_3 NS_31 0 -1.8056402408979944e-01
GC_3_32 b_3 NI_3 NS_32 0 5.8222616453944297e-02
GC_3_33 b_3 NI_3 NS_33 0 -2.5838412793910398e-04
GC_3_34 b_3 NI_3 NS_34 0 8.8719418219103082e-05
GC_3_35 b_3 NI_3 NS_35 0 6.3340938564175147e-08
GC_3_36 b_3 NI_3 NS_36 0 1.5314905031318692e-07
GC_3_37 b_3 NI_3 NS_37 0 -2.9914601800437039e-02
GC_3_38 b_3 NI_3 NS_38 0 -6.1730447422708015e-02
GC_3_39 b_3 NI_3 NS_39 0 7.9867282628517555e-02
GC_3_40 b_3 NI_3 NS_40 0 -1.0211216826739468e-01
GC_3_41 b_3 NI_3 NS_41 0 -7.4453578692055883e-03
GC_3_42 b_3 NI_3 NS_42 0 -4.9122495668140606e-03
GC_3_43 b_3 NI_3 NS_43 0 -1.6828053234393356e-05
GC_3_44 b_3 NI_3 NS_44 0 -2.5005042973138882e-06
GC_3_45 b_3 NI_3 NS_45 0 -2.4057927051444822e-09
GC_3_46 b_3 NI_3 NS_46 0 -4.1381560943654256e-07
GC_3_47 b_3 NI_3 NS_47 0 1.8828664800414126e-03
GC_3_48 b_3 NI_3 NS_48 0 -1.2541806658330386e-02
GC_3_49 b_3 NI_3 NS_49 0 6.8132622328499585e-03
GC_3_50 b_3 NI_3 NS_50 0 1.1344904106816798e-02
GC_3_51 b_3 NI_3 NS_51 0 -1.6930073478816593e-03
GC_3_52 b_3 NI_3 NS_52 0 1.3502364287922241e-03
GC_3_53 b_3 NI_3 NS_53 0 -5.4834376104108819e-06
GC_3_54 b_3 NI_3 NS_54 0 1.1883635424574163e-08
GC_3_55 b_3 NI_3 NS_55 0 2.0709139958615838e-09
GC_3_56 b_3 NI_3 NS_56 0 1.2445061904298917e-07
GC_3_57 b_3 NI_3 NS_57 0 1.8365222464445088e-03
GC_3_58 b_3 NI_3 NS_58 0 -4.4016228950139450e-04
GC_3_59 b_3 NI_3 NS_59 0 -2.0380606253700127e-03
GC_3_60 b_3 NI_3 NS_60 0 -7.6032949324750742e-04
GC_3_61 b_3 NI_3 NS_61 0 -2.3322671330819693e-03
GC_3_62 b_3 NI_3 NS_62 0 -7.3299106530160917e-04
GC_3_63 b_3 NI_3 NS_63 0 -2.1712403229267354e-06
GC_3_64 b_3 NI_3 NS_64 0 7.9797619855397459e-09
GC_3_65 b_3 NI_3 NS_65 0 7.8796782395424921e-11
GC_3_66 b_3 NI_3 NS_66 0 -3.5701773202207393e-08
GC_3_67 b_3 NI_3 NS_67 0 5.4029071943898367e-04
GC_3_68 b_3 NI_3 NS_68 0 -1.1407089600036740e-03
GC_3_69 b_3 NI_3 NS_69 0 1.8427149076859011e-03
GC_3_70 b_3 NI_3 NS_70 0 -1.1617820217932944e-04
GC_3_71 b_3 NI_3 NS_71 0 2.2810331393171546e-04
GC_3_72 b_3 NI_3 NS_72 0 1.9523104902109329e-03
GC_3_73 b_3 NI_3 NS_73 0 2.4668573573564550e-06
GC_3_74 b_3 NI_3 NS_74 0 1.1782357808414174e-07
GC_3_75 b_3 NI_3 NS_75 0 -8.3492749474727398e-11
GC_3_76 b_3 NI_3 NS_76 0 3.2300971650928084e-08
GC_3_77 b_3 NI_3 NS_77 0 3.0095531788116819e-03
GC_3_78 b_3 NI_3 NS_78 0 -1.8743790592256403e-04
GC_3_79 b_3 NI_3 NS_79 0 -5.4033982711598118e-03
GC_3_80 b_3 NI_3 NS_80 0 -5.2386530036741886e-04
GC_3_81 b_3 NI_3 NS_81 0 -1.4365666755094526e-03
GC_3_82 b_3 NI_3 NS_82 0 -5.2555390307240787e-04
GC_3_83 b_3 NI_3 NS_83 0 -1.6806776345275893e-06
GC_3_84 b_3 NI_3 NS_84 0 2.0769026188550992e-07
GC_3_85 b_3 NI_3 NS_85 0 2.2668297248944703e-10
GC_3_86 b_3 NI_3 NS_86 0 -5.5163287780851915e-09
GC_3_87 b_3 NI_3 NS_87 0 3.6567389653507991e-04
GC_3_88 b_3 NI_3 NS_88 0 4.2773835993569132e-04
GC_3_89 b_3 NI_3 NS_89 0 1.4813020334029758e-03
GC_3_90 b_3 NI_3 NS_90 0 -1.7482834881565495e-03
GC_3_91 b_3 NI_3 NS_91 0 8.0853503837957744e-05
GC_3_92 b_3 NI_3 NS_92 0 6.1961854941422609e-04
GC_3_93 b_3 NI_3 NS_93 0 4.5901077523111817e-07
GC_3_94 b_3 NI_3 NS_94 0 1.6709687958626685e-09
GC_3_95 b_3 NI_3 NS_95 0 -2.0540839151132718e-10
GC_3_96 b_3 NI_3 NS_96 0 2.2654604492252261e-09
GC_3_97 b_3 NI_3 NS_97 0 5.4524373557005652e-04
GC_3_98 b_3 NI_3 NS_98 0 8.3637357368031027e-05
GC_3_99 b_3 NI_3 NS_99 0 -1.0621391184145259e-03
GC_3_100 b_3 NI_3 NS_100 0 3.5110894111764761e-04
GC_3_101 b_3 NI_3 NS_101 0 -1.5101101547256504e-04
GC_3_102 b_3 NI_3 NS_102 0 -2.5226873642479234e-04
GC_3_103 b_3 NI_3 NS_103 0 -3.1559083619842678e-07
GC_3_104 b_3 NI_3 NS_104 0 4.4709851055151867e-08
GC_3_105 b_3 NI_3 NS_105 0 1.0763565109496663e-10
GC_3_106 b_3 NI_3 NS_106 0 5.1223218225402046e-11
GC_3_107 b_3 NI_3 NS_107 0 8.6980632206588211e-05
GC_3_108 b_3 NI_3 NS_108 0 1.6471800050515666e-04
GC_3_109 b_3 NI_3 NS_109 0 3.1645865418488691e-04
GC_3_110 b_3 NI_3 NS_110 0 -5.7183067031546487e-04
GC_3_111 b_3 NI_3 NS_111 0 -6.8047032396455873e-05
GC_3_112 b_3 NI_3 NS_112 0 3.4261133561112981e-04
GC_3_113 b_3 NI_3 NS_113 0 -2.0319496336951487e-08
GC_3_114 b_3 NI_3 NS_114 0 1.4268774072850567e-08
GC_3_115 b_3 NI_3 NS_115 0 -1.0175329619432754e-10
GC_3_116 b_3 NI_3 NS_116 0 -9.1092915343631042e-10
GC_3_117 b_3 NI_3 NS_117 0 -5.6817933891895275e-05
GC_3_118 b_3 NI_3 NS_118 0 1.2050288604751119e-04
GC_3_119 b_3 NI_3 NS_119 0 2.1853855541131872e-05
GC_3_120 b_3 NI_3 NS_120 0 5.8520010637099862e-04
GD_3_1 b_3 NI_3 NA_1 0 3.1107304579876829e-02
GD_3_2 b_3 NI_3 NA_2 0 3.7223665651837500e-04
GD_3_3 b_3 NI_3 NA_3 0 -1.9437694054582878e-02
GD_3_4 b_3 NI_3 NA_4 0 2.0560510158963128e-02
GD_3_5 b_3 NI_3 NA_5 0 3.0268489456894625e-02
GD_3_6 b_3 NI_3 NA_6 0 3.6472629992843799e-04
GD_3_7 b_3 NI_3 NA_7 0 3.7468483141920228e-03
GD_3_8 b_3 NI_3 NA_8 0 1.3849076435686723e-04
GD_3_9 b_3 NI_3 NA_9 0 4.2051920717500632e-04
GD_3_10 b_3 NI_3 NA_10 0 -1.3536897167817916e-04
GD_3_11 b_3 NI_3 NA_11 0 3.9286024601949428e-05
GD_3_12 b_3 NI_3 NA_12 0 -1.6521754335559500e-04
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 -1.3064076650635922e-03
GC_4_2 b_4 NI_4 NS_2 0 1.1609671570068636e-03
GC_4_3 b_4 NI_4 NS_3 0 -5.2046701074105827e-06
GC_4_4 b_4 NI_4 NS_4 0 -1.3622416252452102e-07
GC_4_5 b_4 NI_4 NS_5 0 1.8849506907402238e-09
GC_4_6 b_4 NI_4 NS_6 0 1.0944781804581485e-07
GC_4_7 b_4 NI_4 NS_7 0 2.1789912091479606e-03
GC_4_8 b_4 NI_4 NS_8 0 -5.3354771307407233e-04
GC_4_9 b_4 NI_4 NS_9 0 -2.6661110234395880e-03
GC_4_10 b_4 NI_4 NS_10 0 -1.2464190329196801e-03
GC_4_11 b_4 NI_4 NS_11 0 -7.0303330590827115e-03
GC_4_12 b_4 NI_4 NS_12 0 -4.4850017400638060e-03
GC_4_13 b_4 NI_4 NS_13 0 -1.6071362626906194e-05
GC_4_14 b_4 NI_4 NS_14 0 -2.4812561109900059e-06
GC_4_15 b_4 NI_4 NS_15 0 -2.2962509480293271e-09
GC_4_16 b_4 NI_4 NS_16 0 -3.9507715081732348e-07
GC_4_17 b_4 NI_4 NS_17 0 1.7173864573176683e-03
GC_4_18 b_4 NI_4 NS_18 0 -1.3398639507239605e-02
GC_4_19 b_4 NI_4 NS_19 0 5.8796835844652567e-03
GC_4_20 b_4 NI_4 NS_20 0 1.3002224138356774e-02
GC_4_21 b_4 NI_4 NS_21 0 -1.8053477368745591e-01
GC_4_22 b_4 NI_4 NS_22 0 5.8214943362432180e-02
GC_4_23 b_4 NI_4 NS_23 0 -2.5831874125337574e-04
GC_4_24 b_4 NI_4 NS_24 0 8.8703972290716547e-05
GC_4_25 b_4 NI_4 NS_25 0 6.3332061302203367e-08
GC_4_26 b_4 NI_4 NS_26 0 1.5369534788214769e-07
GC_4_27 b_4 NI_4 NS_27 0 -2.9914538229092451e-02
GC_4_28 b_4 NI_4 NS_28 0 -6.1725780150516558e-02
GC_4_29 b_4 NI_4 NS_29 0 7.9857089031509718e-02
GC_4_30 b_4 NI_4 NS_30 0 -1.0210628552638608e-01
GC_4_31 b_4 NI_4 NS_31 0 5.3616779120527064e-02
GC_4_32 b_4 NI_4 NS_32 0 -1.2804945067003930e-02
GC_4_33 b_4 NI_4 NS_33 0 6.3940087657096697e-05
GC_4_34 b_4 NI_4 NS_34 0 -1.3871599455596756e-05
GC_4_35 b_4 NI_4 NS_35 0 -1.0851117673452737e-08
GC_4_36 b_4 NI_4 NS_36 0 -1.2971657354454211e-06
GC_4_37 b_4 NI_4 NS_37 0 -1.9507878599407341e-03
GC_4_38 b_4 NI_4 NS_38 0 7.0862888731600430e-03
GC_4_39 b_4 NI_4 NS_39 0 -1.3281287280820304e-02
GC_4_40 b_4 NI_4 NS_40 0 1.9983224645311447e-02
GC_4_41 b_4 NI_4 NS_41 0 -1.6906647619615888e-03
GC_4_42 b_4 NI_4 NS_42 0 1.3498081337613578e-03
GC_4_43 b_4 NI_4 NS_43 0 -5.4853564407898510e-06
GC_4_44 b_4 NI_4 NS_44 0 1.2354608941308510e-08
GC_4_45 b_4 NI_4 NS_45 0 2.0709613395574615e-09
GC_4_46 b_4 NI_4 NS_46 0 1.2443764671550607e-07
GC_4_47 b_4 NI_4 NS_47 0 1.8367429921158365e-03
GC_4_48 b_4 NI_4 NS_48 0 -4.3939078431075741e-04
GC_4_49 b_4 NI_4 NS_49 0 -2.0386602365681157e-03
GC_4_50 b_4 NI_4 NS_50 0 -7.5963722639747408e-04
GC_4_51 b_4 NI_4 NS_51 0 -7.4378040029148881e-03
GC_4_52 b_4 NI_4 NS_52 0 -4.9141564383269843e-03
GC_4_53 b_4 NI_4 NS_53 0 -1.6815914593756500e-05
GC_4_54 b_4 NI_4 NS_54 0 -2.5025348227531276e-06
GC_4_55 b_4 NI_4 NS_55 0 -2.4059027513451994e-09
GC_4_56 b_4 NI_4 NS_56 0 -4.1378168389794281e-07
GC_4_57 b_4 NI_4 NS_57 0 1.8819564725814338e-03
GC_4_58 b_4 NI_4 NS_58 0 -1.2540693866371440e-02
GC_4_59 b_4 NI_4 NS_59 0 6.8108563693077585e-03
GC_4_60 b_4 NI_4 NS_60 0 1.1346968206311200e-02
GC_4_61 b_4 NI_4 NS_61 0 2.2630995476374629e-04
GC_4_62 b_4 NI_4 NS_62 0 1.9528009480232883e-03
GC_4_63 b_4 NI_4 NS_63 0 2.4633713577156198e-06
GC_4_64 b_4 NI_4 NS_64 0 1.1838736295482264e-07
GC_4_65 b_4 NI_4 NS_65 0 -8.3451289097620632e-11
GC_4_66 b_4 NI_4 NS_66 0 3.2291767275360039e-08
GC_4_67 b_4 NI_4 NS_67 0 3.0097364790043308e-03
GC_4_68 b_4 NI_4 NS_68 0 -1.8752914992742236e-04
GC_4_69 b_4 NI_4 NS_69 0 -5.4027259304871809e-03
GC_4_70 b_4 NI_4 NS_70 0 -5.2429066922317369e-04
GC_4_71 b_4 NI_4 NS_71 0 -2.3327760589818185e-03
GC_4_72 b_4 NI_4 NS_72 0 -7.3280499473649216e-04
GC_4_73 b_4 NI_4 NS_73 0 -2.1736547825694142e-06
GC_4_74 b_4 NI_4 NS_74 0 8.4466433157991678e-09
GC_4_75 b_4 NI_4 NS_75 0 7.8799854867671654e-11
GC_4_76 b_4 NI_4 NS_76 0 -3.5713989682144621e-08
GC_4_77 b_4 NI_4 NS_77 0 5.4021439236045968e-04
GC_4_78 b_4 NI_4 NS_78 0 -1.1406079012404031e-03
GC_4_79 b_4 NI_4 NS_79 0 1.8429926025739906e-03
GC_4_80 b_4 NI_4 NS_80 0 -1.1617592408276236e-04
GC_4_81 b_4 NI_4 NS_81 0 8.1654121462430338e-05
GC_4_82 b_4 NI_4 NS_82 0 6.1942409181479289e-04
GC_4_83 b_4 NI_4 NS_83 0 4.5980700814682754e-07
GC_4_84 b_4 NI_4 NS_84 0 1.5473232055628190e-09
GC_4_85 b_4 NI_4 NS_85 0 -2.0541669074526852e-10
GC_4_86 b_4 NI_4 NS_86 0 2.2671228369173445e-09
GC_4_87 b_4 NI_4 NS_87 0 5.4512433979936878e-04
GC_4_88 b_4 NI_4 NS_88 0 8.3645148241201910e-05
GC_4_89 b_4 NI_4 NS_89 0 -1.0624996024421482e-03
GC_4_90 b_4 NI_4 NS_90 0 3.5134323036855632e-04
GC_4_91 b_4 NI_4 NS_91 0 -1.4365981285533625e-03
GC_4_92 b_4 NI_4 NS_92 0 -5.2554836834912196e-04
GC_4_93 b_4 NI_4 NS_93 0 -1.6806885297593111e-06
GC_4_94 b_4 NI_4 NS_94 0 2.0769313928527144e-07
GC_4_95 b_4 NI_4 NS_95 0 2.2668288943092759e-10
GC_4_96 b_4 NI_4 NS_96 0 -5.5164355151380002e-09
GC_4_97 b_4 NI_4 NS_97 0 3.6567678318688264e-04
GC_4_98 b_4 NI_4 NS_98 0 4.2773342079281218e-04
GC_4_99 b_4 NI_4 NS_99 0 1.4813104413553093e-03
GC_4_100 b_4 NI_4 NS_100 0 -1.7482970824392419e-03
GC_4_101 b_4 NI_4 NS_101 0 -6.8745335049225241e-05
GC_4_102 b_4 NI_4 NS_102 0 3.4274282199370796e-04
GC_4_103 b_4 NI_4 NS_103 0 -2.0454017307283064e-08
GC_4_104 b_4 NI_4 NS_104 0 1.4315479645448529e-08
GC_4_105 b_4 NI_4 NS_105 0 -1.0174599979241521e-10
GC_4_106 b_4 NI_4 NS_106 0 -9.1155877990923631e-10
GC_4_107 b_4 NI_4 NS_107 0 -5.6845318325416464e-05
GC_4_108 b_4 NI_4 NS_108 0 1.2032180497915186e-04
GC_4_109 b_4 NI_4 NS_109 0 2.2055688259251361e-05
GC_4_110 b_4 NI_4 NS_110 0 5.8497488874929653e-04
GC_4_111 b_4 NI_4 NS_111 0 -1.5072974180017139e-04
GC_4_112 b_4 NI_4 NS_112 0 -2.5231601036312034e-04
GC_4_113 b_4 NI_4 NS_113 0 -3.1459273271146477e-07
GC_4_114 b_4 NI_4 NS_114 0 4.4593311782414919e-08
GC_4_115 b_4 NI_4 NS_115 0 1.0762446501307339e-10
GC_4_116 b_4 NI_4 NS_116 0 5.3288867417633135e-11
GC_4_117 b_4 NI_4 NS_117 0 8.6952963580351079e-05
GC_4_118 b_4 NI_4 NS_118 0 1.6486089740420866e-04
GC_4_119 b_4 NI_4 NS_119 0 3.1649716165064063e-04
GC_4_120 b_4 NI_4 NS_120 0 -5.7166537939438609e-04
GD_4_1 b_4 NI_4 NA_1 0 3.7211526732520192e-04
GD_4_2 b_4 NI_4 NA_2 0 3.1099222062001709e-02
GD_4_3 b_4 NI_4 NA_3 0 2.0551875096802001e-02
GD_4_4 b_4 NI_4 NA_4 0 -1.9437694054582878e-02
GD_4_5 b_4 NI_4 NA_5 0 3.6355392340526888e-04
GD_4_6 b_4 NI_4 NA_6 0 3.0267098594982021e-02
GD_4_7 b_4 NI_4 NA_7 0 1.3886656467954533e-04
GD_4_8 b_4 NI_4 NA_8 0 3.7471263744355775e-03
GD_4_9 b_4 NI_4 NA_9 0 -1.3541351404501971e-04
GD_4_10 b_4 NI_4 NA_10 0 4.2053241529844932e-04
GD_4_11 b_4 NI_4 NA_11 0 -1.6492366173784606e-04
GD_4_12 b_4 NI_4 NA_12 0 3.9104219663086600e-05
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 -2.7969920567862752e-03
GC_5_2 b_5 NI_5 NS_2 0 -5.7452506927769273e-04
GC_5_3 b_5 NI_5 NS_3 0 -2.2977364695200834e-06
GC_5_4 b_5 NI_5 NS_4 0 5.4639600786713524e-08
GC_5_5 b_5 NI_5 NS_5 0 1.0754501521530430e-10
GC_5_6 b_5 NI_5 NS_6 0 -3.1810271387062057e-08
GC_5_7 b_5 NI_5 NS_7 0 5.7236763104545954e-04
GC_5_8 b_5 NI_5 NS_8 0 -1.1831822711651785e-03
GC_5_9 b_5 NI_5 NS_9 0 2.0484023784160615e-03
GC_5_10 b_5 NI_5 NS_10 0 -7.4431985879680877e-05
GC_5_11 b_5 NI_5 NS_11 0 4.4879461587188715e-04
GC_5_12 b_5 NI_5 NS_12 0 1.7423941774537904e-03
GC_5_13 b_5 NI_5 NS_13 0 2.5851612781879403e-06
GC_5_14 b_5 NI_5 NS_14 0 6.8465792549908691e-08
GC_5_15 b_5 NI_5 NS_15 0 -1.1309071083045831e-10
GC_5_16 b_5 NI_5 NS_16 0 2.8407691385166663e-08
GC_5_17 b_5 NI_5 NS_17 0 3.2315056701227090e-03
GC_5_18 b_5 NI_5 NS_18 0 -2.7458384256641893e-04
GC_5_19 b_5 NI_5 NS_19 0 -5.7928527581335354e-03
GC_5_20 b_5 NI_5 NS_20 0 -1.0206293933180512e-03
GC_5_21 b_5 NI_5 NS_21 0 -7.4378040029148881e-03
GC_5_22 b_5 NI_5 NS_22 0 -4.9141564383269843e-03
GC_5_23 b_5 NI_5 NS_23 0 -1.6815914593756500e-05
GC_5_24 b_5 NI_5 NS_24 0 -2.5025348227531276e-06
GC_5_25 b_5 NI_5 NS_25 0 -2.4059027513451994e-09
GC_5_26 b_5 NI_5 NS_26 0 -4.1378168389794281e-07
GC_5_27 b_5 NI_5 NS_27 0 1.8819564725814338e-03
GC_5_28 b_5 NI_5 NS_28 0 -1.2540693866371440e-02
GC_5_29 b_5 NI_5 NS_29 0 6.8108563693077585e-03
GC_5_30 b_5 NI_5 NS_30 0 1.1346968206311200e-02
GC_5_31 b_5 NI_5 NS_31 0 -1.6930073478816593e-03
GC_5_32 b_5 NI_5 NS_32 0 1.3502364287922241e-03
GC_5_33 b_5 NI_5 NS_33 0 -5.4834376104108819e-06
GC_5_34 b_5 NI_5 NS_34 0 1.1883635424574163e-08
GC_5_35 b_5 NI_5 NS_35 0 2.0709139958615838e-09
GC_5_36 b_5 NI_5 NS_36 0 1.2445061904298917e-07
GC_5_37 b_5 NI_5 NS_37 0 1.8365222464445088e-03
GC_5_38 b_5 NI_5 NS_38 0 -4.4016228950139450e-04
GC_5_39 b_5 NI_5 NS_39 0 -2.0380606253700127e-03
GC_5_40 b_5 NI_5 NS_40 0 -7.6032949324750742e-04
GC_5_41 b_5 NI_5 NS_41 0 5.4006912402350546e-02
GC_5_42 b_5 NI_5 NS_42 0 -1.2950691146545073e-02
GC_5_43 b_5 NI_5 NS_43 0 6.4022433177070648e-05
GC_5_44 b_5 NI_5 NS_44 0 -1.3923962664081735e-05
GC_5_45 b_5 NI_5 NS_45 0 -1.0941649914308505e-08
GC_5_46 b_5 NI_5 NS_46 0 -1.2992905082218793e-06
GC_5_47 b_5 NI_5 NS_47 0 -1.9794279676321950e-03
GC_5_48 b_5 NI_5 NS_48 0 7.1109620097927701e-03
GC_5_49 b_5 NI_5 NS_49 0 -1.3471842032580358e-02
GC_5_50 b_5 NI_5 NS_50 0 1.9910115330593642e-02
GC_5_51 b_5 NI_5 NS_51 0 -1.8079964333789753e-01
GC_5_52 b_5 NI_5 NS_52 0 5.8436898552091006e-02
GC_5_53 b_5 NI_5 NS_53 0 -2.5852355481785911e-04
GC_5_54 b_5 NI_5 NS_54 0 8.8784818964496231e-05
GC_5_55 b_5 NI_5 NS_55 0 6.3382912203639814e-08
GC_5_56 b_5 NI_5 NS_56 0 1.5614098786017617e-07
GC_5_57 b_5 NI_5 NS_57 0 -3.0132494090102643e-02
GC_5_58 b_5 NI_5 NS_58 0 -6.1641023575303065e-02
GC_5_59 b_5 NI_5 NS_59 0 8.0265196632208782e-02
GC_5_60 b_5 NI_5 NS_60 0 -1.0161816519012962e-01
GC_5_61 b_5 NI_5 NS_61 0 -7.1335350725222563e-03
GC_5_62 b_5 NI_5 NS_62 0 -4.9995367140875154e-03
GC_5_63 b_5 NI_5 NS_63 0 -1.6852299141023232e-05
GC_5_64 b_5 NI_5 NS_64 0 -2.5007847077580000e-06
GC_5_65 b_5 NI_5 NS_65 0 -2.4106580984269951e-09
GC_5_66 b_5 NI_5 NS_66 0 -4.1484901461924044e-07
GC_5_67 b_5 NI_5 NS_67 0 1.8568840199841255e-03
GC_5_68 b_5 NI_5 NS_68 0 -1.2583849639531257e-02
GC_5_69 b_5 NI_5 NS_69 0 6.6065037028949581e-03
GC_5_70 b_5 NI_5 NS_70 0 1.1379025617293689e-02
GC_5_71 b_5 NI_5 NS_71 0 -1.7545021297831079e-03
GC_5_72 b_5 NI_5 NS_72 0 1.3885706843359328e-03
GC_5_73 b_5 NI_5 NS_73 0 -5.3567699787057151e-06
GC_5_74 b_5 NI_5 NS_74 0 -4.8002346001029380e-09
GC_5_75 b_5 NI_5 NS_75 0 2.0762984422569127e-09
GC_5_76 b_5 NI_5 NS_76 0 1.2570450778367722e-07
GC_5_77 b_5 NI_5 NS_77 0 1.8062233681799193e-03
GC_5_78 b_5 NI_5 NS_78 0 -4.1873044973439797e-04
GC_5_79 b_5 NI_5 NS_79 0 -1.9478748151075685e-03
GC_5_80 b_5 NI_5 NS_80 0 -6.8414348926347816e-04
GC_5_81 b_5 NI_5 NS_81 0 -2.3329916798764672e-03
GC_5_82 b_5 NI_5 NS_82 0 -7.3276860499570150e-04
GC_5_83 b_5 NI_5 NS_83 0 -2.1754894548739566e-06
GC_5_84 b_5 NI_5 NS_84 0 8.9813158443094226e-09
GC_5_85 b_5 NI_5 NS_85 0 7.8802453510202652e-11
GC_5_86 b_5 NI_5 NS_86 0 -3.5713227815655763e-08
GC_5_87 b_5 NI_5 NS_87 0 5.4026267907607913e-04
GC_5_88 b_5 NI_5 NS_88 0 -1.1406344561067309e-03
GC_5_89 b_5 NI_5 NS_89 0 1.8430652824974693e-03
GC_5_90 b_5 NI_5 NS_90 0 -1.1628231309278826e-04
GC_5_91 b_5 NI_5 NS_91 0 2.2571822946922183e-04
GC_5_92 b_5 NI_5 NS_92 0 1.9527876275770560e-03
GC_5_93 b_5 NI_5 NS_93 0 2.4667422030195401e-06
GC_5_94 b_5 NI_5 NS_94 0 1.1763930329096830e-07
GC_5_95 b_5 NI_5 NS_95 0 -8.3450274923965756e-11
GC_5_96 b_5 NI_5 NS_96 0 3.2296174829919205e-08
GC_5_97 b_5 NI_5 NS_97 0 3.0097804134294292e-03
GC_5_98 b_5 NI_5 NS_98 0 -1.8781201218584880e-04
GC_5_99 b_5 NI_5 NS_99 0 -5.4027133649887319e-03
GC_5_100 b_5 NI_5 NS_100 0 -5.2475450255814527e-04
GC_5_101 b_5 NI_5 NS_101 0 -1.8102426904621134e-03
GC_5_102 b_5 NI_5 NS_102 0 -4.2556367560624044e-04
GC_5_103 b_5 NI_5 NS_103 0 -1.7767726003691285e-06
GC_5_104 b_5 NI_5 NS_104 0 2.3259814246150690e-07
GC_5_105 b_5 NI_5 NS_105 0 2.3519255691818629e-10
GC_5_106 b_5 NI_5 NS_106 0 -4.8199409832769711e-09
GC_5_107 b_5 NI_5 NS_107 0 3.9578927010691737e-04
GC_5_108 b_5 NI_5 NS_108 0 4.5730820886789983e-04
GC_5_109 b_5 NI_5 NS_109 0 1.7014713360919190e-03
GC_5_110 b_5 NI_5 NS_110 0 -1.8062990478043073e-03
GC_5_111 b_5 NI_5 NS_111 0 1.7713520644807633e-04
GC_5_112 b_5 NI_5 NS_112 0 5.7711503772868910e-04
GC_5_113 b_5 NI_5 NS_113 0 3.8437197205538283e-07
GC_5_114 b_5 NI_5 NS_114 0 5.6131200511718194e-09
GC_5_115 b_5 NI_5 NS_115 0 -2.1142105692611963e-10
GC_5_116 b_5 NI_5 NS_116 0 1.1233157414133004e-09
GC_5_117 b_5 NI_5 NS_117 0 5.7503237530367470e-04
GC_5_118 b_5 NI_5 NS_118 0 7.6072738321982355e-05
GC_5_119 b_5 NI_5 NS_119 0 -1.1522395821956836e-03
GC_5_120 b_5 NI_5 NS_120 0 2.9493613797594543e-04
GD_5_1 b_5 NI_5 NA_1 0 3.8606050553713798e-03
GD_5_2 b_5 NI_5 NA_2 0 2.3520227332051908e-04
GD_5_3 b_5 NI_5 NA_3 0 3.0267098594982021e-02
GD_5_4 b_5 NI_5 NA_4 0 3.6472629992843799e-04
GD_5_5 b_5 NI_5 NA_5 0 -1.9510056231500820e-02
GD_5_6 b_5 NI_5 NA_6 0 2.0461907702647508e-02
GD_5_7 b_5 NI_5 NA_7 0 3.0282091253999912e-02
GD_5_8 b_5 NI_5 NA_8 0 3.3251620337900492e-04
GD_5_9 b_5 NI_5 NA_9 0 3.7471538655471826e-03
GD_5_10 b_5 NI_5 NA_10 0 1.3931914091957427e-04
GD_5_11 b_5 NI_5 NA_11 0 4.3527000620696211e-04
GD_5_12 b_5 NI_5 NA_12 0 -1.3162559052130131e-04
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 4.4221077296529839e-04
GC_6_2 b_6 NI_6 NS_2 0 1.7436489372742686e-03
GC_6_3 b_6 NI_6 NS_3 0 2.5868934374718469e-06
GC_6_4 b_6 NI_6 NS_4 0 6.8132163790513363e-08
GC_6_5 b_6 NI_6 NS_5 0 -1.1317491206945763e-10
GC_6_6 b_6 NI_6 NS_6 0 2.8413703378657205e-08
GC_6_7 b_6 NI_6 NS_7 0 3.2308596094018337e-03
GC_6_8 b_6 NI_6 NS_8 0 -2.7670604659806134e-04
GC_6_9 b_6 NI_6 NS_9 0 -5.7911556532728430e-03
GC_6_10 b_6 NI_6 NS_10 0 -1.0224888052617921e-03
GC_6_11 b_6 NI_6 NS_11 0 -2.7882340457254899e-03
GC_6_12 b_6 NI_6 NS_12 0 -5.7603257060246760e-04
GC_6_13 b_6 NI_6 NS_13 0 -2.2832322525186888e-06
GC_6_14 b_6 NI_6 NS_14 0 5.2509674129389776e-08
GC_6_15 b_6 NI_6 NS_15 0 1.0694927813137638e-10
GC_6_16 b_6 NI_6 NS_16 0 -3.1757470645053139e-08
GC_6_17 b_6 NI_6 NS_17 0 5.7218330748787141e-04
GC_6_18 b_6 NI_6 NS_18 0 -1.1815750180375708e-03
GC_6_19 b_6 NI_6 NS_19 0 2.0454127164122879e-03
GC_6_20 b_6 NI_6 NS_20 0 -7.0599483380387278e-05
GC_6_21 b_6 NI_6 NS_21 0 -1.6906647619615888e-03
GC_6_22 b_6 NI_6 NS_22 0 1.3498081337613578e-03
GC_6_23 b_6 NI_6 NS_23 0 -5.4853564407898510e-06
GC_6_24 b_6 NI_6 NS_24 0 1.2354608941308510e-08
GC_6_25 b_6 NI_6 NS_25 0 2.0709613395574615e-09
GC_6_26 b_6 NI_6 NS_26 0 1.2443764671550607e-07
GC_6_27 b_6 NI_6 NS_27 0 1.8367429921158365e-03
GC_6_28 b_6 NI_6 NS_28 0 -4.3939078431075741e-04
GC_6_29 b_6 NI_6 NS_29 0 -2.0386602365681157e-03
GC_6_30 b_6 NI_6 NS_30 0 -7.5963722639747408e-04
GC_6_31 b_6 NI_6 NS_31 0 -7.4453578692055883e-03
GC_6_32 b_6 NI_6 NS_32 0 -4.9122495668140606e-03
GC_6_33 b_6 NI_6 NS_33 0 -1.6828053234393356e-05
GC_6_34 b_6 NI_6 NS_34 0 -2.5005042973138882e-06
GC_6_35 b_6 NI_6 NS_35 0 -2.4057927051444822e-09
GC_6_36 b_6 NI_6 NS_36 0 -4.1381560943654256e-07
GC_6_37 b_6 NI_6 NS_37 0 1.8828664800414126e-03
GC_6_38 b_6 NI_6 NS_38 0 -1.2541806658330386e-02
GC_6_39 b_6 NI_6 NS_39 0 6.8132622328499585e-03
GC_6_40 b_6 NI_6 NS_40 0 1.1344904106816798e-02
GC_6_41 b_6 NI_6 NS_41 0 -1.8080052518981293e-01
GC_6_42 b_6 NI_6 NS_42 0 5.8437000775994237e-02
GC_6_43 b_6 NI_6 NS_43 0 -2.5852245127656187e-04
GC_6_44 b_6 NI_6 NS_44 0 8.8784467063390699e-05
GC_6_45 b_6 NI_6 NS_45 0 6.3382629439638723e-08
GC_6_46 b_6 NI_6 NS_46 0 1.5615765429789474e-07
GC_6_47 b_6 NI_6 NS_47 0 -3.0132175031306638e-02
GC_6_48 b_6 NI_6 NS_48 0 -6.1641134674318657e-02
GC_6_49 b_6 NI_6 NS_49 0 8.0265403994549123e-02
GC_6_50 b_6 NI_6 NS_50 0 -1.0161874818714424e-01
GC_6_51 b_6 NI_6 NS_51 0 5.4006912402350546e-02
GC_6_52 b_6 NI_6 NS_52 0 -1.2950691146545073e-02
GC_6_53 b_6 NI_6 NS_53 0 6.4022433177070648e-05
GC_6_54 b_6 NI_6 NS_54 0 -1.3923962664081735e-05
GC_6_55 b_6 NI_6 NS_55 0 -1.0941649914308505e-08
GC_6_56 b_6 NI_6 NS_56 0 -1.2992905082218793e-06
GC_6_57 b_6 NI_6 NS_57 0 -1.9794279676321950e-03
GC_6_58 b_6 NI_6 NS_58 0 7.1109620097927701e-03
GC_6_59 b_6 NI_6 NS_59 0 -1.3471842032580358e-02
GC_6_60 b_6 NI_6 NS_60 0 1.9910115330593642e-02
GC_6_61 b_6 NI_6 NS_61 0 -1.7545992716934914e-03
GC_6_62 b_6 NI_6 NS_62 0 1.3886113187470833e-03
GC_6_63 b_6 NI_6 NS_63 0 -5.3570467780378706e-06
GC_6_64 b_6 NI_6 NS_64 0 -4.7668777811152306e-09
GC_6_65 b_6 NI_6 NS_65 0 2.0763013949805005e-09
GC_6_66 b_6 NI_6 NS_66 0 1.2570424061425725e-07
GC_6_67 b_6 NI_6 NS_67 0 1.8063163299997973e-03
GC_6_68 b_6 NI_6 NS_68 0 -4.1865530881807976e-04
GC_6_69 b_6 NI_6 NS_69 0 -1.9477700115534855e-03
GC_6_70 b_6 NI_6 NS_70 0 -6.8416278358347836e-04
GC_6_71 b_6 NI_6 NS_71 0 -7.1335583433311768e-03
GC_6_72 b_6 NI_6 NS_72 0 -4.9995327285223953e-03
GC_6_73 b_6 NI_6 NS_73 0 -1.6852307537586127e-05
GC_6_74 b_6 NI_6 NS_74 0 -2.5007837701117546e-06
GC_6_75 b_6 NI_6 NS_75 0 -2.4106584866412858e-09
GC_6_76 b_6 NI_6 NS_76 0 -4.1484905145946999e-07
GC_6_77 b_6 NI_6 NS_77 0 1.8568853967698838e-03
GC_6_78 b_6 NI_6 NS_78 0 -1.2583855237402349e-02
GC_6_79 b_6 NI_6 NS_79 0 6.6065082787264279e-03
GC_6_80 b_6 NI_6 NS_80 0 1.1379015469041411e-02
GC_6_81 b_6 NI_6 NS_81 0 2.2498716385862400e-04
GC_6_82 b_6 NI_6 NS_82 0 1.9530786948455984e-03
GC_6_83 b_6 NI_6 NS_83 0 2.4631372121652609e-06
GC_6_84 b_6 NI_6 NS_84 0 1.1825817633892398e-07
GC_6_85 b_6 NI_6 NS_85 0 -8.3403319346910024e-11
GC_6_86 b_6 NI_6 NS_86 0 3.2286921814126651e-08
GC_6_87 b_6 NI_6 NS_87 0 3.0098587914049930e-03
GC_6_88 b_6 NI_6 NS_88 0 -1.8773057630928588e-04
GC_6_89 b_6 NI_6 NS_89 0 -5.4023417777550094e-03
GC_6_90 b_6 NI_6 NS_90 0 -5.2475672159504536e-04
GC_6_91 b_6 NI_6 NS_91 0 -2.3329145978155381e-03
GC_6_92 b_6 NI_6 NS_92 0 -7.3285603310363587e-04
GC_6_93 b_6 NI_6 NS_93 0 -2.1737376380831570e-06
GC_6_94 b_6 NI_6 NS_94 0 8.6499861841235125e-09
GC_6_95 b_6 NI_6 NS_95 0 7.8813825396023021e-11
GC_6_96 b_6 NI_6 NS_96 0 -3.5704257177941657e-08
GC_6_97 b_6 NI_6 NS_97 0 5.4038413931800340e-04
GC_6_98 b_6 NI_6 NS_98 0 -1.1407863730068064e-03
GC_6_99 b_6 NI_6 NS_99 0 1.8429279956086277e-03
GC_6_100 b_6 NI_6 NS_100 0 -1.1642622848298793e-04
GC_6_101 b_6 NI_6 NS_101 0 1.7522211295129583e-04
GC_6_102 b_6 NI_6 NS_102 0 5.7756027331900108e-04
GC_6_103 b_6 NI_6 NS_103 0 3.8288848137316545e-07
GC_6_104 b_6 NI_6 NS_104 0 5.8957332192288453e-09
GC_6_105 b_6 NI_6 NS_105 0 -2.1138941227792093e-10
GC_6_106 b_6 NI_6 NS_106 0 1.1214493077146343e-09
GC_6_107 b_6 NI_6 NS_107 0 5.7477864997957143e-04
GC_6_108 b_6 NI_6 NS_108 0 7.5486065024909612e-05
GC_6_109 b_6 NI_6 NS_109 0 -1.1516616088126793e-03
GC_6_110 b_6 NI_6 NS_110 0 2.9458902867056846e-04
GC_6_111 b_6 NI_6 NS_111 0 -1.8082139400216366e-03
GC_6_112 b_6 NI_6 NS_112 0 -4.2594882966600993e-04
GC_6_113 b_6 NI_6 NS_113 0 -1.7706788427184878e-06
GC_6_114 b_6 NI_6 NS_114 0 2.3157148955476831e-07
GC_6_115 b_6 NI_6 NS_115 0 2.3505527812462354e-10
GC_6_116 b_6 NI_6 NS_116 0 -4.7985459397601332e-09
GC_6_117 b_6 NI_6 NS_117 0 3.9569725122428880e-04
GC_6_118 b_6 NI_6 NS_118 0 4.5790575336839251e-04
GC_6_119 b_6 NI_6 NS_119 0 1.7010822969953400e-03
GC_6_120 b_6 NI_6 NS_120 0 -1.8054030035425629e-03
GD_6_1 b_6 NI_6 NA_1 0 2.3853587052750537e-04
GD_6_2 b_6 NI_6 NA_2 0 3.8585855893856912e-03
GD_6_3 b_6 NI_6 NA_3 0 3.6355392340526888e-04
GD_6_4 b_6 NI_6 NA_4 0 3.0268489456894625e-02
GD_6_5 b_6 NI_6 NA_5 0 2.0462026662063738e-02
GD_6_6 b_6 NI_6 NA_6 0 -1.9510056231500820e-02
GD_6_7 b_6 NI_6 NA_7 0 3.3234763115963739e-04
GD_6_8 b_6 NI_6 NA_8 0 3.0282103036456426e-02
GD_6_9 b_6 NI_6 NA_9 0 1.3932018935636532e-04
GD_6_10 b_6 NI_6 NA_10 0 3.7469884696672427e-03
GD_6_11 b_6 NI_6 NA_11 0 -1.3079590950170296e-04
GD_6_12 b_6 NI_6 NA_12 0 4.3459351420468783e-04
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 -1.8103086080908442e-03
GC_7_2 b_7 NI_7 NS_2 0 -4.2554411892932811e-04
GC_7_3 b_7 NI_7 NS_3 0 -1.7770576628909205e-06
GC_7_4 b_7 NI_7 NS_4 0 2.3274736994592285e-07
GC_7_5 b_7 NI_7 NS_5 0 2.3522415508806004e-10
GC_7_6 b_7 NI_7 NS_6 0 -4.8289272699913976e-09
GC_7_7 b_7 NI_7 NS_7 0 3.9578755176589793e-04
GC_7_8 b_7 NI_7 NS_8 0 4.5729849441930533e-04
GC_7_9 b_7 NI_7 NS_9 0 1.7014914530512301e-03
GC_7_10 b_7 NI_7 NS_10 0 -1.8063081690673948e-03
GC_7_11 b_7 NI_7 NS_11 0 1.7726806265213851e-04
GC_7_12 b_7 NI_7 NS_12 0 5.7708080829966266e-04
GC_7_13 b_7 NI_7 NS_13 0 3.8452142880391208e-07
GC_7_14 b_7 NI_7 NS_14 0 5.5176060545675808e-09
GC_7_15 b_7 NI_7 NS_15 0 -2.1149653085821725e-10
GC_7_16 b_7 NI_7 NS_16 0 1.1310143202669461e-09
GC_7_17 b_7 NI_7 NS_17 0 5.7502414607187187e-04
GC_7_18 b_7 NI_7 NS_18 0 7.6086239297994577e-05
GC_7_19 b_7 NI_7 NS_19 0 -1.1522858676960759e-03
GC_7_20 b_7 NI_7 NS_20 0 2.9496670632460673e-04
GC_7_21 b_7 NI_7 NS_21 0 -2.3327760589818185e-03
GC_7_22 b_7 NI_7 NS_22 0 -7.3280499473649216e-04
GC_7_23 b_7 NI_7 NS_23 0 -2.1736547825694142e-06
GC_7_24 b_7 NI_7 NS_24 0 8.4466433157991678e-09
GC_7_25 b_7 NI_7 NS_25 0 7.8799854867671654e-11
GC_7_26 b_7 NI_7 NS_26 0 -3.5713989682144621e-08
GC_7_27 b_7 NI_7 NS_27 0 5.4021439236045968e-04
GC_7_28 b_7 NI_7 NS_28 0 -1.1406079012404031e-03
GC_7_29 b_7 NI_7 NS_29 0 1.8429926025739906e-03
GC_7_30 b_7 NI_7 NS_30 0 -1.1617592408276236e-04
GC_7_31 b_7 NI_7 NS_31 0 2.2810331393171546e-04
GC_7_32 b_7 NI_7 NS_32 0 1.9523104902109329e-03
GC_7_33 b_7 NI_7 NS_33 0 2.4668573573564550e-06
GC_7_34 b_7 NI_7 NS_34 0 1.1782357808414174e-07
GC_7_35 b_7 NI_7 NS_35 0 -8.3492749474727398e-11
GC_7_36 b_7 NI_7 NS_36 0 3.2300971650928084e-08
GC_7_37 b_7 NI_7 NS_37 0 3.0095531788116819e-03
GC_7_38 b_7 NI_7 NS_38 0 -1.8743790592256403e-04
GC_7_39 b_7 NI_7 NS_39 0 -5.4033982711598118e-03
GC_7_40 b_7 NI_7 NS_40 0 -5.2386530036741886e-04
GC_7_41 b_7 NI_7 NS_41 0 -7.1335583433311768e-03
GC_7_42 b_7 NI_7 NS_42 0 -4.9995327285223953e-03
GC_7_43 b_7 NI_7 NS_43 0 -1.6852307537586127e-05
GC_7_44 b_7 NI_7 NS_44 0 -2.5007837701117546e-06
GC_7_45 b_7 NI_7 NS_45 0 -2.4106584866412858e-09
GC_7_46 b_7 NI_7 NS_46 0 -4.1484905145946999e-07
GC_7_47 b_7 NI_7 NS_47 0 1.8568853967698838e-03
GC_7_48 b_7 NI_7 NS_48 0 -1.2583855237402349e-02
GC_7_49 b_7 NI_7 NS_49 0 6.6065082787264279e-03
GC_7_50 b_7 NI_7 NS_50 0 1.1379015469041411e-02
GC_7_51 b_7 NI_7 NS_51 0 -1.7545021297831079e-03
GC_7_52 b_7 NI_7 NS_52 0 1.3885706843359328e-03
GC_7_53 b_7 NI_7 NS_53 0 -5.3567699787057151e-06
GC_7_54 b_7 NI_7 NS_54 0 -4.8002346001029380e-09
GC_7_55 b_7 NI_7 NS_55 0 2.0762984422569127e-09
GC_7_56 b_7 NI_7 NS_56 0 1.2570450778367722e-07
GC_7_57 b_7 NI_7 NS_57 0 1.8062233681799193e-03
GC_7_58 b_7 NI_7 NS_58 0 -4.1873044973439797e-04
GC_7_59 b_7 NI_7 NS_59 0 -1.9478748151075685e-03
GC_7_60 b_7 NI_7 NS_60 0 -6.8414348926347816e-04
GC_7_61 b_7 NI_7 NS_61 0 5.4006195305875582e-02
GC_7_62 b_7 NI_7 NS_62 0 -1.2950685875652967e-02
GC_7_63 b_7 NI_7 NS_63 0 6.4029937987056509e-05
GC_7_64 b_7 NI_7 NS_64 0 -1.3925615523518090e-05
GC_7_65 b_7 NI_7 NS_65 0 -1.0941832731372242e-08
GC_7_66 b_7 NI_7 NS_66 0 -1.2992467142314975e-06
GC_7_67 b_7 NI_7 NS_67 0 -1.9793462077714163e-03
GC_7_68 b_7 NI_7 NS_68 0 7.1107688051664526e-03
GC_7_69 b_7 NI_7 NS_69 0 -1.3471689675817196e-02
GC_7_70 b_7 NI_7 NS_70 0 1.9909622325839892e-02
GC_7_71 b_7 NI_7 NS_71 0 -1.8079962437877359e-01
GC_7_72 b_7 NI_7 NS_72 0 5.8437011537389637e-02
GC_7_73 b_7 NI_7 NS_73 0 -2.5853269315465933e-04
GC_7_74 b_7 NI_7 NS_74 0 8.8787222915376671e-05
GC_7_75 b_7 NI_7 NS_75 0 6.3383867632676292e-08
GC_7_76 b_7 NI_7 NS_76 0 1.5605813858928027e-07
GC_7_77 b_7 NI_7 NS_77 0 -3.0132538012730931e-02
GC_7_78 b_7 NI_7 NS_78 0 -6.1640990378285562e-02
GC_7_79 b_7 NI_7 NS_79 0 8.0265181552842249e-02
GC_7_80 b_7 NI_7 NS_80 0 -1.0161798405703767e-01
GC_7_81 b_7 NI_7 NS_81 0 -7.4389151567008918e-03
GC_7_82 b_7 NI_7 NS_82 0 -4.9138777217378011e-03
GC_7_83 b_7 NI_7 NS_83 0 -1.6817384065761045e-05
GC_7_84 b_7 NI_7 NS_84 0 -2.5022361363910723e-06
GC_7_85 b_7 NI_7 NS_85 0 -2.4058518591219245e-09
GC_7_86 b_7 NI_7 NS_86 0 -4.1377432453105000e-07
GC_7_87 b_7 NI_7 NS_87 0 1.8820577961478513e-03
GC_7_88 b_7 NI_7 NS_88 0 -1.2540780764960473e-02
GC_7_89 b_7 NI_7 NS_89 0 6.8112731294929603e-03
GC_7_90 b_7 NI_7 NS_90 0 1.1346674950468434e-02
GC_7_91 b_7 NI_7 NS_91 0 -1.6924590376648182e-03
GC_7_92 b_7 NI_7 NS_92 0 1.3501145375518274e-03
GC_7_93 b_7 NI_7 NS_93 0 -5.4832940157079633e-06
GC_7_94 b_7 NI_7 NS_94 0 1.1955097696854427e-08
GC_7_95 b_7 NI_7 NS_95 0 2.0709798140686388e-09
GC_7_96 b_7 NI_7 NS_96 0 1.2442755878511398e-07
GC_7_97 b_7 NI_7 NS_97 0 1.8364686691238151e-03
GC_7_98 b_7 NI_7 NS_98 0 -4.4010368481353423e-04
GC_7_99 b_7 NI_7 NS_99 0 -2.0382501866954865e-03
GC_7_100 b_7 NI_7 NS_100 0 -7.6015298818943029e-04
GC_7_101 b_7 NI_7 NS_101 0 -2.7971151411519610e-03
GC_7_102 b_7 NI_7 NS_102 0 -5.7453843688917879e-04
GC_7_103 b_7 NI_7 NS_103 0 -2.2963943578185903e-06
GC_7_104 b_7 NI_7 NS_104 0 5.4353195222753733e-08
GC_7_105 b_7 NI_7 NS_105 0 1.0753259742356695e-10
GC_7_106 b_7 NI_7 NS_106 0 -3.1802393509729266e-08
GC_7_107 b_7 NI_7 NS_107 0 5.7239651384455455e-04
GC_7_108 b_7 NI_7 NS_108 0 -1.1832259322205898e-03
GC_7_109 b_7 NI_7 NS_109 0 2.0484150784670090e-03
GC_7_110 b_7 NI_7 NS_110 0 -7.4558009810014590e-05
GC_7_111 b_7 NI_7 NS_111 0 4.4837993440729763e-04
GC_7_112 b_7 NI_7 NS_112 0 1.7425289508940180e-03
GC_7_113 b_7 NI_7 NS_113 0 2.5838351734011850e-06
GC_7_114 b_7 NI_7 NS_114 0 6.8654595964541843e-08
GC_7_115 b_7 NI_7 NS_115 0 -1.1307784451882576e-10
GC_7_116 b_7 NI_7 NS_116 0 2.8404287293859545e-08
GC_7_117 b_7 NI_7 NS_117 0 3.2315286124498296e-03
GC_7_118 b_7 NI_7 NS_118 0 -2.7458806292783458e-04
GC_7_119 b_7 NI_7 NS_119 0 -5.7926779116929403e-03
GC_7_120 b_7 NI_7 NS_120 0 -1.0206835391601407e-03
GD_7_1 b_7 NI_7 NA_1 0 4.3529775617166675e-04
GD_7_2 b_7 NI_7 NA_2 0 -1.3166542884561320e-04
GD_7_3 b_7 NI_7 NA_3 0 3.7471263744355775e-03
GD_7_4 b_7 NI_7 NA_4 0 1.3849076435686723e-04
GD_7_5 b_7 NI_7 NA_5 0 3.0282103036456426e-02
GD_7_6 b_7 NI_7 NA_6 0 3.3251620337900492e-04
GD_7_7 b_7 NI_7 NA_7 0 -1.9509654583231752e-02
GD_7_8 b_7 NI_7 NA_8 0 2.0461884062731261e-02
GD_7_9 b_7 NI_7 NA_9 0 3.0267336313168261e-02
GD_7_10 b_7 NI_7 NA_10 0 3.6458613786765769e-04
GD_7_11 b_7 NI_7 NA_11 0 3.8606665769386384e-03
GD_7_12 b_7 NI_7 NA_12 0 2.3527094979184168e-04
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 1.7512171572988327e-04
GC_8_2 b_8 NI_8 NS_2 0 5.7758963987158138e-04
GC_8_3 b_8 NI_8 NS_3 0 3.8256035183627728e-07
GC_8_4 b_8 NI_8 NS_4 0 5.8909093128057647e-09
GC_8_5 b_8 NI_8 NS_5 0 -2.1145808913900906e-10
GC_8_6 b_8 NI_8 NS_6 0 1.1273506148340423e-09
GC_8_7 b_8 NI_8 NS_7 0 5.7479252341689562e-04
GC_8_8 b_8 NI_8 NS_8 0 7.5485693406342991e-05
GC_8_9 b_8 NI_8 NS_9 0 -1.1516162709818746e-03
GC_8_10 b_8 NI_8 NS_10 0 2.9456704838688692e-04
GC_8_11 b_8 NI_8 NS_11 0 -1.8083805680269159e-03
GC_8_12 b_8 NI_8 NS_12 0 -4.2589675325296254e-04
GC_8_13 b_8 NI_8 NS_13 0 -1.7713896485539640e-06
GC_8_14 b_8 NI_8 NS_14 0 2.3182273074637414e-07
GC_8_15 b_8 NI_8 NS_15 0 2.3510236112728134e-10
GC_8_16 b_8 NI_8 NS_16 0 -4.8108770705629611e-09
GC_8_17 b_8 NI_8 NS_17 0 3.9570368448633568e-04
GC_8_18 b_8 NI_8 NS_18 0 4.5789574721321875e-04
GC_8_19 b_8 NI_8 NS_19 0 1.7011466517145200e-03
GC_8_20 b_8 NI_8 NS_20 0 -1.8054253450967015e-03
GC_8_21 b_8 NI_8 NS_21 0 2.2630995476374629e-04
GC_8_22 b_8 NI_8 NS_22 0 1.9528009480232883e-03
GC_8_23 b_8 NI_8 NS_23 0 2.4633713577156198e-06
GC_8_24 b_8 NI_8 NS_24 0 1.1838736295482264e-07
GC_8_25 b_8 NI_8 NS_25 0 -8.3451289097620632e-11
GC_8_26 b_8 NI_8 NS_26 0 3.2291767275360039e-08
GC_8_27 b_8 NI_8 NS_27 0 3.0097364790043308e-03
GC_8_28 b_8 NI_8 NS_28 0 -1.8752914992742236e-04
GC_8_29 b_8 NI_8 NS_29 0 -5.4027259304871809e-03
GC_8_30 b_8 NI_8 NS_30 0 -5.2429066922317369e-04
GC_8_31 b_8 NI_8 NS_31 0 -2.3322671330819693e-03
GC_8_32 b_8 NI_8 NS_32 0 -7.3299106530160917e-04
GC_8_33 b_8 NI_8 NS_33 0 -2.1712403229267354e-06
GC_8_34 b_8 NI_8 NS_34 0 7.9797619855397459e-09
GC_8_35 b_8 NI_8 NS_35 0 7.8796782395424921e-11
GC_8_36 b_8 NI_8 NS_36 0 -3.5701773202207393e-08
GC_8_37 b_8 NI_8 NS_37 0 5.4029071943898367e-04
GC_8_38 b_8 NI_8 NS_38 0 -1.1407089600036740e-03
GC_8_39 b_8 NI_8 NS_39 0 1.8427149076859011e-03
GC_8_40 b_8 NI_8 NS_40 0 -1.1617820217932944e-04
GC_8_41 b_8 NI_8 NS_41 0 -1.7545992716934914e-03
GC_8_42 b_8 NI_8 NS_42 0 1.3886113187470833e-03
GC_8_43 b_8 NI_8 NS_43 0 -5.3570467780378706e-06
GC_8_44 b_8 NI_8 NS_44 0 -4.7668777811152306e-09
GC_8_45 b_8 NI_8 NS_45 0 2.0763013949805005e-09
GC_8_46 b_8 NI_8 NS_46 0 1.2570424061425725e-07
GC_8_47 b_8 NI_8 NS_47 0 1.8063163299997973e-03
GC_8_48 b_8 NI_8 NS_48 0 -4.1865530881807976e-04
GC_8_49 b_8 NI_8 NS_49 0 -1.9477700115534855e-03
GC_8_50 b_8 NI_8 NS_50 0 -6.8416278358347836e-04
GC_8_51 b_8 NI_8 NS_51 0 -7.1335350725222563e-03
GC_8_52 b_8 NI_8 NS_52 0 -4.9995367140875154e-03
GC_8_53 b_8 NI_8 NS_53 0 -1.6852299141023232e-05
GC_8_54 b_8 NI_8 NS_54 0 -2.5007847077580000e-06
GC_8_55 b_8 NI_8 NS_55 0 -2.4106580984269951e-09
GC_8_56 b_8 NI_8 NS_56 0 -4.1484901461924044e-07
GC_8_57 b_8 NI_8 NS_57 0 1.8568840199841255e-03
GC_8_58 b_8 NI_8 NS_58 0 -1.2583849639531257e-02
GC_8_59 b_8 NI_8 NS_59 0 6.6065037028949581e-03
GC_8_60 b_8 NI_8 NS_60 0 1.1379025617293689e-02
GC_8_61 b_8 NI_8 NS_61 0 -1.8080058254264517e-01
GC_8_62 b_8 NI_8 NS_62 0 5.8437135541841746e-02
GC_8_63 b_8 NI_8 NS_63 0 -2.5853168604275960e-04
GC_8_64 b_8 NI_8 NS_64 0 8.8786873288582033e-05
GC_8_65 b_8 NI_8 NS_65 0 6.3383578555193156e-08
GC_8_66 b_8 NI_8 NS_66 0 1.5607551915965793e-07
GC_8_67 b_8 NI_8 NS_67 0 -3.0132214468935811e-02
GC_8_68 b_8 NI_8 NS_68 0 -6.1641107205481938e-02
GC_8_69 b_8 NI_8 NS_69 0 8.0265417551285703e-02
GC_8_70 b_8 NI_8 NS_70 0 -1.0161858129957890e-01
GC_8_71 b_8 NI_8 NS_71 0 5.4006195305875582e-02
GC_8_72 b_8 NI_8 NS_72 0 -1.2950685875652967e-02
GC_8_73 b_8 NI_8 NS_73 0 6.4029937987056509e-05
GC_8_74 b_8 NI_8 NS_74 0 -1.3925615523518090e-05
GC_8_75 b_8 NI_8 NS_75 0 -1.0941832731372242e-08
GC_8_76 b_8 NI_8 NS_76 0 -1.2992467142314975e-06
GC_8_77 b_8 NI_8 NS_77 0 -1.9793462077714163e-03
GC_8_78 b_8 NI_8 NS_78 0 7.1107688051664526e-03
GC_8_79 b_8 NI_8 NS_79 0 -1.3471689675817196e-02
GC_8_80 b_8 NI_8 NS_80 0 1.9909622325839892e-02
GC_8_81 b_8 NI_8 NS_81 0 -1.6903764994324194e-03
GC_8_82 b_8 NI_8 NS_82 0 1.3497356703658829e-03
GC_8_83 b_8 NI_8 NS_83 0 -5.4845931134731787e-06
GC_8_84 b_8 NI_8 NS_84 0 1.2152326202624217e-08
GC_8_85 b_8 NI_8 NS_85 0 2.0709716355972255e-09
GC_8_86 b_8 NI_8 NS_86 0 1.2442440059572878e-07
GC_8_87 b_8 NI_8 NS_87 0 1.8367156228869719e-03
GC_8_88 b_8 NI_8 NS_88 0 -4.3936972050341447e-04
GC_8_89 b_8 NI_8 NS_89 0 -2.0387702150236192e-03
GC_8_90 b_8 NI_8 NS_90 0 -7.5956069986714346e-04
GC_8_91 b_8 NI_8 NS_91 0 -7.4460956606887500e-03
GC_8_92 b_8 NI_8 NS_92 0 -4.9120728687247319e-03
GC_8_93 b_8 NI_8 NS_93 0 -1.6829168807819534e-05
GC_8_94 b_8 NI_8 NS_94 0 -2.5002142732340761e-06
GC_8_95 b_8 NI_8 NS_95 0 -2.4057391622560119e-09
GC_8_96 b_8 NI_8 NS_96 0 -4.1381043907329940e-07
GC_8_97 b_8 NI_8 NS_97 0 1.8829292403328706e-03
GC_8_98 b_8 NI_8 NS_98 0 -1.2541882493978097e-02
GC_8_99 b_8 NI_8 NS_99 0 6.8135168116135406e-03
GC_8_100 b_8 NI_8 NS_100 0 1.1344690691195224e-02
GC_8_101 b_8 NI_8 NS_101 0 4.4312076802818063e-04
GC_8_102 b_8 NI_8 NS_102 0 1.7434320196114870e-03
GC_8_103 b_8 NI_8 NS_103 0 2.5874752096212791e-06
GC_8_104 b_8 NI_8 NS_104 0 6.8072367311414042e-08
GC_8_105 b_8 NI_8 NS_105 0 -1.1315508052930240e-10
GC_8_106 b_8 NI_8 NS_106 0 2.8408045874434463e-08
GC_8_107 b_8 NI_8 NS_107 0 3.2307394077003889e-03
GC_8_108 b_8 NI_8 NS_108 0 -2.7665463265152279e-04
GC_8_109 b_8 NI_8 NS_109 0 -5.7915279978725774e-03
GC_8_110 b_8 NI_8 NS_110 0 -1.0222266352664159e-03
GC_8_111 b_8 NI_8 NS_111 0 -2.7874755153256664e-03
GC_8_112 b_8 NI_8 NS_112 0 -5.7624033058046795e-04
GC_8_113 b_8 NI_8 NS_113 0 -2.2810455880852200e-06
GC_8_114 b_8 NI_8 NS_114 0 5.2123773590983789e-08
GC_8_115 b_8 NI_8 NS_115 0 1.0695911914792542e-10
GC_8_116 b_8 NI_8 NS_116 0 -3.1749185512537881e-08
GC_8_117 b_8 NI_8 NS_117 0 5.7212685300815961e-04
GC_8_118 b_8 NI_8 NS_118 0 -1.1815065721432140e-03
GC_8_119 b_8 NI_8 NS_119 0 2.0451472588779804e-03
GC_8_120 b_8 NI_8 NS_120 0 -7.0424879579449208e-05
GD_8_1 b_8 NI_8 NA_1 0 -1.3079564415693494e-04
GD_8_2 b_8 NI_8 NA_2 0 4.3463287813285756e-04
GD_8_3 b_8 NI_8 NA_3 0 1.3886656467954533e-04
GD_8_4 b_8 NI_8 NA_4 0 3.7468483141920228e-03
GD_8_5 b_8 NI_8 NA_5 0 3.3234763115963739e-04
GD_8_6 b_8 NI_8 NA_6 0 3.0282091253999912e-02
GD_8_7 b_8 NI_8 NA_7 0 2.0462020752404206e-02
GD_8_8 b_8 NI_8 NA_8 0 -1.9509654583231752e-02
GD_8_9 b_8 NI_8 NA_9 0 3.6349746612773277e-04
GD_8_10 b_8 NI_8 NA_10 0 3.0268686047503914e-02
GD_8_11 b_8 NI_8 NA_11 0 2.3842103440352533e-04
GD_8_12 b_8 NI_8 NA_12 0 3.8583924691778272e-03
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 -1.5096395792225386e-04
GC_9_2 b_9 NI_9 NS_2 0 -2.5228975229088128e-04
GC_9_3 b_9 NI_9 NS_3 0 -3.1553261516787772e-07
GC_9_4 b_9 NI_9 NS_4 0 4.4725458220605296e-08
GC_9_5 b_9 NI_9 NS_5 0 1.0764361019824762e-10
GC_9_6 b_9 NI_9 NS_6 0 5.1109993696245445e-11
GC_9_7 b_9 NI_9 NS_7 0 8.6978354446912569e-05
GC_9_8 b_9 NI_9 NS_8 0 1.6471009113755645e-04
GC_9_9 b_9 NI_9 NS_9 0 3.1642735768477100e-04
GC_9_10 b_9 NI_9 NS_10 0 -5.7184015220568447e-04
GC_9_11 b_9 NI_9 NS_11 0 -6.8110663934043062e-05
GC_9_12 b_9 NI_9 NS_12 0 3.4263860861849440e-04
GC_9_13 b_9 NI_9 NS_13 0 -2.0423855983249287e-08
GC_9_14 b_9 NI_9 NS_14 0 1.4259177777872977e-08
GC_9_15 b_9 NI_9 NS_15 0 -1.0175926760562784e-10
GC_9_16 b_9 NI_9 NS_16 0 -9.1086072048921074e-10
GC_9_17 b_9 NI_9 NS_17 0 -5.6814754007499051e-05
GC_9_18 b_9 NI_9 NS_18 0 1.2051224837869429e-04
GC_9_19 b_9 NI_9 NS_19 0 2.1893798623872612e-05
GC_9_20 b_9 NI_9 NS_20 0 5.8520957279704835e-04
GC_9_21 b_9 NI_9 NS_21 0 -1.4365981285533625e-03
GC_9_22 b_9 NI_9 NS_22 0 -5.2554836834912196e-04
GC_9_23 b_9 NI_9 NS_23 0 -1.6806885297593111e-06
GC_9_24 b_9 NI_9 NS_24 0 2.0769313928527144e-07
GC_9_25 b_9 NI_9 NS_25 0 2.2668288943092759e-10
GC_9_26 b_9 NI_9 NS_26 0 -5.5164355151380002e-09
GC_9_27 b_9 NI_9 NS_27 0 3.6567678318688264e-04
GC_9_28 b_9 NI_9 NS_28 0 4.2773342079281218e-04
GC_9_29 b_9 NI_9 NS_29 0 1.4813104413553093e-03
GC_9_30 b_9 NI_9 NS_30 0 -1.7482970824392419e-03
GC_9_31 b_9 NI_9 NS_31 0 8.0853503837957744e-05
GC_9_32 b_9 NI_9 NS_32 0 6.1961854941422609e-04
GC_9_33 b_9 NI_9 NS_33 0 4.5901077523111817e-07
GC_9_34 b_9 NI_9 NS_34 0 1.6709687958626685e-09
GC_9_35 b_9 NI_9 NS_35 0 -2.0540839151132718e-10
GC_9_36 b_9 NI_9 NS_36 0 2.2654604492252261e-09
GC_9_37 b_9 NI_9 NS_37 0 5.4524373557005652e-04
GC_9_38 b_9 NI_9 NS_38 0 8.3637357368031027e-05
GC_9_39 b_9 NI_9 NS_39 0 -1.0621391184145259e-03
GC_9_40 b_9 NI_9 NS_40 0 3.5110894111764761e-04
GC_9_41 b_9 NI_9 NS_41 0 -2.3329145978155381e-03
GC_9_42 b_9 NI_9 NS_42 0 -7.3285603310363587e-04
GC_9_43 b_9 NI_9 NS_43 0 -2.1737376380831570e-06
GC_9_44 b_9 NI_9 NS_44 0 8.6499861841235125e-09
GC_9_45 b_9 NI_9 NS_45 0 7.8813825396023021e-11
GC_9_46 b_9 NI_9 NS_46 0 -3.5704257177941657e-08
GC_9_47 b_9 NI_9 NS_47 0 5.4038413931800340e-04
GC_9_48 b_9 NI_9 NS_48 0 -1.1407863730068064e-03
GC_9_49 b_9 NI_9 NS_49 0 1.8429279956086277e-03
GC_9_50 b_9 NI_9 NS_50 0 -1.1642622848298793e-04
GC_9_51 b_9 NI_9 NS_51 0 2.2571822946922183e-04
GC_9_52 b_9 NI_9 NS_52 0 1.9527876275770560e-03
GC_9_53 b_9 NI_9 NS_53 0 2.4667422030195401e-06
GC_9_54 b_9 NI_9 NS_54 0 1.1763930329096830e-07
GC_9_55 b_9 NI_9 NS_55 0 -8.3450274923965756e-11
GC_9_56 b_9 NI_9 NS_56 0 3.2296174829919205e-08
GC_9_57 b_9 NI_9 NS_57 0 3.0097804134294292e-03
GC_9_58 b_9 NI_9 NS_58 0 -1.8781201218584880e-04
GC_9_59 b_9 NI_9 NS_59 0 -5.4027133649887319e-03
GC_9_60 b_9 NI_9 NS_60 0 -5.2475450255814527e-04
GC_9_61 b_9 NI_9 NS_61 0 -7.4460956606887500e-03
GC_9_62 b_9 NI_9 NS_62 0 -4.9120728687247319e-03
GC_9_63 b_9 NI_9 NS_63 0 -1.6829168807819534e-05
GC_9_64 b_9 NI_9 NS_64 0 -2.5002142732340761e-06
GC_9_65 b_9 NI_9 NS_65 0 -2.4057391622560119e-09
GC_9_66 b_9 NI_9 NS_66 0 -4.1381043907329940e-07
GC_9_67 b_9 NI_9 NS_67 0 1.8829292403328706e-03
GC_9_68 b_9 NI_9 NS_68 0 -1.2541882493978097e-02
GC_9_69 b_9 NI_9 NS_69 0 6.8135168116135406e-03
GC_9_70 b_9 NI_9 NS_70 0 1.1344690691195224e-02
GC_9_71 b_9 NI_9 NS_71 0 -1.6924590376648182e-03
GC_9_72 b_9 NI_9 NS_72 0 1.3501145375518274e-03
GC_9_73 b_9 NI_9 NS_73 0 -5.4832940157079633e-06
GC_9_74 b_9 NI_9 NS_74 0 1.1955097696854427e-08
GC_9_75 b_9 NI_9 NS_75 0 2.0709798140686388e-09
GC_9_76 b_9 NI_9 NS_76 0 1.2442755878511398e-07
GC_9_77 b_9 NI_9 NS_77 0 1.8364686691238151e-03
GC_9_78 b_9 NI_9 NS_78 0 -4.4010368481353423e-04
GC_9_79 b_9 NI_9 NS_79 0 -2.0382501866954865e-03
GC_9_80 b_9 NI_9 NS_80 0 -7.6015298818943029e-04
GC_9_81 b_9 NI_9 NS_81 0 5.3616896777345914e-02
GC_9_82 b_9 NI_9 NS_82 0 -1.2804981338122679e-02
GC_9_83 b_9 NI_9 NS_83 0 6.3940330049350603e-05
GC_9_84 b_9 NI_9 NS_84 0 -1.3871628216598860e-05
GC_9_85 b_9 NI_9 NS_85 0 -1.0851120457540901e-08
GC_9_86 b_9 NI_9 NS_86 0 -1.2971656785465817e-06
GC_9_87 b_9 NI_9 NS_87 0 -1.9507989708983128e-03
GC_9_88 b_9 NI_9 NS_88 0 7.0862911648213005e-03
GC_9_89 b_9 NI_9 NS_89 0 -1.3281339308975987e-02
GC_9_90 b_9 NI_9 NS_90 0 1.9983242328530611e-02
GC_9_91 b_9 NI_9 NS_91 0 -1.8056478863254852e-01
GC_9_92 b_9 NI_9 NS_92 0 5.8222882764336167e-02
GC_9_93 b_9 NI_9 NS_93 0 -2.5838659030338906e-04
GC_9_94 b_9 NI_9 NS_94 0 8.8719746021195288e-05
GC_9_95 b_9 NI_9 NS_95 0 6.3340891029122170e-08
GC_9_96 b_9 NI_9 NS_96 0 1.5314824115175121e-07
GC_9_97 b_9 NI_9 NS_97 0 -2.9914530128223038e-02
GC_9_98 b_9 NI_9 NS_98 0 -6.1730431645545744e-02
GC_9_99 b_9 NI_9 NS_99 0 7.9867646357335675e-02
GC_9_100 b_9 NI_9 NS_100 0 -1.0211222722876941e-01
GC_9_101 b_9 NI_9 NS_101 0 -7.0566514973206523e-03
GC_9_102 b_9 NI_9 NS_102 0 -4.4826525389356281e-03
GC_9_103 b_9 NI_9 NS_103 0 -1.6086015613505065e-05
GC_9_104 b_9 NI_9 NS_104 0 -2.4816704104033053e-06
GC_9_105 b_9 NI_9 NS_105 0 -2.2943978362392909e-09
GC_9_106 b_9 NI_9 NS_106 0 -3.9506621399113991e-07
GC_9_107 b_9 NI_9 NS_107 0 1.7173757127493898e-03
GC_9_108 b_9 NI_9 NS_108 0 -1.3406237240908239e-02
GC_9_109 b_9 NI_9 NS_109 0 5.8866758738304733e-03
GC_9_110 b_9 NI_9 NS_110 0 1.2986108939997553e-02
GC_9_111 b_9 NI_9 NS_111 0 -1.3064872164159451e-03
GC_9_112 b_9 NI_9 NS_112 0 1.1610391636487968e-03
GC_9_113 b_9 NI_9 NS_113 0 -5.2056773045755629e-06
GC_9_114 b_9 NI_9 NS_114 0 -1.3609195858071407e-07
GC_9_115 b_9 NI_9 NS_115 0 1.8849426214244058e-09
GC_9_116 b_9 NI_9 NS_116 0 1.0944607695530042e-07
GC_9_117 b_9 NI_9 NS_117 0 2.1790816182797870e-03
GC_9_118 b_9 NI_9 NS_118 0 -5.3341201018435546e-04
GC_9_119 b_9 NI_9 NS_119 0 -2.6659889838270751e-03
GC_9_120 b_9 NI_9 NS_120 0 -1.2463735393863486e-03
GD_9_1 b_9 NI_9 NA_1 0 3.9293699158599537e-05
GD_9_2 b_9 NI_9 NA_2 0 -1.6522435545847635e-04
GD_9_3 b_9 NI_9 NA_3 0 4.2053241529844932e-04
GD_9_4 b_9 NI_9 NA_4 0 -1.3536897167817916e-04
GD_9_5 b_9 NI_9 NA_5 0 3.7469884696672427e-03
GD_9_6 b_9 NI_9 NA_6 0 1.3931914091957427e-04
GD_9_7 b_9 NI_9 NA_7 0 3.0268686047503914e-02
GD_9_8 b_9 NI_9 NA_8 0 3.6458613786765769e-04
GD_9_9 b_9 NI_9 NA_9 0 -1.9437702687596162e-02
GD_9_10 b_9 NI_9 NA_10 0 2.0560518467129904e-02
GD_9_11 b_9 NI_9 NA_11 0 3.1107793494345781e-02
GD_9_12 b_9 NI_9 NA_12 0 3.7194425217160118e-04
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 -6.8799613938542152e-05
GC_10_2 b_10 NI_10 NS_2 0 3.4277166450000614e-04
GC_10_3 b_10 NI_10 NS_3 0 -2.0714519939758428e-08
GC_10_4 b_10 NI_10 NS_4 0 1.4344062583856994e-08
GC_10_5 b_10 NI_10 NS_5 0 -1.0174748616111340e-10
GC_10_6 b_10 NI_10 NS_6 0 -9.1239918190250832e-10
GC_10_7 b_10 NI_10 NS_7 0 -5.6845011500187794e-05
GC_10_8 b_10 NI_10 NS_8 0 1.2033342580408023e-04
GC_10_9 b_10 NI_10 NS_9 0 2.2093533547946310e-05
GC_10_10 b_10 NI_10 NS_10 0 5.8499452995802725e-04
GC_10_11 b_10 NI_10 NS_11 0 -1.5078854548084765e-04
GC_10_12 b_10 NI_10 NS_12 0 -2.5231272645266737e-04
GC_10_13 b_10 NI_10 NS_13 0 -3.1462006780480187e-07
GC_10_14 b_10 NI_10 NS_14 0 4.4620488362912420e-08
GC_10_15 b_10 NI_10 NS_15 0 1.0763234468196428e-10
GC_10_16 b_10 NI_10 NS_16 0 5.2939954377662918e-11
GC_10_17 b_10 NI_10 NS_17 0 8.6961757586850603e-05
GC_10_18 b_10 NI_10 NS_18 0 1.6484274725236408e-04
GC_10_19 b_10 NI_10 NS_19 0 3.1650314601421183e-04
GC_10_20 b_10 NI_10 NS_20 0 -5.7170825778301215e-04
GC_10_21 b_10 NI_10 NS_21 0 8.1654121462430338e-05
GC_10_22 b_10 NI_10 NS_22 0 6.1942409181479289e-04
GC_10_23 b_10 NI_10 NS_23 0 4.5980700814682754e-07
GC_10_24 b_10 NI_10 NS_24 0 1.5473232055628190e-09
GC_10_25 b_10 NI_10 NS_25 0 -2.0541669074526852e-10
GC_10_26 b_10 NI_10 NS_26 0 2.2671228369173445e-09
GC_10_27 b_10 NI_10 NS_27 0 5.4512433979936878e-04
GC_10_28 b_10 NI_10 NS_28 0 8.3645148241201910e-05
GC_10_29 b_10 NI_10 NS_29 0 -1.0624996024421482e-03
GC_10_30 b_10 NI_10 NS_30 0 3.5134323036855632e-04
GC_10_31 b_10 NI_10 NS_31 0 -1.4365666755094526e-03
GC_10_32 b_10 NI_10 NS_32 0 -5.2555390307240787e-04
GC_10_33 b_10 NI_10 NS_33 0 -1.6806776345275893e-06
GC_10_34 b_10 NI_10 NS_34 0 2.0769026188550992e-07
GC_10_35 b_10 NI_10 NS_35 0 2.2668297248944703e-10
GC_10_36 b_10 NI_10 NS_36 0 -5.5163287780851915e-09
GC_10_37 b_10 NI_10 NS_37 0 3.6567389653507991e-04
GC_10_38 b_10 NI_10 NS_38 0 4.2773835993569132e-04
GC_10_39 b_10 NI_10 NS_39 0 1.4813020334029758e-03
GC_10_40 b_10 NI_10 NS_40 0 -1.7482834881565495e-03
GC_10_41 b_10 NI_10 NS_41 0 2.2498716385862400e-04
GC_10_42 b_10 NI_10 NS_42 0 1.9530786948455984e-03
GC_10_43 b_10 NI_10 NS_43 0 2.4631372121652609e-06
GC_10_44 b_10 NI_10 NS_44 0 1.1825817633892398e-07
GC_10_45 b_10 NI_10 NS_45 0 -8.3403319346910024e-11
GC_10_46 b_10 NI_10 NS_46 0 3.2286921814126651e-08
GC_10_47 b_10 NI_10 NS_47 0 3.0098587914049930e-03
GC_10_48 b_10 NI_10 NS_48 0 -1.8773057630928588e-04
GC_10_49 b_10 NI_10 NS_49 0 -5.4023417777550094e-03
GC_10_50 b_10 NI_10 NS_50 0 -5.2475672159504536e-04
GC_10_51 b_10 NI_10 NS_51 0 -2.3329916798764672e-03
GC_10_52 b_10 NI_10 NS_52 0 -7.3276860499570150e-04
GC_10_53 b_10 NI_10 NS_53 0 -2.1754894548739566e-06
GC_10_54 b_10 NI_10 NS_54 0 8.9813158443094226e-09
GC_10_55 b_10 NI_10 NS_55 0 7.8802453510202652e-11
GC_10_56 b_10 NI_10 NS_56 0 -3.5713227815655763e-08
GC_10_57 b_10 NI_10 NS_57 0 5.4026267907607913e-04
GC_10_58 b_10 NI_10 NS_58 0 -1.1406344561067309e-03
GC_10_59 b_10 NI_10 NS_59 0 1.8430652824974693e-03
GC_10_60 b_10 NI_10 NS_60 0 -1.1628231309278826e-04
GC_10_61 b_10 NI_10 NS_61 0 -1.6903764994324194e-03
GC_10_62 b_10 NI_10 NS_62 0 1.3497356703658829e-03
GC_10_63 b_10 NI_10 NS_63 0 -5.4845931134731787e-06
GC_10_64 b_10 NI_10 NS_64 0 1.2152326202624217e-08
GC_10_65 b_10 NI_10 NS_65 0 2.0709716355972255e-09
GC_10_66 b_10 NI_10 NS_66 0 1.2442440059572878e-07
GC_10_67 b_10 NI_10 NS_67 0 1.8367156228869719e-03
GC_10_68 b_10 NI_10 NS_68 0 -4.3936972050341447e-04
GC_10_69 b_10 NI_10 NS_69 0 -2.0387702150236192e-03
GC_10_70 b_10 NI_10 NS_70 0 -7.5956069986714346e-04
GC_10_71 b_10 NI_10 NS_71 0 -7.4389151567008918e-03
GC_10_72 b_10 NI_10 NS_72 0 -4.9138777217378011e-03
GC_10_73 b_10 NI_10 NS_73 0 -1.6817384065761045e-05
GC_10_74 b_10 NI_10 NS_74 0 -2.5022361363910723e-06
GC_10_75 b_10 NI_10 NS_75 0 -2.4058518591219245e-09
GC_10_76 b_10 NI_10 NS_76 0 -4.1377432453105000e-07
GC_10_77 b_10 NI_10 NS_77 0 1.8820577961478513e-03
GC_10_78 b_10 NI_10 NS_78 0 -1.2540780764960473e-02
GC_10_79 b_10 NI_10 NS_79 0 6.8112731294929603e-03
GC_10_80 b_10 NI_10 NS_80 0 1.1346674950468434e-02
GC_10_81 b_10 NI_10 NS_81 0 -1.8053487835711060e-01
GC_10_82 b_10 NI_10 NS_82 0 5.8214972360122470e-02
GC_10_83 b_10 NI_10 NS_83 0 -2.5831896498885434e-04
GC_10_84 b_10 NI_10 NS_84 0 8.8704014865213196e-05
GC_10_85 b_10 NI_10 NS_85 0 6.3332082666254789e-08
GC_10_86 b_10 NI_10 NS_86 0 1.5369414677095390e-07
GC_10_87 b_10 NI_10 NS_87 0 -2.9914529398979435e-02
GC_10_88 b_10 NI_10 NS_88 0 -6.1725786533034108e-02
GC_10_89 b_10 NI_10 NS_89 0 7.9857129787514899e-02
GC_10_90 b_10 NI_10 NS_90 0 -1.0210630810063671e-01
GC_10_91 b_10 NI_10 NS_91 0 5.3616896777345914e-02
GC_10_92 b_10 NI_10 NS_92 0 -1.2804981338122679e-02
GC_10_93 b_10 NI_10 NS_93 0 6.3940330049350603e-05
GC_10_94 b_10 NI_10 NS_94 0 -1.3871628216598860e-05
GC_10_95 b_10 NI_10 NS_95 0 -1.0851120457540901e-08
GC_10_96 b_10 NI_10 NS_96 0 -1.2971656785465817e-06
GC_10_97 b_10 NI_10 NS_97 0 -1.9507989708983128e-03
GC_10_98 b_10 NI_10 NS_98 0 7.0862911648213005e-03
GC_10_99 b_10 NI_10 NS_99 0 -1.3281339308975987e-02
GC_10_100 b_10 NI_10 NS_100 0 1.9983242328530611e-02
GC_10_101 b_10 NI_10 NS_101 0 -1.3061125580791548e-03
GC_10_102 b_10 NI_10 NS_102 0 1.1609039661503548e-03
GC_10_103 b_10 NI_10 NS_103 0 -5.2046723080868838e-06
GC_10_104 b_10 NI_10 NS_104 0 -1.3619515854241348e-07
GC_10_105 b_10 NI_10 NS_105 0 1.8849527256255734e-09
GC_10_106 b_10 NI_10 NS_106 0 1.0944656981071299e-07
GC_10_107 b_10 NI_10 NS_107 0 2.1789648288941632e-03
GC_10_108 b_10 NI_10 NS_108 0 -5.3350899546166777e-04
GC_10_109 b_10 NI_10 NS_109 0 -2.6662046367079903e-03
GC_10_110 b_10 NI_10 NS_110 0 -1.2463188652477935e-03
GC_10_111 b_10 NI_10 NS_111 0 -7.0303427409601120e-03
GC_10_112 b_10 NI_10 NS_112 0 -4.4850612205423511e-03
GC_10_113 b_10 NI_10 NS_113 0 -1.6070237758281345e-05
GC_10_114 b_10 NI_10 NS_114 0 -2.4814686871585115e-06
GC_10_115 b_10 NI_10 NS_115 0 -2.2962574848161942e-09
GC_10_116 b_10 NI_10 NS_116 0 -3.9507264247438605e-07
GC_10_117 b_10 NI_10 NS_117 0 1.7173950787024879e-03
GC_10_118 b_10 NI_10 NS_118 0 -1.3398723896416800e-02
GC_10_119 b_10 NI_10 NS_119 0 5.8795964257928992e-03
GC_10_120 b_10 NI_10 NS_120 0 1.3002086464105812e-02
GD_10_1 b_10 NI_10 NA_1 0 -1.6493460942386661e-04
GD_10_2 b_10 NI_10 NA_2 0 3.9136900122655807e-05
GD_10_3 b_10 NI_10 NA_3 0 -1.3541351404501971e-04
GD_10_4 b_10 NI_10 NA_4 0 4.2051920717500632e-04
GD_10_5 b_10 NI_10 NA_5 0 1.3932018935636532e-04
GD_10_6 b_10 NI_10 NA_6 0 3.7471538655471826e-03
GD_10_7 b_10 NI_10 NA_7 0 3.6349746612773277e-04
GD_10_8 b_10 NI_10 NA_8 0 3.0267336313168261e-02
GD_10_9 b_10 NI_10 NA_9 0 2.0551894646332811e-02
GD_10_10 b_10 NI_10 NA_10 0 -1.9437702687596162e-02
GD_10_11 b_10 NI_10 NA_11 0 3.7202435221328988e-04
GD_10_12 b_10 NI_10 NA_12 0 3.1099351267036241e-02
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 2.9949897747088552e-04
GC_11_2 b_11 NI_11 NS_2 0 -1.6297325967750130e-04
GC_11_3 b_11 NI_11 NS_3 0 3.2141973059138642e-08
GC_11_4 b_11 NI_11 NS_4 0 -1.0197462899819804e-08
GC_11_5 b_11 NI_11 NS_5 0 3.8755308880426955e-11
GC_11_6 b_11 NI_11 NS_6 0 9.2510731016750194e-10
GC_11_7 b_11 NI_11 NS_7 0 -2.7765464681837651e-06
GC_11_8 b_11 NI_11 NS_8 0 1.7958537920894944e-05
GC_11_9 b_11 NI_11 NS_9 0 -1.1314121306781161e-04
GC_11_10 b_11 NI_11 NS_10 0 -1.0759536368278283e-04
GC_11_11 b_11 NI_11 NS_11 0 -9.7220809498346766e-05
GC_11_12 b_11 NI_11 NS_12 0 1.3616955559621417e-04
GC_11_13 b_11 NI_11 NS_13 0 -8.0289895940418349e-09
GC_11_14 b_11 NI_11 NS_14 0 8.0786405512087354e-09
GC_11_15 b_11 NI_11 NS_15 0 -3.8739547827781783e-11
GC_11_16 b_11 NI_11 NS_16 0 -8.7101973761499855e-10
GC_11_17 b_11 NI_11 NS_17 0 -4.7013291556070843e-05
GC_11_18 b_11 NI_11 NS_18 0 4.5272529151951507e-05
GC_11_19 b_11 NI_11 NS_19 0 8.8826450853963002e-05
GC_11_20 b_11 NI_11 NS_20 0 2.2568047343720499e-04
GC_11_21 b_11 NI_11 NS_21 0 -1.5072974180017139e-04
GC_11_22 b_11 NI_11 NS_22 0 -2.5231601036312034e-04
GC_11_23 b_11 NI_11 NS_23 0 -3.1459273271146477e-07
GC_11_24 b_11 NI_11 NS_24 0 4.4593311782414919e-08
GC_11_25 b_11 NI_11 NS_25 0 1.0762446501307339e-10
GC_11_26 b_11 NI_11 NS_26 0 5.3288867417633135e-11
GC_11_27 b_11 NI_11 NS_27 0 8.6952963580351079e-05
GC_11_28 b_11 NI_11 NS_28 0 1.6486089740420866e-04
GC_11_29 b_11 NI_11 NS_29 0 3.1649716165064063e-04
GC_11_30 b_11 NI_11 NS_30 0 -5.7166537939438609e-04
GC_11_31 b_11 NI_11 NS_31 0 -6.8047032396455873e-05
GC_11_32 b_11 NI_11 NS_32 0 3.4261133561112981e-04
GC_11_33 b_11 NI_11 NS_33 0 -2.0319496336951487e-08
GC_11_34 b_11 NI_11 NS_34 0 1.4268774072850567e-08
GC_11_35 b_11 NI_11 NS_35 0 -1.0175329619432754e-10
GC_11_36 b_11 NI_11 NS_36 0 -9.1092915343631042e-10
GC_11_37 b_11 NI_11 NS_37 0 -5.6817933891895275e-05
GC_11_38 b_11 NI_11 NS_38 0 1.2050288604751119e-04
GC_11_39 b_11 NI_11 NS_39 0 2.1853855541131872e-05
GC_11_40 b_11 NI_11 NS_40 0 5.8520010637099862e-04
GC_11_41 b_11 NI_11 NS_41 0 -1.8082139400216366e-03
GC_11_42 b_11 NI_11 NS_42 0 -4.2594882966600993e-04
GC_11_43 b_11 NI_11 NS_43 0 -1.7706788427184878e-06
GC_11_44 b_11 NI_11 NS_44 0 2.3157148955476831e-07
GC_11_45 b_11 NI_11 NS_45 0 2.3505527812462354e-10
GC_11_46 b_11 NI_11 NS_46 0 -4.7985459397601332e-09
GC_11_47 b_11 NI_11 NS_47 0 3.9569725122428880e-04
GC_11_48 b_11 NI_11 NS_48 0 4.5790575336839251e-04
GC_11_49 b_11 NI_11 NS_49 0 1.7010822969953400e-03
GC_11_50 b_11 NI_11 NS_50 0 -1.8054030035425629e-03
GC_11_51 b_11 NI_11 NS_51 0 1.7713520644807633e-04
GC_11_52 b_11 NI_11 NS_52 0 5.7711503772868910e-04
GC_11_53 b_11 NI_11 NS_53 0 3.8437197205538283e-07
GC_11_54 b_11 NI_11 NS_54 0 5.6131200511718194e-09
GC_11_55 b_11 NI_11 NS_55 0 -2.1142105692611963e-10
GC_11_56 b_11 NI_11 NS_56 0 1.1233157414133004e-09
GC_11_57 b_11 NI_11 NS_57 0 5.7503237530367470e-04
GC_11_58 b_11 NI_11 NS_58 0 7.6072738321982355e-05
GC_11_59 b_11 NI_11 NS_59 0 -1.1522395821956836e-03
GC_11_60 b_11 NI_11 NS_60 0 2.9493613797594543e-04
GC_11_61 b_11 NI_11 NS_61 0 -2.7874755153256664e-03
GC_11_62 b_11 NI_11 NS_62 0 -5.7624033058046795e-04
GC_11_63 b_11 NI_11 NS_63 0 -2.2810455880852200e-06
GC_11_64 b_11 NI_11 NS_64 0 5.2123773590983789e-08
GC_11_65 b_11 NI_11 NS_65 0 1.0695911914792542e-10
GC_11_66 b_11 NI_11 NS_66 0 -3.1749185512537881e-08
GC_11_67 b_11 NI_11 NS_67 0 5.7212685300815961e-04
GC_11_68 b_11 NI_11 NS_68 0 -1.1815065721432140e-03
GC_11_69 b_11 NI_11 NS_69 0 2.0451472588779804e-03
GC_11_70 b_11 NI_11 NS_70 0 -7.0424879579449208e-05
GC_11_71 b_11 NI_11 NS_71 0 4.4837993440729763e-04
GC_11_72 b_11 NI_11 NS_72 0 1.7425289508940180e-03
GC_11_73 b_11 NI_11 NS_73 0 2.5838351734011850e-06
GC_11_74 b_11 NI_11 NS_74 0 6.8654595964541843e-08
GC_11_75 b_11 NI_11 NS_75 0 -1.1307784451882576e-10
GC_11_76 b_11 NI_11 NS_76 0 2.8404287293859545e-08
GC_11_77 b_11 NI_11 NS_77 0 3.2315286124498296e-03
GC_11_78 b_11 NI_11 NS_78 0 -2.7458806292783458e-04
GC_11_79 b_11 NI_11 NS_79 0 -5.7926779116929403e-03
GC_11_80 b_11 NI_11 NS_80 0 -1.0206835391601407e-03
GC_11_81 b_11 NI_11 NS_81 0 -7.0303427409601120e-03
GC_11_82 b_11 NI_11 NS_82 0 -4.4850612205423511e-03
GC_11_83 b_11 NI_11 NS_83 0 -1.6070237758281345e-05
GC_11_84 b_11 NI_11 NS_84 0 -2.4814686871585115e-06
GC_11_85 b_11 NI_11 NS_85 0 -2.2962574848161942e-09
GC_11_86 b_11 NI_11 NS_86 0 -3.9507264247438605e-07
GC_11_87 b_11 NI_11 NS_87 0 1.7173950787024879e-03
GC_11_88 b_11 NI_11 NS_88 0 -1.3398723896416800e-02
GC_11_89 b_11 NI_11 NS_89 0 5.8795964257928992e-03
GC_11_90 b_11 NI_11 NS_90 0 1.3002086464105812e-02
GC_11_91 b_11 NI_11 NS_91 0 -1.3064872164159451e-03
GC_11_92 b_11 NI_11 NS_92 0 1.1610391636487968e-03
GC_11_93 b_11 NI_11 NS_93 0 -5.2056773045755629e-06
GC_11_94 b_11 NI_11 NS_94 0 -1.3609195858071407e-07
GC_11_95 b_11 NI_11 NS_95 0 1.8849426214244058e-09
GC_11_96 b_11 NI_11 NS_96 0 1.0944607695530042e-07
GC_11_97 b_11 NI_11 NS_97 0 2.1790816182797870e-03
GC_11_98 b_11 NI_11 NS_98 0 -5.3341201018435546e-04
GC_11_99 b_11 NI_11 NS_99 0 -2.6659889838270751e-03
GC_11_100 b_11 NI_11 NS_100 0 -1.2463735393863486e-03
GC_11_101 b_11 NI_11 NS_101 0 5.2859398508041902e-02
GC_11_102 b_11 NI_11 NS_102 0 -1.3064793307874138e-02
GC_11_103 b_11 NI_11 NS_103 0 5.9279854192276102e-05
GC_11_104 b_11 NI_11 NS_104 0 -1.3381643858258897e-05
GC_11_105 b_11 NI_11 NS_105 0 -8.5088331589078162e-09
GC_11_106 b_11 NI_11 NS_106 0 -1.3098075755340869e-06
GC_11_107 b_11 NI_11 NS_107 0 -1.9013630309753474e-03
GC_11_108 b_11 NI_11 NS_108 0 4.2717618170745328e-03
GC_11_109 b_11 NI_11 NS_109 0 -1.3200571729196761e-02
GC_11_110 b_11 NI_11 NS_110 0 2.3506110531105958e-02
GC_11_111 b_11 NI_11 NS_111 0 -1.7979976521573501e-01
GC_11_112 b_11 NI_11 NS_112 0 5.6387839134505131e-02
GC_11_113 b_11 NI_11 NS_113 0 -2.6203975415478906e-04
GC_11_114 b_11 NI_11 NS_114 0 8.7773995915894961e-05
GC_11_115 b_11 NI_11 NS_115 0 6.1884238521284858e-08
GC_11_116 b_11 NI_11 NS_116 0 6.3199890847947142e-08
GC_11_117 b_11 NI_11 NS_117 0 -3.2557282383069340e-02
GC_11_118 b_11 NI_11 NS_118 0 -6.1488718257204290e-02
GC_11_119 b_11 NI_11 NS_119 0 8.4504622916550420e-02
GC_11_120 b_11 NI_11 NS_120 0 -1.0099258058590413e-01
GD_11_1 b_11 NI_11 NA_1 0 -1.5538174042610196e-06
GD_11_2 b_11 NI_11 NA_2 0 -5.5599313327973641e-05
GD_11_3 b_11 NI_11 NA_3 0 3.9104219663086600e-05
GD_11_4 b_11 NI_11 NA_4 0 -1.6521754335559500e-04
GD_11_5 b_11 NI_11 NA_5 0 4.3459351420468783e-04
GD_11_6 b_11 NI_11 NA_6 0 -1.3162559052130131e-04
GD_11_7 b_11 NI_11 NA_7 0 3.8583924691778272e-03
GD_11_8 b_11 NI_11 NA_8 0 2.3527094979184168e-04
GD_11_9 b_11 NI_11 NA_9 0 3.1099351267036241e-02
GD_11_10 b_11 NI_11 NA_10 0 3.7194425217160118e-04
GD_11_11 b_11 NI_11 NA_11 0 -1.3863806892214475e-02
GD_11_12 b_11 NI_11 NA_12 0 1.9655719725458976e-02
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -9.7681611493678598e-05
GC_12_2 b_12 NI_12 NS_2 0 1.3625652411588271e-04
GC_12_3 b_12 NI_12 NS_3 0 -8.2304077755972315e-09
GC_12_4 b_12 NI_12 NS_4 0 8.1286055351795112e-09
GC_12_5 b_12 NI_12 NS_5 0 -3.8731874586279440e-11
GC_12_6 b_12 NI_12 NS_6 0 -8.7182408139556192e-10
GC_12_7 b_12 NI_12 NS_7 0 -4.6992204407757525e-05
GC_12_8 b_12 NI_12 NS_8 0 4.5214859426022167e-05
GC_12_9 b_12 NI_12 NS_9 0 8.8993848083572329e-05
GC_12_10 b_12 NI_12 NS_10 0 2.2551044614933105e-04
GC_12_11 b_12 NI_12 NS_11 0 2.9950568709309313e-04
GC_12_12 b_12 NI_12 NS_12 0 -1.6297487896081727e-04
GC_12_13 b_12 NI_12 NS_13 0 3.2148093910201142e-08
GC_12_14 b_12 NI_12 NS_14 0 -1.0198415394417565e-08
GC_12_15 b_12 NI_12 NS_15 0 3.8755172796953024e-11
GC_12_16 b_12 NI_12 NS_16 0 9.2512210389744349e-10
GC_12_17 b_12 NI_12 NS_17 0 -2.7773871197578423e-06
GC_12_18 b_12 NI_12 NS_18 0 1.7958982134132495e-05
GC_12_19 b_12 NI_12 NS_19 0 -1.1314384074756495e-04
GC_12_20 b_12 NI_12 NS_20 0 -1.0759340696470801e-04
GC_12_21 b_12 NI_12 NS_21 0 -6.8745335049225241e-05
GC_12_22 b_12 NI_12 NS_22 0 3.4274282199370796e-04
GC_12_23 b_12 NI_12 NS_23 0 -2.0454017307283064e-08
GC_12_24 b_12 NI_12 NS_24 0 1.4315479645448529e-08
GC_12_25 b_12 NI_12 NS_25 0 -1.0174599979241521e-10
GC_12_26 b_12 NI_12 NS_26 0 -9.1155877990923631e-10
GC_12_27 b_12 NI_12 NS_27 0 -5.6845318325416464e-05
GC_12_28 b_12 NI_12 NS_28 0 1.2032180497915186e-04
GC_12_29 b_12 NI_12 NS_29 0 2.2055688259251361e-05
GC_12_30 b_12 NI_12 NS_30 0 5.8497488874929653e-04
GC_12_31 b_12 NI_12 NS_31 0 -1.5101101547256504e-04
GC_12_32 b_12 NI_12 NS_32 0 -2.5226873642479234e-04
GC_12_33 b_12 NI_12 NS_33 0 -3.1559083619842678e-07
GC_12_34 b_12 NI_12 NS_34 0 4.4709851055151867e-08
GC_12_35 b_12 NI_12 NS_35 0 1.0763565109496663e-10
GC_12_36 b_12 NI_12 NS_36 0 5.1223218225402046e-11
GC_12_37 b_12 NI_12 NS_37 0 8.6980632206588211e-05
GC_12_38 b_12 NI_12 NS_38 0 1.6471800050515666e-04
GC_12_39 b_12 NI_12 NS_39 0 3.1645865418488691e-04
GC_12_40 b_12 NI_12 NS_40 0 -5.7183067031546487e-04
GC_12_41 b_12 NI_12 NS_41 0 1.7522211295129583e-04
GC_12_42 b_12 NI_12 NS_42 0 5.7756027331900108e-04
GC_12_43 b_12 NI_12 NS_43 0 3.8288848137316545e-07
GC_12_44 b_12 NI_12 NS_44 0 5.8957332192288453e-09
GC_12_45 b_12 NI_12 NS_45 0 -2.1138941227792093e-10
GC_12_46 b_12 NI_12 NS_46 0 1.1214493077146343e-09
GC_12_47 b_12 NI_12 NS_47 0 5.7477864997957143e-04
GC_12_48 b_12 NI_12 NS_48 0 7.5486065024909612e-05
GC_12_49 b_12 NI_12 NS_49 0 -1.1516616088126793e-03
GC_12_50 b_12 NI_12 NS_50 0 2.9458902867056846e-04
GC_12_51 b_12 NI_12 NS_51 0 -1.8102426904621134e-03
GC_12_52 b_12 NI_12 NS_52 0 -4.2556367560624044e-04
GC_12_53 b_12 NI_12 NS_53 0 -1.7767726003691285e-06
GC_12_54 b_12 NI_12 NS_54 0 2.3259814246150690e-07
GC_12_55 b_12 NI_12 NS_55 0 2.3519255691818629e-10
GC_12_56 b_12 NI_12 NS_56 0 -4.8199409832769711e-09
GC_12_57 b_12 NI_12 NS_57 0 3.9578927010691737e-04
GC_12_58 b_12 NI_12 NS_58 0 4.5730820886789983e-04
GC_12_59 b_12 NI_12 NS_59 0 1.7014713360919190e-03
GC_12_60 b_12 NI_12 NS_60 0 -1.8062990478043073e-03
GC_12_61 b_12 NI_12 NS_61 0 4.4312076802818063e-04
GC_12_62 b_12 NI_12 NS_62 0 1.7434320196114870e-03
GC_12_63 b_12 NI_12 NS_63 0 2.5874752096212791e-06
GC_12_64 b_12 NI_12 NS_64 0 6.8072367311414042e-08
GC_12_65 b_12 NI_12 NS_65 0 -1.1315508052930240e-10
GC_12_66 b_12 NI_12 NS_66 0 2.8408045874434463e-08
GC_12_67 b_12 NI_12 NS_67 0 3.2307394077003889e-03
GC_12_68 b_12 NI_12 NS_68 0 -2.7665463265152279e-04
GC_12_69 b_12 NI_12 NS_69 0 -5.7915279978725774e-03
GC_12_70 b_12 NI_12 NS_70 0 -1.0222266352664159e-03
GC_12_71 b_12 NI_12 NS_71 0 -2.7971151411519610e-03
GC_12_72 b_12 NI_12 NS_72 0 -5.7453843688917879e-04
GC_12_73 b_12 NI_12 NS_73 0 -2.2963943578185903e-06
GC_12_74 b_12 NI_12 NS_74 0 5.4353195222753733e-08
GC_12_75 b_12 NI_12 NS_75 0 1.0753259742356695e-10
GC_12_76 b_12 NI_12 NS_76 0 -3.1802393509729266e-08
GC_12_77 b_12 NI_12 NS_77 0 5.7239651384455455e-04
GC_12_78 b_12 NI_12 NS_78 0 -1.1832259322205898e-03
GC_12_79 b_12 NI_12 NS_79 0 2.0484150784670090e-03
GC_12_80 b_12 NI_12 NS_80 0 -7.4558009810014590e-05
GC_12_81 b_12 NI_12 NS_81 0 -1.3061125580791548e-03
GC_12_82 b_12 NI_12 NS_82 0 1.1609039661503548e-03
GC_12_83 b_12 NI_12 NS_83 0 -5.2046723080868838e-06
GC_12_84 b_12 NI_12 NS_84 0 -1.3619515854241348e-07
GC_12_85 b_12 NI_12 NS_85 0 1.8849527256255734e-09
GC_12_86 b_12 NI_12 NS_86 0 1.0944656981071299e-07
GC_12_87 b_12 NI_12 NS_87 0 2.1789648288941632e-03
GC_12_88 b_12 NI_12 NS_88 0 -5.3350899546166777e-04
GC_12_89 b_12 NI_12 NS_89 0 -2.6662046367079903e-03
GC_12_90 b_12 NI_12 NS_90 0 -1.2463188652477935e-03
GC_12_91 b_12 NI_12 NS_91 0 -7.0566514973206523e-03
GC_12_92 b_12 NI_12 NS_92 0 -4.4826525389356281e-03
GC_12_93 b_12 NI_12 NS_93 0 -1.6086015613505065e-05
GC_12_94 b_12 NI_12 NS_94 0 -2.4816704104033053e-06
GC_12_95 b_12 NI_12 NS_95 0 -2.2943978362392909e-09
GC_12_96 b_12 NI_12 NS_96 0 -3.9506621399113991e-07
GC_12_97 b_12 NI_12 NS_97 0 1.7173757127493898e-03
GC_12_98 b_12 NI_12 NS_98 0 -1.3406237240908239e-02
GC_12_99 b_12 NI_12 NS_99 0 5.8866758738304733e-03
GC_12_100 b_12 NI_12 NS_100 0 1.2986108939997553e-02
GC_12_101 b_12 NI_12 NS_101 0 -1.7980244990755068e-01
GC_12_102 b_12 NI_12 NS_102 0 5.6388736466444656e-02
GC_12_103 b_12 NI_12 NS_103 0 -2.6204708171640540e-04
GC_12_104 b_12 NI_12 NS_104 0 8.7776591566488985e-05
GC_12_105 b_12 NI_12 NS_105 0 6.1886780823697295e-08
GC_12_106 b_12 NI_12 NS_106 0 6.3073454044695431e-08
GC_12_107 b_12 NI_12 NS_107 0 -3.2559836401256544e-02
GC_12_108 b_12 NI_12 NS_108 0 -6.1491335348565879e-02
GC_12_109 b_12 NI_12 NS_109 0 8.4505078097955946e-02
GC_12_110 b_12 NI_12 NS_110 0 -1.0099134515478536e-01
GC_12_111 b_12 NI_12 NS_111 0 5.2859398508041902e-02
GC_12_112 b_12 NI_12 NS_112 0 -1.3064793307874138e-02
GC_12_113 b_12 NI_12 NS_113 0 5.9279854192276102e-05
GC_12_114 b_12 NI_12 NS_114 0 -1.3381643858258897e-05
GC_12_115 b_12 NI_12 NS_115 0 -8.5088331589078162e-09
GC_12_116 b_12 NI_12 NS_116 0 -1.3098075755340869e-06
GC_12_117 b_12 NI_12 NS_117 0 -1.9013630309753474e-03
GC_12_118 b_12 NI_12 NS_118 0 4.2717618170745328e-03
GC_12_119 b_12 NI_12 NS_119 0 -1.3200571729196761e-02
GC_12_120 b_12 NI_12 NS_120 0 2.3506110531105958e-02
GD_12_1 b_12 NI_12 NA_1 0 -5.5459114778578140e-05
GD_12_2 b_12 NI_12 NA_2 0 -1.5547960944828617e-06
GD_12_3 b_12 NI_12 NA_3 0 -1.6492366173784606e-04
GD_12_4 b_12 NI_12 NA_4 0 3.9286024601949428e-05
GD_12_5 b_12 NI_12 NA_5 0 -1.3079590950170296e-04
GD_12_6 b_12 NI_12 NA_6 0 4.3527000620696211e-04
GD_12_7 b_12 NI_12 NA_7 0 2.3842103440352533e-04
GD_12_8 b_12 NI_12 NA_8 0 3.8606665769386384e-03
GD_12_9 b_12 NI_12 NA_9 0 3.7202435221328988e-04
GD_12_10 b_12 NI_12 NA_10 0 3.1107793494345781e-02
GD_12_11 b_12 NI_12 NA_11 0 1.9658445259010188e-02
GD_12_12 b_12 NI_12 NA_12 0 -1.3863806892214475e-02
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 4.0354809530581859e+00
GS_1_1 0 NS_1 NA_1 0 9.2142803748119106e-01
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 6.3411372235753936e+00
GS_2_1 0 NS_2 NA_1 0 9.2142803748119106e-01
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 2.5859585687019660e+01
GS_3_1 0 NS_3 NA_1 0 9.2142803748119106e-01
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 5.0671215210782393e+01
GS_4_1 0 NS_4 NA_1 0 9.2142803748119106e-01
*
* Real pole n. 5
CS_5 NS_5 0 9.9999999999999998e-13
RS_5 NS_5 0 6.2932864196540877e+03
GS_5_1 0 NS_5 NA_1 0 9.2142803748119106e-01
*
* Real pole n. 6
CS_6 NS_6 0 9.9999999999999998e-13
RS_6 NS_6 0 2.5334537631431394e+02
GS_6_1 0 NS_6 NA_1 0 9.2142803748119106e-01
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 6.7467067405495911e+00
RS_8 NS_8 0 6.7467067405495911e+00
GL_7 0 NS_7 NS_8 0 3.3575009023426894e-01
GL_8 0 NS_8 NS_7 0 -3.3575009023426894e-01
GS_7_1 0 NS_7 NA_1 0 9.2142803748119106e-01
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 5.1788602987145635e+00
RS_10 NS_10 0 5.1788602987145627e+00
GL_9 0 NS_9 NS_10 0 1.3722481699036998e-01
GL_10 0 NS_10 NS_9 0 -1.3722481699036998e-01
GS_9_1 0 NS_9 NA_1 0 9.2142803748119106e-01
*
* Real pole n. 11
CS_11 NS_11 0 9.9999999999999998e-13
RS_11 NS_11 0 4.0354809530581859e+00
GS_11_2 0 NS_11 NA_2 0 9.2142803748119106e-01
*
* Real pole n. 12
CS_12 NS_12 0 9.9999999999999998e-13
RS_12 NS_12 0 6.3411372235753936e+00
GS_12_2 0 NS_12 NA_2 0 9.2142803748119106e-01
*
* Real pole n. 13
CS_13 NS_13 0 9.9999999999999998e-13
RS_13 NS_13 0 2.5859585687019660e+01
GS_13_2 0 NS_13 NA_2 0 9.2142803748119106e-01
*
* Real pole n. 14
CS_14 NS_14 0 9.9999999999999998e-13
RS_14 NS_14 0 5.0671215210782393e+01
GS_14_2 0 NS_14 NA_2 0 9.2142803748119106e-01
*
* Real pole n. 15
CS_15 NS_15 0 9.9999999999999998e-13
RS_15 NS_15 0 6.2932864196540877e+03
GS_15_2 0 NS_15 NA_2 0 9.2142803748119106e-01
*
* Real pole n. 16
CS_16 NS_16 0 9.9999999999999998e-13
RS_16 NS_16 0 2.5334537631431394e+02
GS_16_2 0 NS_16 NA_2 0 9.2142803748119106e-01
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 6.7467067405495911e+00
RS_18 NS_18 0 6.7467067405495911e+00
GL_17 0 NS_17 NS_18 0 3.3575009023426894e-01
GL_18 0 NS_18 NS_17 0 -3.3575009023426894e-01
GS_17_2 0 NS_17 NA_2 0 9.2142803748119106e-01
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 5.1788602987145635e+00
RS_20 NS_20 0 5.1788602987145627e+00
GL_19 0 NS_19 NS_20 0 1.3722481699036998e-01
GL_20 0 NS_20 NS_19 0 -1.3722481699036998e-01
GS_19_2 0 NS_19 NA_2 0 9.2142803748119106e-01
*
* Real pole n. 21
CS_21 NS_21 0 9.9999999999999998e-13
RS_21 NS_21 0 4.0354809530581859e+00
GS_21_3 0 NS_21 NA_3 0 9.2142803748119106e-01
*
* Real pole n. 22
CS_22 NS_22 0 9.9999999999999998e-13
RS_22 NS_22 0 6.3411372235753936e+00
GS_22_3 0 NS_22 NA_3 0 9.2142803748119106e-01
*
* Real pole n. 23
CS_23 NS_23 0 9.9999999999999998e-13
RS_23 NS_23 0 2.5859585687019660e+01
GS_23_3 0 NS_23 NA_3 0 9.2142803748119106e-01
*
* Real pole n. 24
CS_24 NS_24 0 9.9999999999999998e-13
RS_24 NS_24 0 5.0671215210782393e+01
GS_24_3 0 NS_24 NA_3 0 9.2142803748119106e-01
*
* Real pole n. 25
CS_25 NS_25 0 9.9999999999999998e-13
RS_25 NS_25 0 6.2932864196540877e+03
GS_25_3 0 NS_25 NA_3 0 9.2142803748119106e-01
*
* Real pole n. 26
CS_26 NS_26 0 9.9999999999999998e-13
RS_26 NS_26 0 2.5334537631431394e+02
GS_26_3 0 NS_26 NA_3 0 9.2142803748119106e-01
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 6.7467067405495911e+00
RS_28 NS_28 0 6.7467067405495911e+00
GL_27 0 NS_27 NS_28 0 3.3575009023426894e-01
GL_28 0 NS_28 NS_27 0 -3.3575009023426894e-01
GS_27_3 0 NS_27 NA_3 0 9.2142803748119106e-01
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 5.1788602987145635e+00
RS_30 NS_30 0 5.1788602987145627e+00
GL_29 0 NS_29 NS_30 0 1.3722481699036998e-01
GL_30 0 NS_30 NS_29 0 -1.3722481699036998e-01
GS_29_3 0 NS_29 NA_3 0 9.2142803748119106e-01
*
* Real pole n. 31
CS_31 NS_31 0 9.9999999999999998e-13
RS_31 NS_31 0 4.0354809530581859e+00
GS_31_4 0 NS_31 NA_4 0 9.2142803748119106e-01
*
* Real pole n. 32
CS_32 NS_32 0 9.9999999999999998e-13
RS_32 NS_32 0 6.3411372235753936e+00
GS_32_4 0 NS_32 NA_4 0 9.2142803748119106e-01
*
* Real pole n. 33
CS_33 NS_33 0 9.9999999999999998e-13
RS_33 NS_33 0 2.5859585687019660e+01
GS_33_4 0 NS_33 NA_4 0 9.2142803748119106e-01
*
* Real pole n. 34
CS_34 NS_34 0 9.9999999999999998e-13
RS_34 NS_34 0 5.0671215210782393e+01
GS_34_4 0 NS_34 NA_4 0 9.2142803748119106e-01
*
* Real pole n. 35
CS_35 NS_35 0 9.9999999999999998e-13
RS_35 NS_35 0 6.2932864196540877e+03
GS_35_4 0 NS_35 NA_4 0 9.2142803748119106e-01
*
* Real pole n. 36
CS_36 NS_36 0 9.9999999999999998e-13
RS_36 NS_36 0 2.5334537631431394e+02
GS_36_4 0 NS_36 NA_4 0 9.2142803748119106e-01
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 6.7467067405495911e+00
RS_38 NS_38 0 6.7467067405495911e+00
GL_37 0 NS_37 NS_38 0 3.3575009023426894e-01
GL_38 0 NS_38 NS_37 0 -3.3575009023426894e-01
GS_37_4 0 NS_37 NA_4 0 9.2142803748119106e-01
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 5.1788602987145635e+00
RS_40 NS_40 0 5.1788602987145627e+00
GL_39 0 NS_39 NS_40 0 1.3722481699036998e-01
GL_40 0 NS_40 NS_39 0 -1.3722481699036998e-01
GS_39_4 0 NS_39 NA_4 0 9.2142803748119106e-01
*
* Real pole n. 41
CS_41 NS_41 0 9.9999999999999998e-13
RS_41 NS_41 0 4.0354809530581859e+00
GS_41_5 0 NS_41 NA_5 0 9.2142803748119106e-01
*
* Real pole n. 42
CS_42 NS_42 0 9.9999999999999998e-13
RS_42 NS_42 0 6.3411372235753936e+00
GS_42_5 0 NS_42 NA_5 0 9.2142803748119106e-01
*
* Real pole n. 43
CS_43 NS_43 0 9.9999999999999998e-13
RS_43 NS_43 0 2.5859585687019660e+01
GS_43_5 0 NS_43 NA_5 0 9.2142803748119106e-01
*
* Real pole n. 44
CS_44 NS_44 0 9.9999999999999998e-13
RS_44 NS_44 0 5.0671215210782393e+01
GS_44_5 0 NS_44 NA_5 0 9.2142803748119106e-01
*
* Real pole n. 45
CS_45 NS_45 0 9.9999999999999998e-13
RS_45 NS_45 0 6.2932864196540877e+03
GS_45_5 0 NS_45 NA_5 0 9.2142803748119106e-01
*
* Real pole n. 46
CS_46 NS_46 0 9.9999999999999998e-13
RS_46 NS_46 0 2.5334537631431394e+02
GS_46_5 0 NS_46 NA_5 0 9.2142803748119106e-01
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 6.7467067405495911e+00
RS_48 NS_48 0 6.7467067405495911e+00
GL_47 0 NS_47 NS_48 0 3.3575009023426894e-01
GL_48 0 NS_48 NS_47 0 -3.3575009023426894e-01
GS_47_5 0 NS_47 NA_5 0 9.2142803748119106e-01
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 5.1788602987145635e+00
RS_50 NS_50 0 5.1788602987145627e+00
GL_49 0 NS_49 NS_50 0 1.3722481699036998e-01
GL_50 0 NS_50 NS_49 0 -1.3722481699036998e-01
GS_49_5 0 NS_49 NA_5 0 9.2142803748119106e-01
*
* Real pole n. 51
CS_51 NS_51 0 9.9999999999999998e-13
RS_51 NS_51 0 4.0354809530581859e+00
GS_51_6 0 NS_51 NA_6 0 9.2142803748119106e-01
*
* Real pole n. 52
CS_52 NS_52 0 9.9999999999999998e-13
RS_52 NS_52 0 6.3411372235753936e+00
GS_52_6 0 NS_52 NA_6 0 9.2142803748119106e-01
*
* Real pole n. 53
CS_53 NS_53 0 9.9999999999999998e-13
RS_53 NS_53 0 2.5859585687019660e+01
GS_53_6 0 NS_53 NA_6 0 9.2142803748119106e-01
*
* Real pole n. 54
CS_54 NS_54 0 9.9999999999999998e-13
RS_54 NS_54 0 5.0671215210782393e+01
GS_54_6 0 NS_54 NA_6 0 9.2142803748119106e-01
*
* Real pole n. 55
CS_55 NS_55 0 9.9999999999999998e-13
RS_55 NS_55 0 6.2932864196540877e+03
GS_55_6 0 NS_55 NA_6 0 9.2142803748119106e-01
*
* Real pole n. 56
CS_56 NS_56 0 9.9999999999999998e-13
RS_56 NS_56 0 2.5334537631431394e+02
GS_56_6 0 NS_56 NA_6 0 9.2142803748119106e-01
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 6.7467067405495911e+00
RS_58 NS_58 0 6.7467067405495911e+00
GL_57 0 NS_57 NS_58 0 3.3575009023426894e-01
GL_58 0 NS_58 NS_57 0 -3.3575009023426894e-01
GS_57_6 0 NS_57 NA_6 0 9.2142803748119106e-01
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 5.1788602987145635e+00
RS_60 NS_60 0 5.1788602987145627e+00
GL_59 0 NS_59 NS_60 0 1.3722481699036998e-01
GL_60 0 NS_60 NS_59 0 -1.3722481699036998e-01
GS_59_6 0 NS_59 NA_6 0 9.2142803748119106e-01
*
* Real pole n. 61
CS_61 NS_61 0 9.9999999999999998e-13
RS_61 NS_61 0 4.0354809530581859e+00
GS_61_7 0 NS_61 NA_7 0 9.2142803748119106e-01
*
* Real pole n. 62
CS_62 NS_62 0 9.9999999999999998e-13
RS_62 NS_62 0 6.3411372235753936e+00
GS_62_7 0 NS_62 NA_7 0 9.2142803748119106e-01
*
* Real pole n. 63
CS_63 NS_63 0 9.9999999999999998e-13
RS_63 NS_63 0 2.5859585687019660e+01
GS_63_7 0 NS_63 NA_7 0 9.2142803748119106e-01
*
* Real pole n. 64
CS_64 NS_64 0 9.9999999999999998e-13
RS_64 NS_64 0 5.0671215210782393e+01
GS_64_7 0 NS_64 NA_7 0 9.2142803748119106e-01
*
* Real pole n. 65
CS_65 NS_65 0 9.9999999999999998e-13
RS_65 NS_65 0 6.2932864196540877e+03
GS_65_7 0 NS_65 NA_7 0 9.2142803748119106e-01
*
* Real pole n. 66
CS_66 NS_66 0 9.9999999999999998e-13
RS_66 NS_66 0 2.5334537631431394e+02
GS_66_7 0 NS_66 NA_7 0 9.2142803748119106e-01
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 6.7467067405495911e+00
RS_68 NS_68 0 6.7467067405495911e+00
GL_67 0 NS_67 NS_68 0 3.3575009023426894e-01
GL_68 0 NS_68 NS_67 0 -3.3575009023426894e-01
GS_67_7 0 NS_67 NA_7 0 9.2142803748119106e-01
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 5.1788602987145635e+00
RS_70 NS_70 0 5.1788602987145627e+00
GL_69 0 NS_69 NS_70 0 1.3722481699036998e-01
GL_70 0 NS_70 NS_69 0 -1.3722481699036998e-01
GS_69_7 0 NS_69 NA_7 0 9.2142803748119106e-01
*
* Real pole n. 71
CS_71 NS_71 0 9.9999999999999998e-13
RS_71 NS_71 0 4.0354809530581859e+00
GS_71_8 0 NS_71 NA_8 0 9.2142803748119106e-01
*
* Real pole n. 72
CS_72 NS_72 0 9.9999999999999998e-13
RS_72 NS_72 0 6.3411372235753936e+00
GS_72_8 0 NS_72 NA_8 0 9.2142803748119106e-01
*
* Real pole n. 73
CS_73 NS_73 0 9.9999999999999998e-13
RS_73 NS_73 0 2.5859585687019660e+01
GS_73_8 0 NS_73 NA_8 0 9.2142803748119106e-01
*
* Real pole n. 74
CS_74 NS_74 0 9.9999999999999998e-13
RS_74 NS_74 0 5.0671215210782393e+01
GS_74_8 0 NS_74 NA_8 0 9.2142803748119106e-01
*
* Real pole n. 75
CS_75 NS_75 0 9.9999999999999998e-13
RS_75 NS_75 0 6.2932864196540877e+03
GS_75_8 0 NS_75 NA_8 0 9.2142803748119106e-01
*
* Real pole n. 76
CS_76 NS_76 0 9.9999999999999998e-13
RS_76 NS_76 0 2.5334537631431394e+02
GS_76_8 0 NS_76 NA_8 0 9.2142803748119106e-01
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 6.7467067405495911e+00
RS_78 NS_78 0 6.7467067405495911e+00
GL_77 0 NS_77 NS_78 0 3.3575009023426894e-01
GL_78 0 NS_78 NS_77 0 -3.3575009023426894e-01
GS_77_8 0 NS_77 NA_8 0 9.2142803748119106e-01
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 5.1788602987145635e+00
RS_80 NS_80 0 5.1788602987145627e+00
GL_79 0 NS_79 NS_80 0 1.3722481699036998e-01
GL_80 0 NS_80 NS_79 0 -1.3722481699036998e-01
GS_79_8 0 NS_79 NA_8 0 9.2142803748119106e-01
*
* Real pole n. 81
CS_81 NS_81 0 9.9999999999999998e-13
RS_81 NS_81 0 4.0354809530581859e+00
GS_81_9 0 NS_81 NA_9 0 9.2142803748119106e-01
*
* Real pole n. 82
CS_82 NS_82 0 9.9999999999999998e-13
RS_82 NS_82 0 6.3411372235753936e+00
GS_82_9 0 NS_82 NA_9 0 9.2142803748119106e-01
*
* Real pole n. 83
CS_83 NS_83 0 9.9999999999999998e-13
RS_83 NS_83 0 2.5859585687019660e+01
GS_83_9 0 NS_83 NA_9 0 9.2142803748119106e-01
*
* Real pole n. 84
CS_84 NS_84 0 9.9999999999999998e-13
RS_84 NS_84 0 5.0671215210782393e+01
GS_84_9 0 NS_84 NA_9 0 9.2142803748119106e-01
*
* Real pole n. 85
CS_85 NS_85 0 9.9999999999999998e-13
RS_85 NS_85 0 6.2932864196540877e+03
GS_85_9 0 NS_85 NA_9 0 9.2142803748119106e-01
*
* Real pole n. 86
CS_86 NS_86 0 9.9999999999999998e-13
RS_86 NS_86 0 2.5334537631431394e+02
GS_86_9 0 NS_86 NA_9 0 9.2142803748119106e-01
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 6.7467067405495911e+00
RS_88 NS_88 0 6.7467067405495911e+00
GL_87 0 NS_87 NS_88 0 3.3575009023426894e-01
GL_88 0 NS_88 NS_87 0 -3.3575009023426894e-01
GS_87_9 0 NS_87 NA_9 0 9.2142803748119106e-01
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 5.1788602987145635e+00
RS_90 NS_90 0 5.1788602987145627e+00
GL_89 0 NS_89 NS_90 0 1.3722481699036998e-01
GL_90 0 NS_90 NS_89 0 -1.3722481699036998e-01
GS_89_9 0 NS_89 NA_9 0 9.2142803748119106e-01
*
* Real pole n. 91
CS_91 NS_91 0 9.9999999999999998e-13
RS_91 NS_91 0 4.0354809530581859e+00
GS_91_10 0 NS_91 NA_10 0 9.2142803748119106e-01
*
* Real pole n. 92
CS_92 NS_92 0 9.9999999999999998e-13
RS_92 NS_92 0 6.3411372235753936e+00
GS_92_10 0 NS_92 NA_10 0 9.2142803748119106e-01
*
* Real pole n. 93
CS_93 NS_93 0 9.9999999999999998e-13
RS_93 NS_93 0 2.5859585687019660e+01
GS_93_10 0 NS_93 NA_10 0 9.2142803748119106e-01
*
* Real pole n. 94
CS_94 NS_94 0 9.9999999999999998e-13
RS_94 NS_94 0 5.0671215210782393e+01
GS_94_10 0 NS_94 NA_10 0 9.2142803748119106e-01
*
* Real pole n. 95
CS_95 NS_95 0 9.9999999999999998e-13
RS_95 NS_95 0 6.2932864196540877e+03
GS_95_10 0 NS_95 NA_10 0 9.2142803748119106e-01
*
* Real pole n. 96
CS_96 NS_96 0 9.9999999999999998e-13
RS_96 NS_96 0 2.5334537631431394e+02
GS_96_10 0 NS_96 NA_10 0 9.2142803748119106e-01
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 6.7467067405495911e+00
RS_98 NS_98 0 6.7467067405495911e+00
GL_97 0 NS_97 NS_98 0 3.3575009023426894e-01
GL_98 0 NS_98 NS_97 0 -3.3575009023426894e-01
GS_97_10 0 NS_97 NA_10 0 9.2142803748119106e-01
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 5.1788602987145635e+00
RS_100 NS_100 0 5.1788602987145627e+00
GL_99 0 NS_99 NS_100 0 1.3722481699036998e-01
GL_100 0 NS_100 NS_99 0 -1.3722481699036998e-01
GS_99_10 0 NS_99 NA_10 0 9.2142803748119106e-01
*
* Real pole n. 101
CS_101 NS_101 0 9.9999999999999998e-13
RS_101 NS_101 0 4.0354809530581859e+00
GS_101_11 0 NS_101 NA_11 0 9.2142803748119106e-01
*
* Real pole n. 102
CS_102 NS_102 0 9.9999999999999998e-13
RS_102 NS_102 0 6.3411372235753936e+00
GS_102_11 0 NS_102 NA_11 0 9.2142803748119106e-01
*
* Real pole n. 103
CS_103 NS_103 0 9.9999999999999998e-13
RS_103 NS_103 0 2.5859585687019660e+01
GS_103_11 0 NS_103 NA_11 0 9.2142803748119106e-01
*
* Real pole n. 104
CS_104 NS_104 0 9.9999999999999998e-13
RS_104 NS_104 0 5.0671215210782393e+01
GS_104_11 0 NS_104 NA_11 0 9.2142803748119106e-01
*
* Real pole n. 105
CS_105 NS_105 0 9.9999999999999998e-13
RS_105 NS_105 0 6.2932864196540877e+03
GS_105_11 0 NS_105 NA_11 0 9.2142803748119106e-01
*
* Real pole n. 106
CS_106 NS_106 0 9.9999999999999998e-13
RS_106 NS_106 0 2.5334537631431394e+02
GS_106_11 0 NS_106 NA_11 0 9.2142803748119106e-01
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 6.7467067405495911e+00
RS_108 NS_108 0 6.7467067405495911e+00
GL_107 0 NS_107 NS_108 0 3.3575009023426894e-01
GL_108 0 NS_108 NS_107 0 -3.3575009023426894e-01
GS_107_11 0 NS_107 NA_11 0 9.2142803748119106e-01
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 5.1788602987145635e+00
RS_110 NS_110 0 5.1788602987145627e+00
GL_109 0 NS_109 NS_110 0 1.3722481699036998e-01
GL_110 0 NS_110 NS_109 0 -1.3722481699036998e-01
GS_109_11 0 NS_109 NA_11 0 9.2142803748119106e-01
*
* Real pole n. 111
CS_111 NS_111 0 9.9999999999999998e-13
RS_111 NS_111 0 4.0354809530581859e+00
GS_111_12 0 NS_111 NA_12 0 9.2142803748119106e-01
*
* Real pole n. 112
CS_112 NS_112 0 9.9999999999999998e-13
RS_112 NS_112 0 6.3411372235753936e+00
GS_112_12 0 NS_112 NA_12 0 9.2142803748119106e-01
*
* Real pole n. 113
CS_113 NS_113 0 9.9999999999999998e-13
RS_113 NS_113 0 2.5859585687019660e+01
GS_113_12 0 NS_113 NA_12 0 9.2142803748119106e-01
*
* Real pole n. 114
CS_114 NS_114 0 9.9999999999999998e-13
RS_114 NS_114 0 5.0671215210782393e+01
GS_114_12 0 NS_114 NA_12 0 9.2142803748119106e-01
*
* Real pole n. 115
CS_115 NS_115 0 9.9999999999999998e-13
RS_115 NS_115 0 6.2932864196540877e+03
GS_115_12 0 NS_115 NA_12 0 9.2142803748119106e-01
*
* Real pole n. 116
CS_116 NS_116 0 9.9999999999999998e-13
RS_116 NS_116 0 2.5334537631431394e+02
GS_116_12 0 NS_116 NA_12 0 9.2142803748119106e-01
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 6.7467067405495911e+00
RS_118 NS_118 0 6.7467067405495911e+00
GL_117 0 NS_117 NS_118 0 3.3575009023426894e-01
GL_118 0 NS_118 NS_117 0 -3.3575009023426894e-01
GS_117_12 0 NS_117 NA_12 0 9.2142803748119106e-01
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 5.1788602987145635e+00
RS_120 NS_120 0 5.1788602987145627e+00
GL_119 0 NS_119 NS_120 0 1.3722481699036998e-01
GL_120 0 NS_120 NS_119 0 -1.3722481699036998e-01
GS_119_12 0 NS_119 NA_12 0 9.2142803748119106e-01
*
******************************


.ends
*******************
* End of subcircuit
*******************
