**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [6 2 22] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** n/a - passivity was not enforced
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_13_PCB_wire_0p25inch_lowloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 -1.5427134833671494e-05
GC_1_2 b_1 NI_1 NS_2 0 -3.7324314463545671e-06
GC_1_3 b_1 NI_1 NS_3 0 -2.3081208574539930e-08
GC_1_4 b_1 NI_1 NS_4 0 -3.8674152015124863e-07
GC_1_5 b_1 NI_1 NS_5 0 4.5760065321819544e-03
GC_1_6 b_1 NI_1 NS_6 0 3.7993286796473413e-03
GC_1_7 b_1 NI_1 NS_7 0 1.3872401175672972e-02
GC_1_8 b_1 NI_1 NS_8 0 -2.1406272364670791e-02
GC_1_9 b_1 NI_1 NS_9 0 -2.2493840945157238e-02
GC_1_10 b_1 NI_1 NS_10 0 2.6058892826137971e-02
GC_1_11 b_1 NI_1 NS_11 0 3.8337056193939845e-02
GC_1_12 b_1 NI_1 NS_12 0 -3.0181707170744618e-02
GC_1_13 b_1 NI_1 NS_13 0 -4.8685823011493726e-02
GC_1_14 b_1 NI_1 NS_14 0 1.9831379205208496e-02
GC_1_15 b_1 NI_1 NS_15 0 2.6967890308017876e-02
GC_1_16 b_1 NI_1 NS_16 0 -1.5945601193033111e-02
GC_1_17 b_1 NI_1 NS_17 0 -1.4394992250511156e-02
GC_1_18 b_1 NI_1 NS_18 0 6.8900418217842071e-03
GC_1_19 b_1 NI_1 NS_19 0 -4.8273798048062144e-03
GC_1_20 b_1 NI_1 NS_20 0 -1.6678597174271628e-02
GC_1_21 b_1 NI_1 NS_21 0 8.9998734551854876e-05
GC_1_22 b_1 NI_1 NS_22 0 3.6211869169675083e-06
GC_1_23 b_1 NI_1 NS_23 0 5.9682354758434722e-09
GC_1_24 b_1 NI_1 NS_24 0 5.9667522902359863e-07
GC_1_25 b_1 NI_1 NS_25 0 4.7508861022456356e-02
GC_1_26 b_1 NI_1 NS_26 0 -9.6471124299470808e-03
GC_1_27 b_1 NI_1 NS_27 0 -4.5582916284812439e-02
GC_1_28 b_1 NI_1 NS_28 0 2.0552301948532230e-02
GC_1_29 b_1 NI_1 NS_29 0 -5.7696873069333687e-02
GC_1_30 b_1 NI_1 NS_30 0 -6.7350307522222236e-02
GC_1_31 b_1 NI_1 NS_31 0 6.3862086522426101e-02
GC_1_32 b_1 NI_1 NS_32 0 -2.2063737480482501e-02
GC_1_33 b_1 NI_1 NS_33 0 2.8382271166397396e-02
GC_1_34 b_1 NI_1 NS_34 0 8.9387912540108805e-02
GC_1_35 b_1 NI_1 NS_35 0 -5.4366407764440933e-02
GC_1_36 b_1 NI_1 NS_36 0 2.7979863436566029e-03
GC_1_37 b_1 NI_1 NS_37 0 -1.3847775043581515e-02
GC_1_38 b_1 NI_1 NS_38 0 -4.7095073864144334e-02
GC_1_39 b_1 NI_1 NS_39 0 1.6380424383275735e-02
GC_1_40 b_1 NI_1 NS_40 0 -3.9016261579912184e-02
GC_1_41 b_1 NI_1 NS_41 0 -1.0356264848364811e-05
GC_1_42 b_1 NI_1 NS_42 0 -2.1272069476427938e-07
GC_1_43 b_1 NI_1 NS_43 0 -1.2831320148494259e-09
GC_1_44 b_1 NI_1 NS_44 0 -2.5390347645538870e-08
GC_1_45 b_1 NI_1 NS_45 0 -4.2497281814668159e-03
GC_1_46 b_1 NI_1 NS_46 0 -3.4927766090990550e-03
GC_1_47 b_1 NI_1 NS_47 0 -1.2922365127891406e-02
GC_1_48 b_1 NI_1 NS_48 0 1.7065796230691491e-02
GC_1_49 b_1 NI_1 NS_49 0 1.7371354225988563e-02
GC_1_50 b_1 NI_1 NS_50 0 -1.9447062637168996e-02
GC_1_51 b_1 NI_1 NS_51 0 -3.3168706678817890e-02
GC_1_52 b_1 NI_1 NS_52 0 2.5454421766033537e-02
GC_1_53 b_1 NI_1 NS_53 0 4.0789606058407438e-02
GC_1_54 b_1 NI_1 NS_54 0 -1.1433470437631330e-02
GC_1_55 b_1 NI_1 NS_55 0 -2.1059355346524658e-02
GC_1_56 b_1 NI_1 NS_56 0 1.5315260733975060e-02
GC_1_57 b_1 NI_1 NS_57 0 1.4123842664329858e-02
GC_1_58 b_1 NI_1 NS_58 0 -3.7538561739732805e-03
GC_1_59 b_1 NI_1 NS_59 0 7.0868353733450707e-03
GC_1_60 b_1 NI_1 NS_60 0 1.3573780074925436e-02
GC_1_61 b_1 NI_1 NS_61 0 -1.8490439615139437e-06
GC_1_62 b_1 NI_1 NS_62 0 2.5677074933392194e-07
GC_1_63 b_1 NI_1 NS_63 0 1.6912981785828298e-09
GC_1_64 b_1 NI_1 NS_64 0 1.3611966266223569e-08
GC_1_65 b_1 NI_1 NS_65 0 1.1406458022347574e-03
GC_1_66 b_1 NI_1 NS_66 0 -2.1726047860165824e-03
GC_1_67 b_1 NI_1 NS_67 0 3.4952390932754688e-03
GC_1_68 b_1 NI_1 NS_68 0 -1.3003077579089521e-02
GC_1_69 b_1 NI_1 NS_69 0 -3.9401362279387793e-02
GC_1_70 b_1 NI_1 NS_70 0 -3.6438011076934138e-04
GC_1_71 b_1 NI_1 NS_71 0 -2.6247364897834035e-02
GC_1_72 b_1 NI_1 NS_72 0 2.8990158213005355e-02
GC_1_73 b_1 NI_1 NS_73 0 5.2202631372588425e-02
GC_1_74 b_1 NI_1 NS_74 0 3.8208679971992614e-02
GC_1_75 b_1 NI_1 NS_75 0 1.7572267408916771e-02
GC_1_76 b_1 NI_1 NS_76 0 -1.4394059888813116e-02
GC_1_77 b_1 NI_1 NS_77 0 -9.1651297154559906e-03
GC_1_78 b_1 NI_1 NS_78 0 -3.7458099504316571e-03
GC_1_79 b_1 NI_1 NS_79 0 8.0623393298334071e-03
GC_1_80 b_1 NI_1 NS_80 0 5.8595893515523386e-03
GC_1_81 b_1 NI_1 NS_81 0 -2.8092440288425173e-08
GC_1_82 b_1 NI_1 NS_82 0 1.2625337474215857e-09
GC_1_83 b_1 NI_1 NS_83 0 -9.9117586587806565e-12
GC_1_84 b_1 NI_1 NS_84 0 2.2550558458697022e-11
GC_1_85 b_1 NI_1 NS_85 0 4.4972689419318870e-06
GC_1_86 b_1 NI_1 NS_86 0 2.2387586722816038e-06
GC_1_87 b_1 NI_1 NS_87 0 9.9893573540610767e-06
GC_1_88 b_1 NI_1 NS_88 0 9.6249760329734133e-06
GC_1_89 b_1 NI_1 NS_89 0 1.8703103400856396e-05
GC_1_90 b_1 NI_1 NS_90 0 -2.3516915801382316e-05
GC_1_91 b_1 NI_1 NS_91 0 1.1345871735913158e-05
GC_1_92 b_1 NI_1 NS_92 0 -3.3422993560431516e-06
GC_1_93 b_1 NI_1 NS_93 0 -6.9544968254494872e-06
GC_1_94 b_1 NI_1 NS_94 0 -5.3248456054245464e-05
GC_1_95 b_1 NI_1 NS_95 0 -1.4962316211438840e-05
GC_1_96 b_1 NI_1 NS_96 0 -1.7861800586854711e-05
GC_1_97 b_1 NI_1 NS_97 0 -2.7583405432856385e-05
GC_1_98 b_1 NI_1 NS_98 0 -1.2422759826088116e-05
GC_1_99 b_1 NI_1 NS_99 0 -1.9191335618816399e-05
GC_1_100 b_1 NI_1 NS_100 0 5.8309121447318445e-06
GC_1_101 b_1 NI_1 NS_101 0 1.9598946470227410e-09
GC_1_102 b_1 NI_1 NS_102 0 -2.0086874360900031e-10
GC_1_103 b_1 NI_1 NS_103 0 1.6947995157649516e-11
GC_1_104 b_1 NI_1 NS_104 0 -8.9403567446646518e-11
GC_1_105 b_1 NI_1 NS_105 0 -1.5359112189243393e-06
GC_1_106 b_1 NI_1 NS_106 0 -1.4180235571302273e-06
GC_1_107 b_1 NI_1 NS_107 0 -5.6310779670129126e-06
GC_1_108 b_1 NI_1 NS_108 0 1.3500611750431549e-05
GC_1_109 b_1 NI_1 NS_109 0 3.5171791665529070e-05
GC_1_110 b_1 NI_1 NS_110 0 1.0738187807399045e-05
GC_1_111 b_1 NI_1 NS_111 0 3.2592497147550180e-05
GC_1_112 b_1 NI_1 NS_112 0 -2.6153534908048104e-05
GC_1_113 b_1 NI_1 NS_113 0 -4.0881138315577420e-05
GC_1_114 b_1 NI_1 NS_114 0 -5.0758189819292667e-05
GC_1_115 b_1 NI_1 NS_115 0 -2.0190319845236130e-05
GC_1_116 b_1 NI_1 NS_116 0 9.6138439711589819e-06
GC_1_117 b_1 NI_1 NS_117 0 3.9348241833565739e-06
GC_1_118 b_1 NI_1 NS_118 0 1.2590336294826159e-07
GC_1_119 b_1 NI_1 NS_119 0 -1.3016787727210123e-05
GC_1_120 b_1 NI_1 NS_120 0 -6.9640822669126007e-06
GC_1_121 b_1 NI_1 NS_121 0 2.0299546140481705e-08
GC_1_122 b_1 NI_1 NS_122 0 -1.0034002686525121e-09
GC_1_123 b_1 NI_1 NS_123 0 -1.9109342675463624e-11
GC_1_124 b_1 NI_1 NS_124 0 1.5480761836615813e-10
GC_1_125 b_1 NI_1 NS_125 0 -1.0725434622452993e-06
GC_1_126 b_1 NI_1 NS_126 0 -8.5344075162897932e-07
GC_1_127 b_1 NI_1 NS_127 0 -1.9513310892946869e-06
GC_1_128 b_1 NI_1 NS_128 0 -1.3188138025883565e-08
GC_1_129 b_1 NI_1 NS_129 0 -3.0922827393656368e-06
GC_1_130 b_1 NI_1 NS_130 0 7.4413712648172044e-07
GC_1_131 b_1 NI_1 NS_131 0 -4.1341886827109643e-06
GC_1_132 b_1 NI_1 NS_132 0 4.2201126647395223e-06
GC_1_133 b_1 NI_1 NS_133 0 3.1590338887411926e-06
GC_1_134 b_1 NI_1 NS_134 0 5.3423798158732478e-06
GC_1_135 b_1 NI_1 NS_135 0 -9.0664820051612160e-07
GC_1_136 b_1 NI_1 NS_136 0 5.9322125548371897e-06
GC_1_137 b_1 NI_1 NS_137 0 5.9750664309987333e-06
GC_1_138 b_1 NI_1 NS_138 0 3.2312446526880142e-06
GC_1_139 b_1 NI_1 NS_139 0 5.7326862601811489e-06
GC_1_140 b_1 NI_1 NS_140 0 1.6824495324711960e-06
GC_1_141 b_1 NI_1 NS_141 0 -2.3936347645166899e-08
GC_1_142 b_1 NI_1 NS_142 0 1.2234640188227060e-09
GC_1_143 b_1 NI_1 NS_143 0 2.1495916698099719e-11
GC_1_144 b_1 NI_1 NS_144 0 -1.7598162135548903e-10
GC_1_145 b_1 NI_1 NS_145 0 1.8751005647204246e-06
GC_1_146 b_1 NI_1 NS_146 0 -4.2198207591646423e-06
GC_1_147 b_1 NI_1 NS_147 0 2.4962608508731053e-06
GC_1_148 b_1 NI_1 NS_148 0 3.3570575042169042e-08
GC_1_149 b_1 NI_1 NS_149 0 -1.6539764370095475e-06
GC_1_150 b_1 NI_1 NS_150 0 -4.5468556956447017e-06
GC_1_151 b_1 NI_1 NS_151 0 9.6538947329780083e-07
GC_1_152 b_1 NI_1 NS_152 0 -7.3307017335965299e-06
GC_1_153 b_1 NI_1 NS_153 0 -8.9355030981749736e-06
GC_1_154 b_1 NI_1 NS_154 0 -4.6687538325722228e-06
GC_1_155 b_1 NI_1 NS_155 0 -3.3134578113383491e-06
GC_1_156 b_1 NI_1 NS_156 0 1.4348150263421389e-06
GC_1_157 b_1 NI_1 NS_157 0 -1.9277165976358564e-06
GC_1_158 b_1 NI_1 NS_158 0 -4.7310371470009925e-07
GC_1_159 b_1 NI_1 NS_159 0 -3.2465968730777669e-06
GC_1_160 b_1 NI_1 NS_160 0 -1.4929324878008046e-06
GC_1_161 b_1 NI_1 NS_161 0 1.2106842237884703e-08
GC_1_162 b_1 NI_1 NS_162 0 -8.1571298811555564e-10
GC_1_163 b_1 NI_1 NS_163 0 -1.6071023418781674e-11
GC_1_164 b_1 NI_1 NS_164 0 1.3071903269525911e-10
GC_1_165 b_1 NI_1 NS_165 0 7.0579052575455553e-08
GC_1_166 b_1 NI_1 NS_166 0 -1.7341292851143489e-08
GC_1_167 b_1 NI_1 NS_167 0 -5.8731127869909124e-07
GC_1_168 b_1 NI_1 NS_168 0 5.5956805176833051e-07
GC_1_169 b_1 NI_1 NS_169 0 1.6811068744447512e-06
GC_1_170 b_1 NI_1 NS_170 0 -5.0795584588021045e-07
GC_1_171 b_1 NI_1 NS_171 0 -9.8095867614861980e-07
GC_1_172 b_1 NI_1 NS_172 0 1.0424098484702523e-07
GC_1_173 b_1 NI_1 NS_173 0 1.6471580138523334e-06
GC_1_174 b_1 NI_1 NS_174 0 -1.1441251756289331e-06
GC_1_175 b_1 NI_1 NS_175 0 -9.0813493777810186e-07
GC_1_176 b_1 NI_1 NS_176 0 -8.6585062111804777e-07
GC_1_177 b_1 NI_1 NS_177 0 -1.1417346081240492e-06
GC_1_178 b_1 NI_1 NS_178 0 -2.4697843848620396e-07
GC_1_179 b_1 NI_1 NS_179 0 8.7317971471414561e-08
GC_1_180 b_1 NI_1 NS_180 0 1.1733539946370222e-06
GC_1_181 b_1 NI_1 NS_181 0 -8.0862450612965640e-09
GC_1_182 b_1 NI_1 NS_182 0 6.7986866325640429e-10
GC_1_183 b_1 NI_1 NS_183 0 1.5646924258080400e-11
GC_1_184 b_1 NI_1 NS_184 0 -1.2067900853629605e-10
GC_1_185 b_1 NI_1 NS_185 0 -2.1903688072239168e-06
GC_1_186 b_1 NI_1 NS_186 0 2.1886429252156328e-07
GC_1_187 b_1 NI_1 NS_187 0 -2.1895702693708999e-06
GC_1_188 b_1 NI_1 NS_188 0 2.7884235005604448e-06
GC_1_189 b_1 NI_1 NS_189 0 -1.1327115041868474e-06
GC_1_190 b_1 NI_1 NS_190 0 6.5773615222719144e-06
GC_1_191 b_1 NI_1 NS_191 0 -4.1803954700632813e-07
GC_1_192 b_1 NI_1 NS_192 0 2.1422267847399631e-06
GC_1_193 b_1 NI_1 NS_193 0 7.2190705524395957e-06
GC_1_194 b_1 NI_1 NS_194 0 5.1224416474795141e-06
GC_1_195 b_1 NI_1 NS_195 0 1.6120534398522007e-06
GC_1_196 b_1 NI_1 NS_196 0 3.1394760665465149e-06
GC_1_197 b_1 NI_1 NS_197 0 4.8357385644198927e-06
GC_1_198 b_1 NI_1 NS_198 0 1.1501568808445245e-06
GC_1_199 b_1 NI_1 NS_199 0 2.9137147537947708e-06
GC_1_200 b_1 NI_1 NS_200 0 -1.3217648486956743e-06
GC_1_201 b_1 NI_1 NS_201 0 2.2396157452627350e-09
GC_1_202 b_1 NI_1 NS_202 0 -6.1561076042089695e-11
GC_1_203 b_1 NI_1 NS_203 0 -1.4862050536700992e-12
GC_1_204 b_1 NI_1 NS_204 0 1.6503533637686690e-11
GC_1_205 b_1 NI_1 NS_205 0 -5.6364933938874718e-07
GC_1_206 b_1 NI_1 NS_206 0 4.0935838158504715e-07
GC_1_207 b_1 NI_1 NS_207 0 -2.8795952928024670e-07
GC_1_208 b_1 NI_1 NS_208 0 1.5345503807726983e-06
GC_1_209 b_1 NI_1 NS_209 0 7.1636298814122615e-07
GC_1_210 b_1 NI_1 NS_210 0 -5.3800515958739559e-07
GC_1_211 b_1 NI_1 NS_211 0 -5.0824258465736391e-07
GC_1_212 b_1 NI_1 NS_212 0 2.2104028450888111e-06
GC_1_213 b_1 NI_1 NS_213 0 2.2909990647961379e-06
GC_1_214 b_1 NI_1 NS_214 0 -1.4800226174704842e-06
GC_1_215 b_1 NI_1 NS_215 0 -7.8890914683715793e-07
GC_1_216 b_1 NI_1 NS_216 0 9.3935833472566150e-07
GC_1_217 b_1 NI_1 NS_217 0 8.4704636416236091e-07
GC_1_218 b_1 NI_1 NS_218 0 7.6970617360841139e-08
GC_1_219 b_1 NI_1 NS_219 0 7.2184154615945984e-07
GC_1_220 b_1 NI_1 NS_220 0 5.7000023822011174e-07
GC_1_221 b_1 NI_1 NS_221 0 -1.1015629863834296e-09
GC_1_222 b_1 NI_1 NS_222 0 -2.6549958891719780e-11
GC_1_223 b_1 NI_1 NS_223 0 -5.3034840223828454e-13
GC_1_224 b_1 NI_1 NS_224 0 -6.8049665643590616e-12
GC_1_225 b_1 NI_1 NS_225 0 -5.8840398742393816e-08
GC_1_226 b_1 NI_1 NS_226 0 -6.1578144303334940e-07
GC_1_227 b_1 NI_1 NS_227 0 -3.4130228134294928e-07
GC_1_228 b_1 NI_1 NS_228 0 -1.0123465797124970e-07
GC_1_229 b_1 NI_1 NS_229 0 -1.1029923849319420e-06
GC_1_230 b_1 NI_1 NS_230 0 1.5334423106785697e-06
GC_1_231 b_1 NI_1 NS_231 0 6.9658928443120067e-07
GC_1_232 b_1 NI_1 NS_232 0 8.5933513051534568e-07
GC_1_233 b_1 NI_1 NS_233 0 2.1615730602530171e-06
GC_1_234 b_1 NI_1 NS_234 0 -1.4800255934375675e-06
GC_1_235 b_1 NI_1 NS_235 0 -1.9795094232726746e-07
GC_1_236 b_1 NI_1 NS_236 0 -9.9053906696821745e-07
GC_1_237 b_1 NI_1 NS_237 0 -1.0678574077154779e-06
GC_1_238 b_1 NI_1 NS_238 0 -4.1564960536129056e-07
GC_1_239 b_1 NI_1 NS_239 0 -4.0950187893463552e-07
GC_1_240 b_1 NI_1 NS_240 0 1.2021646057613325e-07
GD_1_1 b_1 NI_1 NA_1 0 -9.5068692159427804e-03
GD_1_2 b_1 NI_1 NA_2 0 5.5525392089087145e-03
GD_1_3 b_1 NI_1 NA_3 0 6.7730081992907008e-03
GD_1_4 b_1 NI_1 NA_4 0 -3.3302468896282736e-03
GD_1_5 b_1 NI_1 NA_5 0 1.5200615815968786e-05
GD_1_6 b_1 NI_1 NA_6 0 4.8447122923810510e-06
GD_1_7 b_1 NI_1 NA_7 0 -9.6392316489659132e-07
GD_1_8 b_1 NI_1 NA_8 0 1.0239339079594321e-05
GD_1_9 b_1 NI_1 NA_9 0 3.3803651775093737e-07
GD_1_10 b_1 NI_1 NA_10 0 -7.7230341037443803e-06
GD_1_11 b_1 NI_1 NA_11 0 -1.5460728728675082e-06
GD_1_12 b_1 NI_1 NA_12 0 3.4772174162415355e-07
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 8.9999190166085749e-05
GC_2_2 b_2 NI_2 NS_2 0 3.6211572619918142e-06
GC_2_3 b_2 NI_2 NS_3 0 5.9678538713479614e-09
GC_2_4 b_2 NI_2 NS_4 0 5.9667815251363812e-07
GC_2_5 b_2 NI_2 NS_5 0 4.7508813598207855e-02
GC_2_6 b_2 NI_2 NS_6 0 -9.6471254307658356e-03
GC_2_7 b_2 NI_2 NS_7 0 -4.5582968010781183e-02
GC_2_8 b_2 NI_2 NS_8 0 2.0552255624712346e-02
GC_2_9 b_2 NI_2 NS_9 0 -5.7696971352543966e-02
GC_2_10 b_2 NI_2 NS_10 0 -6.7350096687222555e-02
GC_2_11 b_2 NI_2 NS_11 0 6.3862106477352409e-02
GC_2_12 b_2 NI_2 NS_12 0 -2.2063600411148052e-02
GC_2_13 b_2 NI_2 NS_13 0 2.8382466276717130e-02
GC_2_14 b_2 NI_2 NS_14 0 8.9387906610425297e-02
GC_2_15 b_2 NI_2 NS_15 0 -5.4366402609714828e-02
GC_2_16 b_2 NI_2 NS_16 0 2.7979807087300688e-03
GC_2_17 b_2 NI_2 NS_17 0 -1.3847752516525336e-02
GC_2_18 b_2 NI_2 NS_18 0 -4.7095021041774848e-02
GC_2_19 b_2 NI_2 NS_19 0 1.6380501998999319e-02
GC_2_20 b_2 NI_2 NS_20 0 -3.9016241061821062e-02
GC_2_21 b_2 NI_2 NS_21 0 -1.5427134833673530e-05
GC_2_22 b_2 NI_2 NS_22 0 -3.7324314463540962e-06
GC_2_23 b_2 NI_2 NS_23 0 -2.3081208574536304e-08
GC_2_24 b_2 NI_2 NS_24 0 -3.8674152015128616e-07
GC_2_25 b_2 NI_2 NS_25 0 4.5760065321819726e-03
GC_2_26 b_2 NI_2 NS_26 0 3.7993286796473577e-03
GC_2_27 b_2 NI_2 NS_27 0 1.3872401175673038e-02
GC_2_28 b_2 NI_2 NS_28 0 -2.1406272364670773e-02
GC_2_29 b_2 NI_2 NS_29 0 -2.2493840945157176e-02
GC_2_30 b_2 NI_2 NS_30 0 2.6058892826137880e-02
GC_2_31 b_2 NI_2 NS_31 0 3.8337056193939921e-02
GC_2_32 b_2 NI_2 NS_32 0 -3.0181707170744677e-02
GC_2_33 b_2 NI_2 NS_33 0 -4.8685823011493809e-02
GC_2_34 b_2 NI_2 NS_34 0 1.9831379205208298e-02
GC_2_35 b_2 NI_2 NS_35 0 2.6967890308017828e-02
GC_2_36 b_2 NI_2 NS_36 0 -1.5945601193033197e-02
GC_2_37 b_2 NI_2 NS_37 0 -1.4394992250511275e-02
GC_2_38 b_2 NI_2 NS_38 0 6.8900418217841585e-03
GC_2_39 b_2 NI_2 NS_39 0 -4.8273798048063124e-03
GC_2_40 b_2 NI_2 NS_40 0 -1.6678597174271628e-02
GC_2_41 b_2 NI_2 NS_41 0 -1.8490432689311067e-06
GC_2_42 b_2 NI_2 NS_42 0 2.5677072774764679e-07
GC_2_43 b_2 NI_2 NS_43 0 1.6912981353217913e-09
GC_2_44 b_2 NI_2 NS_44 0 1.3611967492200204e-08
GC_2_45 b_2 NI_2 NS_45 0 1.1406455708583255e-03
GC_2_46 b_2 NI_2 NS_46 0 -2.1726046512128218e-03
GC_2_47 b_2 NI_2 NS_47 0 3.4952388385406201e-03
GC_2_48 b_2 NI_2 NS_48 0 -1.3003077419957746e-02
GC_2_49 b_2 NI_2 NS_49 0 -3.9401362309773112e-02
GC_2_50 b_2 NI_2 NS_50 0 -3.6437957861373019e-04
GC_2_51 b_2 NI_2 NS_51 0 -2.6247365013333229e-02
GC_2_52 b_2 NI_2 NS_52 0 2.8990158552302144e-02
GC_2_53 b_2 NI_2 NS_53 0 5.2202631961657302e-02
GC_2_54 b_2 NI_2 NS_54 0 3.8208680679658859e-02
GC_2_55 b_2 NI_2 NS_55 0 1.7572267735017501e-02
GC_2_56 b_2 NI_2 NS_56 0 -1.4394059592167791e-02
GC_2_57 b_2 NI_2 NS_57 0 -9.1651292323489640e-03
GC_2_58 b_2 NI_2 NS_58 0 -3.7458099120903140e-03
GC_2_59 b_2 NI_2 NS_59 0 8.0623396411401340e-03
GC_2_60 b_2 NI_2 NS_60 0 5.8595893032171754e-03
GC_2_61 b_2 NI_2 NS_61 0 -1.0355529880404218e-05
GC_2_62 b_2 NI_2 NS_62 0 -2.1274256833402216e-07
GC_2_63 b_2 NI_2 NS_63 0 -1.2832450400108521e-09
GC_2_64 b_2 NI_2 NS_64 0 -2.5390014001036675e-08
GC_2_65 b_2 NI_2 NS_65 0 -4.2497323834282267e-03
GC_2_66 b_2 NI_2 NS_66 0 -3.4927923471721749e-03
GC_2_67 b_2 NI_2 NS_67 0 -1.2922477450098393e-02
GC_2_68 b_2 NI_2 NS_68 0 1.7065692973002193e-02
GC_2_69 b_2 NI_2 NS_69 0 1.7371378752297752e-02
GC_2_70 b_2 NI_2 NS_70 0 -1.9446861927124425e-02
GC_2_71 b_2 NI_2 NS_71 0 -3.3168754752004551e-02
GC_2_72 b_2 NI_2 NS_72 0 2.5454292399461884e-02
GC_2_73 b_2 NI_2 NS_73 0 4.0789565934951817e-02
GC_2_74 b_2 NI_2 NS_74 0 -1.1433260033183347e-02
GC_2_75 b_2 NI_2 NS_75 0 -2.1059403287576946e-02
GC_2_76 b_2 NI_2 NS_76 0 1.5315262372466762e-02
GC_2_77 b_2 NI_2 NS_77 0 1.4123880964770012e-02
GC_2_78 b_2 NI_2 NS_78 0 -3.7536569665759900e-03
GC_2_79 b_2 NI_2 NS_79 0 7.0870158476398458e-03
GC_2_80 b_2 NI_2 NS_80 0 1.3573831644007557e-02
GC_2_81 b_2 NI_2 NS_81 0 1.9604852788726349e-09
GC_2_82 b_2 NI_2 NS_82 0 -2.0091526388615055e-10
GC_2_83 b_2 NI_2 NS_83 0 1.6947532415274508e-11
GC_2_84 b_2 NI_2 NS_84 0 -8.9399790297473540e-11
GC_2_85 b_2 NI_2 NS_85 0 -1.5357424455689392e-06
GC_2_86 b_2 NI_2 NS_86 0 -1.4180438831206701e-06
GC_2_87 b_2 NI_2 NS_87 0 -5.6306080906594459e-06
GC_2_88 b_2 NI_2 NS_88 0 1.3500657748422429e-05
GC_2_89 b_2 NI_2 NS_89 0 3.5171687032293902e-05
GC_2_90 b_2 NI_2 NS_90 0 1.0737047668327977e-05
GC_2_91 b_2 NI_2 NS_91 0 3.2592131103119838e-05
GC_2_92 b_2 NI_2 NS_92 0 -2.6154287044429459e-05
GC_2_93 b_2 NI_2 NS_93 0 -4.0882398407775127e-05
GC_2_94 b_2 NI_2 NS_94 0 -5.0757256993609718e-05
GC_2_95 b_2 NI_2 NS_95 0 -2.0190237784648093e-05
GC_2_96 b_2 NI_2 NS_96 0 9.6142443525415032e-06
GC_2_97 b_2 NI_2 NS_97 0 3.9350711279937617e-06
GC_2_98 b_2 NI_2 NS_98 0 1.2601215998924943e-07
GC_2_99 b_2 NI_2 NS_99 0 -1.3016677197569990e-05
GC_2_100 b_2 NI_2 NS_100 0 -6.9640875432022361e-06
GC_2_101 b_2 NI_2 NS_101 0 -2.7923125774226328e-08
GC_2_102 b_2 NI_2 NS_102 0 1.2536813934649216e-09
GC_2_103 b_2 NI_2 NS_103 0 -9.9739505539133315e-12
GC_2_104 b_2 NI_2 NS_104 0 2.3134353988249122e-11
GC_2_105 b_2 NI_2 NS_105 0 4.4587604978169435e-06
GC_2_106 b_2 NI_2 NS_106 0 2.3149763989935091e-06
GC_2_107 b_2 NI_2 NS_107 0 9.9868190898202963e-06
GC_2_108 b_2 NI_2 NS_108 0 9.7173874939187713e-06
GC_2_109 b_2 NI_2 NS_109 0 1.8696326367134671e-05
GC_2_110 b_2 NI_2 NS_110 0 -2.3425383884676492e-05
GC_2_111 b_2 NI_2 NS_111 0 1.1422717757635607e-05
GC_2_112 b_2 NI_2 NS_112 0 -3.1566161289885828e-06
GC_2_113 b_2 NI_2 NS_113 0 -6.8037249938342225e-06
GC_2_114 b_2 NI_2 NS_114 0 -5.3300295458185595e-05
GC_2_115 b_2 NI_2 NS_115 0 -1.4916969153581901e-05
GC_2_116 b_2 NI_2 NS_116 0 -1.7768778399842951e-05
GC_2_117 b_2 NI_2 NS_117 0 -2.7486796157655815e-05
GC_2_118 b_2 NI_2 NS_118 0 -1.2413931710816263e-05
GC_2_119 b_2 NI_2 NS_119 0 -1.9106840008349110e-05
GC_2_120 b_2 NI_2 NS_120 0 5.8361989575897929e-06
GC_2_121 b_2 NI_2 NS_121 0 -2.3908523234125537e-08
GC_2_122 b_2 NI_2 NS_122 0 1.2224989733165013e-09
GC_2_123 b_2 NI_2 NS_123 0 2.1485254456742414e-11
GC_2_124 b_2 NI_2 NS_124 0 -1.7590194319704380e-10
GC_2_125 b_2 NI_2 NS_125 0 1.8930936224716691e-06
GC_2_126 b_2 NI_2 NS_126 0 -4.2142294530380668e-06
GC_2_127 b_2 NI_2 NS_127 0 2.5243760144951360e-06
GC_2_128 b_2 NI_2 NS_128 0 5.0918948835923102e-08
GC_2_129 b_2 NI_2 NS_129 0 -1.6404747600687275e-06
GC_2_130 b_2 NI_2 NS_130 0 -4.6526885821658506e-06
GC_2_131 b_2 NI_2 NS_131 0 9.2496762166540442e-07
GC_2_132 b_2 NI_2 NS_132 0 -7.3960095786705500e-06
GC_2_133 b_2 NI_2 NS_133 0 -9.0332921936587167e-06
GC_2_134 b_2 NI_2 NS_134 0 -4.5741787561415314e-06
GC_2_135 b_2 NI_2 NS_135 0 -3.2971986365740275e-06
GC_2_136 b_2 NI_2 NS_136 0 1.4734746772318877e-06
GC_2_137 b_2 NI_2 NS_137 0 -1.9003383982323848e-06
GC_2_138 b_2 NI_2 NS_138 0 -4.7685587262859305e-07
GC_2_139 b_2 NI_2 NS_139 0 -3.2417996388603735e-06
GC_2_140 b_2 NI_2 NS_140 0 -1.4954314330784851e-06
GC_2_141 b_2 NI_2 NS_141 0 2.0308403902655277e-08
GC_2_142 b_2 NI_2 NS_142 0 -1.0039751858470065e-09
GC_2_143 b_2 NI_2 NS_143 0 -1.9110577895048245e-11
GC_2_144 b_2 NI_2 NS_144 0 1.5484026839687705e-10
GC_2_145 b_2 NI_2 NS_145 0 -1.0722359562227930e-06
GC_2_146 b_2 NI_2 NS_146 0 -8.5235515144468894e-07
GC_2_147 b_2 NI_2 NS_147 0 -1.9506686830661488e-06
GC_2_148 b_2 NI_2 NS_148 0 -1.2482927928276412e-08
GC_2_149 b_2 NI_2 NS_149 0 -3.0919926703168450e-06
GC_2_150 b_2 NI_2 NS_150 0 7.4445421550881869e-07
GC_2_151 b_2 NI_2 NS_151 0 -4.1324093158809334e-06
GC_2_152 b_2 NI_2 NS_152 0 4.2217629535418763e-06
GC_2_153 b_2 NI_2 NS_153 0 3.1598677310450003e-06
GC_2_154 b_2 NI_2 NS_154 0 5.3390135227791481e-06
GC_2_155 b_2 NI_2 NS_155 0 -9.0731364395962377e-07
GC_2_156 b_2 NI_2 NS_156 0 5.9324207748569021e-06
GC_2_157 b_2 NI_2 NS_157 0 5.9750962457929427e-06
GC_2_158 b_2 NI_2 NS_158 0 3.2313789873680945e-06
GC_2_159 b_2 NI_2 NS_159 0 5.7328775981044180e-06
GC_2_160 b_2 NI_2 NS_160 0 1.6826699780220596e-06
GC_2_161 b_2 NI_2 NS_161 0 -8.0862417481882517e-09
GC_2_162 b_2 NI_2 NS_162 0 6.7986839486542468e-10
GC_2_163 b_2 NI_2 NS_163 0 1.5646920700517975e-11
GC_2_164 b_2 NI_2 NS_164 0 -1.2067897764148527e-10
GC_2_165 b_2 NI_2 NS_165 0 -2.1903678985632206e-06
GC_2_166 b_2 NI_2 NS_166 0 2.1886701232454442e-07
GC_2_167 b_2 NI_2 NS_167 0 -2.1895685047983085e-06
GC_2_168 b_2 NI_2 NS_168 0 2.7884235887420626e-06
GC_2_169 b_2 NI_2 NS_169 0 -1.1327165606225950e-06
GC_2_170 b_2 NI_2 NS_170 0 6.5773529509389916e-06
GC_2_171 b_2 NI_2 NS_171 0 -4.1805363041955437e-07
GC_2_172 b_2 NI_2 NS_172 0 2.1422233725341662e-06
GC_2_173 b_2 NI_2 NS_173 0 7.2190734551721315e-06
GC_2_174 b_2 NI_2 NS_174 0 5.1224751283217904e-06
GC_2_175 b_2 NI_2 NS_175 0 1.6120647361843836e-06
GC_2_176 b_2 NI_2 NS_176 0 3.1394830292940118e-06
GC_2_177 b_2 NI_2 NS_177 0 4.8357482425744014e-06
GC_2_178 b_2 NI_2 NS_178 0 1.1501519105330648e-06
GC_2_179 b_2 NI_2 NS_179 0 2.9137167102917309e-06
GC_2_180 b_2 NI_2 NS_180 0 -1.3217668035907330e-06
GC_2_181 b_2 NI_2 NS_181 0 1.2088122144263996e-08
GC_2_182 b_2 NI_2 NS_182 0 -8.1496960457312789e-10
GC_2_183 b_2 NI_2 NS_183 0 -1.6058676906252965e-11
GC_2_184 b_2 NI_2 NS_184 0 1.3065452190541024e-10
GC_2_185 b_2 NI_2 NS_185 0 6.7658987941781301e-08
GC_2_186 b_2 NI_2 NS_186 0 -1.2554500534109858e-08
GC_2_187 b_2 NI_2 NS_187 0 -5.8630537147780822e-07
GC_2_188 b_2 NI_2 NS_188 0 5.6735526469643323e-07
GC_2_189 b_2 NI_2 NS_189 0 1.6812066593347299e-06
GC_2_190 b_2 NI_2 NS_190 0 -5.0520102910590609e-07
GC_2_191 b_2 NI_2 NS_191 0 -9.7641441693587768e-07
GC_2_192 b_2 NI_2 NS_192 0 1.1750298519143401e-07
GC_2_193 b_2 NI_2 NS_193 0 1.6591569763562076e-06
GC_2_194 b_2 NI_2 NS_194 0 -1.1492634252151207e-06
GC_2_195 b_2 NI_2 NS_195 0 -9.0302151436305048e-07
GC_2_196 b_2 NI_2 NS_196 0 -8.6140223471503724e-07
GC_2_197 b_2 NI_2 NS_197 0 -1.1367785483040083e-06
GC_2_198 b_2 NI_2 NS_198 0 -2.5235764802674883e-07
GC_2_199 b_2 NI_2 NS_199 0 8.6997582195573543e-08
GC_2_200 b_2 NI_2 NS_200 0 1.1717149430683317e-06
GC_2_201 b_2 NI_2 NS_201 0 -1.1046897993113746e-09
GC_2_202 b_2 NI_2 NS_202 0 -2.6299903039481296e-11
GC_2_203 b_2 NI_2 NS_203 0 -5.2637224831364711e-13
GC_2_204 b_2 NI_2 NS_204 0 -6.8308769529236783e-12
GC_2_205 b_2 NI_2 NS_205 0 -5.6995941193330348e-08
GC_2_206 b_2 NI_2 NS_206 0 -6.1544892377173382e-07
GC_2_207 b_2 NI_2 NS_207 0 -3.3915795639183863e-07
GC_2_208 b_2 NI_2 NS_208 0 -9.9907671104722794e-08
GC_2_209 b_2 NI_2 NS_209 0 -1.1012111807461664e-06
GC_2_210 b_2 NI_2 NS_210 0 1.5244120090490377e-06
GC_2_211 b_2 NI_2 NS_211 0 6.9375560335145676e-07
GC_2_212 b_2 NI_2 NS_212 0 8.5371679391019377e-07
GC_2_213 b_2 NI_2 NS_213 0 2.1527501889350394e-06
GC_2_214 b_2 NI_2 NS_214 0 -1.4741002469637863e-06
GC_2_215 b_2 NI_2 NS_215 0 -1.9736984512668063e-07
GC_2_216 b_2 NI_2 NS_216 0 -9.8761908922844942e-07
GC_2_217 b_2 NI_2 NS_217 0 -1.0659946076328012e-06
GC_2_218 b_2 NI_2 NS_218 0 -4.1594105812968707e-07
GC_2_219 b_2 NI_2 NS_219 0 -4.0970882085670685e-07
GC_2_220 b_2 NI_2 NS_220 0 1.1981977083908726e-07
GC_2_221 b_2 NI_2 NS_221 0 2.2395748087674939e-09
GC_2_222 b_2 NI_2 NS_222 0 -6.1558498738993909e-11
GC_2_223 b_2 NI_2 NS_223 0 -1.4861569372661307e-12
GC_2_224 b_2 NI_2 NS_224 0 1.6503232506218042e-11
GC_2_225 b_2 NI_2 NS_225 0 -5.6363581950771241e-07
GC_2_226 b_2 NI_2 NS_226 0 4.0935471619371628e-07
GC_2_227 b_2 NI_2 NS_227 0 -2.8794739183938974e-07
GC_2_228 b_2 NI_2 NS_228 0 1.5345560781331815e-06
GC_2_229 b_2 NI_2 NS_229 0 7.1637550141177257e-07
GC_2_230 b_2 NI_2 NS_230 0 -5.3803637853951479e-07
GC_2_231 b_2 NI_2 NS_231 0 -5.0822717986590916e-07
GC_2_232 b_2 NI_2 NS_232 0 2.2103913046970427e-06
GC_2_233 b_2 NI_2 NS_233 0 2.2909579048656214e-06
GC_2_234 b_2 NI_2 NS_234 0 -1.4800634842362092e-06
GC_2_235 b_2 NI_2 NS_235 0 -7.8891777831041268e-07
GC_2_236 b_2 NI_2 NS_236 0 9.3936142405522612e-07
GC_2_237 b_2 NI_2 NS_237 0 8.4703261567315227e-07
GC_2_238 b_2 NI_2 NS_238 0 7.6963614072742491e-08
GC_2_239 b_2 NI_2 NS_239 0 7.2183075636571366e-07
GC_2_240 b_2 NI_2 NS_240 0 5.7000291858870880e-07
GD_2_1 b_2 NI_2 NA_1 0 5.5524724040559364e-03
GD_2_2 b_2 NI_2 NA_2 0 -9.5068692159426971e-03
GD_2_3 b_2 NI_2 NA_3 0 -3.3302476158489414e-03
GD_2_4 b_2 NI_2 NA_4 0 6.7731249295636129e-03
GD_2_5 b_2 NI_2 NA_5 0 4.8451604085130311e-06
GD_2_6 b_2 NI_2 NA_6 0 1.4811101802870812e-05
GD_2_7 b_2 NI_2 NA_7 0 1.0254584292221343e-05
GD_2_8 b_2 NI_2 NA_8 0 -9.6795235974316782e-07
GD_2_9 b_2 NI_2 NA_9 0 -7.7230413691639899e-06
GD_2_10 b_2 NI_2 NA_10 0 3.1367551797316232e-07
GD_2_11 b_2 NI_2 NA_11 0 3.4974454918927533e-07
GD_2_12 b_2 NI_2 NA_12 0 -1.5460811361145363e-06
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 -1.0355529880404518e-05
GC_3_2 b_3 NI_3 NS_2 0 -2.1274256833408915e-07
GC_3_3 b_3 NI_3 NS_3 0 -1.2832450400069960e-09
GC_3_4 b_3 NI_3 NS_4 0 -2.5390014001067446e-08
GC_3_5 b_3 NI_3 NS_5 0 -4.2497323834282119e-03
GC_3_6 b_3 NI_3 NS_6 0 -3.4927923471721836e-03
GC_3_7 b_3 NI_3 NS_7 0 -1.2922477450098379e-02
GC_3_8 b_3 NI_3 NS_8 0 1.7065692973002162e-02
GC_3_9 b_3 NI_3 NS_9 0 1.7371378752297724e-02
GC_3_10 b_3 NI_3 NS_10 0 -1.9446861927124429e-02
GC_3_11 b_3 NI_3 NS_11 0 -3.3168754752004571e-02
GC_3_12 b_3 NI_3 NS_12 0 2.5454292399461891e-02
GC_3_13 b_3 NI_3 NS_13 0 4.0789565934951831e-02
GC_3_14 b_3 NI_3 NS_14 0 -1.1433260033183327e-02
GC_3_15 b_3 NI_3 NS_15 0 -2.1059403287576946e-02
GC_3_16 b_3 NI_3 NS_16 0 1.5315262372466762e-02
GC_3_17 b_3 NI_3 NS_17 0 1.4123880964770019e-02
GC_3_18 b_3 NI_3 NS_18 0 -3.7536569665759900e-03
GC_3_19 b_3 NI_3 NS_19 0 7.0870158476398467e-03
GC_3_20 b_3 NI_3 NS_20 0 1.3573831644007557e-02
GC_3_21 b_3 NI_3 NS_21 0 -1.8490438988644939e-06
GC_3_22 b_3 NI_3 NS_22 0 2.5677074680421776e-07
GC_3_23 b_3 NI_3 NS_23 0 1.6912981705721218e-09
GC_3_24 b_3 NI_3 NS_24 0 1.3611966370737097e-08
GC_3_25 b_3 NI_3 NS_25 0 1.1406457930701562e-03
GC_3_26 b_3 NI_3 NS_26 0 -2.1726047917648996e-03
GC_3_27 b_3 NI_3 NS_27 0 3.4952390751082796e-03
GC_3_28 b_3 NI_3 NS_28 0 -1.3003077589556929e-02
GC_3_29 b_3 NI_3 NS_29 0 -3.9401362309484780e-02
GC_3_30 b_3 NI_3 NS_30 0 -3.6438007419600717e-04
GC_3_31 b_3 NI_3 NS_31 0 -2.6247364909958073e-02
GC_3_32 b_3 NI_3 NS_32 0 2.8990158240220401e-02
GC_3_33 b_3 NI_3 NS_33 0 5.2202631407155385e-02
GC_3_34 b_3 NI_3 NS_34 0 3.8208680017635860e-02
GC_3_35 b_3 NI_3 NS_35 0 1.7572267423582623e-02
GC_3_36 b_3 NI_3 NS_36 0 -1.4394059869843325e-02
GC_3_37 b_3 NI_3 NS_37 0 -9.1651296869080055e-03
GC_3_38 b_3 NI_3 NS_38 0 -3.7458099411661243e-03
GC_3_39 b_3 NI_3 NS_39 0 8.0623393527399188e-03
GC_3_40 b_3 NI_3 NS_40 0 5.8595893506551335e-03
GC_3_41 b_3 NI_3 NS_41 0 -1.6276376083511130e-05
GC_3_42 b_3 NI_3 NS_42 0 -3.6835869480387372e-06
GC_3_43 b_3 NI_3 NS_43 0 -2.2928932972614377e-08
GC_3_44 b_3 NI_3 NS_44 0 -3.8914239402373816e-07
GC_3_45 b_3 NI_3 NS_45 0 4.5530397110479254e-03
GC_3_46 b_3 NI_3 NS_46 0 3.8169600042903522e-03
GC_3_47 b_3 NI_3 NS_47 0 1.3858626071957416e-02
GC_3_48 b_3 NI_3 NS_48 0 -2.1367083698543090e-02
GC_3_49 b_3 NI_3 NS_49 0 -2.2487121350575304e-02
GC_3_50 b_3 NI_3 NS_50 0 2.6079640325127895e-02
GC_3_51 b_3 NI_3 NS_51 0 3.8329043046791994e-02
GC_3_52 b_3 NI_3 NS_52 0 -3.0114597187179827e-02
GC_3_53 b_3 NI_3 NS_53 0 -4.8600025534500116e-02
GC_3_54 b_3 NI_3 NS_54 0 1.9841748148375499e-02
GC_3_55 b_3 NI_3 NS_55 0 2.6998114871042304e-02
GC_3_56 b_3 NI_3 NS_56 0 -1.5909282696620272e-02
GC_3_57 b_3 NI_3 NS_57 0 -1.4330190300066270e-02
GC_3_58 b_3 NI_3 NS_58 0 6.8408592040238494e-03
GC_3_59 b_3 NI_3 NS_59 0 -4.8601515355699071e-03
GC_3_60 b_3 NI_3 NS_60 0 -1.6721195153551638e-02
GC_3_61 b_3 NI_3 NS_61 0 8.9222503585804791e-05
GC_3_62 b_3 NI_3 NS_62 0 3.6749061774156831e-06
GC_3_63 b_3 NI_3 NS_63 0 6.5785472494238862e-09
GC_3_64 b_3 NI_3 NS_64 0 5.9211960324826194e-07
GC_3_65 b_3 NI_3 NS_65 0 4.7462853332893865e-02
GC_3_66 b_3 NI_3 NS_66 0 -9.5881597164119946e-03
GC_3_67 b_3 NI_3 NS_67 0 -4.5650675707979649e-02
GC_3_68 b_3 NI_3 NS_68 0 2.0563547184382663e-02
GC_3_69 b_3 NI_3 NS_69 0 -5.7680587918086536e-02
GC_3_70 b_3 NI_3 NS_70 0 -6.7211174157165571e-02
GC_3_71 b_3 NI_3 NS_71 0 6.3843296160758525e-02
GC_3_72 b_3 NI_3 NS_72 0 -2.1942062128457153e-02
GC_3_73 b_3 NI_3 NS_73 0 2.8542719293894115e-02
GC_3_74 b_3 NI_3 NS_74 0 8.9518926126440732e-02
GC_3_75 b_3 NI_3 NS_75 0 -5.4297956932849931e-02
GC_3_76 b_3 NI_3 NS_76 0 2.8478266776892974e-03
GC_3_77 b_3 NI_3 NS_77 0 -1.3713164323650252e-02
GC_3_78 b_3 NI_3 NS_78 0 -4.7078862498526913e-02
GC_3_79 b_3 NI_3 NS_79 0 1.6430654705521061e-02
GC_3_80 b_3 NI_3 NS_80 0 -3.9060974829509716e-02
GC_3_81 b_3 NI_3 NS_81 0 -5.4549210608330184e-08
GC_3_82 b_3 NI_3 NS_82 0 -2.0955089589676602e-09
GC_3_83 b_3 NI_3 NS_83 0 -1.0056422574831398e-10
GC_3_84 b_3 NI_3 NS_84 0 3.2111226395797933e-10
GC_3_85 b_3 NI_3 NS_85 0 -1.3498608773630498e-05
GC_3_86 b_3 NI_3 NS_86 0 -1.1749813954730540e-05
GC_3_87 b_3 NI_3 NS_87 0 -4.4778893554938589e-05
GC_3_88 b_3 NI_3 NS_88 0 4.2451447189743566e-05
GC_3_89 b_3 NI_3 NS_89 0 4.9954079145832937e-05
GC_3_90 b_3 NI_3 NS_90 0 -4.4097075711862196e-05
GC_3_91 b_3 NI_3 NS_91 0 -1.0686413605100913e-04
GC_3_92 b_3 NI_3 NS_92 0 6.6403484143851292e-05
GC_3_93 b_3 NI_3 NS_93 0 1.2727377646230102e-04
GC_3_94 b_3 NI_3 NS_94 0 -7.6158834385833419e-06
GC_3_95 b_3 NI_3 NS_95 0 -5.8523906738008992e-05
GC_3_96 b_3 NI_3 NS_96 0 4.1104294135137665e-05
GC_3_97 b_3 NI_3 NS_97 0 4.5420874071449214e-05
GC_3_98 b_3 NI_3 NS_98 0 -5.0322590373786632e-06
GC_3_99 b_3 NI_3 NS_99 0 2.5831324828247464e-05
GC_3_100 b_3 NI_3 NS_100 0 3.8190405596921607e-05
GC_3_101 b_3 NI_3 NS_101 0 6.1704204611500170e-08
GC_3_102 b_3 NI_3 NS_102 0 1.2660808026659556e-09
GC_3_103 b_3 NI_3 NS_103 0 1.6398710172210104e-10
GC_3_104 b_3 NI_3 NS_104 0 -6.8655449777241208e-10
GC_3_105 b_3 NI_3 NS_105 0 -1.0004015498735078e-05
GC_3_106 b_3 NI_3 NS_106 0 -5.4826723330268039e-06
GC_3_107 b_3 NI_3 NS_107 0 1.5174730675954420e-06
GC_3_108 b_3 NI_3 NS_108 0 -1.4462000377827409e-05
GC_3_109 b_3 NI_3 NS_109 0 -1.1184072756880178e-04
GC_3_110 b_3 NI_3 NS_110 0 3.9184477241259155e-05
GC_3_111 b_3 NI_3 NS_111 0 -7.9769108318366932e-05
GC_3_112 b_3 NI_3 NS_112 0 7.8276874556310719e-05
GC_3_113 b_3 NI_3 NS_113 0 1.9275207558602618e-04
GC_3_114 b_3 NI_3 NS_114 0 1.3386994113989069e-04
GC_3_115 b_3 NI_3 NS_115 0 5.7427660497060864e-05
GC_3_116 b_3 NI_3 NS_116 0 -1.9414654753774555e-05
GC_3_117 b_3 NI_3 NS_117 0 -4.7733075781125739e-06
GC_3_118 b_3 NI_3 NS_118 0 -8.4252422978962683e-06
GC_3_119 b_3 NI_3 NS_119 0 3.7519337703540680e-05
GC_3_120 b_3 NI_3 NS_120 0 9.6450131856198730e-06
GC_3_121 b_3 NI_3 NS_121 0 -2.8873926576664789e-08
GC_3_122 b_3 NI_3 NS_122 0 8.6794397828226697e-10
GC_3_123 b_3 NI_3 NS_123 0 -1.4875501391169310e-11
GC_3_124 b_3 NI_3 NS_124 0 6.7611109103727131e-11
GC_3_125 b_3 NI_3 NS_125 0 4.0217078483307668e-06
GC_3_126 b_3 NI_3 NS_126 0 2.7674566954845836e-06
GC_3_127 b_3 NI_3 NS_127 0 9.4641818359249975e-06
GC_3_128 b_3 NI_3 NS_128 0 1.0309426283756137e-05
GC_3_129 b_3 NI_3 NS_129 0 1.9370375353955013e-05
GC_3_130 b_3 NI_3 NS_130 0 -2.2294981716770753e-05
GC_3_131 b_3 NI_3 NS_131 0 1.1424263074155789e-05
GC_3_132 b_3 NI_3 NS_132 0 -2.5122773266785977e-06
GC_3_133 b_3 NI_3 NS_133 0 -4.9910962902228301e-06
GC_3_134 b_3 NI_3 NS_134 0 -5.2807265709480471e-05
GC_3_135 b_3 NI_3 NS_135 0 -1.4282076751128546e-05
GC_3_136 b_3 NI_3 NS_136 0 -1.7913591378453619e-05
GC_3_137 b_3 NI_3 NS_137 0 -2.7057560633672118e-05
GC_3_138 b_3 NI_3 NS_138 0 -1.2982227856194106e-05
GC_3_139 b_3 NI_3 NS_139 0 -1.9361092732665781e-05
GC_3_140 b_3 NI_3 NS_140 0 5.4944462469671546e-06
GC_3_141 b_3 NI_3 NS_141 0 8.5556734467643192e-09
GC_3_142 b_3 NI_3 NS_142 0 -6.8782359327380786e-11
GC_3_143 b_3 NI_3 NS_143 0 1.9395383795071008e-11
GC_3_144 b_3 NI_3 NS_144 0 -1.1529159218652285e-10
GC_3_145 b_3 NI_3 NS_145 0 -2.0028562967330632e-06
GC_3_146 b_3 NI_3 NS_146 0 -1.3631238950097677e-06
GC_3_147 b_3 NI_3 NS_147 0 -6.1770683286078986e-06
GC_3_148 b_3 NI_3 NS_148 0 1.3444025449663790e-05
GC_3_149 b_3 NI_3 NS_149 0 3.4355390258455108e-05
GC_3_150 b_3 NI_3 NS_150 0 1.2051900647873328e-05
GC_3_151 b_3 NI_3 NS_151 0 3.1744499708276636e-05
GC_3_152 b_3 NI_3 NS_152 0 -2.5606784189652760e-05
GC_3_153 b_3 NI_3 NS_153 0 -3.9672992449617925e-05
GC_3_154 b_3 NI_3 NS_154 0 -4.8329186141366939e-05
GC_3_155 b_3 NI_3 NS_155 0 -2.0078434701598177e-05
GC_3_156 b_3 NI_3 NS_156 0 1.0823486275999271e-05
GC_3_157 b_3 NI_3 NS_157 0 5.4292695568741710e-06
GC_3_158 b_3 NI_3 NS_158 0 1.5199028266985819e-06
GC_3_159 b_3 NI_3 NS_159 0 -1.0987725731552888e-05
GC_3_160 b_3 NI_3 NS_160 0 -6.5992097941249840e-06
GC_3_161 b_3 NI_3 NS_161 0 -3.3864674725516121e-10
GC_3_162 b_3 NI_3 NS_162 0 2.4529398445319242e-10
GC_3_163 b_3 NI_3 NS_163 0 5.1902615261627132e-12
GC_3_164 b_3 NI_3 NS_164 0 -1.2433846629163551e-11
GC_3_165 b_3 NI_3 NS_165 0 -1.5827626811463050e-06
GC_3_166 b_3 NI_3 NS_166 0 7.4475369069846336e-07
GC_3_167 b_3 NI_3 NS_167 0 -2.4991303745999922e-06
GC_3_168 b_3 NI_3 NS_168 0 1.5671831500026475e-06
GC_3_169 b_3 NI_3 NS_169 0 6.6684087571416742e-07
GC_3_170 b_3 NI_3 NS_170 0 3.1009811081154088e-06
GC_3_171 b_3 NI_3 NS_171 0 -2.4062952858700963e-06
GC_3_172 b_3 NI_3 NS_172 0 3.2308237351507997e-06
GC_3_173 b_3 NI_3 NS_173 0 5.2075167856537086e-06
GC_3_174 b_3 NI_3 NS_174 0 4.2312117262503590e-06
GC_3_175 b_3 NI_3 NS_175 0 -6.0809239945553697e-08
GC_3_176 b_3 NI_3 NS_176 0 3.4339391251201637e-06
GC_3_177 b_3 NI_3 NS_177 0 5.0339041861181077e-06
GC_3_178 b_3 NI_3 NS_178 0 2.2607893496869355e-06
GC_3_179 b_3 NI_3 NS_179 0 3.8677360878047681e-06
GC_3_180 b_3 NI_3 NS_180 0 2.0110295890484790e-07
GC_3_181 b_3 NI_3 NS_181 0 -5.4833814467484070e-09
GC_3_182 b_3 NI_3 NS_182 0 -1.1889748466481436e-10
GC_3_183 b_3 NI_3 NS_183 0 -8.7976138207791731e-12
GC_3_184 b_3 NI_3 NS_184 0 1.2303218485222241e-11
GC_3_185 b_3 NI_3 NS_185 0 2.8877995719496378e-06
GC_3_186 b_3 NI_3 NS_186 0 -3.3700212519888746e-06
GC_3_187 b_3 NI_3 NS_187 0 3.9433199743612119e-06
GC_3_188 b_3 NI_3 NS_188 0 -1.1977393726373229e-06
GC_3_189 b_3 NI_3 NS_189 0 -1.9626918729766032e-06
GC_3_190 b_3 NI_3 NS_190 0 -6.4897711656872423e-06
GC_3_191 b_3 NI_3 NS_191 0 1.2536646758761601e-06
GC_3_192 b_3 NI_3 NS_192 0 -5.0193344574078501e-06
GC_3_193 b_3 NI_3 NS_193 0 -3.5332533464715268e-06
GC_3_194 b_3 NI_3 NS_194 0 -9.5121434827749131e-06
GC_3_195 b_3 NI_3 NS_195 0 -2.5204736747884079e-06
GC_3_196 b_3 NI_3 NS_196 0 -6.0280721378257165e-06
GC_3_197 b_3 NI_3 NS_197 0 -9.7106992562458986e-06
GC_3_198 b_3 NI_3 NS_198 0 -4.8418374803948609e-06
GC_3_199 b_3 NI_3 NS_199 0 -7.2832410780474679e-06
GC_3_200 b_3 NI_3 NS_200 0 5.3200546492472691e-07
GC_3_201 b_3 NI_3 NS_201 0 1.2106006956954586e-08
GC_3_202 b_3 NI_3 NS_202 0 -8.1607725955684340e-10
GC_3_203 b_3 NI_3 NS_203 0 -1.6069712823546570e-11
GC_3_204 b_3 NI_3 NS_204 0 1.3075628238106635e-10
GC_3_205 b_3 NI_3 NS_205 0 6.7316822588730167e-08
GC_3_206 b_3 NI_3 NS_206 0 -1.0258733780435687e-08
GC_3_207 b_3 NI_3 NS_207 0 -5.8672885351322148e-07
GC_3_208 b_3 NI_3 NS_208 0 5.6507220738065023e-07
GC_3_209 b_3 NI_3 NS_209 0 1.6793028872568002e-06
GC_3_210 b_3 NI_3 NS_210 0 -4.9707775017724074e-07
GC_3_211 b_3 NI_3 NS_211 0 -9.7352485421797951e-07
GC_3_212 b_3 NI_3 NS_212 0 1.1756511766500204e-07
GC_3_213 b_3 NI_3 NS_213 0 1.6616849728960241e-06
GC_3_214 b_3 NI_3 NS_214 0 -1.1455584703510304e-06
GC_3_215 b_3 NI_3 NS_215 0 -9.0102798840054306e-07
GC_3_216 b_3 NI_3 NS_216 0 -8.6217891943433918e-07
GC_3_217 b_3 NI_3 NS_217 0 -1.1351757070676733e-06
GC_3_218 b_3 NI_3 NS_218 0 -2.5009878316923763e-07
GC_3_219 b_3 NI_3 NS_219 0 8.9211369333922681e-08
GC_3_220 b_3 NI_3 NS_220 0 1.1707706689430232e-06
GC_3_221 b_3 NI_3 NS_221 0 -8.0831890802940624e-09
GC_3_222 b_3 NI_3 NS_222 0 6.7951711470364199e-10
GC_3_223 b_3 NI_3 NS_223 0 1.5642915009344743e-11
GC_3_224 b_3 NI_3 NS_224 0 -1.2064088754624331e-10
GC_3_225 b_3 NI_3 NS_225 0 -2.1882725635612118e-06
GC_3_226 b_3 NI_3 NS_226 0 2.1734553743875468e-07
GC_3_227 b_3 NI_3 NS_227 0 -2.1912528558260467e-06
GC_3_228 b_3 NI_3 NS_228 0 2.7906333776331638e-06
GC_3_229 b_3 NI_3 NS_229 0 -1.1302477192788392e-06
GC_3_230 b_3 NI_3 NS_230 0 6.5760336575148070e-06
GC_3_231 b_3 NI_3 NS_231 0 -4.1809920509408275e-07
GC_3_232 b_3 NI_3 NS_232 0 2.1387821923278500e-06
GC_3_233 b_3 NI_3 NS_233 0 7.2163468082858510e-06
GC_3_234 b_3 NI_3 NS_234 0 5.1185253122720565e-06
GC_3_235 b_3 NI_3 NS_235 0 1.6097745885896683e-06
GC_3_236 b_3 NI_3 NS_236 0 3.1433821168253118e-06
GC_3_237 b_3 NI_3 NS_237 0 4.8364254637692954e-06
GC_3_238 b_3 NI_3 NS_238 0 1.1505222941834284e-06
GC_3_239 b_3 NI_3 NS_239 0 2.9136130509841236e-06
GC_3_240 b_3 NI_3 NS_240 0 -1.3226685510506915e-06
GD_3_1 b_3 NI_3 NA_1 0 6.7731249295635886e-03
GD_3_2 b_3 NI_3 NA_2 0 -3.3302469036985542e-03
GD_3_3 b_3 NI_3 NA_3 0 -9.5852748204677332e-03
GD_3_4 b_3 NI_3 NA_4 0 5.3317577349758878e-03
GD_3_5 b_3 NI_3 NA_5 0 2.2411103750888878e-05
GD_3_6 b_3 NI_3 NA_6 0 -5.5822644697282615e-05
GD_3_7 b_3 NI_3 NA_7 0 1.3060694789158776e-05
GD_3_8 b_3 NI_3 NA_8 0 3.5140059858188311e-06
GD_3_9 b_3 NI_3 NA_9 0 -5.2908402367067881e-06
GD_3_10 b_3 NI_3 NA_10 0 1.2166293037161280e-05
GD_3_11 b_3 NI_3 NA_11 0 3.0621156193219034e-07
GD_3_12 b_3 NI_3 NA_12 0 -7.7232171148659777e-06
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 -1.8490432701957148e-06
GC_4_2 b_4 NI_4 NS_2 0 2.5677072811178663e-07
GC_4_3 b_4 NI_4 NS_3 0 1.6912978303957608e-09
GC_4_4 b_4 NI_4 NS_4 0 1.3611967604735484e-08
GC_4_5 b_4 NI_4 NS_5 0 1.1406455706463846e-03
GC_4_6 b_4 NI_4 NS_6 0 -2.1726046514023395e-03
GC_4_7 b_4 NI_4 NS_7 0 3.4952388382647509e-03
GC_4_8 b_4 NI_4 NS_8 0 -1.3003077420434843e-02
GC_4_9 b_4 NI_4 NS_9 0 -3.9401362311358497e-02
GC_4_10 b_4 NI_4 NS_10 0 -3.6437957826918277e-04
GC_4_11 b_4 NI_4 NS_11 0 -2.6247365014822440e-02
GC_4_12 b_4 NI_4 NS_12 0 2.8990158553066792e-02
GC_4_13 b_4 NI_4 NS_13 0 5.2202631962548061e-02
GC_4_14 b_4 NI_4 NS_14 0 3.8208680683020892e-02
GC_4_15 b_4 NI_4 NS_15 0 1.7572267735831874e-02
GC_4_16 b_4 NI_4 NS_16 0 -1.4394059590820482e-02
GC_4_17 b_4 NI_4 NS_17 0 -9.1651292305929867e-03
GC_4_18 b_4 NI_4 NS_18 0 -3.7458099115582405e-03
GC_4_19 b_4 NI_4 NS_19 0 8.0623396423227956e-03
GC_4_20 b_4 NI_4 NS_20 0 5.8595893030517938e-03
GC_4_21 b_4 NI_4 NS_21 0 -1.0356264848365143e-05
GC_4_22 b_4 NI_4 NS_22 0 -2.1272069476427758e-07
GC_4_23 b_4 NI_4 NS_23 0 -1.2831320148477391e-09
GC_4_24 b_4 NI_4 NS_24 0 -2.5390347645561548e-08
GC_4_25 b_4 NI_4 NS_25 0 -4.2497281814668263e-03
GC_4_26 b_4 NI_4 NS_26 0 -3.4927766090990351e-03
GC_4_27 b_4 NI_4 NS_27 0 -1.2922365127891394e-02
GC_4_28 b_4 NI_4 NS_28 0 1.7065796230691495e-02
GC_4_29 b_4 NI_4 NS_29 0 1.7371354225988570e-02
GC_4_30 b_4 NI_4 NS_30 0 -1.9447062637169003e-02
GC_4_31 b_4 NI_4 NS_31 0 -3.3168706678817911e-02
GC_4_32 b_4 NI_4 NS_32 0 2.5454421766033526e-02
GC_4_33 b_4 NI_4 NS_33 0 4.0789606058407431e-02
GC_4_34 b_4 NI_4 NS_34 0 -1.1433470437631318e-02
GC_4_35 b_4 NI_4 NS_35 0 -2.1059355346524665e-02
GC_4_36 b_4 NI_4 NS_36 0 1.5315260733975079e-02
GC_4_37 b_4 NI_4 NS_37 0 1.4123842664329872e-02
GC_4_38 b_4 NI_4 NS_38 0 -3.7538561739732593e-03
GC_4_39 b_4 NI_4 NS_39 0 7.0868353733450958e-03
GC_4_40 b_4 NI_4 NS_40 0 1.3573780074925441e-02
GC_4_41 b_4 NI_4 NS_41 0 8.9222419501535527e-05
GC_4_42 b_4 NI_4 NS_42 0 3.6749132353070791e-06
GC_4_43 b_4 NI_4 NS_43 0 6.5786641838421933e-09
GC_4_44 b_4 NI_4 NS_44 0 5.9211884765179745e-07
GC_4_45 b_4 NI_4 NS_45 0 4.7462887092685216e-02
GC_4_46 b_4 NI_4 NS_46 0 -9.5881529940481589e-03
GC_4_47 b_4 NI_4 NS_47 0 -4.5650645617307077e-02
GC_4_48 b_4 NI_4 NS_48 0 2.0563576716745340e-02
GC_4_49 b_4 NI_4 NS_49 0 -5.7680546160371965e-02
GC_4_50 b_4 NI_4 NS_50 0 -6.7211347487177803e-02
GC_4_51 b_4 NI_4 NS_51 0 6.3843233987005477e-02
GC_4_52 b_4 NI_4 NS_52 0 -2.1942170418654840e-02
GC_4_53 b_4 NI_4 NS_53 0 2.8542538099582470e-02
GC_4_54 b_4 NI_4 NS_54 0 8.9519055461347030e-02
GC_4_55 b_4 NI_4 NS_55 0 -5.4297952568354707e-02
GC_4_56 b_4 NI_4 NS_56 0 2.8479060360913334e-03
GC_4_57 b_4 NI_4 NS_57 0 -1.3713101282009938e-02
GC_4_58 b_4 NI_4 NS_58 0 -4.7078848688976119e-02
GC_4_59 b_4 NI_4 NS_59 0 1.6430668105227891e-02
GC_4_60 b_4 NI_4 NS_60 0 -3.9060986405084652e-02
GC_4_61 b_4 NI_4 NS_61 0 -1.6276376083510920e-05
GC_4_62 b_4 NI_4 NS_62 0 -3.6835869480389367e-06
GC_4_63 b_4 NI_4 NS_63 0 -2.2928932972616687e-08
GC_4_64 b_4 NI_4 NS_64 0 -3.8914239402371439e-07
GC_4_65 b_4 NI_4 NS_65 0 4.5530397110479098e-03
GC_4_66 b_4 NI_4 NS_66 0 3.8169600042903635e-03
GC_4_67 b_4 NI_4 NS_67 0 1.3858626071957382e-02
GC_4_68 b_4 NI_4 NS_68 0 -2.1367083698543059e-02
GC_4_69 b_4 NI_4 NS_69 0 -2.2487121350575259e-02
GC_4_70 b_4 NI_4 NS_70 0 2.6079640325127912e-02
GC_4_71 b_4 NI_4 NS_71 0 3.8329043046791959e-02
GC_4_72 b_4 NI_4 NS_72 0 -3.0114597187179806e-02
GC_4_73 b_4 NI_4 NS_73 0 -4.8600025534500046e-02
GC_4_74 b_4 NI_4 NS_74 0 1.9841748148375554e-02
GC_4_75 b_4 NI_4 NS_75 0 2.6998114871042325e-02
GC_4_76 b_4 NI_4 NS_76 0 -1.5909282696620251e-02
GC_4_77 b_4 NI_4 NS_77 0 -1.4330190300066234e-02
GC_4_78 b_4 NI_4 NS_78 0 6.8408592040238433e-03
GC_4_79 b_4 NI_4 NS_79 0 -4.8601515355698923e-03
GC_4_80 b_4 NI_4 NS_80 0 -1.6721195153551641e-02
GC_4_81 b_4 NI_4 NS_81 0 6.1677766343849838e-08
GC_4_82 b_4 NI_4 NS_82 0 1.2669494224174599e-09
GC_4_83 b_4 NI_4 NS_83 0 1.6399362866972895e-10
GC_4_84 b_4 NI_4 NS_84 0 -6.8660941723314503e-10
GC_4_85 b_4 NI_4 NS_85 0 -1.0021558047793940e-05
GC_4_86 b_4 NI_4 NS_86 0 -5.4883439806934467e-06
GC_4_87 b_4 NI_4 NS_87 0 1.4900704373333057e-06
GC_4_88 b_4 NI_4 NS_88 0 -1.4479541823707826e-05
GC_4_89 b_4 NI_4 NS_89 0 -1.1185421230508268e-04
GC_4_90 b_4 NI_4 NS_90 0 3.9288817160982158e-05
GC_4_91 b_4 NI_4 NS_91 0 -7.9728855875448563e-05
GC_4_92 b_4 NI_4 NS_92 0 7.8341206766294489e-05
GC_4_93 b_4 NI_4 NS_93 0 1.9284808419524834e-04
GC_4_94 b_4 NI_4 NS_94 0 1.3377504041656453e-04
GC_4_95 b_4 NI_4 NS_95 0 5.7410792430328639e-05
GC_4_96 b_4 NI_4 NS_96 0 -1.9453200939423888e-05
GC_4_97 b_4 NI_4 NS_97 0 -4.8009480197536796e-06
GC_4_98 b_4 NI_4 NS_98 0 -8.4210384618054360e-06
GC_4_99 b_4 NI_4 NS_99 0 3.7514588743837150e-05
GC_4_100 b_4 NI_4 NS_100 0 9.6476630184289767e-06
GC_4_101 b_4 NI_4 NS_101 0 -5.4561561068293565e-08
GC_4_102 b_4 NI_4 NS_102 0 -2.0950021925183736e-09
GC_4_103 b_4 NI_4 NS_103 0 -1.0056334578832291e-10
GC_4_104 b_4 NI_4 NS_104 0 3.2108262567304042e-10
GC_4_105 b_4 NI_4 NS_105 0 -1.3498690865487997e-05
GC_4_106 b_4 NI_4 NS_106 0 -1.1750814233770695e-05
GC_4_107 b_4 NI_4 NS_107 0 -4.4779272935724558e-05
GC_4_108 b_4 NI_4 NS_108 0 4.2450788885289540e-05
GC_4_109 b_4 NI_4 NS_109 0 4.9954070167012760e-05
GC_4_110 b_4 NI_4 NS_110 0 -4.4097729395530223e-05
GC_4_111 b_4 NI_4 NS_111 0 -1.0686547177891550e-04
GC_4_112 b_4 NI_4 NS_112 0 6.6401822178292926e-05
GC_4_113 b_4 NI_4 NS_113 0 1.2727304651976258e-04
GC_4_114 b_4 NI_4 NS_114 0 -7.6138314080397109e-06
GC_4_115 b_4 NI_4 NS_115 0 -5.8523238301711753e-05
GC_4_116 b_4 NI_4 NS_116 0 4.1103429169409825e-05
GC_4_117 b_4 NI_4 NS_117 0 4.5420168059158734e-05
GC_4_118 b_4 NI_4 NS_118 0 -5.0333340820386233e-06
GC_4_119 b_4 NI_4 NS_119 0 2.5829953018934378e-05
GC_4_120 b_4 NI_4 NS_120 0 3.8189923677398833e-05
GC_4_121 b_4 NI_4 NS_121 0 8.5552374072510627e-09
GC_4_122 b_4 NI_4 NS_122 0 -6.8743751083017320e-11
GC_4_123 b_4 NI_4 NS_123 0 1.9395779480082281e-11
GC_4_124 b_4 NI_4 NS_124 0 -1.1529477964491152e-10
GC_4_125 b_4 NI_4 NS_125 0 -2.0030697019467825e-06
GC_4_126 b_4 NI_4 NS_126 0 -1.3631112372404010e-06
GC_4_127 b_4 NI_4 NS_127 0 -6.1775750385786398e-06
GC_4_128 b_4 NI_4 NS_128 0 1.3443933038774419e-05
GC_4_129 b_4 NI_4 NS_129 0 3.4355404835467198e-05
GC_4_130 b_4 NI_4 NS_130 0 1.2053255053106789e-05
GC_4_131 b_4 NI_4 NS_131 0 3.1744906971074869e-05
GC_4_132 b_4 NI_4 NS_132 0 -2.5605882951053705e-05
GC_4_133 b_4 NI_4 NS_133 0 -3.9671497342349534e-05
GC_4_134 b_4 NI_4 NS_134 0 -4.8330196162698599e-05
GC_4_135 b_4 NI_4 NS_135 0 -2.0078507057459110e-05
GC_4_136 b_4 NI_4 NS_136 0 1.0823027997846755e-05
GC_4_137 b_4 NI_4 NS_137 0 5.4289939198273120e-06
GC_4_138 b_4 NI_4 NS_138 0 1.5197978448762857e-06
GC_4_139 b_4 NI_4 NS_139 0 -1.0987816924257252e-05
GC_4_140 b_4 NI_4 NS_140 0 -6.5991928129225256e-06
GC_4_141 b_4 NI_4 NS_141 0 -2.9031622171304460e-08
GC_4_142 b_4 NI_4 NS_142 0 8.7636030709564117e-10
GC_4_143 b_4 NI_4 NS_143 0 -1.4816261998091007e-11
GC_4_144 b_4 NI_4 NS_144 0 6.7054218521014788e-11
GC_4_145 b_4 NI_4 NS_145 0 4.0592951735025578e-06
GC_4_146 b_4 NI_4 NS_146 0 2.6907844350418541e-06
GC_4_147 b_4 NI_4 NS_147 0 9.4653612161286075e-06
GC_4_148 b_4 NI_4 NS_148 0 1.0215857384098309e-05
GC_4_149 b_4 NI_4 NS_149 0 1.9372833183751840e-05
GC_4_150 b_4 NI_4 NS_150 0 -2.2384281659024826e-05
GC_4_151 b_4 NI_4 NS_151 0 1.1343539511849331e-05
GC_4_152 b_4 NI_4 NS_152 0 -2.6952227890324833e-06
GC_4_153 b_4 NI_4 NS_153 0 -5.1382559186932719e-06
GC_4_154 b_4 NI_4 NS_154 0 -5.2745958064313502e-05
GC_4_155 b_4 NI_4 NS_155 0 -1.4325005209326608e-05
GC_4_156 b_4 NI_4 NS_156 0 -1.8002955613140436e-05
GC_4_157 b_4 NI_4 NS_157 0 -2.7149276257855480e-05
GC_4_158 b_4 NI_4 NS_158 0 -1.2989279815600287e-05
GC_4_159 b_4 NI_4 NS_159 0 -1.9441644717617884e-05
GC_4_160 b_4 NI_4 NS_160 0 5.4890785512462912e-06
GC_4_161 b_4 NI_4 NS_161 0 -5.4818371649066236e-09
GC_4_162 b_4 NI_4 NS_162 0 -1.1901796049475389e-10
GC_4_163 b_4 NI_4 NS_163 0 -8.7994518695916208e-12
GC_4_164 b_4 NI_4 NS_164 0 1.2315142963664801e-11
GC_4_165 b_4 NI_4 NS_165 0 2.8858211537417031e-06
GC_4_166 b_4 NI_4 NS_166 0 -3.3702242116261308e-06
GC_4_167 b_4 NI_4 NS_167 0 3.9410259368147069e-06
GC_4_168 b_4 NI_4 NS_168 0 -1.1989223234137028e-06
GC_4_169 b_4 NI_4 NS_169 0 -1.9642433880287631e-06
GC_4_170 b_4 NI_4 NS_170 0 -6.4802158723046093e-06
GC_4_171 b_4 NI_4 NS_171 0 1.2567716824085263e-06
GC_4_172 b_4 NI_4 NS_172 0 -5.0134050233295088e-06
GC_4_173 b_4 NI_4 NS_173 0 -3.5237885585713972e-06
GC_4_174 b_4 NI_4 NS_174 0 -9.5185281593917652e-06
GC_4_175 b_4 NI_4 NS_175 0 -2.5209703585581226e-06
GC_4_176 b_4 NI_4 NS_176 0 -6.0312525650058470e-06
GC_4_177 b_4 NI_4 NS_177 0 -9.7127123453665514e-06
GC_4_178 b_4 NI_4 NS_178 0 -4.8417688883052603e-06
GC_4_179 b_4 NI_4 NS_179 0 -7.2832299507205544e-06
GC_4_180 b_4 NI_4 NS_180 0 5.3233994989961372e-07
GC_4_181 b_4 NI_4 NS_181 0 -3.3859883087635165e-10
GC_4_182 b_4 NI_4 NS_182 0 2.4529151661449522e-10
GC_4_183 b_4 NI_4 NS_183 0 5.1902204304678520e-12
GC_4_184 b_4 NI_4 NS_184 0 -1.2433599528851051e-11
GC_4_185 b_4 NI_4 NS_185 0 -1.5827743464796938e-06
GC_4_186 b_4 NI_4 NS_186 0 7.4475466439671627e-07
GC_4_187 b_4 NI_4 NS_187 0 -2.4991417266455317e-06
GC_4_188 b_4 NI_4 NS_188 0 1.5671735056923162e-06
GC_4_189 b_4 NI_4 NS_189 0 6.6682294953050091e-07
GC_4_190 b_4 NI_4 NS_190 0 3.1010091667621887e-06
GC_4_191 b_4 NI_4 NS_191 0 -2.4063142448289807e-06
GC_4_192 b_4 NI_4 NS_192 0 3.2308341364502626e-06
GC_4_193 b_4 NI_4 NS_193 0 5.2075548560408698e-06
GC_4_194 b_4 NI_4 NS_194 0 4.2312570220811752e-06
GC_4_195 b_4 NI_4 NS_195 0 -6.0801452312503040e-08
GC_4_196 b_4 NI_4 NS_196 0 3.4339368915667544e-06
GC_4_197 b_4 NI_4 NS_197 0 5.0339180689199024e-06
GC_4_198 b_4 NI_4 NS_198 0 2.2607987292745665e-06
GC_4_199 b_4 NI_4 NS_199 0 3.8677487007284419e-06
GC_4_200 b_4 NI_4 NS_200 0 2.0110103386488468e-07
GC_4_201 b_4 NI_4 NS_201 0 -8.0831953789018070e-09
GC_4_202 b_4 NI_4 NS_202 0 6.7951732942200894e-10
GC_4_203 b_4 NI_4 NS_203 0 1.5642916247863941e-11
GC_4_204 b_4 NI_4 NS_204 0 -1.2064090575273783e-10
GC_4_205 b_4 NI_4 NS_205 0 -2.1882729742021485e-06
GC_4_206 b_4 NI_4 NS_206 0 2.1734096249892573e-07
GC_4_207 b_4 NI_4 NS_207 0 -2.1912511733562971e-06
GC_4_208 b_4 NI_4 NS_208 0 2.7906294964400894e-06
GC_4_209 b_4 NI_4 NS_209 0 -1.1302628992833111e-06
GC_4_210 b_4 NI_4 NS_210 0 6.5760377685747830e-06
GC_4_211 b_4 NI_4 NS_211 0 -4.1810170942281865e-07
GC_4_212 b_4 NI_4 NS_212 0 2.1387920953709941e-06
GC_4_213 b_4 NI_4 NS_213 0 7.2163592441393801e-06
GC_4_214 b_4 NI_4 NS_214 0 5.1185248820630036e-06
GC_4_215 b_4 NI_4 NS_215 0 1.6097744637809077e-06
GC_4_216 b_4 NI_4 NS_216 0 3.1433799468975925e-06
GC_4_217 b_4 NI_4 NS_217 0 4.8364246709907083e-06
GC_4_218 b_4 NI_4 NS_218 0 1.1505236042177926e-06
GC_4_219 b_4 NI_4 NS_219 0 2.9136141097550729e-06
GC_4_220 b_4 NI_4 NS_220 0 -1.3226685779113845e-06
GC_4_221 b_4 NI_4 NS_221 0 1.2124744748315953e-08
GC_4_222 b_4 NI_4 NS_222 0 -8.1682181925457122e-10
GC_4_223 b_4 NI_4 NS_223 0 -1.6082078493818995e-11
GC_4_224 b_4 NI_4 NS_224 0 1.3082088836440345e-10
GC_4_225 b_4 NI_4 NS_225 0 7.0237137154054835e-08
GC_4_226 b_4 NI_4 NS_226 0 -1.5046100602807478e-08
GC_4_227 b_4 NI_4 NS_227 0 -5.8773516479748986e-07
GC_4_228 b_4 NI_4 NS_228 0 5.5728451311275108e-07
GC_4_229 b_4 NI_4 NS_229 0 1.6792028015234382e-06
GC_4_230 b_4 NI_4 NS_230 0 -4.9983190161395739e-07
GC_4_231 b_4 NI_4 NS_231 0 -9.7806812458105507e-07
GC_4_232 b_4 NI_4 NS_232 0 1.0430328669730802e-07
GC_4_233 b_4 NI_4 NS_233 0 1.6496852836970744e-06
GC_4_234 b_4 NI_4 NS_234 0 -1.1404220659832494e-06
GC_4_235 b_4 NI_4 NS_235 0 -9.0614256642167145e-07
GC_4_236 b_4 NI_4 NS_236 0 -8.6662744441435901e-07
GC_4_237 b_4 NI_4 NS_237 0 -1.1401322789173552e-06
GC_4_238 b_4 NI_4 NS_238 0 -2.4471838474591632e-07
GC_4_239 b_4 NI_4 NS_239 0 8.9532567616223394e-08
GC_4_240 b_4 NI_4 NS_240 0 1.1724103873260396e-06
GD_4_1 b_4 NI_4 NA_1 0 -3.3302476163286280e-03
GD_4_2 b_4 NI_4 NA_2 0 6.7730081992907224e-03
GD_4_3 b_4 NI_4 NA_3 0 5.3317895465105972e-03
GD_4_4 b_4 NI_4 NA_4 0 -9.5852748204678200e-03
GD_4_5 b_4 NI_4 NA_5 0 -5.5836870580439680e-05
GD_4_6 b_4 NI_4 NA_6 0 2.2415266044034365e-05
GD_4_7 b_4 NI_4 NA_7 0 3.5134970198040297e-06
GD_4_8 b_4 NI_4 NA_8 0 1.3447892212093689e-05
GD_4_9 b_4 NI_4 NA_9 0 1.2163792536105277e-05
GD_4_10 b_4 NI_4 NA_10 0 -5.2908253082863328e-06
GD_4_11 b_4 NI_4 NA_11 0 -7.7232130318499107e-06
GD_4_12 b_4 NI_4 NA_12 0 3.3057303322647529e-07
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 -2.7923124691350910e-08
GC_5_2 b_5 NI_5 NS_2 0 1.2536815712132948e-09
GC_5_3 b_5 NI_5 NS_3 0 -9.9739487076124692e-12
GC_5_4 b_5 NI_5 NS_4 0 2.3134321425664088e-11
GC_5_5 b_5 NI_5 NS_5 0 4.4587604533018080e-06
GC_5_6 b_5 NI_5 NS_6 0 2.3149763981336355e-06
GC_5_7 b_5 NI_5 NS_7 0 9.9868190271577679e-06
GC_5_8 b_5 NI_5 NS_8 0 9.7173874857916071e-06
GC_5_9 b_5 NI_5 NS_9 0 1.8696326294226554e-05
GC_5_10 b_5 NI_5 NS_10 0 -2.3425383782450823e-05
GC_5_11 b_5 NI_5 NS_11 0 1.1422717685310508e-05
GC_5_12 b_5 NI_5 NS_12 0 -3.1566160935719605e-06
GC_5_13 b_5 NI_5 NS_13 0 -6.8037250224544765e-06
GC_5_14 b_5 NI_5 NS_14 0 -5.3300295188769093e-05
GC_5_15 b_5 NI_5 NS_15 0 -1.4916969173799026e-05
GC_5_16 b_5 NI_5 NS_16 0 -1.7768778202809616e-05
GC_5_17 b_5 NI_5 NS_17 0 -2.7486795951589168e-05
GC_5_18 b_5 NI_5 NS_18 0 -1.2413931464518155e-05
GC_5_19 b_5 NI_5 NS_19 0 -1.9106839705044043e-05
GC_5_20 b_5 NI_5 NS_20 0 5.8361990204607296e-06
GC_5_21 b_5 NI_5 NS_21 0 1.9598934763184864e-09
GC_5_22 b_5 NI_5 NS_22 0 -2.0086832472399546e-10
GC_5_23 b_5 NI_5 NS_23 0 1.6948014982972321e-11
GC_5_24 b_5 NI_5 NS_24 0 -8.9403656119748818e-11
GC_5_25 b_5 NI_5 NS_25 0 -1.5359113827957648e-06
GC_5_26 b_5 NI_5 NS_26 0 -1.4180233990432019e-06
GC_5_27 b_5 NI_5 NS_27 0 -5.6310781471521074e-06
GC_5_28 b_5 NI_5 NS_28 0 1.3500611931389617e-05
GC_5_29 b_5 NI_5 NS_29 0 3.5171791823724562e-05
GC_5_30 b_5 NI_5 NS_30 0 1.0738188299303173e-05
GC_5_31 b_5 NI_5 NS_31 0 3.2592497296194610e-05
GC_5_32 b_5 NI_5 NS_32 0 -2.6153534597446313e-05
GC_5_33 b_5 NI_5 NS_33 0 -4.0881137715698488e-05
GC_5_34 b_5 NI_5 NS_34 0 -5.0758189867169578e-05
GC_5_35 b_5 NI_5 NS_35 0 -2.0190319739241903e-05
GC_5_36 b_5 NI_5 NS_36 0 9.6138438963685323e-06
GC_5_37 b_5 NI_5 NS_37 0 3.9348242489290908e-06
GC_5_38 b_5 NI_5 NS_38 0 1.2590336015284537e-07
GC_5_39 b_5 NI_5 NS_39 0 -1.3016787634257337e-05
GC_5_40 b_5 NI_5 NS_40 0 -6.9640822807283620e-06
GC_5_41 b_5 NI_5 NS_41 0 -5.4561569564327847e-08
GC_5_42 b_5 NI_5 NS_42 0 -2.0950014170457977e-09
GC_5_43 b_5 NI_5 NS_43 0 -1.0056334028213010e-10
GC_5_44 b_5 NI_5 NS_44 0 3.2108259609170147e-10
GC_5_45 b_5 NI_5 NS_45 0 -1.3498690817229335e-05
GC_5_46 b_5 NI_5 NS_46 0 -1.1750814225702265e-05
GC_5_47 b_5 NI_5 NS_47 0 -4.4779272850936404e-05
GC_5_48 b_5 NI_5 NS_48 0 4.2450788856547733e-05
GC_5_49 b_5 NI_5 NS_49 0 4.9954070089977282e-05
GC_5_50 b_5 NI_5 NS_50 0 -4.4097729568267773e-05
GC_5_51 b_5 NI_5 NS_51 0 -1.0686547194669208e-04
GC_5_52 b_5 NI_5 NS_52 0 6.6401822130587271e-05
GC_5_53 b_5 NI_5 NS_53 0 1.2727304655689204e-04
GC_5_54 b_5 NI_5 NS_54 0 -7.6138310814273877e-06
GC_5_55 b_5 NI_5 NS_55 0 -5.8523238024984612e-05
GC_5_56 b_5 NI_5 NS_56 0 4.1103429217737743e-05
GC_5_57 b_5 NI_5 NS_57 0 4.5420168203443201e-05
GC_5_58 b_5 NI_5 NS_58 0 -5.0333344890631766e-06
GC_5_59 b_5 NI_5 NS_59 0 2.5829952628643368e-05
GC_5_60 b_5 NI_5 NS_60 0 3.8189923382862363e-05
GC_5_61 b_5 NI_5 NS_61 0 6.1704202984796410e-08
GC_5_62 b_5 NI_5 NS_62 0 1.2660808754303996e-09
GC_5_63 b_5 NI_5 NS_63 0 1.6398710151821976e-10
GC_5_64 b_5 NI_5 NS_64 0 -6.8655450263965292e-10
GC_5_65 b_5 NI_5 NS_65 0 -1.0004015465445989e-05
GC_5_66 b_5 NI_5 NS_66 0 -5.4826721762471929e-06
GC_5_67 b_5 NI_5 NS_67 0 1.5174731402820260e-06
GC_5_68 b_5 NI_5 NS_68 0 -1.4462000067996589e-05
GC_5_69 b_5 NI_5 NS_69 0 -1.1184072675492020e-04
GC_5_70 b_5 NI_5 NS_70 0 3.9184477224405538e-05
GC_5_71 b_5 NI_5 NS_71 0 -7.9769107629553979e-05
GC_5_72 b_5 NI_5 NS_72 0 7.8276874305719342e-05
GC_5_73 b_5 NI_5 NS_73 0 1.9275207550530950e-04
GC_5_74 b_5 NI_5 NS_74 0 1.3386993970600984e-04
GC_5_75 b_5 NI_5 NS_75 0 5.7427660373365126e-05
GC_5_76 b_5 NI_5 NS_76 0 -1.9414655481526226e-05
GC_5_77 b_5 NI_5 NS_77 0 -4.7733084209288887e-06
GC_5_78 b_5 NI_5 NS_78 0 -8.4252428590257904e-06
GC_5_79 b_5 NI_5 NS_79 0 3.7519336943135385e-05
GC_5_80 b_5 NI_5 NS_80 0 9.6450131727861820e-06
GC_5_81 b_5 NI_5 NS_81 0 -1.5463093138223280e-05
GC_5_82 b_5 NI_5 NS_82 0 -3.7113235284201742e-06
GC_5_83 b_5 NI_5 NS_83 0 -2.3018576090338935e-08
GC_5_84 b_5 NI_5 NS_84 0 -3.8858820771317450e-07
GC_5_85 b_5 NI_5 NS_85 0 4.5345249190916715e-03
GC_5_86 b_5 NI_5 NS_86 0 3.8285450979865204e-03
GC_5_87 b_5 NI_5 NS_87 0 1.3835635390211187e-02
GC_5_88 b_5 NI_5 NS_88 0 -2.1353740646470533e-02
GC_5_89 b_5 NI_5 NS_89 0 -2.2486096743710830e-02
GC_5_90 b_5 NI_5 NS_90 0 2.6120598454944879e-02
GC_5_91 b_5 NI_5 NS_91 0 3.8309154981649995e-02
GC_5_92 b_5 NI_5 NS_92 0 -3.0087483472848890e-02
GC_5_93 b_5 NI_5 NS_93 0 -4.8554176284704466e-02
GC_5_94 b_5 NI_5 NS_94 0 1.9895869176736150e-02
GC_5_95 b_5 NI_5 NS_95 0 2.6986020389083123e-02
GC_5_96 b_5 NI_5 NS_96 0 -1.5889694902449677e-02
GC_5_97 b_5 NI_5 NS_97 0 -1.4309121714042727e-02
GC_5_98 b_5 NI_5 NS_98 0 6.9209609955556512e-03
GC_5_99 b_5 NI_5 NS_99 0 -4.7570098518152238e-03
GC_5_100 b_5 NI_5 NS_100 0 -1.6677668433030920e-02
GC_5_101 b_5 NI_5 NS_101 0 9.0218498673363110e-05
GC_5_102 b_5 NI_5 NS_102 0 3.5894574595358378e-06
GC_5_103 b_5 NI_5 NS_103 0 5.3419368460603899e-09
GC_5_104 b_5 NI_5 NS_104 0 6.0135185111483185e-07
GC_5_105 b_5 NI_5 NS_105 0 4.7513062286576813e-02
GC_5_106 b_5 NI_5 NS_106 0 -9.6277234691041526e-03
GC_5_107 b_5 NI_5 NS_107 0 -4.5583690652245219e-02
GC_5_108 b_5 NI_5 NS_108 0 2.0520639180749756e-02
GC_5_109 b_5 NI_5 NS_109 0 -5.7692165395681401e-02
GC_5_110 b_5 NI_5 NS_110 0 -6.7344965287313222e-02
GC_5_111 b_5 NI_5 NS_111 0 6.3851924086485393e-02
GC_5_112 b_5 NI_5 NS_112 0 -2.2031911241825644e-02
GC_5_113 b_5 NI_5 NS_113 0 2.8432494601250025e-02
GC_5_114 b_5 NI_5 NS_114 0 8.9369942471789712e-02
GC_5_115 b_5 NI_5 NS_115 0 -5.4359628001037358e-02
GC_5_116 b_5 NI_5 NS_116 0 2.7514733172397093e-03
GC_5_117 b_5 NI_5 NS_117 0 -1.3881473517597189e-02
GC_5_118 b_5 NI_5 NS_118 0 -4.7121694833386497e-02
GC_5_119 b_5 NI_5 NS_119 0 1.6357842588927106e-02
GC_5_120 b_5 NI_5 NS_120 0 -3.9002013699552154e-02
GC_5_121 b_5 NI_5 NS_121 0 -1.0349953958275891e-05
GC_5_122 b_5 NI_5 NS_122 0 -2.1316754009336968e-07
GC_5_123 b_5 NI_5 NS_123 0 -1.2660235834400570e-09
GC_5_124 b_5 NI_5 NS_124 0 -2.5543420737476787e-08
GC_5_125 b_5 NI_5 NS_125 0 -4.2480397462394803e-03
GC_5_126 b_5 NI_5 NS_126 0 -3.4907699650810410e-03
GC_5_127 b_5 NI_5 NS_127 0 -1.2926398897791642e-02
GC_5_128 b_5 NI_5 NS_128 0 1.7064707780997578e-02
GC_5_129 b_5 NI_5 NS_129 0 1.7381905686225656e-02
GC_5_130 b_5 NI_5 NS_130 0 -1.9436891295307211e-02
GC_5_131 b_5 NI_5 NS_131 0 -3.3160398510843646e-02
GC_5_132 b_5 NI_5 NS_132 0 2.5454388828446247e-02
GC_5_133 b_5 NI_5 NS_133 0 4.0799770165464516e-02
GC_5_134 b_5 NI_5 NS_134 0 -1.1454429797341452e-02
GC_5_135 b_5 NI_5 NS_135 0 -2.1063045481597327e-02
GC_5_136 b_5 NI_5 NS_136 0 1.5303540864951387e-02
GC_5_137 b_5 NI_5 NS_137 0 1.4115522372272005e-02
GC_5_138 b_5 NI_5 NS_138 0 -3.7637543500676045e-03
GC_5_139 b_5 NI_5 NS_139 0 7.0728043525807938e-03
GC_5_140 b_5 NI_5 NS_140 0 1.3571593783590505e-02
GC_5_141 b_5 NI_5 NS_141 0 -1.8513493899295285e-06
GC_5_142 b_5 NI_5 NS_142 0 2.5575445312156877e-07
GC_5_143 b_5 NI_5 NS_143 0 1.6675703226009014e-09
GC_5_144 b_5 NI_5 NS_144 0 1.3815226234037955e-08
GC_5_145 b_5 NI_5 NS_145 0 1.1369543036640721e-03
GC_5_146 b_5 NI_5 NS_146 0 -2.1664743213213279e-03
GC_5_147 b_5 NI_5 NS_147 0 3.4943906453732310e-03
GC_5_148 b_5 NI_5 NS_148 0 -1.2990553284985176e-02
GC_5_149 b_5 NI_5 NS_149 0 -3.9378869909784474e-02
GC_5_150 b_5 NI_5 NS_150 0 -3.6054851395279669e-04
GC_5_151 b_5 NI_5 NS_151 0 -2.6238831230157907e-02
GC_5_152 b_5 NI_5 NS_152 0 2.8978927054347653e-02
GC_5_153 b_5 NI_5 NS_153 0 5.2196790950131008e-02
GC_5_154 b_5 NI_5 NS_154 0 3.8196066069323777e-02
GC_5_155 b_5 NI_5 NS_155 0 1.7566178593046489e-02
GC_5_156 b_5 NI_5 NS_156 0 -1.4392572455005484e-02
GC_5_157 b_5 NI_5 NS_157 0 -9.1635687513091282e-03
GC_5_158 b_5 NI_5 NS_158 0 -3.7446291391962723e-03
GC_5_159 b_5 NI_5 NS_159 0 8.0613894069748015e-03
GC_5_160 b_5 NI_5 NS_160 0 5.8589432140919440e-03
GC_5_161 b_5 NI_5 NS_161 0 -2.7807364352481097e-08
GC_5_162 b_5 NI_5 NS_162 0 8.0981225233898658e-10
GC_5_163 b_5 NI_5 NS_163 0 -1.5187365283490889e-11
GC_5_164 b_5 NI_5 NS_164 0 7.2084391797050138e-11
GC_5_165 b_5 NI_5 NS_165 0 4.1642275850109524e-06
GC_5_166 b_5 NI_5 NS_166 0 2.5912863085221852e-06
GC_5_167 b_5 NI_5 NS_167 0 9.5706833326626421e-06
GC_5_168 b_5 NI_5 NS_168 0 1.0122654107189798e-05
GC_5_169 b_5 NI_5 NS_169 0 1.9377846290706080e-05
GC_5_170 b_5 NI_5 NS_170 0 -2.2684105905676801e-05
GC_5_171 b_5 NI_5 NS_171 0 1.1294700522921069e-05
GC_5_172 b_5 NI_5 NS_172 0 -2.9403257986622225e-06
GC_5_173 b_5 NI_5 NS_173 0 -5.4388631518847627e-06
GC_5_174 b_5 NI_5 NS_174 0 -5.2854993937379103e-05
GC_5_175 b_5 NI_5 NS_175 0 -1.4373071972407834e-05
GC_5_176 b_5 NI_5 NS_176 0 -1.8172894657484738e-05
GC_5_177 b_5 NI_5 NS_177 0 -2.7456964330486272e-05
GC_5_178 b_5 NI_5 NS_178 0 -1.3076036408659439e-05
GC_5_179 b_5 NI_5 NS_179 0 -1.9571260205948100e-05
GC_5_180 b_5 NI_5 NS_180 0 5.5880008509162627e-06
GC_5_181 b_5 NI_5 NS_181 0 7.1854199516570721e-09
GC_5_182 b_5 NI_5 NS_182 0 2.2463982532401806e-11
GC_5_183 b_5 NI_5 NS_183 0 2.0136528402966687e-11
GC_5_184 b_5 NI_5 NS_184 0 -1.2273056645649860e-10
GC_5_185 b_5 NI_5 NS_185 0 -2.1095037643416079e-06
GC_5_186 b_5 NI_5 NS_186 0 -1.2999236650784924e-06
GC_5_187 b_5 NI_5 NS_187 0 -6.2931078936699155e-06
GC_5_188 b_5 NI_5 NS_188 0 1.3497473245167949e-05
GC_5_189 b_5 NI_5 NS_189 0 3.4249418972078463e-05
GC_5_190 b_5 NI_5 NS_190 0 1.2262045703420404e-05
GC_5_191 b_5 NI_5 NS_191 0 3.1603969976309555e-05
GC_5_192 b_5 NI_5 NS_192 0 -2.5423271129533440e-05
GC_5_193 b_5 NI_5 NS_193 0 -3.9478418815785943e-05
GC_5_194 b_5 NI_5 NS_194 0 -4.7737604930462616e-05
GC_5_195 b_5 NI_5 NS_195 0 -1.9905276024478461e-05
GC_5_196 b_5 NI_5 NS_196 0 1.1122842176561719e-05
GC_5_197 b_5 NI_5 NS_197 0 5.8928629382809743e-06
GC_5_198 b_5 NI_5 NS_198 0 1.6678091834620214e-06
GC_5_199 b_5 NI_5 NS_199 0 -1.0738280350499075e-05
GC_5_200 b_5 NI_5 NS_200 0 -6.7127708104186512e-06
GC_5_201 b_5 NI_5 NS_201 0 2.0778195936989297e-08
GC_5_202 b_5 NI_5 NS_202 0 -1.0272255302554099e-09
GC_5_203 b_5 NI_5 NS_203 0 -1.9428689757195630e-11
GC_5_204 b_5 NI_5 NS_204 0 1.5753099575968302e-10
GC_5_205 b_5 NI_5 NS_205 0 -1.1217624880046448e-06
GC_5_206 b_5 NI_5 NS_206 0 -8.0925816984924033e-07
GC_5_207 b_5 NI_5 NS_207 0 -2.0036364579880455e-06
GC_5_208 b_5 NI_5 NS_208 0 3.6547330537952460e-08
GC_5_209 b_5 NI_5 NS_209 0 -3.0739377035217024e-06
GC_5_210 b_5 NI_5 NS_210 0 8.6266627408548295e-07
GC_5_211 b_5 NI_5 NS_211 0 -4.1492024228943606e-06
GC_5_212 b_5 NI_5 NS_212 0 4.3129834150431052e-06
GC_5_213 b_5 NI_5 NS_213 0 3.3149237246716839e-06
GC_5_214 b_5 NI_5 NS_214 0 5.4267708388420411e-06
GC_5_215 b_5 NI_5 NS_215 0 -8.9973918604331059e-07
GC_5_216 b_5 NI_5 NS_216 0 5.9728357018210710e-06
GC_5_217 b_5 NI_5 NS_217 0 6.0574025209169526e-06
GC_5_218 b_5 NI_5 NS_218 0 3.3263249260727735e-06
GC_5_219 b_5 NI_5 NS_219 0 5.8642833348653532e-06
GC_5_220 b_5 NI_5 NS_220 0 1.7030941970030566e-06
GC_5_221 b_5 NI_5 NS_221 0 -2.4099530210314082e-08
GC_5_222 b_5 NI_5 NS_222 0 1.2312870981145740e-09
GC_5_223 b_5 NI_5 NS_223 0 2.1599265978424943e-11
GC_5_224 b_5 NI_5 NS_224 0 -1.7722969548801152e-10
GC_5_225 b_5 NI_5 NS_225 0 1.8333073269437817e-06
GC_5_226 b_5 NI_5 NS_226 0 -4.1855575088977378e-06
GC_5_227 b_5 NI_5 NS_227 0 2.4443899379798524e-06
GC_5_228 b_5 NI_5 NS_228 0 7.5715587036162879e-08
GC_5_229 b_5 NI_5 NS_229 0 -1.6176202535224682e-06
GC_5_230 b_5 NI_5 NS_230 0 -4.3834845702583308e-06
GC_5_231 b_5 NI_5 NS_231 0 1.0020626084563424e-06
GC_5_232 b_5 NI_5 NS_232 0 -7.2532092352636712e-06
GC_5_233 b_5 NI_5 NS_233 0 -8.7087205385327074e-06
GC_5_234 b_5 NI_5 NS_234 0 -4.7028288919249329e-06
GC_5_235 b_5 NI_5 NS_235 0 -3.2786364418600656e-06
GC_5_236 b_5 NI_5 NS_236 0 1.3949522064841812e-06
GC_5_237 b_5 NI_5 NS_237 0 -1.9194178681185603e-06
GC_5_238 b_5 NI_5 NS_238 0 -5.4219324937889567e-07
GC_5_239 b_5 NI_5 NS_239 0 -3.2888266602591204e-06
GC_5_240 b_5 NI_5 NS_240 0 -1.5163216469431046e-06
GD_5_1 b_5 NI_5 NA_1 0 1.4811101677325513e-05
GD_5_2 b_5 NI_5 NA_2 0 4.8447116803312470e-06
GD_5_3 b_5 NI_5 NA_3 0 2.2415266046305738e-05
GD_5_4 b_5 NI_5 NA_4 0 -5.5822644692711185e-05
GD_5_5 b_5 NI_5 NA_5 0 -9.6518867068792636e-03
GD_5_6 b_5 NI_5 NA_6 0 5.5541233396464319e-03
GD_5_7 b_5 NI_5 NA_7 0 6.7712145109744713e-03
GD_5_8 b_5 NI_5 NA_8 0 -3.3437475323618415e-03
GD_5_9 b_5 NI_5 NA_9 0 1.3910657017617279e-05
GD_5_10 b_5 NI_5 NA_10 0 3.0880584766365765e-06
GD_5_11 b_5 NI_5 NA_11 0 -1.1680798973691237e-06
GD_5_12 b_5 NI_5 NA_12 0 1.0083329928954350e-05
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 1.9604827830782515e-09
GC_6_2 b_6 NI_6 NS_2 0 -2.0091514800021308e-10
GC_6_3 b_6 NI_6 NS_3 0 1.6947532319169950e-11
GC_6_4 b_6 NI_6 NS_4 0 -8.9399793521601689e-11
GC_6_5 b_6 NI_6 NS_5 0 -1.5357422933152633e-06
GC_6_6 b_6 NI_6 NS_6 0 -1.4180437166354096e-06
GC_6_7 b_6 NI_6 NS_7 0 -5.6306077416537357e-06
GC_6_8 b_6 NI_6 NS_8 0 1.3500657911951440e-05
GC_6_9 b_6 NI_6 NS_9 0 3.5171687454704517e-05
GC_6_10 b_6 NI_6 NS_10 0 1.0737047101803751e-05
GC_6_11 b_6 NI_6 NS_11 0 3.2592131254318384e-05
GC_6_12 b_6 NI_6 NS_12 0 -2.6154287337496831e-05
GC_6_13 b_6 NI_6 NS_13 0 -4.0882398560458643e-05
GC_6_14 b_6 NI_6 NS_14 0 -5.0757257704051900e-05
GC_6_15 b_6 NI_6 NS_15 0 -2.0190237823403160e-05
GC_6_16 b_6 NI_6 NS_16 0 9.6142438172427980e-06
GC_6_17 b_6 NI_6 NS_17 0 3.9350704921754933e-06
GC_6_18 b_6 NI_6 NS_18 0 1.2601171458113056e-07
GC_6_19 b_6 NI_6 NS_19 0 -1.3016677802276930e-05
GC_6_20 b_6 NI_6 NS_20 0 -6.9640875839880075e-06
GC_6_21 b_6 NI_6 NS_21 0 -2.8092440361794687e-08
GC_6_22 b_6 NI_6 NS_22 0 1.2625336458669506e-09
GC_6_23 b_6 NI_6 NS_23 0 -9.9117772157191163e-12
GC_6_24 b_6 NI_6 NS_24 0 2.2550619963543961e-11
GC_6_25 b_6 NI_6 NS_25 0 4.4972689470959310e-06
GC_6_26 b_6 NI_6 NS_26 0 2.2387586862493406e-06
GC_6_27 b_6 NI_6 NS_27 0 9.9893573699537052e-06
GC_6_28 b_6 NI_6 NS_28 0 9.6249760574098784e-06
GC_6_29 b_6 NI_6 NS_29 0 1.8703103456593553e-05
GC_6_30 b_6 NI_6 NS_30 0 -2.3516915830969245e-05
GC_6_31 b_6 NI_6 NS_31 0 1.1345871762316627e-05
GC_6_32 b_6 NI_6 NS_32 0 -3.3422993870302998e-06
GC_6_33 b_6 NI_6 NS_33 0 -6.9544968558510616e-06
GC_6_34 b_6 NI_6 NS_34 0 -5.3248456117640947e-05
GC_6_35 b_6 NI_6 NS_35 0 -1.4962316214552076e-05
GC_6_36 b_6 NI_6 NS_36 0 -1.7861800609159752e-05
GC_6_37 b_6 NI_6 NS_37 0 -2.7583405459367039e-05
GC_6_38 b_6 NI_6 NS_38 0 -1.2422759868052168e-05
GC_6_39 b_6 NI_6 NS_39 0 -1.9191335674622318e-05
GC_6_40 b_6 NI_6 NS_40 0 5.8309121307191929e-06
GC_6_41 b_6 NI_6 NS_41 0 6.1677766459094732e-08
GC_6_42 b_6 NI_6 NS_42 0 1.2669495478499282e-09
GC_6_43 b_6 NI_6 NS_43 0 1.6399362489482193e-10
GC_6_44 b_6 NI_6 NS_44 0 -6.8660944025229873e-10
GC_6_45 b_6 NI_6 NS_45 0 -1.0021558735457105e-05
GC_6_46 b_6 NI_6 NS_46 0 -5.4883440367866527e-06
GC_6_47 b_6 NI_6 NS_47 0 1.4900690210184307e-06
GC_6_48 b_6 NI_6 NS_48 0 -1.4479541704894820e-05
GC_6_49 b_6 NI_6 NS_49 0 -1.1185421245698944e-04
GC_6_50 b_6 NI_6 NS_50 0 3.9288819923528026e-05
GC_6_51 b_6 NI_6 NS_51 0 -7.9728855551602850e-05
GC_6_52 b_6 NI_6 NS_52 0 7.8341208257694904e-05
GC_6_53 b_6 NI_6 NS_53 0 1.9284808673156843e-04
GC_6_54 b_6 NI_6 NS_54 0 1.3377504115888111e-04
GC_6_55 b_6 NI_6 NS_55 0 5.7410793278272214e-05
GC_6_56 b_6 NI_6 NS_56 0 -1.9453200790137479e-05
GC_6_57 b_6 NI_6 NS_57 0 -4.8009473033744608e-06
GC_6_58 b_6 NI_6 NS_58 0 -8.4210387803408596e-06
GC_6_59 b_6 NI_6 NS_59 0 3.7514589085846781e-05
GC_6_60 b_6 NI_6 NS_60 0 9.6476628665192894e-06
GC_6_61 b_6 NI_6 NS_61 0 -5.4549211238926692e-08
GC_6_62 b_6 NI_6 NS_62 0 -2.0955088690325817e-09
GC_6_63 b_6 NI_6 NS_63 0 -1.0056422443866788e-10
GC_6_64 b_6 NI_6 NS_64 0 3.2111225146416855e-10
GC_6_65 b_6 NI_6 NS_65 0 -1.3498608767791119e-05
GC_6_66 b_6 NI_6 NS_66 0 -1.1749813932926006e-05
GC_6_67 b_6 NI_6 NS_67 0 -4.4778893550487295e-05
GC_6_68 b_6 NI_6 NS_68 0 4.2451447230670165e-05
GC_6_69 b_6 NI_6 NS_69 0 4.9954079253378359e-05
GC_6_70 b_6 NI_6 NS_70 0 -4.4097075684274855e-05
GC_6_71 b_6 NI_6 NS_71 0 -1.0686413593653601e-04
GC_6_72 b_6 NI_6 NS_72 0 6.6403484170360631e-05
GC_6_73 b_6 NI_6 NS_73 0 1.2727377659504002e-04
GC_6_74 b_6 NI_6 NS_74 0 -7.6158837192898895e-06
GC_6_75 b_6 NI_6 NS_75 0 -5.8523906708703590e-05
GC_6_76 b_6 NI_6 NS_76 0 4.1104293931107492e-05
GC_6_77 b_6 NI_6 NS_77 0 4.5420873863384692e-05
GC_6_78 b_6 NI_6 NS_78 0 -5.0322592430726497e-06
GC_6_79 b_6 NI_6 NS_79 0 2.5831324603454427e-05
GC_6_80 b_6 NI_6 NS_80 0 3.8190405578631550e-05
GC_6_81 b_6 NI_6 NS_81 0 9.0218499688407347e-05
GC_6_82 b_6 NI_6 NS_82 0 3.5894574033663602e-06
GC_6_83 b_6 NI_6 NS_83 0 5.3419361839614819e-09
GC_6_84 b_6 NI_6 NS_84 0 6.0135185639577056e-07
GC_6_85 b_6 NI_6 NS_85 0 4.7513062011700448e-02
GC_6_86 b_6 NI_6 NS_86 0 -9.6277234593040613e-03
GC_6_87 b_6 NI_6 NS_87 0 -4.5583691085500568e-02
GC_6_88 b_6 NI_6 NS_88 0 2.0520639159310738e-02
GC_6_89 b_6 NI_6 NS_89 0 -5.7692165766263639e-02
GC_6_90 b_6 NI_6 NS_90 0 -6.7344964383529077e-02
GC_6_91 b_6 NI_6 NS_91 0 6.3851923941562333e-02
GC_6_92 b_6 NI_6 NS_92 0 -2.2031910559920331e-02
GC_6_93 b_6 NI_6 NS_93 0 2.8432495618086751e-02
GC_6_94 b_6 NI_6 NS_94 0 8.9369943252157358e-02
GC_6_95 b_6 NI_6 NS_95 0 -5.4359627623583401e-02
GC_6_96 b_6 NI_6 NS_96 0 2.7514735995811880e-03
GC_6_97 b_6 NI_6 NS_97 0 -1.3881472979163034e-02
GC_6_98 b_6 NI_6 NS_98 0 -4.7121694776249737e-02
GC_6_99 b_6 NI_6 NS_99 0 1.6357842969523112e-02
GC_6_100 b_6 NI_6 NS_100 0 -3.9002013745733449e-02
GC_6_101 b_6 NI_6 NS_101 0 -1.5463093138225740e-05
GC_6_102 b_6 NI_6 NS_102 0 -3.7113235284196241e-06
GC_6_103 b_6 NI_6 NS_103 0 -2.3018576090332437e-08
GC_6_104 b_6 NI_6 NS_104 0 -3.8858820771322548e-07
GC_6_105 b_6 NI_6 NS_105 0 4.5345249190916585e-03
GC_6_106 b_6 NI_6 NS_106 0 3.8285450979865161e-03
GC_6_107 b_6 NI_6 NS_107 0 1.3835635390211164e-02
GC_6_108 b_6 NI_6 NS_108 0 -2.1353740646470554e-02
GC_6_109 b_6 NI_6 NS_109 0 -2.2486096743710875e-02
GC_6_110 b_6 NI_6 NS_110 0 2.6120598454944924e-02
GC_6_111 b_6 NI_6 NS_111 0 3.8309154981649968e-02
GC_6_112 b_6 NI_6 NS_112 0 -3.0087483472848838e-02
GC_6_113 b_6 NI_6 NS_113 0 -4.8554176284704383e-02
GC_6_114 b_6 NI_6 NS_114 0 1.9895869176736209e-02
GC_6_115 b_6 NI_6 NS_115 0 2.6986020389083137e-02
GC_6_116 b_6 NI_6 NS_116 0 -1.5889694902449663e-02
GC_6_117 b_6 NI_6 NS_117 0 -1.4309121714042691e-02
GC_6_118 b_6 NI_6 NS_118 0 6.9209609955556591e-03
GC_6_119 b_6 NI_6 NS_119 0 -4.7570098518151978e-03
GC_6_120 b_6 NI_6 NS_120 0 -1.6677668433030916e-02
GC_6_121 b_6 NI_6 NS_121 0 -1.8513499671640072e-06
GC_6_122 b_6 NI_6 NS_122 0 2.5575447761234043e-07
GC_6_123 b_6 NI_6 NS_123 0 1.6675703955056872e-09
GC_6_124 b_6 NI_6 NS_124 0 1.3815225133691497e-08
GC_6_125 b_6 NI_6 NS_125 0 1.1369543523702614e-03
GC_6_126 b_6 NI_6 NS_126 0 -2.1664743002109054e-03
GC_6_127 b_6 NI_6 NS_127 0 3.4943906894775627e-03
GC_6_128 b_6 NI_6 NS_128 0 -1.2990553244954826e-02
GC_6_129 b_6 NI_6 NS_129 0 -3.9378869866403161e-02
GC_6_130 b_6 NI_6 NS_130 0 -3.6054868580326886e-04
GC_6_131 b_6 NI_6 NS_131 0 -2.6238831259690898e-02
GC_6_132 b_6 NI_6 NS_132 0 2.8978926982025113e-02
GC_6_133 b_6 NI_6 NS_133 0 5.2196790921335993e-02
GC_6_134 b_6 NI_6 NS_134 0 3.8196066152359855e-02
GC_6_135 b_6 NI_6 NS_135 0 1.7566178694236975e-02
GC_6_136 b_6 NI_6 NS_136 0 -1.4392572524268841e-02
GC_6_137 b_6 NI_6 NS_137 0 -9.1635688226028873e-03
GC_6_138 b_6 NI_6 NS_138 0 -3.7446293230960583e-03
GC_6_139 b_6 NI_6 NS_139 0 8.0613892485741391e-03
GC_6_140 b_6 NI_6 NS_140 0 5.8589431802656723e-03
GC_6_141 b_6 NI_6 NS_141 0 -1.0349953947742934e-05
GC_6_142 b_6 NI_6 NS_142 0 -2.1316754054524233e-07
GC_6_143 b_6 NI_6 NS_143 0 -1.2660235847175938e-09
GC_6_144 b_6 NI_6 NS_144 0 -2.5543420716095991e-08
GC_6_145 b_6 NI_6 NS_145 0 -4.2480397441673617e-03
GC_6_146 b_6 NI_6 NS_146 0 -3.4907699661083235e-03
GC_6_147 b_6 NI_6 NS_147 0 -1.2926398894721185e-02
GC_6_148 b_6 NI_6 NS_148 0 1.7064707778669249e-02
GC_6_149 b_6 NI_6 NS_149 0 1.7381905682377952e-02
GC_6_150 b_6 NI_6 NS_150 0 -1.9436891301835096e-02
GC_6_151 b_6 NI_6 NS_151 0 -3.3160398514071744e-02
GC_6_152 b_6 NI_6 NS_152 0 2.5454388825887866e-02
GC_6_153 b_6 NI_6 NS_153 0 4.0799770158819450e-02
GC_6_154 b_6 NI_6 NS_154 0 -1.1454429793721573e-02
GC_6_155 b_6 NI_6 NS_155 0 -2.1063045483320952e-02
GC_6_156 b_6 NI_6 NS_156 0 1.5303540867818198e-02
GC_6_157 b_6 NI_6 NS_157 0 1.4115522373870227e-02
GC_6_158 b_6 NI_6 NS_158 0 -3.7637543469367083e-03
GC_6_159 b_6 NI_6 NS_159 0 7.0728043549368085e-03
GC_6_160 b_6 NI_6 NS_160 0 1.3571593784218749e-02
GC_6_161 b_6 NI_6 NS_161 0 7.1854881813297068e-09
GC_6_162 b_6 NI_6 NS_162 0 2.2479995654004664e-11
GC_6_163 b_6 NI_6 NS_163 0 2.0136715087475737e-11
GC_6_164 b_6 NI_6 NS_164 0 -1.2273214753647510e-10
GC_6_165 b_6 NI_6 NS_165 0 -2.1096709923798715e-06
GC_6_166 b_6 NI_6 NS_166 0 -1.2998928360082714e-06
GC_6_167 b_6 NI_6 NS_167 0 -6.2934656757459617e-06
GC_6_168 b_6 NI_6 NS_168 0 1.3497434132054178e-05
GC_6_169 b_6 NI_6 NS_169 0 3.4249374886744684e-05
GC_6_170 b_6 NI_6 NS_170 0 1.2262958998267503e-05
GC_6_171 b_6 NI_6 NS_171 0 3.1604141179292504e-05
GC_6_172 b_6 NI_6 NS_172 0 -2.5422645117072160e-05
GC_6_173 b_6 NI_6 NS_173 0 -3.9477361308842852e-05
GC_6_174 b_6 NI_6 NS_174 0 -4.7737993528208787e-05
GC_6_175 b_6 NI_6 NS_175 0 -1.9905263437515359e-05
GC_6_176 b_6 NI_6 NS_176 0 1.1122633918341686e-05
GC_6_177 b_6 NI_6 NS_177 0 5.8928106945511438e-06
GC_6_178 b_6 NI_6 NS_178 0 1.6678145791323972e-06
GC_6_179 b_6 NI_6 NS_179 0 -1.0738206877000946e-05
GC_6_180 b_6 NI_6 NS_180 0 -6.7127512475465279e-06
GC_6_181 b_6 NI_6 NS_181 0 -2.7643468422334792e-08
GC_6_182 b_6 NI_6 NS_182 0 8.0098526232942438e-10
GC_6_183 b_6 NI_6 NS_183 0 -1.5252017746931417e-11
GC_6_184 b_6 NI_6 NS_184 0 7.2677014517694059e-11
GC_6_185 b_6 NI_6 NS_185 0 4.1256396025753677e-06
GC_6_186 b_6 NI_6 NS_186 0 2.6677180412753289e-06
GC_6_187 b_6 NI_6 NS_187 0 9.5682087516342433e-06
GC_6_188 b_6 NI_6 NS_188 0 1.0216481061170554e-05
GC_6_189 b_6 NI_6 NS_189 0 1.9376033425933281e-05
GC_6_190 b_6 NI_6 NS_190 0 -2.2593580530887805e-05
GC_6_191 b_6 NI_6 NS_191 0 1.1373791657047345e-05
GC_6_192 b_6 NI_6 NS_192 0 -2.7583655380216521e-06
GC_6_193 b_6 NI_6 NS_193 0 -5.2913335843761499e-06
GC_6_194 b_6 NI_6 NS_194 0 -5.2911831798658552e-05
GC_6_195 b_6 NI_6 NS_195 0 -1.4329145239331920e-05
GC_6_196 b_6 NI_6 NS_196 0 -1.8082861952609308e-05
GC_6_197 b_6 NI_6 NS_197 0 -2.7364161700548423e-05
GC_6_198 b_6 NI_6 NS_198 0 -1.3068178053941816e-05
GC_6_199 b_6 NI_6 NS_199 0 -1.9489167007288623e-05
GC_6_200 b_6 NI_6 NS_200 0 5.5936316671906848e-06
GC_6_201 b_6 NI_6 NS_201 0 -2.4072623166394023e-08
GC_6_202 b_6 NI_6 NS_202 0 1.2303582292995059e-09
GC_6_203 b_6 NI_6 NS_203 0 2.1589039811450104e-11
GC_6_204 b_6 NI_6 NS_204 0 -1.7715315527549914e-10
GC_6_205 b_6 NI_6 NS_205 0 1.8511908287664064e-06
GC_6_206 b_6 NI_6 NS_206 0 -4.1799796137779077e-06
GC_6_207 b_6 NI_6 NS_207 0 2.4721017975487148e-06
GC_6_208 b_6 NI_6 NS_208 0 9.2956239740711766e-08
GC_6_209 b_6 NI_6 NS_209 0 -1.6039211287656701e-06
GC_6_210 b_6 NI_6 NS_210 0 -4.4881546093933058e-06
GC_6_211 b_6 NI_6 NS_211 0 9.6225859519559063e-07
GC_6_212 b_6 NI_6 NS_212 0 -7.3177751128954375e-06
GC_6_213 b_6 NI_6 NS_213 0 -8.8052555665384768e-06
GC_6_214 b_6 NI_6 NS_214 0 -4.6098776432908940e-06
GC_6_215 b_6 NI_6 NS_215 0 -3.2625429725014267e-06
GC_6_216 b_6 NI_6 NS_216 0 1.4328971487351356e-06
GC_6_217 b_6 NI_6 NS_217 0 -1.8926888690737559e-06
GC_6_218 b_6 NI_6 NS_218 0 -5.4632541315331183e-07
GC_6_219 b_6 NI_6 NS_219 0 -3.2845052668505904e-06
GC_6_220 b_6 NI_6 NS_220 0 -1.5188068225328758e-06
GC_6_221 b_6 NI_6 NS_221 0 2.0768895948580851e-08
GC_6_222 b_6 NI_6 NS_222 0 -1.0266108896198756e-09
GC_6_223 b_6 NI_6 NS_223 0 -1.9426118057760797e-11
GC_6_224 b_6 NI_6 NS_224 0 1.5749233684995178e-10
GC_6_225 b_6 NI_6 NS_225 0 -1.1217130528244135e-06
GC_6_226 b_6 NI_6 NS_226 0 -8.1021153889261965e-07
GC_6_227 b_6 NI_6 NS_227 0 -2.0037374167279018e-06
GC_6_228 b_6 NI_6 NS_228 0 3.5848983956333890e-08
GC_6_229 b_6 NI_6 NS_229 0 -3.0743117932636520e-06
GC_6_230 b_6 NI_6 NS_230 0 8.6171738066585947e-07
GC_6_231 b_6 NI_6 NS_231 0 -4.1502959904431947e-06
GC_6_232 b_6 NI_6 NS_232 0 4.3114704609334525e-06
GC_6_233 b_6 NI_6 NS_233 0 3.3134004765228827e-06
GC_6_234 b_6 NI_6 NS_234 0 5.4284203752211894e-06
GC_6_235 b_6 NI_6 NS_235 0 -8.9968142481886455e-07
GC_6_236 b_6 NI_6 NS_236 0 5.9726067064414733e-06
GC_6_237 b_6 NI_6 NS_237 0 6.0570612608695188e-06
GC_6_238 b_6 NI_6 NS_238 0 3.3263267320167050e-06
GC_6_239 b_6 NI_6 NS_239 0 5.8639217402273652e-06
GC_6_240 b_6 NI_6 NS_240 0 1.7029363024306995e-06
GD_6_1 b_6 NI_6 NA_1 0 4.8451604984338582e-06
GD_6_2 b_6 NI_6 NA_2 0 1.5200615813122763e-05
GD_6_3 b_6 NI_6 NA_3 0 -5.5836872143735613e-05
GD_6_4 b_6 NI_6 NA_4 0 2.2411103753543215e-05
GD_6_5 b_6 NI_6 NA_5 0 5.5541226909173414e-03
GD_6_6 b_6 NI_6 NA_6 0 -9.6518867068792896e-03
GD_6_7 b_6 NI_6 NA_7 0 -3.3437475291103330e-03
GD_6_8 b_6 NI_6 NA_8 0 6.7712145152012118e-03
GD_6_9 b_6 NI_6 NA_9 0 3.0875897660319961e-06
GD_6_10 b_6 NI_6 NA_10 0 1.3524373889132782e-05
GD_6_11 b_6 NI_6 NA_11 0 1.0098377215587846e-05
GD_6_12 b_6 NI_6 NA_12 0 -1.1644152985624877e-06
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 2.0308402598486642e-08
GC_7_2 b_7 NI_7 NS_2 0 -1.0039750939935007e-09
GC_7_3 b_7 NI_7 NS_3 0 -1.9110575435930744e-11
GC_7_4 b_7 NI_7 NS_4 0 1.5484024294356069e-10
GC_7_5 b_7 NI_7 NS_5 0 -1.0722359773115095e-06
GC_7_6 b_7 NI_7 NS_6 0 -8.5235517903430253e-07
GC_7_7 b_7 NI_7 NS_7 0 -1.9506687511606466e-06
GC_7_8 b_7 NI_7 NS_8 0 -1.2482950387529962e-08
GC_7_9 b_7 NI_7 NS_9 0 -3.0919927235436234e-06
GC_7_10 b_7 NI_7 NS_10 0 7.4445433475246381e-07
GC_7_11 b_7 NI_7 NS_11 0 -4.1324093293388241e-06
GC_7_12 b_7 NI_7 NS_12 0 4.2217630317936244e-06
GC_7_13 b_7 NI_7 NS_13 0 3.1598678701574386e-06
GC_7_14 b_7 NI_7 NS_14 0 5.3390136116707116e-06
GC_7_15 b_7 NI_7 NS_15 0 -9.0731354704219589e-07
GC_7_16 b_7 NI_7 NS_16 0 5.9324207974835424e-06
GC_7_17 b_7 NI_7 NS_17 0 5.9750963306107842e-06
GC_7_18 b_7 NI_7 NS_18 0 3.2313788606390890e-06
GC_7_19 b_7 NI_7 NS_19 0 5.7328774923184436e-06
GC_7_20 b_7 NI_7 NS_20 0 1.6826698841534174e-06
GC_7_21 b_7 NI_7 NS_21 0 -2.3936347149078703e-08
GC_7_22 b_7 NI_7 NS_22 0 1.2234639228557475e-09
GC_7_23 b_7 NI_7 NS_23 0 2.1495912135450298e-11
GC_7_24 b_7 NI_7 NS_24 0 -1.7598159666021412e-10
GC_7_25 b_7 NI_7 NS_25 0 1.8751008390970340e-06
GC_7_26 b_7 NI_7 NS_26 0 -4.2198207235496843e-06
GC_7_27 b_7 NI_7 NS_27 0 2.4962612760178384e-06
GC_7_28 b_7 NI_7 NS_28 0 3.3570514187435951e-08
GC_7_29 b_7 NI_7 NS_29 0 -1.6539763328507257e-06
GC_7_30 b_7 NI_7 NS_30 0 -4.5468564695944350e-06
GC_7_31 b_7 NI_7 NS_31 0 9.6538948992990325e-07
GC_7_32 b_7 NI_7 NS_32 0 -7.3307021692487106e-06
GC_7_33 b_7 NI_7 NS_33 0 -8.9355038128141216e-06
GC_7_34 b_7 NI_7 NS_34 0 -4.6687543392506300e-06
GC_7_35 b_7 NI_7 NS_35 0 -3.3134581965229515e-06
GC_7_36 b_7 NI_7 NS_36 0 1.4348148238389367e-06
GC_7_37 b_7 NI_7 NS_37 0 -1.9277169841723072e-06
GC_7_38 b_7 NI_7 NS_38 0 -4.7310350609293157e-07
GC_7_39 b_7 NI_7 NS_39 0 -3.2465969303585123e-06
GC_7_40 b_7 NI_7 NS_40 0 -1.4929323717757760e-06
GC_7_41 b_7 NI_7 NS_41 0 -2.9031620960743867e-08
GC_7_42 b_7 NI_7 NS_42 0 8.7636027093703715e-10
GC_7_43 b_7 NI_7 NS_43 0 -1.4816280151215723e-11
GC_7_44 b_7 NI_7 NS_44 0 6.7054246600502079e-11
GC_7_45 b_7 NI_7 NS_45 0 4.0592950908727557e-06
GC_7_46 b_7 NI_7 NS_46 0 2.6907844646426563e-06
GC_7_47 b_7 NI_7 NS_47 0 9.4653610952736620e-06
GC_7_48 b_7 NI_7 NS_48 0 1.0215857407310115e-05
GC_7_49 b_7 NI_7 NS_49 0 1.9372833128320083e-05
GC_7_50 b_7 NI_7 NS_50 0 -2.2384281389530957e-05
GC_7_51 b_7 NI_7 NS_51 0 1.1343539513129804e-05
GC_7_52 b_7 NI_7 NS_52 0 -2.6952226034522639e-06
GC_7_53 b_7 NI_7 NS_53 0 -5.1382556721611020e-06
GC_7_54 b_7 NI_7 NS_54 0 -5.2745957926989898e-05
GC_7_55 b_7 NI_7 NS_55 0 -1.4325005217061793e-05
GC_7_56 b_7 NI_7 NS_56 0 -1.8002955538546896e-05
GC_7_57 b_7 NI_7 NS_57 0 -2.7149276126787048e-05
GC_7_58 b_7 NI_7 NS_58 0 -1.2989279596568725e-05
GC_7_59 b_7 NI_7 NS_59 0 -1.9441644438439541e-05
GC_7_60 b_7 NI_7 NS_60 0 5.4890786149537805e-06
GC_7_61 b_7 NI_7 NS_61 0 8.5556714407722106e-09
GC_7_62 b_7 NI_7 NS_62 0 -6.8782371264959805e-11
GC_7_63 b_7 NI_7 NS_63 0 1.9395402785764801e-11
GC_7_64 b_7 NI_7 NS_64 0 -1.1529163919598110e-10
GC_7_65 b_7 NI_7 NS_65 0 -2.0028560946062559e-06
GC_7_66 b_7 NI_7 NS_66 0 -1.3631238314291123e-06
GC_7_67 b_7 NI_7 NS_67 0 -6.1770680038347812e-06
GC_7_68 b_7 NI_7 NS_68 0 1.3444025569354297e-05
GC_7_69 b_7 NI_7 NS_69 0 3.4355390717192790e-05
GC_7_70 b_7 NI_7 NS_70 0 1.2051900028178313e-05
GC_7_71 b_7 NI_7 NS_71 0 3.1744499942199238e-05
GC_7_72 b_7 NI_7 NS_72 0 -2.5606784604828128e-05
GC_7_73 b_7 NI_7 NS_73 0 -3.9672992881193003e-05
GC_7_74 b_7 NI_7 NS_74 0 -4.8329187031210138e-05
GC_7_75 b_7 NI_7 NS_75 0 -2.0078434807717822e-05
GC_7_76 b_7 NI_7 NS_76 0 1.0823485809187198e-05
GC_7_77 b_7 NI_7 NS_77 0 5.4292689603850797e-06
GC_7_78 b_7 NI_7 NS_78 0 1.5199022833234827e-06
GC_7_79 b_7 NI_7 NS_79 0 -1.0987726510998054e-05
GC_7_80 b_7 NI_7 NS_80 0 -6.5992099095698996e-06
GC_7_81 b_7 NI_7 NS_81 0 -1.0349953947744301e-05
GC_7_82 b_7 NI_7 NS_82 0 -2.1316754054514227e-07
GC_7_83 b_7 NI_7 NS_83 0 -1.2660235847172915e-09
GC_7_84 b_7 NI_7 NS_84 0 -2.5543420716107330e-08
GC_7_85 b_7 NI_7 NS_85 0 -4.2480397441673574e-03
GC_7_86 b_7 NI_7 NS_86 0 -3.4907699661083031e-03
GC_7_87 b_7 NI_7 NS_87 0 -1.2926398894721150e-02
GC_7_88 b_7 NI_7 NS_88 0 1.7064707778669270e-02
GC_7_89 b_7 NI_7 NS_89 0 1.7381905682378011e-02
GC_7_90 b_7 NI_7 NS_90 0 -1.9436891301835148e-02
GC_7_91 b_7 NI_7 NS_91 0 -3.3160398514071696e-02
GC_7_92 b_7 NI_7 NS_92 0 2.5454388825887825e-02
GC_7_93 b_7 NI_7 NS_93 0 4.0799770158819408e-02
GC_7_94 b_7 NI_7 NS_94 0 -1.1454429793721684e-02
GC_7_95 b_7 NI_7 NS_95 0 -2.1063045483320990e-02
GC_7_96 b_7 NI_7 NS_96 0 1.5303540867818164e-02
GC_7_97 b_7 NI_7 NS_97 0 1.4115522373870178e-02
GC_7_98 b_7 NI_7 NS_98 0 -3.7637543469367252e-03
GC_7_99 b_7 NI_7 NS_99 0 7.0728043549367625e-03
GC_7_100 b_7 NI_7 NS_100 0 1.3571593784218745e-02
GC_7_101 b_7 NI_7 NS_101 0 -1.8513494007626723e-06
GC_7_102 b_7 NI_7 NS_102 0 2.5575445489220321e-07
GC_7_103 b_7 NI_7 NS_103 0 1.6675703264204748e-09
GC_7_104 b_7 NI_7 NS_104 0 1.3815226051981620e-08
GC_7_105 b_7 NI_7 NS_105 0 1.1369543036031022e-03
GC_7_106 b_7 NI_7 NS_106 0 -2.1664743216562102e-03
GC_7_107 b_7 NI_7 NS_107 0 3.4943906451710693e-03
GC_7_108 b_7 NI_7 NS_108 0 -1.2990553285539714e-02
GC_7_109 b_7 NI_7 NS_109 0 -3.9378869911133207e-02
GC_7_110 b_7 NI_7 NS_110 0 -3.6054851366724804e-04
GC_7_111 b_7 NI_7 NS_111 0 -2.6238831231058937e-02
GC_7_112 b_7 NI_7 NS_112 0 2.8978927055115893e-02
GC_7_113 b_7 NI_7 NS_113 0 5.2196790951274809e-02
GC_7_114 b_7 NI_7 NS_114 0 3.8196066071054524e-02
GC_7_115 b_7 NI_7 NS_115 0 1.7566178593826341e-02
GC_7_116 b_7 NI_7 NS_116 0 -1.4392572454675156e-02
GC_7_117 b_7 NI_7 NS_117 0 -9.1635687506150358e-03
GC_7_118 b_7 NI_7 NS_118 0 -3.7446291397158428e-03
GC_7_119 b_7 NI_7 NS_119 0 8.0613894067779780e-03
GC_7_120 b_7 NI_7 NS_120 0 5.8589432136555040e-03
GC_7_121 b_7 NI_7 NS_121 0 -1.5463085782081824e-05
GC_7_122 b_7 NI_7 NS_122 0 -3.7113238203608699e-06
GC_7_123 b_7 NI_7 NS_123 0 -2.3018577090184498e-08
GC_7_124 b_7 NI_7 NS_124 0 -3.8858819412814409e-07
GC_7_125 b_7 NI_7 NS_125 0 4.5345248115713985e-03
GC_7_126 b_7 NI_7 NS_126 0 3.8285448816379906e-03
GC_7_127 b_7 NI_7 NS_127 0 1.3835635213407260e-02
GC_7_128 b_7 NI_7 NS_128 0 -2.1353741124443226e-02
GC_7_129 b_7 NI_7 NS_129 0 -2.2486098121026522e-02
GC_7_130 b_7 NI_7 NS_130 0 2.6120598049385206e-02
GC_7_131 b_7 NI_7 NS_131 0 3.8309152499632501e-02
GC_7_132 b_7 NI_7 NS_132 0 -3.0087483901807922e-02
GC_7_133 b_7 NI_7 NS_133 0 -4.8554176854155272e-02
GC_7_134 b_7 NI_7 NS_134 0 1.9895874892674990e-02
GC_7_135 b_7 NI_7 NS_135 0 2.6986021369989413e-02
GC_7_136 b_7 NI_7 NS_136 0 -1.5889692568148695e-02
GC_7_137 b_7 NI_7 NS_137 0 -1.4309119112052000e-02
GC_7_138 b_7 NI_7 NS_138 0 6.9209623898226474e-03
GC_7_139 b_7 NI_7 NS_139 0 -4.7570075546656152e-03
GC_7_140 b_7 NI_7 NS_140 0 -1.6677668350921087e-02
GC_7_141 b_7 NI_7 NS_141 0 9.0218499076511396e-05
GC_7_142 b_7 NI_7 NS_142 0 3.5894574940617367e-06
GC_7_143 b_7 NI_7 NS_143 0 5.3419378208384192e-09
GC_7_144 b_7 NI_7 NS_144 0 6.0135184560224317e-07
GC_7_145 b_7 NI_7 NS_145 0 4.7513059778792360e-02
GC_7_146 b_7 NI_7 NS_146 0 -9.6277217005798759e-03
GC_7_147 b_7 NI_7 NS_147 0 -4.5583693078616185e-02
GC_7_148 b_7 NI_7 NS_148 0 2.0520641397986247e-02
GC_7_149 b_7 NI_7 NS_149 0 -5.7692164632266209e-02
GC_7_150 b_7 NI_7 NS_150 0 -6.7344959227193024e-02
GC_7_151 b_7 NI_7 NS_151 0 6.3851924366771756e-02
GC_7_152 b_7 NI_7 NS_152 0 -2.2031906852666681e-02
GC_7_153 b_7 NI_7 NS_153 0 2.8432503096589755e-02
GC_7_154 b_7 NI_7 NS_154 0 8.9369945454574190e-02
GC_7_155 b_7 NI_7 NS_155 0 -5.4359625111176590e-02
GC_7_156 b_7 NI_7 NS_156 0 2.7514735049838975e-03
GC_7_157 b_7 NI_7 NS_157 0 -1.3881471252999364e-02
GC_7_158 b_7 NI_7 NS_158 0 -4.7121695848641960e-02
GC_7_159 b_7 NI_7 NS_159 0 1.6357843729325555e-02
GC_7_160 b_7 NI_7 NS_160 0 -3.9002014227731578e-02
GC_7_161 b_7 NI_7 NS_161 0 -5.5372266664983193e-08
GC_7_162 b_7 NI_7 NS_162 0 -2.0698404009485823e-09
GC_7_163 b_7 NI_7 NS_163 0 -1.0036912891436134e-10
GC_7_164 b_7 NI_7 NS_164 0 3.2118675203965048e-10
GC_7_165 b_7 NI_7 NS_165 0 -1.3057976893899547e-05
GC_7_166 b_7 NI_7 NS_166 0 -1.2121355214976902e-05
GC_7_167 b_7 NI_7 NS_167 0 -4.4199162038479153e-05
GC_7_168 b_7 NI_7 NS_168 0 4.2015911154331553e-05
GC_7_169 b_7 NI_7 NS_169 0 4.9655942344418255e-05
GC_7_170 b_7 NI_7 NS_170 0 -4.5267462596750191e-05
GC_7_171 b_7 NI_7 NS_171 0 -1.0660547764705324e-04
GC_7_172 b_7 NI_7 NS_172 0 6.5657554186562090e-05
GC_7_173 b_7 NI_7 NS_173 0 1.2561071361605848e-04
GC_7_174 b_7 NI_7 NS_174 0 -8.6598583089383844e-06
GC_7_175 b_7 NI_7 NS_175 0 -5.8946727833178148e-05
GC_7_176 b_7 NI_7 NS_176 0 4.0869752558371764e-05
GC_7_177 b_7 NI_7 NS_177 0 4.4689149851088784e-05
GC_7_178 b_7 NI_7 NS_178 0 -5.2904252762722482e-06
GC_7_179 b_7 NI_7 NS_179 0 2.5177397457381439e-05
GC_7_180 b_7 NI_7 NS_180 0 3.8246853472087470e-05
GC_7_181 b_7 NI_7 NS_181 0 5.9928607787127386e-08
GC_7_182 b_7 NI_7 NS_182 0 1.3687395134155103e-09
GC_7_183 b_7 NI_7 NS_183 0 1.6472083144839028e-10
GC_7_184 b_7 NI_7 NS_184 0 -6.9445082709331730e-10
GC_7_185 b_7 NI_7 NS_185 0 -9.5337281204900740e-06
GC_7_186 b_7 NI_7 NS_186 0 -5.9434691484757439e-06
GC_7_187 b_7 NI_7 NS_187 0 1.9546602872675080e-06
GC_7_188 b_7 NI_7 NS_188 0 -1.4939358952878093e-05
GC_7_189 b_7 NI_7 NS_189 0 -1.1210929150737505e-04
GC_7_190 b_7 NI_7 NS_190 0 3.7775222383628991e-05
GC_7_191 b_7 NI_7 NS_191 0 -7.9681739295999783e-05
GC_7_192 b_7 NI_7 NS_192 0 7.7640564228990958e-05
GC_7_193 b_7 NI_7 NS_193 0 1.9081247283508868e-04
GC_7_194 b_7 NI_7 NS_194 0 1.3314012857386484e-04
GC_7_195 b_7 NI_7 NS_195 0 5.7036572023150067e-05
GC_7_196 b_7 NI_7 NS_196 0 -1.9615088201760255e-05
GC_7_197 b_7 NI_7 NS_197 0 -5.4481406855992492e-06
GC_7_198 b_7 NI_7 NS_198 0 -8.3263834426774030e-06
GC_7_199 b_7 NI_7 NS_199 0 3.7160520039688663e-05
GC_7_200 b_7 NI_7 NS_200 0 9.7251560104406765e-06
GC_7_201 b_7 NI_7 NS_201 0 -2.5754064648857980e-08
GC_7_202 b_7 NI_7 NS_202 0 1.1438284879377590e-09
GC_7_203 b_7 NI_7 NS_203 0 -1.1059887723800844e-11
GC_7_204 b_7 NI_7 NS_204 0 3.1894463353368207e-11
GC_7_205 b_7 NI_7 NS_205 0 4.4269009498271563e-06
GC_7_206 b_7 NI_7 NS_206 0 2.3386907252314359e-06
GC_7_207 b_7 NI_7 NS_207 0 9.9199540048149036e-06
GC_7_208 b_7 NI_7 NS_208 0 9.7652561060266453e-06
GC_7_209 b_7 NI_7 NS_209 0 1.8817727602255084e-05
GC_7_210 b_7 NI_7 NS_210 0 -2.3372956456713281e-05
GC_7_211 b_7 NI_7 NS_211 0 1.1289948438730449e-05
GC_7_212 b_7 NI_7 NS_212 0 -3.2013245051689467e-06
GC_7_213 b_7 NI_7 NS_213 0 -6.5988113720183717e-06
GC_7_214 b_7 NI_7 NS_214 0 -5.3073158508640626e-05
GC_7_215 b_7 NI_7 NS_215 0 -1.4827253649678679e-05
GC_7_216 b_7 NI_7 NS_216 0 -1.7892238087596487e-05
GC_7_217 b_7 NI_7 NS_217 0 -2.7603790063017063e-05
GC_7_218 b_7 NI_7 NS_218 0 -1.2421187980035711e-05
GC_7_219 b_7 NI_7 NS_219 0 -1.9027359143531106e-05
GC_7_220 b_7 NI_7 NS_220 0 5.9411137870301416e-06
GC_7_221 b_7 NI_7 NS_221 0 1.1016516164503194e-09
GC_7_222 b_7 NI_7 NS_222 0 -1.2971137923553618e-10
GC_7_223 b_7 NI_7 NS_223 0 1.7862402132351913e-11
GC_7_224 b_7 NI_7 NS_224 0 -9.6106651331500777e-11
GC_7_225 b_7 NI_7 NS_225 0 -1.9128837492933734e-06
GC_7_226 b_7 NI_7 NS_226 0 -1.1371208177488090e-06
GC_7_227 b_7 NI_7 NS_227 0 -6.0331197681405545e-06
GC_7_228 b_7 NI_7 NS_228 0 1.3796847544603874e-05
GC_7_229 b_7 NI_7 NS_229 0 3.5155088846427304e-05
GC_7_230 b_7 NI_7 NS_230 0 1.1739874225946811e-05
GC_7_231 b_7 NI_7 NS_231 0 3.2374480861564711e-05
GC_7_232 b_7 NI_7 NS_232 0 -2.5607924418786508e-05
GC_7_233 b_7 NI_7 NS_233 0 -3.9768424611497577e-05
GC_7_234 b_7 NI_7 NS_234 0 -4.9607873062286408e-05
GC_7_235 b_7 NI_7 NS_235 0 -1.9812838165824242e-05
GC_7_236 b_7 NI_7 NS_236 0 1.0190725397008221e-05
GC_7_237 b_7 NI_7 NS_237 0 4.9362496595826359e-06
GC_7_238 b_7 NI_7 NS_238 0 3.9503206173261735e-07
GC_7_239 b_7 NI_7 NS_239 0 -1.2398818543469652e-05
GC_7_240 b_7 NI_7 NS_240 0 -7.1395544494296740e-06
GD_7_1 b_7 NI_7 NA_1 0 -9.6795238849265317e-07
GD_7_2 b_7 NI_7 NA_2 0 1.0239339449112561e-05
GD_7_3 b_7 NI_7 NA_3 0 1.3447891948918530e-05
GD_7_4 b_7 NI_7 NA_4 0 3.5140063146195559e-06
GD_7_5 b_7 NI_7 NA_5 0 6.7712145152012647e-03
GD_7_6 b_7 NI_7 NA_6 0 -3.3437475320033105e-03
GD_7_7 b_7 NI_7 NA_7 0 -9.6518873014063492e-03
GD_7_8 b_7 NI_7 NA_8 0 5.5541158591456887e-03
GD_7_9 b_7 NI_7 NA_9 0 2.4227205234474679e-05
GD_7_10 b_7 NI_7 NA_10 0 -5.3839434842203685e-05
GD_7_11 b_7 NI_7 NA_11 0 1.4712435961715527e-05
GD_7_12 b_7 NI_7 NA_12 0 3.3225507489141470e-06
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 -2.3908523376360200e-08
GC_8_2 b_8 NI_8 NS_2 0 1.2224990530175730e-09
GC_8_3 b_8 NI_8 NS_3 0 2.1485244883925260e-11
GC_8_4 b_8 NI_8 NS_4 0 -1.7590191201697083e-10
GC_8_5 b_8 NI_8 NS_5 0 1.8930935618405023e-06
GC_8_6 b_8 NI_8 NS_6 0 -4.2142295402140277e-06
GC_8_7 b_8 NI_8 NS_7 0 2.5243758763162093e-06
GC_8_8 b_8 NI_8 NS_8 0 5.0918793191389289e-08
GC_8_9 b_8 NI_8 NS_9 0 -1.6404752179600091e-06
GC_8_10 b_8 NI_8 NS_10 0 -4.6526884260699409e-06
GC_8_11 b_8 NI_8 NS_11 0 9.2496720811147026e-07
GC_8_12 b_8 NI_8 NS_12 0 -7.3960094374648206e-06
GC_8_13 b_8 NI_8 NS_13 0 -9.0332922200943151e-06
GC_8_14 b_8 NI_8 NS_14 0 -4.5741776910452687e-06
GC_8_15 b_8 NI_8 NS_15 0 -3.2971985659804730e-06
GC_8_16 b_8 NI_8 NS_16 0 1.4734753333752264e-06
GC_8_17 b_8 NI_8 NS_17 0 -1.9003376107287650e-06
GC_8_18 b_8 NI_8 NS_18 0 -4.7685538269711010e-07
GC_8_19 b_8 NI_8 NS_19 0 -3.2417990197473164e-06
GC_8_20 b_8 NI_8 NS_20 0 -1.4954314827063772e-06
GC_8_21 b_8 NI_8 NS_21 0 2.0299545770449321e-08
GC_8_22 b_8 NI_8 NS_22 0 -1.0034002210460646e-09
GC_8_23 b_8 NI_8 NS_23 0 -1.9109341689581415e-11
GC_8_24 b_8 NI_8 NS_24 0 1.5480761937531662e-10
GC_8_25 b_8 NI_8 NS_25 0 -1.0725434548538138e-06
GC_8_26 b_8 NI_8 NS_26 0 -8.5344072598230112e-07
GC_8_27 b_8 NI_8 NS_27 0 -1.9513310564582947e-06
GC_8_28 b_8 NI_8 NS_28 0 -1.3188102615803828e-08
GC_8_29 b_8 NI_8 NS_29 0 -3.0922826700100027e-06
GC_8_30 b_8 NI_8 NS_30 0 7.4413707336782746e-07
GC_8_31 b_8 NI_8 NS_31 0 -4.1341886516126113e-06
GC_8_32 b_8 NI_8 NS_32 0 4.2201126273883127e-06
GC_8_33 b_8 NI_8 NS_33 0 3.1590338509409375e-06
GC_8_34 b_8 NI_8 NS_34 0 5.3423797236740300e-06
GC_8_35 b_8 NI_8 NS_35 0 -9.0664822714762075e-07
GC_8_36 b_8 NI_8 NS_36 0 5.9322125158233579e-06
GC_8_37 b_8 NI_8 NS_37 0 5.9750663833850115e-06
GC_8_38 b_8 NI_8 NS_38 0 3.2312446396819881e-06
GC_8_39 b_8 NI_8 NS_39 0 5.7326862226021451e-06
GC_8_40 b_8 NI_8 NS_40 0 1.6824495306353415e-06
GC_8_41 b_8 NI_8 NS_41 0 8.5552414657857903e-09
GC_8_42 b_8 NI_8 NS_42 0 -6.8743886753121097e-11
GC_8_43 b_8 NI_8 NS_43 0 1.9395794000963330e-11
GC_8_44 b_8 NI_8 NS_44 0 -1.1529482108751473e-10
GC_8_45 b_8 NI_8 NS_45 0 -2.0030699890984852e-06
GC_8_46 b_8 NI_8 NS_46 0 -1.3631111479816519e-06
GC_8_47 b_8 NI_8 NS_47 0 -6.1775754697539286e-06
GC_8_48 b_8 NI_8 NS_48 0 1.3443933064859785e-05
GC_8_49 b_8 NI_8 NS_49 0 3.4355404529504172e-05
GC_8_50 b_8 NI_8 NS_50 0 1.2053255983872879e-05
GC_8_51 b_8 NI_8 NS_51 0 3.1744906799396686e-05
GC_8_52 b_8 NI_8 NS_52 0 -2.5605882352139866e-05
GC_8_53 b_8 NI_8 NS_53 0 -3.9671496519268456e-05
GC_8_54 b_8 NI_8 NS_54 0 -4.8330195180565401e-05
GC_8_55 b_8 NI_8 NS_55 0 -2.0078506796946053e-05
GC_8_56 b_8 NI_8 NS_56 0 1.0823028506417180e-05
GC_8_57 b_8 NI_8 NS_57 0 5.4289946730006231e-06
GC_8_58 b_8 NI_8 NS_58 0 1.5197982943230366e-06
GC_8_59 b_8 NI_8 NS_59 0 -1.0987816131006844e-05
GC_8_60 b_8 NI_8 NS_60 0 -6.5991927488239113e-06
GC_8_61 b_8 NI_8 NS_61 0 -2.8873926808889625e-08
GC_8_62 b_8 NI_8 NS_62 0 8.6794416700660869e-10
GC_8_63 b_8 NI_8 NS_63 0 -1.4875514101685988e-11
GC_8_64 b_8 NI_8 NS_64 0 6.7611104861018029e-11
GC_8_65 b_8 NI_8 NS_65 0 4.0217078753580034e-06
GC_8_66 b_8 NI_8 NS_66 0 2.7674566952151132e-06
GC_8_67 b_8 NI_8 NS_67 0 9.4641818825118519e-06
GC_8_68 b_8 NI_8 NS_68 0 1.0309426271287153e-05
GC_8_69 b_8 NI_8 NS_69 0 1.9370375339903224e-05
GC_8_70 b_8 NI_8 NS_70 0 -2.2294981830877045e-05
GC_8_71 b_8 NI_8 NS_71 0 1.1424263010993573e-05
GC_8_72 b_8 NI_8 NS_72 0 -2.5122774186767328e-06
GC_8_73 b_8 NI_8 NS_73 0 -4.9910964781205054e-06
GC_8_74 b_8 NI_8 NS_74 0 -5.2807265593622214e-05
GC_8_75 b_8 NI_8 NS_75 0 -1.4282076805887971e-05
GC_8_76 b_8 NI_8 NS_76 0 -1.7913591270644068e-05
GC_8_77 b_8 NI_8 NS_77 0 -2.7057560551645508e-05
GC_8_78 b_8 NI_8 NS_78 0 -1.2982227715911269e-05
GC_8_79 b_8 NI_8 NS_79 0 -1.9361092604084692e-05
GC_8_80 b_8 NI_8 NS_80 0 5.4944462731053547e-06
GC_8_81 b_8 NI_8 NS_81 0 -1.8513499671749782e-06
GC_8_82 b_8 NI_8 NS_82 0 2.5575447761495729e-07
GC_8_83 b_8 NI_8 NS_83 0 1.6675703954548088e-09
GC_8_84 b_8 NI_8 NS_84 0 1.3815225133507906e-08
GC_8_85 b_8 NI_8 NS_85 0 1.1369543523708770e-03
GC_8_86 b_8 NI_8 NS_86 0 -2.1664743002075145e-03
GC_8_87 b_8 NI_8 NS_87 0 3.4943906894795147e-03
GC_8_88 b_8 NI_8 NS_88 0 -1.2990553244949939e-02
GC_8_89 b_8 NI_8 NS_89 0 -3.9378869866391206e-02
GC_8_90 b_8 NI_8 NS_90 0 -3.6054868580438900e-04
GC_8_91 b_8 NI_8 NS_91 0 -2.6238831259680944e-02
GC_8_92 b_8 NI_8 NS_92 0 2.8978926982022462e-02
GC_8_93 b_8 NI_8 NS_93 0 5.2196790921334897e-02
GC_8_94 b_8 NI_8 NS_94 0 3.8196066152336956e-02
GC_8_95 b_8 NI_8 NS_95 0 1.7566178694232281e-02
GC_8_96 b_8 NI_8 NS_96 0 -1.4392572524278668e-02
GC_8_97 b_8 NI_8 NS_97 0 -9.1635688226141473e-03
GC_8_98 b_8 NI_8 NS_98 0 -3.7446293231003414e-03
GC_8_99 b_8 NI_8 NS_99 0 8.0613892485659738e-03
GC_8_100 b_8 NI_8 NS_100 0 5.8589431802663332e-03
GC_8_101 b_8 NI_8 NS_101 0 -1.0349953958273454e-05
GC_8_102 b_8 NI_8 NS_102 0 -2.1316754009410218e-07
GC_8_103 b_8 NI_8 NS_103 0 -1.2660235834495063e-09
GC_8_104 b_8 NI_8 NS_104 0 -2.5543420737366643e-08
GC_8_105 b_8 NI_8 NS_105 0 -4.2480397462394638e-03
GC_8_106 b_8 NI_8 NS_106 0 -3.4907699650810575e-03
GC_8_107 b_8 NI_8 NS_107 0 -1.2926398897791656e-02
GC_8_108 b_8 NI_8 NS_108 0 1.7064707780997539e-02
GC_8_109 b_8 NI_8 NS_109 0 1.7381905686225566e-02
GC_8_110 b_8 NI_8 NS_110 0 -1.9436891295307176e-02
GC_8_111 b_8 NI_8 NS_111 0 -3.3160398510843715e-02
GC_8_112 b_8 NI_8 NS_112 0 2.5454388828446313e-02
GC_8_113 b_8 NI_8 NS_113 0 4.0799770165464627e-02
GC_8_114 b_8 NI_8 NS_114 0 -1.1454429797341313e-02
GC_8_115 b_8 NI_8 NS_115 0 -2.1063045481597271e-02
GC_8_116 b_8 NI_8 NS_116 0 1.5303540864951413e-02
GC_8_117 b_8 NI_8 NS_117 0 1.4115522372272054e-02
GC_8_118 b_8 NI_8 NS_118 0 -3.7637543500676149e-03
GC_8_119 b_8 NI_8 NS_119 0 7.0728043525808224e-03
GC_8_120 b_8 NI_8 NS_120 0 1.3571593783590505e-02
GC_8_121 b_8 NI_8 NS_121 0 9.0218498754969571e-05
GC_8_122 b_8 NI_8 NS_122 0 3.5894575141347713e-06
GC_8_123 b_8 NI_8 NS_123 0 5.3419380499845483e-09
GC_8_124 b_8 NI_8 NS_124 0 6.0135184366276081e-07
GC_8_125 b_8 NI_8 NS_125 0 4.7513059791977751e-02
GC_8_126 b_8 NI_8 NS_126 0 -9.6277216961446373e-03
GC_8_127 b_8 NI_8 NS_127 0 -4.5583693056558745e-02
GC_8_128 b_8 NI_8 NS_128 0 2.0520641417564475e-02
GC_8_129 b_8 NI_8 NS_129 0 -5.7692164564510214e-02
GC_8_130 b_8 NI_8 NS_130 0 -6.7344959263317850e-02
GC_8_131 b_8 NI_8 NS_131 0 6.3851924433093260e-02
GC_8_132 b_8 NI_8 NS_132 0 -2.2031906886441049e-02
GC_8_133 b_8 NI_8 NS_133 0 2.8432503060880094e-02
GC_8_134 b_8 NI_8 NS_134 0 8.9369945281271110e-02
GC_8_135 b_8 NI_8 NS_135 0 -5.4359625146366587e-02
GC_8_136 b_8 NI_8 NS_136 0 2.7514734238907896e-03
GC_8_137 b_8 NI_8 NS_137 0 -1.3881471352158836e-02
GC_8_138 b_8 NI_8 NS_138 0 -4.7121695896976283e-02
GC_8_139 b_8 NI_8 NS_139 0 1.6357843643316688e-02
GC_8_140 b_8 NI_8 NS_140 0 -3.9002014229856073e-02
GC_8_141 b_8 NI_8 NS_141 0 -1.5463085782082915e-05
GC_8_142 b_8 NI_8 NS_142 0 -3.7113238203605209e-06
GC_8_143 b_8 NI_8 NS_143 0 -2.3018577090181689e-08
GC_8_144 b_8 NI_8 NS_144 0 -3.8858819412816617e-07
GC_8_145 b_8 NI_8 NS_145 0 4.5345248115714358e-03
GC_8_146 b_8 NI_8 NS_146 0 3.8285448816379780e-03
GC_8_147 b_8 NI_8 NS_147 0 1.3835635213407272e-02
GC_8_148 b_8 NI_8 NS_148 0 -2.1353741124443271e-02
GC_8_149 b_8 NI_8 NS_149 0 -2.2486098121026591e-02
GC_8_150 b_8 NI_8 NS_150 0 2.6120598049385192e-02
GC_8_151 b_8 NI_8 NS_151 0 3.8309152499632466e-02
GC_8_152 b_8 NI_8 NS_152 0 -3.0087483901807904e-02
GC_8_153 b_8 NI_8 NS_153 0 -4.8554176854155230e-02
GC_8_154 b_8 NI_8 NS_154 0 1.9895874892675001e-02
GC_8_155 b_8 NI_8 NS_155 0 2.6986021369989413e-02
GC_8_156 b_8 NI_8 NS_156 0 -1.5889692568148716e-02
GC_8_157 b_8 NI_8 NS_157 0 -1.4309119112052010e-02
GC_8_158 b_8 NI_8 NS_158 0 6.9209623898226283e-03
GC_8_159 b_8 NI_8 NS_159 0 -4.7570075546656343e-03
GC_8_160 b_8 NI_8 NS_160 0 -1.6677668350921087e-02
GC_8_161 b_8 NI_8 NS_161 0 5.9902842863302531e-08
GC_8_162 b_8 NI_8 NS_162 0 1.3695849204786296e-09
GC_8_163 b_8 NI_8 NS_163 0 1.6472719001903974e-10
GC_8_164 b_8 NI_8 NS_164 0 -6.9450434269704248e-10
GC_8_165 b_8 NI_8 NS_165 0 -9.5511617838509243e-06
GC_8_166 b_8 NI_8 NS_166 0 -5.9491244241203354e-06
GC_8_167 b_8 NI_8 NS_167 0 1.9276576281713021e-06
GC_8_168 b_8 NI_8 NS_168 0 -1.4956781608311702e-05
GC_8_169 b_8 NI_8 NS_169 0 -1.1212294648190245e-04
GC_8_170 b_8 NI_8 NS_170 0 3.7878411785785902e-05
GC_8_171 b_8 NI_8 NS_171 0 -7.9642075961477310e-05
GC_8_172 b_8 NI_8 NS_172 0 7.7704165831143061e-05
GC_8_173 b_8 NI_8 NS_173 0 1.9090727074380369e-04
GC_8_174 b_8 NI_8 NS_174 0 1.3304677911219376e-04
GC_8_175 b_8 NI_8 NS_175 0 5.7019878415249709e-05
GC_8_176 b_8 NI_8 NS_176 0 -1.9652975331635071e-05
GC_8_177 b_8 NI_8 NS_177 0 -5.4751856196237679e-06
GC_8_178 b_8 NI_8 NS_178 0 -8.3218542127282402e-06
GC_8_179 b_8 NI_8 NS_179 0 3.7156186010252443e-05
GC_8_180 b_8 NI_8 NS_180 0 9.7277837983443741e-06
GC_8_181 b_8 NI_8 NS_181 0 -5.5359599424378504e-08
GC_8_182 b_8 NI_8 NS_182 0 -2.0704056517732812e-09
GC_8_183 b_8 NI_8 NS_183 0 -1.0037045945726831e-10
GC_8_184 b_8 NI_8 NS_184 0 3.2121630299065353e-10
GC_8_185 b_8 NI_8 NS_185 0 -1.3058224327566672e-05
GC_8_186 b_8 NI_8 NS_186 0 -1.2120478538255689e-05
GC_8_187 b_8 NI_8 NS_187 0 -4.4199314341231065e-05
GC_8_188 b_8 NI_8 NS_188 0 4.2016566232179795e-05
GC_8_189 b_8 NI_8 NS_189 0 4.9656079253780703e-05
GC_8_190 b_8 NI_8 NS_190 0 -4.5266201048751713e-05
GC_8_191 b_8 NI_8 NS_191 0 -1.0660475212441537e-04
GC_8_192 b_8 NI_8 NS_192 0 6.5659091562060752e-05
GC_8_193 b_8 NI_8 NS_193 0 1.2561218753332507e-04
GC_8_194 b_8 NI_8 NS_194 0 -8.6604311644105561e-06
GC_8_195 b_8 NI_8 NS_195 0 -5.8946835085473599e-05
GC_8_196 b_8 NI_8 NS_196 0 4.0870477952169338e-05
GC_8_197 b_8 NI_8 NS_197 0 4.4689994150164994e-05
GC_8_198 b_8 NI_8 NS_198 0 -5.2895347108169919e-06
GC_8_199 b_8 NI_8 NS_199 0 2.5178844363802749e-05
GC_8_200 b_8 NI_8 NS_200 0 3.8247291133897129e-05
GC_8_201 b_8 NI_8 NS_201 0 1.1017305163556556e-09
GC_8_202 b_8 NI_8 NS_202 0 -1.2973356084544113e-10
GC_8_203 b_8 NI_8 NS_203 0 1.7862140539337658e-11
GC_8_204 b_8 NI_8 NS_204 0 -9.6104624647440653e-11
GC_8_205 b_8 NI_8 NS_205 0 -1.9127610684637098e-06
GC_8_206 b_8 NI_8 NS_206 0 -1.1371602954370355e-06
GC_8_207 b_8 NI_8 NS_207 0 -6.0327984341615081e-06
GC_8_208 b_8 NI_8 NS_208 0 1.3796838394416037e-05
GC_8_209 b_8 NI_8 NS_209 0 3.5155038201109612e-05
GC_8_210 b_8 NI_8 NS_210 0 1.1739173831793734e-05
GC_8_211 b_8 NI_8 NS_211 0 3.2374347249562897e-05
GC_8_212 b_8 NI_8 NS_212 0 -2.5608400564646464e-05
GC_8_213 b_8 NI_8 NS_213 0 -3.9769248107332664e-05
GC_8_214 b_8 NI_8 NS_214 0 -4.9607554737818210e-05
GC_8_215 b_8 NI_8 NS_215 0 -1.9812840984530885e-05
GC_8_216 b_8 NI_8 NS_216 0 1.0190879443117163e-05
GC_8_217 b_8 NI_8 NS_217 0 4.9362771498468141e-06
GC_8_218 b_8 NI_8 NS_218 0 3.9503380476092955e-07
GC_8_219 b_8 NI_8 NS_219 0 -1.2398868750962824e-05
GC_8_220 b_8 NI_8 NS_220 0 -7.1395621963900314e-06
GC_8_221 b_8 NI_8 NS_221 0 -2.5925743947527895e-08
GC_8_222 b_8 NI_8 NS_222 0 1.1529333622976366e-09
GC_8_223 b_8 NI_8 NS_223 0 -1.0993201109843437e-11
GC_8_224 b_8 NI_8 NS_224 0 3.1284473599936635e-11
GC_8_225 b_8 NI_8 NS_225 0 4.4658843764132860e-06
GC_8_226 b_8 NI_8 NS_226 0 2.2626211872327774e-06
GC_8_227 b_8 NI_8 NS_227 0 9.9229977550412083e-06
GC_8_228 b_8 NI_8 NS_228 0 9.6721828705981198e-06
GC_8_229 b_8 NI_8 NS_229 0 1.8821990088643682e-05
GC_8_230 b_8 NI_8 NS_230 0 -2.3464206870715885e-05
GC_8_231 b_8 NI_8 NS_231 0 1.1213140551861190e-05
GC_8_232 b_8 NI_8 NS_232 0 -3.3843357992134624e-06
GC_8_233 b_8 NI_8 NS_233 0 -6.7473936959766888e-06
GC_8_234 b_8 NI_8 NS_234 0 -5.3021724352220091e-05
GC_8_235 b_8 NI_8 NS_235 0 -1.4872212717022044e-05
GC_8_236 b_8 NI_8 NS_236 0 -1.7984609360484102e-05
GC_8_237 b_8 NI_8 NS_237 0 -2.7699452931528875e-05
GC_8_238 b_8 NI_8 NS_238 0 -1.2430480263581680e-05
GC_8_239 b_8 NI_8 NS_239 0 -1.9111947280303820e-05
GC_8_240 b_8 NI_8 NS_240 0 5.9354257008595398e-06
GD_8_1 b_8 NI_8 NA_1 0 1.0254584098881482e-05
GD_8_2 b_8 NI_8 NA_2 0 -9.6392317503807296e-07
GD_8_3 b_8 NI_8 NA_3 0 3.5134960645226050e-06
GD_8_4 b_8 NI_8 NA_4 0 1.3060694799291506e-05
GD_8_5 b_8 NI_8 NA_5 0 -3.3437475291121354e-03
GD_8_6 b_8 NI_8 NA_6 0 6.7712145109744158e-03
GD_8_7 b_8 NI_8 NA_7 0 5.5541159113289638e-03
GD_8_8 b_8 NI_8 NA_8 0 -9.6518873014063335e-03
GD_8_9 b_8 NI_8 NA_9 0 -5.3853460106419274e-05
GD_8_10 b_8 NI_8 NA_10 0 2.4223441825095968e-05
GD_8_11 b_8 NI_8 NA_11 0 3.3229601080506427e-06
GD_8_12 b_8 NI_8 NA_12 0 1.5099444127781766e-05
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 1.2088123459337427e-08
GC_9_2 b_9 NI_9 NS_2 0 -8.1496970130157824e-10
GC_9_3 b_9 NI_9 NS_3 0 -1.6058681327176953e-11
GC_9_4 b_9 NI_9 NS_4 0 1.3065453480248421e-10
GC_9_5 b_9 NI_9 NS_5 0 6.7658967692906657e-08
GC_9_6 b_9 NI_9 NS_6 0 -1.2554508018271056e-08
GC_9_7 b_9 NI_9 NS_7 0 -5.8630541163050299e-07
GC_9_8 b_9 NI_9 NS_8 0 5.6735525770875182e-07
GC_9_9 b_9 NI_9 NS_9 0 1.6812066328390143e-06
GC_9_10 b_9 NI_9 NS_10 0 -5.0520096791566311e-07
GC_9_11 b_9 NI_9 NS_11 0 -9.7641443665908538e-07
GC_9_12 b_9 NI_9 NS_12 0 1.1750300024974223e-07
GC_9_13 b_9 NI_9 NS_13 0 1.6591569524997925e-06
GC_9_14 b_9 NI_9 NS_14 0 -1.1492633357344439e-06
GC_9_15 b_9 NI_9 NS_15 0 -9.0302156088360417e-07
GC_9_16 b_9 NI_9 NS_16 0 -8.6140215593144392e-07
GC_9_17 b_9 NI_9 NS_17 0 -1.1367784787962444e-06
GC_9_18 b_9 NI_9 NS_18 0 -2.5235747715113701e-07
GC_9_19 b_9 NI_9 NS_19 0 8.6997773625294326e-08
GC_9_20 b_9 NI_9 NS_20 0 1.1717150089213943e-06
GC_9_21 b_9 NI_9 NS_21 0 -8.0862474117938583e-09
GC_9_22 b_9 NI_9 NS_22 0 6.7986876039155784e-10
GC_9_23 b_9 NI_9 NS_23 0 1.5646929769061646e-11
GC_9_24 b_9 NI_9 NS_24 0 -1.2067902589302462e-10
GC_9_25 b_9 NI_9 NS_25 0 -2.1903687640893429e-06
GC_9_26 b_9 NI_9 NS_26 0 2.1886446261441094e-07
GC_9_27 b_9 NI_9 NS_27 0 -2.1895701238172224e-06
GC_9_28 b_9 NI_9 NS_28 0 2.7884237644963512e-06
GC_9_29 b_9 NI_9 NS_29 0 -1.1327109188332638e-06
GC_9_30 b_9 NI_9 NS_30 0 6.5773613987983140e-06
GC_9_31 b_9 NI_9 NS_31 0 -4.1803908124301069e-07
GC_9_32 b_9 NI_9 NS_32 0 2.1422267230030422e-06
GC_9_33 b_9 NI_9 NS_33 0 7.2190707962389696e-06
GC_9_34 b_9 NI_9 NS_34 0 5.1224404333900628e-06
GC_9_35 b_9 NI_9 NS_35 0 1.6120533390669766e-06
GC_9_36 b_9 NI_9 NS_36 0 3.1394752839629968e-06
GC_9_37 b_9 NI_9 NS_37 0 4.8357377515413603e-06
GC_9_38 b_9 NI_9 NS_38 0 1.1501563862083032e-06
GC_9_39 b_9 NI_9 NS_39 0 2.9137140609115429e-06
GC_9_40 b_9 NI_9 NS_40 0 -1.3217648764209678e-06
GC_9_41 b_9 NI_9 NS_41 0 -3.3859863904254525e-10
GC_9_42 b_9 NI_9 NS_42 0 2.4529145269220358e-10
GC_9_43 b_9 NI_9 NS_43 0 5.1902229666319652e-12
GC_9_44 b_9 NI_9 NS_44 0 -1.2433590070472335e-11
GC_9_45 b_9 NI_9 NS_45 0 -1.5827743636708918e-06
GC_9_46 b_9 NI_9 NS_46 0 7.4475468121840055e-07
GC_9_47 b_9 NI_9 NS_47 0 -2.4991417335532137e-06
GC_9_48 b_9 NI_9 NS_48 0 1.5671735100594544e-06
GC_9_49 b_9 NI_9 NS_49 0 6.6682291141731250e-07
GC_9_50 b_9 NI_9 NS_50 0 3.1010091849612044e-06
GC_9_51 b_9 NI_9 NS_51 0 -2.4063142968841994e-06
GC_9_52 b_9 NI_9 NS_52 0 3.2308341548225504e-06
GC_9_53 b_9 NI_9 NS_53 0 5.2075548500172518e-06
GC_9_54 b_9 NI_9 NS_54 0 4.2312571753700278e-06
GC_9_55 b_9 NI_9 NS_55 0 -6.0801449677925113e-08
GC_9_56 b_9 NI_9 NS_56 0 3.4339369967366203e-06
GC_9_57 b_9 NI_9 NS_57 0 5.0339181939226489e-06
GC_9_58 b_9 NI_9 NS_58 0 2.2607988292484626e-06
GC_9_59 b_9 NI_9 NS_59 0 3.8677488225692439e-06
GC_9_60 b_9 NI_9 NS_60 0 2.0110103523571253e-07
GC_9_61 b_9 NI_9 NS_61 0 -5.4833829822955736e-09
GC_9_62 b_9 NI_9 NS_62 0 -1.1889739531692169e-10
GC_9_63 b_9 NI_9 NS_63 0 -8.7976089162406984e-12
GC_9_64 b_9 NI_9 NS_64 0 1.2303198140108776e-11
GC_9_65 b_9 NI_9 NS_65 0 2.8877995215041497e-06
GC_9_66 b_9 NI_9 NS_66 0 -3.3700211751688477e-06
GC_9_67 b_9 NI_9 NS_67 0 3.9433199517964702e-06
GC_9_68 b_9 NI_9 NS_68 0 -1.1977393394484600e-06
GC_9_69 b_9 NI_9 NS_69 0 -1.9626919454646774e-06
GC_9_70 b_9 NI_9 NS_70 0 -6.4897710475789265e-06
GC_9_71 b_9 NI_9 NS_71 0 1.2536645771166293e-06
GC_9_72 b_9 NI_9 NS_72 0 -5.0193343188160694e-06
GC_9_73 b_9 NI_9 NS_73 0 -3.5332530761102703e-06
GC_9_74 b_9 NI_9 NS_74 0 -9.5121431503138647e-06
GC_9_75 b_9 NI_9 NS_75 0 -2.5204734656598353e-06
GC_9_76 b_9 NI_9 NS_76 0 -6.0280720261952257e-06
GC_9_77 b_9 NI_9 NS_77 0 -9.7106990318218545e-06
GC_9_78 b_9 NI_9 NS_78 0 -4.8418376319791716e-06
GC_9_79 b_9 NI_9 NS_79 0 -7.2832411310277787e-06
GC_9_80 b_9 NI_9 NS_80 0 5.3200533983852105e-07
GC_9_81 b_9 NI_9 NS_81 0 -2.7643471420272211e-08
GC_9_82 b_9 NI_9 NS_82 0 8.0098552561472182e-10
GC_9_83 b_9 NI_9 NS_83 0 -1.5252025686165523e-11
GC_9_84 b_9 NI_9 NS_84 0 7.2677023337438917e-11
GC_9_85 b_9 NI_9 NS_85 0 4.1256396360657731e-06
GC_9_86 b_9 NI_9 NS_86 0 2.6677180504402813e-06
GC_9_87 b_9 NI_9 NS_87 0 9.5682087960191221e-06
GC_9_88 b_9 NI_9 NS_88 0 1.0216481086741431e-05
GC_9_89 b_9 NI_9 NS_89 0 1.9376033536868980e-05
GC_9_90 b_9 NI_9 NS_90 0 -2.2593580598893458e-05
GC_9_91 b_9 NI_9 NS_91 0 1.1373791753991274e-05
GC_9_92 b_9 NI_9 NS_92 0 -2.7583655875270399e-06
GC_9_93 b_9 NI_9 NS_93 0 -5.2913335796614383e-06
GC_9_94 b_9 NI_9 NS_94 0 -5.2911832072160727e-05
GC_9_95 b_9 NI_9 NS_95 0 -1.4329145221574527e-05
GC_9_96 b_9 NI_9 NS_96 0 -1.8082862119734448e-05
GC_9_97 b_9 NI_9 NS_97 0 -2.7364161860539553e-05
GC_9_98 b_9 NI_9 NS_98 0 -1.3068178294104021e-05
GC_9_99 b_9 NI_9 NS_99 0 -1.9489167315248817e-05
GC_9_100 b_9 NI_9 NS_100 0 5.5936315706487113e-06
GC_9_101 b_9 NI_9 NS_101 0 7.1854157299091598e-09
GC_9_102 b_9 NI_9 NS_102 0 2.2464234729853902e-11
GC_9_103 b_9 NI_9 NS_103 0 2.0136508811792832e-11
GC_9_104 b_9 NI_9 NS_104 0 -1.2273053865240682e-10
GC_9_105 b_9 NI_9 NS_105 0 -2.1095036109939568e-06
GC_9_106 b_9 NI_9 NS_106 0 -1.2999235739844057e-06
GC_9_107 b_9 NI_9 NS_107 0 -6.2931075777899012e-06
GC_9_108 b_9 NI_9 NS_108 0 1.3497473419153023e-05
GC_9_109 b_9 NI_9 NS_109 0 3.4249419478038199e-05
GC_9_110 b_9 NI_9 NS_110 0 1.2262045131326663e-05
GC_9_111 b_9 NI_9 NS_111 0 3.1603970270400573e-05
GC_9_112 b_9 NI_9 NS_112 0 -2.5423271516891107e-05
GC_9_113 b_9 NI_9 NS_113 0 -3.9478419220890421e-05
GC_9_114 b_9 NI_9 NS_114 0 -4.7737605894194924e-05
GC_9_115 b_9 NI_9 NS_115 0 -1.9905276143987593e-05
GC_9_116 b_9 NI_9 NS_116 0 1.1122841702354280e-05
GC_9_117 b_9 NI_9 NS_117 0 5.8928623430032139e-06
GC_9_118 b_9 NI_9 NS_118 0 1.6678086547024906e-06
GC_9_119 b_9 NI_9 NS_119 0 -1.0738281121528716e-05
GC_9_120 b_9 NI_9 NS_120 0 -6.7127709387204716e-06
GC_9_121 b_9 NI_9 NS_121 0 -5.5359599791114455e-08
GC_9_122 b_9 NI_9 NS_122 0 -2.0704057398251863e-09
GC_9_123 b_9 NI_9 NS_123 0 -1.0037046304438618e-10
GC_9_124 b_9 NI_9 NS_124 0 3.2121632988503290e-10
GC_9_125 b_9 NI_9 NS_125 0 -1.3058224220505718e-05
GC_9_126 b_9 NI_9 NS_126 0 -1.2120478520087456e-05
GC_9_127 b_9 NI_9 NS_127 0 -4.4199314182585291e-05
GC_9_128 b_9 NI_9 NS_128 0 4.2016566311888570e-05
GC_9_129 b_9 NI_9 NS_129 0 4.9656079589274285e-05
GC_9_130 b_9 NI_9 NS_130 0 -4.5266201309794318e-05
GC_9_131 b_9 NI_9 NS_131 0 -1.0660475181430455e-04
GC_9_132 b_9 NI_9 NS_132 0 6.5659091404509479e-05
GC_9_133 b_9 NI_9 NS_133 0 1.2561218749265551e-04
GC_9_134 b_9 NI_9 NS_134 0 -8.6604321284077216e-06
GC_9_135 b_9 NI_9 NS_135 0 -5.8946835208946736e-05
GC_9_136 b_9 NI_9 NS_136 0 4.0870477336001732e-05
GC_9_137 b_9 NI_9 NS_137 0 4.4689993412846754e-05
GC_9_138 b_9 NI_9 NS_138 0 -5.2895351090532065e-06
GC_9_139 b_9 NI_9 NS_139 0 2.5178843789635272e-05
GC_9_140 b_9 NI_9 NS_140 0 3.8247291166327853e-05
GC_9_141 b_9 NI_9 NS_141 0 5.9928608547547549e-08
GC_9_142 b_9 NI_9 NS_142 0 1.3687394720631383e-09
GC_9_143 b_9 NI_9 NS_143 0 1.6472082433167449e-10
GC_9_144 b_9 NI_9 NS_144 0 -6.9445080854302796e-10
GC_9_145 b_9 NI_9 NS_145 0 -9.5337283939971872e-06
GC_9_146 b_9 NI_9 NS_146 0 -5.9434688778598219e-06
GC_9_147 b_9 NI_9 NS_147 0 1.9546600520512794e-06
GC_9_148 b_9 NI_9 NS_148 0 -1.4939358042743400e-05
GC_9_149 b_9 NI_9 NS_149 0 -1.1210928952594424e-04
GC_9_150 b_9 NI_9 NS_150 0 3.7775222738267632e-05
GC_9_151 b_9 NI_9 NS_151 0 -7.9681737954587396e-05
GC_9_152 b_9 NI_9 NS_152 0 7.7640563676732659e-05
GC_9_153 b_9 NI_9 NS_153 0 1.9081247246732487e-04
GC_9_154 b_9 NI_9 NS_154 0 1.3314012598281971e-04
GC_9_155 b_9 NI_9 NS_155 0 5.7036571384641120e-05
GC_9_156 b_9 NI_9 NS_156 0 -1.9615089216589243e-05
GC_9_157 b_9 NI_9 NS_157 0 -5.4481419343213027e-06
GC_9_158 b_9 NI_9 NS_158 0 -8.3263835394805787e-06
GC_9_159 b_9 NI_9 NS_159 0 3.7160519546687136e-05
GC_9_160 b_9 NI_9 NS_160 0 9.7251562597782957e-06
GC_9_161 b_9 NI_9 NS_161 0 -1.6276376620293364e-05
GC_9_162 b_9 NI_9 NS_162 0 -3.6835869170720415e-06
GC_9_163 b_9 NI_9 NS_163 0 -2.2928932851337686e-08
GC_9_164 b_9 NI_9 NS_164 0 -3.8914239545499710e-07
GC_9_165 b_9 NI_9 NS_165 0 4.5530395277775023e-03
GC_9_166 b_9 NI_9 NS_166 0 3.8169598798565539e-03
GC_9_167 b_9 NI_9 NS_167 0 1.3858625682191395e-02
GC_9_168 b_9 NI_9 NS_168 0 -2.1367083898151652e-02
GC_9_169 b_9 NI_9 NS_169 0 -2.2487121893657022e-02
GC_9_170 b_9 NI_9 NS_170 0 2.6079640738487106e-02
GC_9_171 b_9 NI_9 NS_171 0 3.8329041774220064e-02
GC_9_172 b_9 NI_9 NS_172 0 -3.0114596950807260e-02
GC_9_173 b_9 NI_9 NS_173 0 -4.8600024054157434e-02
GC_9_174 b_9 NI_9 NS_174 0 1.9841750849277237e-02
GC_9_175 b_9 NI_9 NS_175 0 2.6998116012690629e-02
GC_9_176 b_9 NI_9 NS_176 0 -1.5909282707089543e-02
GC_9_177 b_9 NI_9 NS_177 0 -1.4330189877374923e-02
GC_9_178 b_9 NI_9 NS_178 0 6.8408587009178463e-03
GC_9_179 b_9 NI_9 NS_179 0 -4.8601514556090011e-03
GC_9_180 b_9 NI_9 NS_180 0 -1.6721195306677868e-02
GC_9_181 b_9 NI_9 NS_181 0 8.9222515767978884e-05
GC_9_182 b_9 NI_9 NS_182 0 3.6749054305357087e-06
GC_9_183 b_9 NI_9 NS_183 0 6.5785375774819149e-09
GC_9_184 b_9 NI_9 NS_184 0 5.9211967668965912e-07
GC_9_185 b_9 NI_9 NS_185 0 4.7462852297715630e-02
GC_9_186 b_9 NI_9 NS_186 0 -9.5881604591076686e-03
GC_9_187 b_9 NI_9 NS_187 0 -4.5650677633938978e-02
GC_9_188 b_9 NI_9 NS_188 0 2.0563545412997535e-02
GC_9_189 b_9 NI_9 NS_189 0 -5.7680593181111878e-02
GC_9_190 b_9 NI_9 NS_190 0 -6.7211170247604049e-02
GC_9_191 b_9 NI_9 NS_191 0 6.3843292984651259e-02
GC_9_192 b_9 NI_9 NS_192 0 -2.1942058420593546e-02
GC_9_193 b_9 NI_9 NS_193 0 2.8542724300669418e-02
GC_9_194 b_9 NI_9 NS_194 0 8.9518934996959440e-02
GC_9_195 b_9 NI_9 NS_195 0 -5.4297954280909277e-02
GC_9_196 b_9 NI_9 NS_196 0 2.8478297858244069e-03
GC_9_197 b_9 NI_9 NS_197 0 -1.3713159769321300e-02
GC_9_198 b_9 NI_9 NS_198 0 -4.7078861173502455e-02
GC_9_199 b_9 NI_9 NS_199 0 1.6430658303161417e-02
GC_9_200 b_9 NI_9 NS_200 0 -3.9060974951704200e-02
GC_9_201 b_9 NI_9 NS_201 0 -1.0355529015791051e-05
GC_9_202 b_9 NI_9 NS_202 0 -2.1274259819667828e-07
GC_9_203 b_9 NI_9 NS_203 0 -1.2832451361410014e-09
GC_9_204 b_9 NI_9 NS_204 0 -2.5390012878609004e-08
GC_9_205 b_9 NI_9 NS_205 0 -4.2497322965482434e-03
GC_9_206 b_9 NI_9 NS_206 0 -3.4927923626545533e-03
GC_9_207 b_9 NI_9 NS_207 0 -1.2922477265220869e-02
GC_9_208 b_9 NI_9 NS_208 0 1.7065692851498011e-02
GC_9_209 b_9 NI_9 NS_209 0 1.7371378434938835e-02
GC_9_210 b_9 NI_9 NS_210 0 -1.9446862252898930e-02
GC_9_211 b_9 NI_9 NS_211 0 -3.3168754961407691e-02
GC_9_212 b_9 NI_9 NS_212 0 2.5454292393380304e-02
GC_9_213 b_9 NI_9 NS_213 0 4.0789565682369619e-02
GC_9_214 b_9 NI_9 NS_214 0 -1.1433259751476585e-02
GC_9_215 b_9 NI_9 NS_215 0 -2.1059403379134214e-02
GC_9_216 b_9 NI_9 NS_216 0 1.5315262612977363e-02
GC_9_217 b_9 NI_9 NS_217 0 1.4123881158377607e-02
GC_9_218 b_9 NI_9 NS_218 0 -3.7536567067230223e-03
GC_9_219 b_9 NI_9 NS_219 0 7.0870161015161538e-03
GC_9_220 b_9 NI_9 NS_220 0 1.3573831691721272e-02
GC_9_221 b_9 NI_9 NS_221 0 -1.8490444357835950e-06
GC_9_222 b_9 NI_9 NS_222 0 2.5677075981751627e-07
GC_9_223 b_9 NI_9 NS_223 0 1.6912982074270045e-09
GC_9_224 b_9 NI_9 NS_224 0 1.3611965998209290e-08
GC_9_225 b_9 NI_9 NS_225 0 1.1406457287261131e-03
GC_9_226 b_9 NI_9 NS_226 0 -2.1726047766020876e-03
GC_9_227 b_9 NI_9 NS_227 0 3.4952389071990068e-03
GC_9_228 b_9 NI_9 NS_228 0 -1.3003077534147438e-02
GC_9_229 b_9 NI_9 NS_229 0 -3.9401362133573800e-02
GC_9_230 b_9 NI_9 NS_230 0 -3.6437965189726785e-04
GC_9_231 b_9 NI_9 NS_231 0 -2.6247364552274215e-02
GC_9_232 b_9 NI_9 NS_232 0 2.8990158451350057e-02
GC_9_233 b_9 NI_9 NS_233 0 5.2202631798501667e-02
GC_9_234 b_9 NI_9 NS_234 0 3.8208679384923068e-02
GC_9_235 b_9 NI_9 NS_235 0 1.7572267409945871e-02
GC_9_236 b_9 NI_9 NS_236 0 -1.4394060190426484e-02
GC_9_237 b_9 NI_9 NS_237 0 -9.1651299739626008e-03
GC_9_238 b_9 NI_9 NS_238 0 -3.7458101634088663e-03
GC_9_239 b_9 NI_9 NS_239 0 8.0623390969349965e-03
GC_9_240 b_9 NI_9 NS_240 0 5.8595893376968784e-03
GD_9_1 b_9 NI_9 NA_1 0 3.1367547041557106e-07
GD_9_2 b_9 NI_9 NA_2 0 -7.7230341600206242e-06
GD_9_3 b_9 NI_9 NA_3 0 -5.2908253988354390e-06
GD_9_4 b_9 NI_9 NA_4 0 1.2166292731830236e-05
GD_9_5 b_9 NI_9 NA_5 0 1.3524373978260853e-05
GD_9_6 b_9 NI_9 NA_6 0 3.0880587850413712e-06
GD_9_7 b_9 NI_9 NA_7 0 2.4223442152152600e-05
GD_9_8 b_9 NI_9 NA_8 0 -5.3839434947247229e-05
GD_9_9 b_9 NI_9 NA_9 0 -9.5852751720691132e-03
GD_9_10 b_9 NI_9 NA_10 0 5.3317556315548775e-03
GD_9_11 b_9 NI_9 NA_11 0 6.7731250245859206e-03
GD_9_12 b_9 NI_9 NA_12 0 -3.3302470009204236e-03
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 -8.0862429425631542e-09
GC_10_2 b_10 NI_10 NS_2 0 6.7986853628853092e-10
GC_10_3 b_10 NI_10 NS_3 0 1.5646926565497410e-11
GC_10_4 b_10 NI_10 NS_4 0 -1.2067899612524435e-10
GC_10_5 b_10 NI_10 NS_5 0 -2.1903676063695700e-06
GC_10_6 b_10 NI_10 NS_6 0 2.1886699250466421e-07
GC_10_7 b_10 NI_10 NS_7 0 -2.1895680331061825e-06
GC_10_8 b_10 NI_10 NS_8 0 2.7884236398782645e-06
GC_10_9 b_10 NI_10 NS_9 0 -1.1327160790076451e-06
GC_10_10 b_10 NI_10 NS_10 0 6.5773519729230505e-06
GC_10_11 b_10 NI_10 NS_11 0 -4.1805333405201739e-07
GC_10_12 b_10 NI_10 NS_12 0 2.1422226419866412e-06
GC_10_13 b_10 NI_10 NS_13 0 7.2190723247341023e-06
GC_10_14 b_10 NI_10 NS_14 0 5.1224739287487711e-06
GC_10_15 b_10 NI_10 NS_15 0 1.6120642164153096e-06
GC_10_16 b_10 NI_10 NS_16 0 3.1394825979609483e-06
GC_10_17 b_10 NI_10 NS_17 0 4.8357474811900809e-06
GC_10_18 b_10 NI_10 NS_18 0 1.1501518584872333e-06
GC_10_19 b_10 NI_10 NS_19 0 2.9137162497862428e-06
GC_10_20 b_10 NI_10 NS_20 0 -1.3217667056904295e-06
GC_10_21 b_10 NI_10 NS_21 0 1.2106842905142488e-08
GC_10_22 b_10 NI_10 NS_22 0 -8.1571308952176727e-10
GC_10_23 b_10 NI_10 NS_23 0 -1.6071025340007973e-11
GC_10_24 b_10 NI_10 NS_24 0 1.3071904809656657e-10
GC_10_25 b_10 NI_10 NS_25 0 7.0579025090415643e-08
GC_10_26 b_10 NI_10 NS_26 0 -1.7341315485362095e-08
GC_10_27 b_10 NI_10 NS_27 0 -5.8731133393872786e-07
GC_10_28 b_10 NI_10 NS_28 0 5.5956800275594364e-07
GC_10_29 b_10 NI_10 NS_29 0 1.6811067354598341e-06
GC_10_30 b_10 NI_10 NS_30 0 -5.0795573744212536e-07
GC_10_31 b_10 NI_10 NS_31 0 -9.8095875690495444e-07
GC_10_32 b_10 NI_10 NS_32 0 1.0424108306403679e-07
GC_10_33 b_10 NI_10 NS_33 0 1.6471581389013903e-06
GC_10_34 b_10 NI_10 NS_34 0 -1.1441249430947431e-06
GC_10_35 b_10 NI_10 NS_35 0 -9.0813486808954271e-07
GC_10_36 b_10 NI_10 NS_36 0 -8.6585053648909310e-07
GC_10_37 b_10 NI_10 NS_37 0 -1.1417344897309673e-06
GC_10_38 b_10 NI_10 NS_38 0 -2.4697839840979059e-07
GC_10_39 b_10 NI_10 NS_39 0 8.7318073965828909e-08
GC_10_40 b_10 NI_10 NS_40 0 1.1733539979702182e-06
GC_10_41 b_10 NI_10 NS_41 0 -5.4818324424450644e-09
GC_10_42 b_10 NI_10 NS_42 0 -1.1901835741469128e-10
GC_10_43 b_10 NI_10 NS_43 0 -8.7994515202676744e-12
GC_10_44 b_10 NI_10 NS_44 0 1.2315176722815721e-11
GC_10_45 b_10 NI_10 NS_45 0 2.8858209527946445e-06
GC_10_46 b_10 NI_10 NS_46 0 -3.3702241853339397e-06
GC_10_47 b_10 NI_10 NS_47 0 3.9410256489470293e-06
GC_10_48 b_10 NI_10 NS_48 0 -1.1989223610866349e-06
GC_10_49 b_10 NI_10 NS_49 0 -1.9642437738130119e-06
GC_10_50 b_10 NI_10 NS_50 0 -6.4802153682235693e-06
GC_10_51 b_10 NI_10 NS_51 0 1.2567712838821434e-06
GC_10_52 b_10 NI_10 NS_52 0 -5.0134047537357725e-06
GC_10_53 b_10 NI_10 NS_53 0 -3.5237884466218855e-06
GC_10_54 b_10 NI_10 NS_54 0 -9.5185268064895474e-06
GC_10_55 b_10 NI_10 NS_55 0 -2.5209703165457264e-06
GC_10_56 b_10 NI_10 NS_56 0 -6.0312516466059491e-06
GC_10_57 b_10 NI_10 NS_57 0 -9.7127112443458909e-06
GC_10_58 b_10 NI_10 NS_58 0 -4.8417680116899474e-06
GC_10_59 b_10 NI_10 NS_59 0 -7.2832288177636864e-06
GC_10_60 b_10 NI_10 NS_60 0 5.3234003849588913e-07
GC_10_61 b_10 NI_10 NS_61 0 -3.3864652711196353e-10
GC_10_62 b_10 NI_10 NS_62 0 2.4529395010533287e-10
GC_10_63 b_10 NI_10 NS_63 0 5.1902605450978487e-12
GC_10_64 b_10 NI_10 NS_64 0 -1.2433837194779225e-11
GC_10_65 b_10 NI_10 NS_65 0 -1.5827626835614125e-06
GC_10_66 b_10 NI_10 NS_66 0 7.4475369233895886e-07
GC_10_67 b_10 NI_10 NS_67 0 -2.4991303777528208e-06
GC_10_68 b_10 NI_10 NS_68 0 1.5671831489314346e-06
GC_10_69 b_10 NI_10 NS_69 0 6.6684086788187250e-07
GC_10_70 b_10 NI_10 NS_70 0 3.1009811147786875e-06
GC_10_71 b_10 NI_10 NS_71 0 -2.4062952941829602e-06
GC_10_72 b_10 NI_10 NS_72 0 3.2308237399731522e-06
GC_10_73 b_10 NI_10 NS_73 0 5.2075167889360714e-06
GC_10_74 b_10 NI_10 NS_74 0 4.2312117521726851e-06
GC_10_75 b_10 NI_10 NS_75 0 -6.0809236297035762e-08
GC_10_76 b_10 NI_10 NS_76 0 3.4339391390181084e-06
GC_10_77 b_10 NI_10 NS_77 0 5.0339042001961214e-06
GC_10_78 b_10 NI_10 NS_78 0 2.2607893633775146e-06
GC_10_79 b_10 NI_10 NS_79 0 3.8677361095028935e-06
GC_10_80 b_10 NI_10 NS_80 0 2.0110296499558791e-07
GC_10_81 b_10 NI_10 NS_81 0 7.1854928984595203e-09
GC_10_82 b_10 NI_10 NS_82 0 2.2479657377056623e-11
GC_10_83 b_10 NI_10 NS_83 0 2.0136707547946319e-11
GC_10_84 b_10 NI_10 NS_84 0 -1.2273208181719761e-10
GC_10_85 b_10 NI_10 NS_85 0 -2.1096712486059104e-06
GC_10_86 b_10 NI_10 NS_86 0 -1.2998927811752803e-06
GC_10_87 b_10 NI_10 NS_87 0 -6.2934660538879975e-06
GC_10_88 b_10 NI_10 NS_88 0 1.3497434156992927e-05
GC_10_89 b_10 NI_10 NS_89 0 3.4249374585142340e-05
GC_10_90 b_10 NI_10 NS_90 0 1.2262959746333759e-05
GC_10_91 b_10 NI_10 NS_91 0 3.1604140904388727e-05
GC_10_92 b_10 NI_10 NS_92 0 -2.5422644597209839e-05
GC_10_93 b_10 NI_10 NS_93 0 -3.9477360525499071e-05
GC_10_94 b_10 NI_10 NS_94 0 -4.7737992460718595e-05
GC_10_95 b_10 NI_10 NS_95 0 -1.9905263090725417e-05
GC_10_96 b_10 NI_10 NS_96 0 1.1122634355785685e-05
GC_10_97 b_10 NI_10 NS_97 0 5.8928113277687483e-06
GC_10_98 b_10 NI_10 NS_98 0 1.6678148716154533e-06
GC_10_99 b_10 NI_10 NS_99 0 -1.0738206206862035e-05
GC_10_100 b_10 NI_10 NS_100 0 -6.7127511662373408e-06
GC_10_101 b_10 NI_10 NS_101 0 -2.7807365128967029e-08
GC_10_102 b_10 NI_10 NS_102 0 8.0981223177863883e-10
GC_10_103 b_10 NI_10 NS_103 0 -1.5187385029306241e-11
GC_10_104 b_10 NI_10 NS_104 0 7.2084451894071040e-11
GC_10_105 b_10 NI_10 NS_105 0 4.1642274389458009e-06
GC_10_106 b_10 NI_10 NS_106 0 2.5912863178490564e-06
GC_10_107 b_10 NI_10 NS_107 0 9.5706831032568584e-06
GC_10_108 b_10 NI_10 NS_108 0 1.0122654099038685e-05
GC_10_109 b_10 NI_10 NS_109 0 1.9377846095135266e-05
GC_10_110 b_10 NI_10 NS_110 0 -2.2684105418625281e-05
GC_10_111 b_10 NI_10 NS_111 0 1.1294700433726763e-05
GC_10_112 b_10 NI_10 NS_112 0 -2.9403254197072107e-06
GC_10_113 b_10 NI_10 NS_113 0 -5.4388625196974942e-06
GC_10_114 b_10 NI_10 NS_114 0 -5.2854993492073391e-05
GC_10_115 b_10 NI_10 NS_115 0 -1.4373071668690942e-05
GC_10_116 b_10 NI_10 NS_116 0 -1.8172894557346663e-05
GC_10_117 b_10 NI_10 NS_117 0 -2.7456964069959592e-05
GC_10_118 b_10 NI_10 NS_118 0 -1.3076036553376653e-05
GC_10_119 b_10 NI_10 NS_119 0 -1.9571260158777062e-05
GC_10_120 b_10 NI_10 NS_120 0 5.5880007596961506e-06
GC_10_121 b_10 NI_10 NS_121 0 5.9902836314631399e-08
GC_10_122 b_10 NI_10 NS_122 0 1.3695854086778263e-09
GC_10_123 b_10 NI_10 NS_123 0 1.6472719510125378e-10
GC_10_124 b_10 NI_10 NS_124 0 -6.9450440199314813e-10
GC_10_125 b_10 NI_10 NS_125 0 -9.5511611120860599e-06
GC_10_126 b_10 NI_10 NS_126 0 -5.9491244688905109e-06
GC_10_127 b_10 NI_10 NS_127 0 1.9276587029548481e-06
GC_10_128 b_10 NI_10 NS_128 0 -1.4956781516650164e-05
GC_10_129 b_10 NI_10 NS_129 0 -1.1212294553213076e-04
GC_10_130 b_10 NI_10 NS_130 0 3.7878409671072394e-05
GC_10_131 b_10 NI_10 NS_131 0 -7.9642075310816429e-05
GC_10_132 b_10 NI_10 NS_132 0 7.7704164508358270e-05
GC_10_133 b_10 NI_10 NS_133 0 1.9090726902570764e-04
GC_10_134 b_10 NI_10 NS_134 0 1.3304677632984438e-04
GC_10_135 b_10 NI_10 NS_135 0 5.7019877806471301e-05
GC_10_136 b_10 NI_10 NS_136 0 -1.9652976749049302e-05
GC_10_137 b_10 NI_10 NS_137 0 -5.4751876055237403e-06
GC_10_138 b_10 NI_10 NS_138 0 -8.3218554711010356e-06
GC_10_139 b_10 NI_10 NS_139 0 3.7156183936561682e-05
GC_10_140 b_10 NI_10 NS_140 0 9.7277836656017786e-06
GC_10_141 b_10 NI_10 NS_141 0 -5.5372264074574203e-08
GC_10_142 b_10 NI_10 NS_142 0 -2.0698405003956447e-09
GC_10_143 b_10 NI_10 NS_143 0 -1.0036913013043493e-10
GC_10_144 b_10 NI_10 NS_144 0 3.2118675094755313e-10
GC_10_145 b_10 NI_10 NS_145 0 -1.3057977126047742e-05
GC_10_146 b_10 NI_10 NS_146 0 -1.2121355181200021e-05
GC_10_147 b_10 NI_10 NS_147 0 -4.4199162340438443e-05
GC_10_148 b_10 NI_10 NS_148 0 4.2015911170957170e-05
GC_10_149 b_10 NI_10 NS_149 0 4.9655942058050381e-05
GC_10_150 b_10 NI_10 NS_150 0 -4.5267462078757824e-05
GC_10_151 b_10 NI_10 NS_151 0 -1.0660547794756488e-04
GC_10_152 b_10 NI_10 NS_152 0 6.5657554411257732e-05
GC_10_153 b_10 NI_10 NS_153 0 1.2561071358901135e-04
GC_10_154 b_10 NI_10 NS_154 0 -8.6598571144387529e-06
GC_10_155 b_10 NI_10 NS_155 0 -5.8946727886662037e-05
GC_10_156 b_10 NI_10 NS_156 0 4.0869753509480727e-05
GC_10_157 b_10 NI_10 NS_157 0 4.4689150976666890e-05
GC_10_158 b_10 NI_10 NS_158 0 -5.2904242922244085e-06
GC_10_159 b_10 NI_10 NS_159 0 2.5177398627135203e-05
GC_10_160 b_10 NI_10 NS_160 0 3.8246853529692717e-05
GC_10_161 b_10 NI_10 NS_161 0 8.9222421995792891e-05
GC_10_162 b_10 NI_10 NS_162 0 3.6749130943961404e-06
GC_10_163 b_10 NI_10 NS_163 0 6.5786627378165616e-09
GC_10_164 b_10 NI_10 NS_164 0 5.9211886052560896e-07
GC_10_165 b_10 NI_10 NS_165 0 4.7462886305466585e-02
GC_10_166 b_10 NI_10 NS_166 0 -9.5881530848590107e-03
GC_10_167 b_10 NI_10 NS_167 0 -4.5650646954405197e-02
GC_10_168 b_10 NI_10 NS_168 0 2.0563576409542247e-02
GC_10_169 b_10 NI_10 NS_169 0 -5.7680547906318907e-02
GC_10_170 b_10 NI_10 NS_170 0 -6.7211344845207646e-02
GC_10_171 b_10 NI_10 NS_171 0 6.3843232630716604e-02
GC_10_172 b_10 NI_10 NS_172 0 -2.1942168262716683e-02
GC_10_173 b_10 NI_10 NS_173 0 2.8542542012470567e-02
GC_10_174 b_10 NI_10 NS_174 0 8.9519059621235186e-02
GC_10_175 b_10 NI_10 NS_175 0 -5.4297950706615382e-02
GC_10_176 b_10 NI_10 NS_176 0 2.8479068636053937e-03
GC_10_177 b_10 NI_10 NS_177 0 -1.3713099434847276e-02
GC_10_178 b_10 NI_10 NS_178 0 -4.7078848912118477e-02
GC_10_179 b_10 NI_10 NS_179 0 1.6430669201775220e-02
GC_10_180 b_10 NI_10 NS_180 0 -3.9060986660119278e-02
GC_10_181 b_10 NI_10 NS_181 0 -1.6276376620293679e-05
GC_10_182 b_10 NI_10 NS_182 0 -3.6835869170718272e-06
GC_10_183 b_10 NI_10 NS_183 0 -2.2928932851337957e-08
GC_10_184 b_10 NI_10 NS_184 0 -3.8914239545499371e-07
GC_10_185 b_10 NI_10 NS_185 0 4.5530395277774659e-03
GC_10_186 b_10 NI_10 NS_186 0 3.8169598798565448e-03
GC_10_187 b_10 NI_10 NS_187 0 1.3858625682191388e-02
GC_10_188 b_10 NI_10 NS_188 0 -2.1367083898151652e-02
GC_10_189 b_10 NI_10 NS_189 0 -2.2487121893657057e-02
GC_10_190 b_10 NI_10 NS_190 0 2.6079640738487151e-02
GC_10_191 b_10 NI_10 NS_191 0 3.8329041774220071e-02
GC_10_192 b_10 NI_10 NS_192 0 -3.0114596950807253e-02
GC_10_193 b_10 NI_10 NS_193 0 -4.8600024054157420e-02
GC_10_194 b_10 NI_10 NS_194 0 1.9841750849277275e-02
GC_10_195 b_10 NI_10 NS_195 0 2.6998116012690646e-02
GC_10_196 b_10 NI_10 NS_196 0 -1.5909282707089547e-02
GC_10_197 b_10 NI_10 NS_197 0 -1.4330189877374916e-02
GC_10_198 b_10 NI_10 NS_198 0 6.8408587009178515e-03
GC_10_199 b_10 NI_10 NS_199 0 -4.8601514556089881e-03
GC_10_200 b_10 NI_10 NS_200 0 -1.6721195306677868e-02
GC_10_201 b_10 NI_10 NS_201 0 -1.8490440325849337e-06
GC_10_202 b_10 NI_10 NS_202 0 2.5677074895948616e-07
GC_10_203 b_10 NI_10 NS_203 0 1.6912978857590798e-09
GC_10_204 b_10 NI_10 NS_204 0 1.3611966836481582e-08
GC_10_205 b_10 NI_10 NS_205 0 1.1406456014744885e-03
GC_10_206 b_10 NI_10 NS_206 0 -2.1726046681587005e-03
GC_10_207 b_10 NI_10 NS_207 0 3.4952388266333233e-03
GC_10_208 b_10 NI_10 NS_208 0 -1.3003077401551761e-02
GC_10_209 b_10 NI_10 NS_209 0 -3.9401362128267073e-02
GC_10_210 b_10 NI_10 NS_210 0 -3.6437949506928485e-04
GC_10_211 b_10 NI_10 NS_211 0 -2.6247364684288919e-02
GC_10_212 b_10 NI_10 NS_212 0 2.8990158567300840e-02
GC_10_213 b_10 NI_10 NS_213 0 5.2202632001435427e-02
GC_10_214 b_10 NI_10 NS_214 0 3.8208679920845603e-02
GC_10_215 b_10 NI_10 NS_215 0 1.7572267604284250e-02
GC_10_216 b_10 NI_10 NS_216 0 -1.4394059928293807e-02
GC_10_217 b_10 NI_10 NS_217 0 -9.1651296143751542e-03
GC_10_218 b_10 NI_10 NS_218 0 -3.7458101137161429e-03
GC_10_219 b_10 NI_10 NS_219 0 8.0623393113781906e-03
GC_10_220 b_10 NI_10 NS_220 0 5.8595892994051293e-03
GC_10_221 b_10 NI_10 NS_221 0 -1.0356264724050639e-05
GC_10_222 b_10 NI_10 NS_222 0 -2.1272066910781319e-07
GC_10_223 b_10 NI_10 NS_223 0 -1.2831318769616312e-09
GC_10_224 b_10 NI_10 NS_224 0 -2.5390349103913194e-08
GC_10_225 b_10 NI_10 NS_225 0 -4.2497282974039595e-03
GC_10_226 b_10 NI_10 NS_226 0 -3.4927765861530180e-03
GC_10_227 b_10 NI_10 NS_227 0 -1.2922365284355081e-02
GC_10_228 b_10 NI_10 NS_228 0 1.7065796242937883e-02
GC_10_229 b_10 NI_10 NS_229 0 1.7371354068310418e-02
GC_10_230 b_10 NI_10 NS_230 0 -1.9447062281415850e-02
GC_10_231 b_10 NI_10 NS_231 0 -3.3168706673441066e-02
GC_10_232 b_10 NI_10 NS_232 0 2.5454422060204401e-02
GC_10_233 b_10 NI_10 NS_233 0 4.0789606324396155e-02
GC_10_234 b_10 NI_10 NS_234 0 -1.1433470216096055e-02
GC_10_235 b_10 NI_10 NS_235 0 -2.1059355324638526e-02
GC_10_236 b_10 NI_10 NS_236 0 1.5315260980555735e-02
GC_10_237 b_10 NI_10 NS_237 0 1.4123842999471408e-02
GC_10_238 b_10 NI_10 NS_238 0 -3.7538559430493365e-03
GC_10_239 b_10 NI_10 NS_239 0 7.0868356914228353e-03
GC_10_240 b_10 NI_10 NS_240 0 1.3573780069431456e-02
GD_10_1 b_10 NI_10 NA_1 0 -7.7230405332677081e-06
GD_10_2 b_10 NI_10 NA_2 0 3.3803646505013203e-07
GD_10_3 b_10 NI_10 NA_3 0 1.2163791812448901e-05
GD_10_4 b_10 NI_10 NA_4 0 -5.2908402516629234e-06
GD_10_5 b_10 NI_10 NA_5 0 3.0875889695450648e-06
GD_10_6 b_10 NI_10 NA_6 0 1.3910656666057643e-05
GD_10_7 b_10 NI_10 NA_7 0 -5.3853458210282143e-05
GD_10_8 b_10 NI_10 NA_8 0 2.4227204553939678e-05
GD_10_9 b_10 NI_10 NA_9 0 5.3317874208177818e-03
GD_10_10 b_10 NI_10 NA_10 0 -9.5852751720690212e-03
GD_10_11 b_10 NI_10 NA_11 0 -3.3302474407708280e-03
GD_10_12 b_10 NI_10 NA_12 0 6.7730078664015488e-03
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 2.2395738343677488e-09
GC_11_2 b_11 NI_11 NS_2 0 -6.1558476047547845e-11
GC_11_3 b_11 NI_11 NS_3 0 -1.4861658374094376e-12
GC_11_4 b_11 NI_11 NS_4 0 1.6503249921698269e-11
GC_11_5 b_11 NI_11 NS_5 0 -5.6363583213756244e-07
GC_11_6 b_11 NI_11 NS_6 0 4.0935474549865688e-07
GC_11_7 b_11 NI_11 NS_7 0 -2.8794740970991849e-07
GC_11_8 b_11 NI_11 NS_8 0 1.5345561224319849e-06
GC_11_9 b_11 NI_11 NS_9 0 7.1637558426986786e-07
GC_11_10 b_11 NI_11 NS_10 0 -5.3803630323437651e-07
GC_11_11 b_11 NI_11 NS_11 0 -5.0822709272192711e-07
GC_11_12 b_11 NI_11 NS_12 0 2.2103913740334615e-06
GC_11_13 b_11 NI_11 NS_13 0 2.2909581102689927e-06
GC_11_14 b_11 NI_11 NS_14 0 -1.4800636805869496e-06
GC_11_15 b_11 NI_11 NS_15 0 -7.8891771318784974e-07
GC_11_16 b_11 NI_11 NS_16 0 9.3936125386882881e-07
GC_11_17 b_11 NI_11 NS_17 0 8.4703247342769325e-07
GC_11_18 b_11 NI_11 NS_18 0 7.6963402416810992e-08
GC_11_19 b_11 NI_11 NS_19 0 7.2183054273667128e-07
GC_11_20 b_11 NI_11 NS_20 0 5.7000287097420042e-07
GC_11_21 b_11 NI_11 NS_21 0 -1.1015623704594474e-09
GC_11_22 b_11 NI_11 NS_22 0 -2.6549909328046467e-11
GC_11_23 b_11 NI_11 NS_23 0 -5.3034250402839469e-13
GC_11_24 b_11 NI_11 NS_24 0 -6.8049911445173450e-12
GC_11_25 b_11 NI_11 NS_25 0 -5.8840407325761900e-08
GC_11_26 b_11 NI_11 NS_26 0 -6.1578153394293002e-07
GC_11_27 b_11 NI_11 NS_27 0 -3.4130239288733140e-07
GC_11_28 b_11 NI_11 NS_28 0 -1.0123479225734651e-07
GC_11_29 b_11 NI_11 NS_29 0 -1.1029926730503831e-06
GC_11_30 b_11 NI_11 NS_30 0 1.5334424956307699e-06
GC_11_31 b_11 NI_11 NS_31 0 6.9658915384646699e-07
GC_11_32 b_11 NI_11 NS_32 0 8.5933532703793078e-07
GC_11_33 b_11 NI_11 NS_33 0 2.1615732983857669e-06
GC_11_34 b_11 NI_11 NS_34 0 -1.4800253009785432e-06
GC_11_35 b_11 NI_11 NS_35 0 -1.9795090989705576e-07
GC_11_36 b_11 NI_11 NS_36 0 -9.9053898808474952e-07
GC_11_37 b_11 NI_11 NS_37 0 -1.0678572701212045e-06
GC_11_38 b_11 NI_11 NS_38 0 -4.1564945858280948e-07
GC_11_39 b_11 NI_11 NS_39 0 -4.0950167754025826e-07
GC_11_40 b_11 NI_11 NS_40 0 1.2021649037414041e-07
GC_11_41 b_11 NI_11 NS_41 0 1.2124745556995733e-08
GC_11_42 b_11 NI_11 NS_42 0 -8.1682186850862606e-10
GC_11_43 b_11 NI_11 NS_43 0 -1.6082074221028918e-11
GC_11_44 b_11 NI_11 NS_44 0 1.3082088109253331e-10
GC_11_45 b_11 NI_11 NS_45 0 7.0237185005250259e-08
GC_11_46 b_11 NI_11 NS_46 0 -1.5046103959732042e-08
GC_11_47 b_11 NI_11 NS_47 0 -5.8773509465538331e-07
GC_11_48 b_11 NI_11 NS_48 0 5.5728452394883659e-07
GC_11_49 b_11 NI_11 NS_49 0 1.6792028947161364e-06
GC_11_50 b_11 NI_11 NS_50 0 -4.9983203933124169e-07
GC_11_51 b_11 NI_11 NS_51 0 -9.7806804612696847e-07
GC_11_52 b_11 NI_11 NS_52 0 1.0430318477577697e-07
GC_11_53 b_11 NI_11 NS_53 0 1.6496851442707612e-06
GC_11_54 b_11 NI_11 NS_54 0 -1.1404223409920525e-06
GC_11_55 b_11 NI_11 NS_55 0 -9.0614266959089292e-07
GC_11_56 b_11 NI_11 NS_56 0 -8.6662758942946901e-07
GC_11_57 b_11 NI_11 NS_57 0 -1.1401325009421186e-06
GC_11_58 b_11 NI_11 NS_58 0 -2.4471837740874721e-07
GC_11_59 b_11 NI_11 NS_59 0 8.9532514154139703e-08
GC_11_60 b_11 NI_11 NS_60 0 1.1724104597568607e-06
GC_11_61 b_11 NI_11 NS_61 0 -8.0831916955979319e-09
GC_11_62 b_11 NI_11 NS_62 0 6.7951718459366812e-10
GC_11_63 b_11 NI_11 NS_63 0 1.5642918129532941e-11
GC_11_64 b_11 NI_11 NS_64 0 -1.2064089991393890e-10
GC_11_65 b_11 NI_11 NS_65 0 -2.1882725000884367e-06
GC_11_66 b_11 NI_11 NS_66 0 2.1734556172316175e-07
GC_11_67 b_11 NI_11 NS_67 0 -2.1912527686827508e-06
GC_11_68 b_11 NI_11 NS_68 0 2.7906333782337800e-06
GC_11_69 b_11 NI_11 NS_69 0 -1.1302476646992286e-06
GC_11_70 b_11 NI_11 NS_70 0 6.5760335640018249e-06
GC_11_71 b_11 NI_11 NS_71 0 -4.1809912937988589e-07
GC_11_72 b_11 NI_11 NS_72 0 2.1387822117820339e-06
GC_11_73 b_11 NI_11 NS_73 0 7.2163470227411025e-06
GC_11_74 b_11 NI_11 NS_74 0 5.1185250623867466e-06
GC_11_75 b_11 NI_11 NS_75 0 1.6097748600473306e-06
GC_11_76 b_11 NI_11 NS_76 0 3.1433818307163161e-06
GC_11_77 b_11 NI_11 NS_77 0 4.8364251853179645e-06
GC_11_78 b_11 NI_11 NS_78 0 1.1505215892388850e-06
GC_11_79 b_11 NI_11 NS_79 0 2.9136123734502448e-06
GC_11_80 b_11 NI_11 NS_80 0 -1.3226687332598515e-06
GC_11_81 b_11 NI_11 NS_81 0 2.0768895667569918e-08
GC_11_82 b_11 NI_11 NS_82 0 -1.0266109490189834e-09
GC_11_83 b_11 NI_11 NS_83 0 -1.9426111434699114e-11
GC_11_84 b_11 NI_11 NS_84 0 1.5749234171268774e-10
GC_11_85 b_11 NI_11 NS_85 0 -1.1217130347970750e-06
GC_11_86 b_11 NI_11 NS_86 0 -8.1021153432838907e-07
GC_11_87 b_11 NI_11 NS_87 0 -2.0037373811811460e-06
GC_11_88 b_11 NI_11 NS_88 0 3.5848970353834649e-08
GC_11_89 b_11 NI_11 NS_89 0 -3.0743118329312175e-06
GC_11_90 b_11 NI_11 NS_90 0 8.6171731281222673e-07
GC_11_91 b_11 NI_11 NS_91 0 -4.1502960449123667e-06
GC_11_92 b_11 NI_11 NS_92 0 4.3114704550708062e-06
GC_11_93 b_11 NI_11 NS_93 0 3.3134004680986720e-06
GC_11_94 b_11 NI_11 NS_94 0 5.4284204535535411e-06
GC_11_95 b_11 NI_11 NS_95 0 -8.9968139539892171e-07
GC_11_96 b_11 NI_11 NS_96 0 5.9726067275538619e-06
GC_11_97 b_11 NI_11 NS_97 0 6.0570612853233583e-06
GC_11_98 b_11 NI_11 NS_98 0 3.3263267045521445e-06
GC_11_99 b_11 NI_11 NS_99 0 5.8639217214175510e-06
GC_11_100 b_11 NI_11 NS_100 0 1.7029362831189067e-06
GC_11_101 b_11 NI_11 NS_101 0 -2.4099524019331689e-08
GC_11_102 b_11 NI_11 NS_102 0 1.2312867652762508e-09
GC_11_103 b_11 NI_11 NS_103 0 2.1599268163163194e-11
GC_11_104 b_11 NI_11 NS_104 0 -1.7722969911922579e-10
GC_11_105 b_11 NI_11 NS_105 0 1.8333069647984085e-06
GC_11_106 b_11 NI_11 NS_106 0 -4.1855572864766310e-06
GC_11_107 b_11 NI_11 NS_107 0 2.4443895867784114e-06
GC_11_108 b_11 NI_11 NS_108 0 7.5715890058606818e-08
GC_11_109 b_11 NI_11 NS_109 0 -1.6176201312295375e-06
GC_11_110 b_11 NI_11 NS_110 0 -4.3834838139503211e-06
GC_11_111 b_11 NI_11 NS_111 0 1.0020625871023608e-06
GC_11_112 b_11 NI_11 NS_112 0 -7.2532088098346539e-06
GC_11_113 b_11 NI_11 NS_113 0 -8.7087199478208018e-06
GC_11_114 b_11 NI_11 NS_114 0 -4.7028282904740683e-06
GC_11_115 b_11 NI_11 NS_115 0 -3.2786364004082251e-06
GC_11_116 b_11 NI_11 NS_116 0 1.3949526537140679e-06
GC_11_117 b_11 NI_11 NS_117 0 -1.9194172549351789e-06
GC_11_118 b_11 NI_11 NS_118 0 -5.4219261060331632e-07
GC_11_119 b_11 NI_11 NS_119 0 -3.2888257473440780e-06
GC_11_120 b_11 NI_11 NS_120 0 -1.5163214527416041e-06
GC_11_121 b_11 NI_11 NS_121 0 -2.5925745127603500e-08
GC_11_122 b_11 NI_11 NS_122 0 1.1529335398274651e-09
GC_11_123 b_11 NI_11 NS_123 0 -1.0993192444707395e-11
GC_11_124 b_11 NI_11 NS_124 0 3.1284423661570616e-11
GC_11_125 b_11 NI_11 NS_125 0 4.4658844035384920e-06
GC_11_126 b_11 NI_11 NS_126 0 2.2626212029459831e-06
GC_11_127 b_11 NI_11 NS_127 0 9.9229978114461097e-06
GC_11_128 b_11 NI_11 NS_128 0 9.6721828936730693e-06
GC_11_129 b_11 NI_11 NS_129 0 1.8821990151604254e-05
GC_11_130 b_11 NI_11 NS_130 0 -2.3464206978695570e-05
GC_11_131 b_11 NI_11 NS_131 0 1.1213140567439407e-05
GC_11_132 b_11 NI_11 NS_132 0 -3.3843358572877514e-06
GC_11_133 b_11 NI_11 NS_133 0 -6.7473937484409067e-06
GC_11_134 b_11 NI_11 NS_134 0 -5.3021724455831431e-05
GC_11_135 b_11 NI_11 NS_135 0 -1.4872212726895500e-05
GC_11_136 b_11 NI_11 NS_136 0 -1.7984609424269335e-05
GC_11_137 b_11 NI_11 NS_137 0 -2.7699453003828182e-05
GC_11_138 b_11 NI_11 NS_138 0 -1.2430480343366660e-05
GC_11_139 b_11 NI_11 NS_139 0 -1.9111947397054776e-05
GC_11_140 b_11 NI_11 NS_140 0 5.9354256697731410e-06
GC_11_141 b_11 NI_11 NS_141 0 1.1016561122603096e-09
GC_11_142 b_11 NI_11 NS_142 0 -1.2971191919709161e-10
GC_11_143 b_11 NI_11 NS_143 0 1.7862379697115573e-11
GC_11_144 b_11 NI_11 NS_144 0 -9.6106570732850838e-11
GC_11_145 b_11 NI_11 NS_145 0 -1.9128838357417402e-06
GC_11_146 b_11 NI_11 NS_146 0 -1.1371208884424316e-06
GC_11_147 b_11 NI_11 NS_147 0 -6.0331199268242744e-06
GC_11_148 b_11 NI_11 NS_148 0 1.3796847501518855e-05
GC_11_149 b_11 NI_11 NS_149 0 3.5155088732053217e-05
GC_11_150 b_11 NI_11 NS_150 0 1.1739874487382219e-05
GC_11_151 b_11 NI_11 NS_151 0 3.2374480867563567e-05
GC_11_152 b_11 NI_11 NS_152 0 -2.5607924312700215e-05
GC_11_153 b_11 NI_11 NS_153 0 -3.9768424582202082e-05
GC_11_154 b_11 NI_11 NS_154 0 -4.9607872925322454e-05
GC_11_155 b_11 NI_11 NS_155 0 -1.9812838261914891e-05
GC_11_156 b_11 NI_11 NS_156 0 1.0190725540275987e-05
GC_11_157 b_11 NI_11 NS_157 0 4.9362497903320495e-06
GC_11_158 b_11 NI_11 NS_158 0 3.9503240476232038e-07
GC_11_159 b_11 NI_11 NS_159 0 -1.2398818152153722e-05
GC_11_160 b_11 NI_11 NS_160 0 -7.1395543002243443e-06
GC_11_161 b_11 NI_11 NS_161 0 -1.0356264724048311e-05
GC_11_162 b_11 NI_11 NS_162 0 -2.1272066910863974e-07
GC_11_163 b_11 NI_11 NS_163 0 -1.2831318769650057e-09
GC_11_164 b_11 NI_11 NS_164 0 -2.5390349103888902e-08
GC_11_165 b_11 NI_11 NS_165 0 -4.2497282974039464e-03
GC_11_166 b_11 NI_11 NS_166 0 -3.4927765861530367e-03
GC_11_167 b_11 NI_11 NS_167 0 -1.2922365284355097e-02
GC_11_168 b_11 NI_11 NS_168 0 1.7065796242937876e-02
GC_11_169 b_11 NI_11 NS_169 0 1.7371354068310436e-02
GC_11_170 b_11 NI_11 NS_170 0 -1.9447062281415871e-02
GC_11_171 b_11 NI_11 NS_171 0 -3.3168706673441066e-02
GC_11_172 b_11 NI_11 NS_172 0 2.5454422060204387e-02
GC_11_173 b_11 NI_11 NS_173 0 4.0789606324396113e-02
GC_11_174 b_11 NI_11 NS_174 0 -1.1433470216096073e-02
GC_11_175 b_11 NI_11 NS_175 0 -2.1059355324638523e-02
GC_11_176 b_11 NI_11 NS_176 0 1.5315260980555714e-02
GC_11_177 b_11 NI_11 NS_177 0 1.4123842999471371e-02
GC_11_178 b_11 NI_11 NS_178 0 -3.7538559430493530e-03
GC_11_179 b_11 NI_11 NS_179 0 7.0868356914228110e-03
GC_11_180 b_11 NI_11 NS_180 0 1.3573780069431454e-02
GC_11_181 b_11 NI_11 NS_181 0 -1.8490444358048100e-06
GC_11_182 b_11 NI_11 NS_182 0 2.5677075982013329e-07
GC_11_183 b_11 NI_11 NS_183 0 1.6912982073973982e-09
GC_11_184 b_11 NI_11 NS_184 0 1.3611965998259831e-08
GC_11_185 b_11 NI_11 NS_185 0 1.1406457287262612e-03
GC_11_186 b_11 NI_11 NS_186 0 -2.1726047766017975e-03
GC_11_187 b_11 NI_11 NS_187 0 3.4952389072004774e-03
GC_11_188 b_11 NI_11 NS_188 0 -1.3003077534147230e-02
GC_11_189 b_11 NI_11 NS_189 0 -3.9401362133573939e-02
GC_11_190 b_11 NI_11 NS_190 0 -3.6437965189990332e-04
GC_11_191 b_11 NI_11 NS_191 0 -2.6247364552274995e-02
GC_11_192 b_11 NI_11 NS_192 0 2.8990158451349730e-02
GC_11_193 b_11 NI_11 NS_193 0 5.2202631798501424e-02
GC_11_194 b_11 NI_11 NS_194 0 3.8208679384921937e-02
GC_11_195 b_11 NI_11 NS_195 0 1.7572267409945067e-02
GC_11_196 b_11 NI_11 NS_196 0 -1.4394060190427067e-02
GC_11_197 b_11 NI_11 NS_197 0 -9.1651299739631872e-03
GC_11_198 b_11 NI_11 NS_198 0 -3.7458101634095698e-03
GC_11_199 b_11 NI_11 NS_199 0 8.0623390969336746e-03
GC_11_200 b_11 NI_11 NS_200 0 5.8595893376966234e-03
GC_11_201 b_11 NI_11 NS_201 0 -1.5427135100829775e-05
GC_11_202 b_11 NI_11 NS_202 0 -3.7324314362845172e-06
GC_11_203 b_11 NI_11 NS_203 0 -2.3081208540648690e-08
GC_11_204 b_11 NI_11 NS_204 0 -3.8674152064337953e-07
GC_11_205 b_11 NI_11 NS_205 0 4.5760065486724890e-03
GC_11_206 b_11 NI_11 NS_206 0 3.7993286749984792e-03
GC_11_207 b_11 NI_11 NS_207 0 1.3872401194724840e-02
GC_11_208 b_11 NI_11 NS_208 0 -2.1406272357366678e-02
GC_11_209 b_11 NI_11 NS_209 0 -2.2493840892053685e-02
GC_11_210 b_11 NI_11 NS_210 0 2.6058892794354329e-02
GC_11_211 b_11 NI_11 NS_211 0 3.8337056260354004e-02
GC_11_212 b_11 NI_11 NS_212 0 -3.0181707200149149e-02
GC_11_213 b_11 NI_11 NS_213 0 -4.8685823046150975e-02
GC_11_214 b_11 NI_11 NS_214 0 1.9831379025888919e-02
GC_11_215 b_11 NI_11 NS_215 0 2.6967890269789584e-02
GC_11_216 b_11 NI_11 NS_216 0 -1.5945601277777981e-02
GC_11_217 b_11 NI_11 NS_217 0 -1.4394992355179019e-02
GC_11_218 b_11 NI_11 NS_218 0 6.8900417725550646e-03
GC_11_219 b_11 NI_11 NS_219 0 -4.8273798937391614e-03
GC_11_220 b_11 NI_11 NS_220 0 -1.6678597174828426e-02
GC_11_221 b_11 NI_11 NS_221 0 8.9998716174948435e-05
GC_11_222 b_11 NI_11 NS_222 0 3.6211880582123379e-06
GC_11_223 b_11 NI_11 NS_223 0 5.9682499092563400e-09
GC_11_224 b_11 NI_11 NS_224 0 5.9667511698087758e-07
GC_11_225 b_11 NI_11 NS_225 0 4.7508862642063471e-02
GC_11_226 b_11 NI_11 NS_226 0 -9.6471114695072090e-03
GC_11_227 b_11 NI_11 NS_227 0 -4.5582913306079817e-02
GC_11_228 b_11 NI_11 NS_228 0 2.0552304035070239e-02
GC_11_229 b_11 NI_11 NS_229 0 -5.7696866703446030e-02
GC_11_230 b_11 NI_11 NS_230 0 -6.7350313493443684e-02
GC_11_231 b_11 NI_11 NS_231 0 6.3862089875377726e-02
GC_11_232 b_11 NI_11 NS_232 0 -2.2063742598215173e-02
GC_11_233 b_11 NI_11 NS_233 0 2.8382264866129117e-02
GC_11_234 b_11 NI_11 NS_234 0 8.9387902159478241e-02
GC_11_235 b_11 NI_11 NS_235 0 -5.4366410708933430e-02
GC_11_236 b_11 NI_11 NS_236 0 2.7979819975819244e-03
GC_11_237 b_11 NI_11 NS_237 0 -1.3847781195743720e-02
GC_11_238 b_11 NI_11 NS_238 0 -4.7095076153860223e-02
GC_11_239 b_11 NI_11 NS_239 0 1.6380419252626524e-02
GC_11_240 b_11 NI_11 NS_240 0 -3.9016261544321161e-02
GD_11_1 b_11 NI_11 NA_1 0 -1.5460811934903774e-06
GD_11_2 b_11 NI_11 NA_2 0 3.4772172746934404e-07
GD_11_3 b_11 NI_11 NA_3 0 3.3057317500745035e-07
GD_11_4 b_11 NI_11 NA_4 0 -7.7232170305271223e-06
GD_11_5 b_11 NI_11 NA_5 0 -1.1644152972350560e-06
GD_11_6 b_11 NI_11 NA_6 0 1.0083328886852959e-05
GD_11_7 b_11 NI_11 NA_7 0 1.5099444170113518e-05
GD_11_8 b_11 NI_11 NA_8 0 3.3225507644304590e-06
GD_11_9 b_11 NI_11 NA_9 0 6.7730078664016286e-03
GD_11_10 b_11 NI_11 NA_10 0 -3.3302470009183077e-03
GD_11_11 b_11 NI_11 NA_11 0 -9.5068691426405533e-03
GD_11_12 b_11 NI_11 NA_12 0 5.5525421417793874e-03
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -1.1046906440981123e-09
GC_12_2 b_12 NI_12 NS_2 0 -2.6299755093010511e-11
GC_12_3 b_12 NI_12 NS_3 0 -5.2636187210249694e-13
GC_12_4 b_12 NI_12 NS_4 0 -6.8309082363625461e-12
GC_12_5 b_12 NI_12 NS_5 0 -5.6996025020906859e-08
GC_12_6 b_12 NI_12 NS_6 0 -6.1544886072464830e-07
GC_12_7 b_12 NI_12 NS_7 0 -3.3915803365226771e-07
GC_12_8 b_12 NI_12 NS_8 0 -9.9907673970843927e-08
GC_12_9 b_12 NI_12 NS_9 0 -1.1012113680797633e-06
GC_12_10 b_12 NI_12 NS_10 0 1.5244122405969686e-06
GC_12_11 b_12 NI_12 NS_11 0 6.9375546872322093e-07
GC_12_12 b_12 NI_12 NS_12 0 8.5371702533888434e-07
GC_12_13 b_12 NI_12 NS_13 0 2.1527505059997690e-06
GC_12_14 b_12 NI_12 NS_14 0 -1.4740997862130439e-06
GC_12_15 b_12 NI_12 NS_15 0 -1.9736969920695288e-07
GC_12_16 b_12 NI_12 NS_16 0 -9.8761886623425301e-07
GC_12_17 b_12 NI_12 NS_17 0 -1.0659942557986130e-06
GC_12_18 b_12 NI_12 NS_18 0 -4.1594097543504030e-07
GC_12_19 b_12 NI_12 NS_19 0 -4.0970861873034791e-07
GC_12_20 b_12 NI_12 NS_20 0 1.1981970866248892e-07
GC_12_21 b_12 NI_12 NS_21 0 2.2396167113473174e-09
GC_12_22 b_12 NI_12 NS_22 0 -6.1561128763768491e-11
GC_12_23 b_12 NI_12 NS_23 0 -1.4862083830941954e-12
GC_12_24 b_12 NI_12 NS_24 0 1.6503540031658315e-11
GC_12_25 b_12 NI_12 NS_25 0 -5.6364936760525864e-07
GC_12_26 b_12 NI_12 NS_26 0 4.0935839248077542e-07
GC_12_27 b_12 NI_12 NS_27 0 -2.8795956868861392e-07
GC_12_28 b_12 NI_12 NS_28 0 1.5345503766143033e-06
GC_12_29 b_12 NI_12 NS_29 0 7.1636293599735773e-07
GC_12_30 b_12 NI_12 NS_30 0 -5.3800506682514607e-07
GC_12_31 b_12 NI_12 NS_31 0 -5.0824261669073087e-07
GC_12_32 b_12 NI_12 NS_32 0 2.2104029143316395e-06
GC_12_33 b_12 NI_12 NS_33 0 2.2909991570676821e-06
GC_12_34 b_12 NI_12 NS_34 0 -1.4800224857008827e-06
GC_12_35 b_12 NI_12 NS_35 0 -7.8890911287081858e-07
GC_12_36 b_12 NI_12 NS_36 0 9.3935839661420669e-07
GC_12_37 b_12 NI_12 NS_37 0 8.4704644890086722e-07
GC_12_38 b_12 NI_12 NS_38 0 7.6970670324237981e-08
GC_12_39 b_12 NI_12 NS_39 0 7.2184164606210784e-07
GC_12_40 b_12 NI_12 NS_40 0 5.7000025669550418e-07
GC_12_41 b_12 NI_12 NS_41 0 -8.0831969364444200e-09
GC_12_42 b_12 NI_12 NS_42 0 6.7951745087779999e-10
GC_12_43 b_12 NI_12 NS_43 0 1.5642919002214455e-11
GC_12_44 b_12 NI_12 NS_44 0 -1.2064091411708442e-10
GC_12_45 b_12 NI_12 NS_45 0 -2.1882726311756117e-06
GC_12_46 b_12 NI_12 NS_46 0 2.1734101965580886e-07
GC_12_47 b_12 NI_12 NS_47 0 -2.1912506480021271e-06
GC_12_48 b_12 NI_12 NS_48 0 2.7906296105152532e-06
GC_12_49 b_12 NI_12 NS_49 0 -1.1302622064664544e-06
GC_12_50 b_12 NI_12 NS_50 0 6.5760368578741155e-06
GC_12_51 b_12 NI_12 NS_51 0 -4.1810107968636913e-07
GC_12_52 b_12 NI_12 NS_52 0 2.1387914932411373e-06
GC_12_53 b_12 NI_12 NS_53 0 7.2163585024804401e-06
GC_12_54 b_12 NI_12 NS_54 0 5.1185228015276619e-06
GC_12_55 b_12 NI_12 NS_55 0 1.6097738392966683e-06
GC_12_56 b_12 NI_12 NS_56 0 3.1433788916466673e-06
GC_12_57 b_12 NI_12 NS_57 0 4.8364232917524590e-06
GC_12_58 b_12 NI_12 NS_58 0 1.1505232861193836e-06
GC_12_59 b_12 NI_12 NS_59 0 2.9136132480920116e-06
GC_12_60 b_12 NI_12 NS_60 0 -1.3226684409065287e-06
GC_12_61 b_12 NI_12 NS_61 0 1.2106007700698675e-08
GC_12_62 b_12 NI_12 NS_62 0 -8.1607724473917441e-10
GC_12_63 b_12 NI_12 NS_63 0 -1.6069712447068123e-11
GC_12_64 b_12 NI_12 NS_64 0 1.3075627944756318e-10
GC_12_65 b_12 NI_12 NS_65 0 6.7316804626362200e-08
GC_12_66 b_12 NI_12 NS_66 0 -1.0258734476238071e-08
GC_12_67 b_12 NI_12 NS_67 0 -5.8672887394209879e-07
GC_12_68 b_12 NI_12 NS_68 0 5.6507219275813845e-07
GC_12_69 b_12 NI_12 NS_69 0 1.6793028172713135e-06
GC_12_70 b_12 NI_12 NS_70 0 -4.9707772017475448e-07
GC_12_71 b_12 NI_12 NS_71 0 -9.7352492628771473e-07
GC_12_72 b_12 NI_12 NS_72 0 1.1756514757272984e-07
GC_12_73 b_12 NI_12 NS_73 0 1.6616849787553703e-06
GC_12_74 b_12 NI_12 NS_74 0 -1.1455582813553621e-06
GC_12_75 b_12 NI_12 NS_75 0 -9.0102798366742374e-07
GC_12_76 b_12 NI_12 NS_76 0 -8.6217881073158520e-07
GC_12_77 b_12 NI_12 NS_77 0 -1.1351755872321114e-06
GC_12_78 b_12 NI_12 NS_78 0 -2.5009866294180292e-07
GC_12_79 b_12 NI_12 NS_79 0 8.9211526006683745e-08
GC_12_80 b_12 NI_12 NS_80 0 1.1707706966858266e-06
GC_12_81 b_12 NI_12 NS_81 0 -2.4072625796988510e-08
GC_12_82 b_12 NI_12 NS_82 0 1.2303584415501799e-09
GC_12_83 b_12 NI_12 NS_83 0 2.1589039643871709e-11
GC_12_84 b_12 NI_12 NS_84 0 -1.7715317255558408e-10
GC_12_85 b_12 NI_12 NS_85 0 1.8511907218037083e-06
GC_12_86 b_12 NI_12 NS_86 0 -4.1799796668254263e-06
GC_12_87 b_12 NI_12 NS_87 0 2.4721015583538056e-06
GC_12_88 b_12 NI_12 NS_88 0 9.2956230577807551e-08
GC_12_89 b_12 NI_12 NS_89 0 -1.6039211486997497e-06
GC_12_90 b_12 NI_12 NS_90 0 -4.4881541102459727e-06
GC_12_91 b_12 NI_12 NS_91 0 9.6225879227102122e-07
GC_12_92 b_12 NI_12 NS_92 0 -7.3177748083844976e-06
GC_12_93 b_12 NI_12 NS_93 0 -8.8052550289210104e-06
GC_12_94 b_12 NI_12 NS_94 0 -4.6098778630091865e-06
GC_12_95 b_12 NI_12 NS_95 0 -3.2625427767199931e-06
GC_12_96 b_12 NI_12 NS_96 0 1.4328969672693819e-06
GC_12_97 b_12 NI_12 NS_97 0 -1.8926889321340110e-06
GC_12_98 b_12 NI_12 NS_98 0 -5.4632580839357924e-07
GC_12_99 b_12 NI_12 NS_99 0 -3.2845056178010501e-06
GC_12_100 b_12 NI_12 NS_100 0 -1.5188069760774799e-06
GC_12_101 b_12 NI_12 NS_101 0 2.0778198330531370e-08
GC_12_102 b_12 NI_12 NS_102 0 -1.0272256493056005e-09
GC_12_103 b_12 NI_12 NS_103 0 -1.9428684944092260e-11
GC_12_104 b_12 NI_12 NS_104 0 1.5753100077666516e-10
GC_12_105 b_12 NI_12 NS_105 0 -1.1217624682380167e-06
GC_12_106 b_12 NI_12 NS_106 0 -8.0925817113875196e-07
GC_12_107 b_12 NI_12 NS_107 0 -2.0036364271147203e-06
GC_12_108 b_12 NI_12 NS_108 0 3.6547335154770767e-08
GC_12_109 b_12 NI_12 NS_109 0 -3.0739376635560486e-06
GC_12_110 b_12 NI_12 NS_110 0 8.6266621104533135e-07
GC_12_111 b_12 NI_12 NS_111 0 -4.1492023864912274e-06
GC_12_112 b_12 NI_12 NS_112 0 4.3129833637817266e-06
GC_12_113 b_12 NI_12 NS_113 0 3.3149236285788492e-06
GC_12_114 b_12 NI_12 NS_114 0 5.4267707069496117e-06
GC_12_115 b_12 NI_12 NS_115 0 -8.9973928816588690e-07
GC_12_116 b_12 NI_12 NS_116 0 5.9728356453656474e-06
GC_12_117 b_12 NI_12 NS_117 0 6.0574023997706786e-06
GC_12_118 b_12 NI_12 NS_118 0 3.3263250418503469e-06
GC_12_119 b_12 NI_12 NS_119 0 5.8642834330265700e-06
GC_12_120 b_12 NI_12 NS_120 0 1.7030943136346586e-06
GC_12_121 b_12 NI_12 NS_121 0 1.1017192562109760e-09
GC_12_122 b_12 NI_12 NS_122 0 -1.2973268727606295e-10
GC_12_123 b_12 NI_12 NS_123 0 1.7862164751323448e-11
GC_12_124 b_12 NI_12 NS_124 0 -9.6104739320483837e-11
GC_12_125 b_12 NI_12 NS_125 0 -1.9127609136197165e-06
GC_12_126 b_12 NI_12 NS_126 0 -1.1371603682902866e-06
GC_12_127 b_12 NI_12 NS_127 0 -6.0327982251055266e-06
GC_12_128 b_12 NI_12 NS_128 0 1.3796838375104208e-05
GC_12_129 b_12 NI_12 NS_129 0 3.5155038418529905e-05
GC_12_130 b_12 NI_12 NS_130 0 1.1739173386579375e-05
GC_12_131 b_12 NI_12 NS_131 0 3.2374347428810980e-05
GC_12_132 b_12 NI_12 NS_132 0 -2.5608400859484606e-05
GC_12_133 b_12 NI_12 NS_133 0 -3.9769248371542705e-05
GC_12_134 b_12 NI_12 NS_134 0 -4.9607555460096675e-05
GC_12_135 b_12 NI_12 NS_135 0 -1.9812840964574548e-05
GC_12_136 b_12 NI_12 NS_136 0 1.0190878968906249e-05
GC_12_137 b_12 NI_12 NS_137 0 4.9362766377343271e-06
GC_12_138 b_12 NI_12 NS_138 0 3.9503311961443643e-07
GC_12_139 b_12 NI_12 NS_139 0 -1.2398869698488733e-05
GC_12_140 b_12 NI_12 NS_140 0 -7.1395625148057625e-06
GC_12_141 b_12 NI_12 NS_141 0 -2.5754063776220947e-08
GC_12_142 b_12 NI_12 NS_142 0 1.1438284551779549e-09
GC_12_143 b_12 NI_12 NS_143 0 -1.1059886470990824e-11
GC_12_144 b_12 NI_12 NS_144 0 3.1894465303223854e-11
GC_12_145 b_12 NI_12 NS_145 0 4.4269009274707093e-06
GC_12_146 b_12 NI_12 NS_146 0 2.3386907249128186e-06
GC_12_147 b_12 NI_12 NS_147 0 9.9199539753604205e-06
GC_12_148 b_12 NI_12 NS_148 0 9.7652561005697354e-06
GC_12_149 b_12 NI_12 NS_149 0 1.8817727558306793e-05
GC_12_150 b_12 NI_12 NS_150 0 -2.3372956409274537e-05
GC_12_151 b_12 NI_12 NS_151 0 1.1289948395455642e-05
GC_12_152 b_12 NI_12 NS_152 0 -3.2013244823291166e-06
GC_12_153 b_12 NI_12 NS_153 0 -6.5988113817069921e-06
GC_12_154 b_12 NI_12 NS_154 0 -5.3073158368814812e-05
GC_12_155 b_12 NI_12 NS_155 0 -1.4827253670180887e-05
GC_12_156 b_12 NI_12 NS_156 0 -1.7892237989297917e-05
GC_12_157 b_12 NI_12 NS_157 0 -2.7603789960950623e-05
GC_12_158 b_12 NI_12 NS_158 0 -1.2421187832311726e-05
GC_12_159 b_12 NI_12 NS_159 0 -1.9027358968843341e-05
GC_12_160 b_12 NI_12 NS_160 0 5.9411138282685284e-06
GC_12_161 b_12 NI_12 NS_161 0 -1.8490440641954348e-06
GC_12_162 b_12 NI_12 NS_162 0 2.5677075147041633e-07
GC_12_163 b_12 NI_12 NS_163 0 1.6912978920197489e-09
GC_12_164 b_12 NI_12 NS_164 0 1.3611966760933655e-08
GC_12_165 b_12 NI_12 NS_165 0 1.1406456016643991e-03
GC_12_166 b_12 NI_12 NS_166 0 -2.1726046680037923e-03
GC_12_167 b_12 NI_12 NS_167 0 3.4952388269267648e-03
GC_12_168 b_12 NI_12 NS_168 0 -1.3003077401248245e-02
GC_12_169 b_12 NI_12 NS_169 0 -3.9401362127337594e-02
GC_12_170 b_12 NI_12 NS_170 0 -3.6437949542473440e-04
GC_12_171 b_12 NI_12 NS_171 0 -2.6247364683507662e-02
GC_12_172 b_12 NI_12 NS_172 0 2.8990158567117112e-02
GC_12_173 b_12 NI_12 NS_173 0 5.2202632001945491e-02
GC_12_174 b_12 NI_12 NS_174 0 3.8208679918731628e-02
GC_12_175 b_12 NI_12 NS_175 0 1.7572267604685811e-02
GC_12_176 b_12 NI_12 NS_176 0 -1.4394059929725983e-02
GC_12_177 b_12 NI_12 NS_177 0 -9.1651296156218011e-03
GC_12_178 b_12 NI_12 NS_178 0 -3.7458101159816241e-03
GC_12_179 b_12 NI_12 NS_179 0 8.0623393086459733e-03
GC_12_180 b_12 NI_12 NS_180 0 5.8595892984327214e-03
GC_12_181 b_12 NI_12 NS_181 0 -1.0355529015791468e-05
GC_12_182 b_12 NI_12 NS_182 0 -2.1274259819609918e-07
GC_12_183 b_12 NI_12 NS_183 0 -1.2832451361373878e-09
GC_12_184 b_12 NI_12 NS_184 0 -2.5390012878643017e-08
GC_12_185 b_12 NI_12 NS_185 0 -4.2497322965482408e-03
GC_12_186 b_12 NI_12 NS_186 0 -3.4927923626545312e-03
GC_12_187 b_12 NI_12 NS_187 0 -1.2922477265220875e-02
GC_12_188 b_12 NI_12 NS_188 0 1.7065692851498025e-02
GC_12_189 b_12 NI_12 NS_189 0 1.7371378434938866e-02
GC_12_190 b_12 NI_12 NS_190 0 -1.9446862252898902e-02
GC_12_191 b_12 NI_12 NS_191 0 -3.3168754961407691e-02
GC_12_192 b_12 NI_12 NS_192 0 2.5454292393380318e-02
GC_12_193 b_12 NI_12 NS_193 0 4.0789565682369668e-02
GC_12_194 b_12 NI_12 NS_194 0 -1.1433259751476599e-02
GC_12_195 b_12 NI_12 NS_195 0 -2.1059403379134214e-02
GC_12_196 b_12 NI_12 NS_196 0 1.5315262612977363e-02
GC_12_197 b_12 NI_12 NS_197 0 1.4123881158377621e-02
GC_12_198 b_12 NI_12 NS_198 0 -3.7536567067230223e-03
GC_12_199 b_12 NI_12 NS_199 0 7.0870161015161642e-03
GC_12_200 b_12 NI_12 NS_200 0 1.3573831691721277e-02
GC_12_201 b_12 NI_12 NS_201 0 8.9999191136949723e-05
GC_12_202 b_12 NI_12 NS_202 0 3.6211572001889603e-06
GC_12_203 b_12 NI_12 NS_203 0 5.9678531418353555e-09
GC_12_204 b_12 NI_12 NS_204 0 5.9667815859358460e-07
GC_12_205 b_12 NI_12 NS_205 0 4.7508813473330587e-02
GC_12_206 b_12 NI_12 NS_206 0 -9.6471254253403787e-03
GC_12_207 b_12 NI_12 NS_207 0 -4.5582968181618368e-02
GC_12_208 b_12 NI_12 NS_208 0 2.0552255656018408e-02
GC_12_209 b_12 NI_12 NS_209 0 -5.7696971420534350e-02
GC_12_210 b_12 NI_12 NS_210 0 -6.7350096396171621e-02
GC_12_211 b_12 NI_12 NS_211 0 6.3862106370389721e-02
GC_12_212 b_12 NI_12 NS_212 0 -2.2063600270370499e-02
GC_12_213 b_12 NI_12 NS_213 0 2.8382466453299202e-02
GC_12_214 b_12 NI_12 NS_214 0 8.9387907056920748e-02
GC_12_215 b_12 NI_12 NS_215 0 -5.4366402503193280e-02
GC_12_216 b_12 NI_12 NS_216 0 2.7979809770003854e-03
GC_12_217 b_12 NI_12 NS_217 0 -1.3847752170212951e-02
GC_12_218 b_12 NI_12 NS_218 0 -4.7095020884852339e-02
GC_12_219 b_12 NI_12 NS_219 0 1.6380502283893608e-02
GC_12_220 b_12 NI_12 NS_220 0 -3.9016241064613558e-02
GC_12_221 b_12 NI_12 NS_221 0 -1.5427135100830025e-05
GC_12_222 b_12 NI_12 NS_222 0 -3.7324314362848548e-06
GC_12_223 b_12 NI_12 NS_223 0 -2.3081208540649659e-08
GC_12_224 b_12 NI_12 NS_224 0 -3.8674152064337271e-07
GC_12_225 b_12 NI_12 NS_225 0 4.5760065486724934e-03
GC_12_226 b_12 NI_12 NS_226 0 3.7993286749984554e-03
GC_12_227 b_12 NI_12 NS_227 0 1.3872401194724821e-02
GC_12_228 b_12 NI_12 NS_228 0 -2.1406272357366692e-02
GC_12_229 b_12 NI_12 NS_229 0 -2.2493840892053685e-02
GC_12_230 b_12 NI_12 NS_230 0 2.6058892794354339e-02
GC_12_231 b_12 NI_12 NS_231 0 3.8337056260354004e-02
GC_12_232 b_12 NI_12 NS_232 0 -3.0181707200149149e-02
GC_12_233 b_12 NI_12 NS_233 0 -4.8685823046150968e-02
GC_12_234 b_12 NI_12 NS_234 0 1.9831379025888881e-02
GC_12_235 b_12 NI_12 NS_235 0 2.6967890269789570e-02
GC_12_236 b_12 NI_12 NS_236 0 -1.5945601277778002e-02
GC_12_237 b_12 NI_12 NS_237 0 -1.4394992355179034e-02
GC_12_238 b_12 NI_12 NS_238 0 6.8900417725550351e-03
GC_12_239 b_12 NI_12 NS_239 0 -4.8273798937392039e-03
GC_12_240 b_12 NI_12 NS_240 0 -1.6678597174828440e-02
GD_12_1 b_12 NI_12 NA_1 0 3.4974418709710693e-07
GD_12_2 b_12 NI_12 NA_2 0 -1.5460729796501311e-06
GD_12_3 b_12 NI_12 NA_3 0 -7.7232122284489841e-06
GD_12_4 b_12 NI_12 NA_4 0 3.0621149873090703e-07
GD_12_5 b_12 NI_12 NA_5 0 1.0098377175198105e-05
GD_12_6 b_12 NI_12 NA_6 0 -1.1680798391685690e-06
GD_12_7 b_12 NI_12 NA_7 0 3.3229607739967262e-06
GD_12_8 b_12 NI_12 NA_8 0 1.4712435896906739e-05
GD_12_9 b_12 NI_12 NA_9 0 -3.3302474403628201e-03
GD_12_10 b_12 NI_12 NA_10 0 6.7731250245857870e-03
GD_12_11 b_12 NI_12 NA_11 0 5.5524721466031516e-03
GD_12_12 b_12 NI_12 NA_12 0 -9.5068691426404475e-03
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 6.8759459879260660e+01
GS_1_1 0 NS_1 NA_1 0 6.0286980150450964e-01
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 2.4827714035206478e+02
GS_2_1 0 NS_2 NA_1 0 6.0286980150450964e-01
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 5.8935503054175797e+03
GS_3_1 0 NS_3 NA_1 0 6.0286980150450964e-01
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 1.2841015484081297e+03
GS_4_1 0 NS_4 NA_1 0 6.0286980150450964e-01
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 2.8319423052259118e+01
RS_6 NS_6 0 2.8319423052259115e+01
GL_5 0 NS_5 NS_6 0 3.0726343572183612e-01
GL_6 0 NS_6 NS_5 0 -3.0726343572183612e-01
GS_5_1 0 NS_5 NA_1 0 6.0286980150450964e-01
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 1.8367949753848961e+01
RS_8 NS_8 0 1.8367949753848965e+01
GL_7 0 NS_7 NS_8 0 2.4584800021674161e-01
GL_8 0 NS_8 NS_7 0 -2.4584800021674161e-01
GS_7_1 0 NS_7 NA_1 0 6.0286980150450964e-01
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 1.4690910804179261e+01
RS_10 NS_10 0 1.4690910804179261e+01
GL_9 0 NS_9 NS_10 0 2.1320637363820186e-01
GL_10 0 NS_10 NS_9 0 -2.1320637363820186e-01
GS_9_1 0 NS_9 NA_1 0 6.0286980150450964e-01
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 1.6315799932686236e+01
RS_12 NS_12 0 1.6315799932686236e+01
GL_11 0 NS_11 NS_12 0 1.6372677698710228e-01
GL_12 0 NS_12 NS_11 0 -1.6372677698710228e-01
GS_11_1 0 NS_11 NA_1 0 6.0286980150450964e-01
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 1.3805021583364081e+01
RS_14 NS_14 0 1.3805021583364081e+01
GL_13 0 NS_13 NS_14 0 1.3053652152390091e-01
GL_14 0 NS_14 NS_13 0 -1.3053652152390091e-01
GS_13_1 0 NS_13 NA_1 0 6.0286980150450964e-01
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 1.7453012154519879e+01
RS_16 NS_16 0 1.7453012154519879e+01
GL_15 0 NS_15 NS_16 0 8.4170507635427994e-02
GL_16 0 NS_16 NS_15 0 -8.4170507635427994e-02
GS_15_1 0 NS_15 NA_1 0 6.0286980150450964e-01
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 1.7836078439168801e+01
RS_18 NS_18 0 1.7836078439168805e+01
GL_17 0 NS_17 NS_18 0 5.3586142573527437e-02
GL_18 0 NS_18 NS_17 0 -5.3586142573527437e-02
GS_17_1 0 NS_17 NA_1 0 6.0286980150450964e-01
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 1.9366404748437819e+01
RS_20 NS_20 0 1.9366404748437819e+01
GL_19 0 NS_19 NS_20 0 2.0213646406074141e-02
GL_20 0 NS_20 NS_19 0 -2.0213646406074141e-02
GS_19_1 0 NS_19 NA_1 0 6.0286980150450964e-01
*
* Real pole n. 21
CS_21 NS_21 0 9.9999999999999998e-13
RS_21 NS_21 0 6.8759459879260660e+01
GS_21_2 0 NS_21 NA_2 0 6.0286980150450964e-01
*
* Real pole n. 22
CS_22 NS_22 0 9.9999999999999998e-13
RS_22 NS_22 0 2.4827714035206478e+02
GS_22_2 0 NS_22 NA_2 0 6.0286980150450964e-01
*
* Real pole n. 23
CS_23 NS_23 0 9.9999999999999998e-13
RS_23 NS_23 0 5.8935503054175797e+03
GS_23_2 0 NS_23 NA_2 0 6.0286980150450964e-01
*
* Real pole n. 24
CS_24 NS_24 0 9.9999999999999998e-13
RS_24 NS_24 0 1.2841015484081297e+03
GS_24_2 0 NS_24 NA_2 0 6.0286980150450964e-01
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 2.8319423052259118e+01
RS_26 NS_26 0 2.8319423052259115e+01
GL_25 0 NS_25 NS_26 0 3.0726343572183612e-01
GL_26 0 NS_26 NS_25 0 -3.0726343572183612e-01
GS_25_2 0 NS_25 NA_2 0 6.0286980150450964e-01
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 1.8367949753848961e+01
RS_28 NS_28 0 1.8367949753848965e+01
GL_27 0 NS_27 NS_28 0 2.4584800021674161e-01
GL_28 0 NS_28 NS_27 0 -2.4584800021674161e-01
GS_27_2 0 NS_27 NA_2 0 6.0286980150450964e-01
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 1.4690910804179261e+01
RS_30 NS_30 0 1.4690910804179261e+01
GL_29 0 NS_29 NS_30 0 2.1320637363820186e-01
GL_30 0 NS_30 NS_29 0 -2.1320637363820186e-01
GS_29_2 0 NS_29 NA_2 0 6.0286980150450964e-01
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 1.6315799932686236e+01
RS_32 NS_32 0 1.6315799932686236e+01
GL_31 0 NS_31 NS_32 0 1.6372677698710228e-01
GL_32 0 NS_32 NS_31 0 -1.6372677698710228e-01
GS_31_2 0 NS_31 NA_2 0 6.0286980150450964e-01
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 1.3805021583364081e+01
RS_34 NS_34 0 1.3805021583364081e+01
GL_33 0 NS_33 NS_34 0 1.3053652152390091e-01
GL_34 0 NS_34 NS_33 0 -1.3053652152390091e-01
GS_33_2 0 NS_33 NA_2 0 6.0286980150450964e-01
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 1.7453012154519879e+01
RS_36 NS_36 0 1.7453012154519879e+01
GL_35 0 NS_35 NS_36 0 8.4170507635427994e-02
GL_36 0 NS_36 NS_35 0 -8.4170507635427994e-02
GS_35_2 0 NS_35 NA_2 0 6.0286980150450964e-01
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 1.7836078439168801e+01
RS_38 NS_38 0 1.7836078439168805e+01
GL_37 0 NS_37 NS_38 0 5.3586142573527437e-02
GL_38 0 NS_38 NS_37 0 -5.3586142573527437e-02
GS_37_2 0 NS_37 NA_2 0 6.0286980150450964e-01
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 1.9366404748437819e+01
RS_40 NS_40 0 1.9366404748437819e+01
GL_39 0 NS_39 NS_40 0 2.0213646406074141e-02
GL_40 0 NS_40 NS_39 0 -2.0213646406074141e-02
GS_39_2 0 NS_39 NA_2 0 6.0286980150450964e-01
*
* Real pole n. 41
CS_41 NS_41 0 9.9999999999999998e-13
RS_41 NS_41 0 6.8759459879260660e+01
GS_41_3 0 NS_41 NA_3 0 6.0286980150450964e-01
*
* Real pole n. 42
CS_42 NS_42 0 9.9999999999999998e-13
RS_42 NS_42 0 2.4827714035206478e+02
GS_42_3 0 NS_42 NA_3 0 6.0286980150450964e-01
*
* Real pole n. 43
CS_43 NS_43 0 9.9999999999999998e-13
RS_43 NS_43 0 5.8935503054175797e+03
GS_43_3 0 NS_43 NA_3 0 6.0286980150450964e-01
*
* Real pole n. 44
CS_44 NS_44 0 9.9999999999999998e-13
RS_44 NS_44 0 1.2841015484081297e+03
GS_44_3 0 NS_44 NA_3 0 6.0286980150450964e-01
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 2.8319423052259118e+01
RS_46 NS_46 0 2.8319423052259115e+01
GL_45 0 NS_45 NS_46 0 3.0726343572183612e-01
GL_46 0 NS_46 NS_45 0 -3.0726343572183612e-01
GS_45_3 0 NS_45 NA_3 0 6.0286980150450964e-01
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 1.8367949753848961e+01
RS_48 NS_48 0 1.8367949753848965e+01
GL_47 0 NS_47 NS_48 0 2.4584800021674161e-01
GL_48 0 NS_48 NS_47 0 -2.4584800021674161e-01
GS_47_3 0 NS_47 NA_3 0 6.0286980150450964e-01
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 1.4690910804179261e+01
RS_50 NS_50 0 1.4690910804179261e+01
GL_49 0 NS_49 NS_50 0 2.1320637363820186e-01
GL_50 0 NS_50 NS_49 0 -2.1320637363820186e-01
GS_49_3 0 NS_49 NA_3 0 6.0286980150450964e-01
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 1.6315799932686236e+01
RS_52 NS_52 0 1.6315799932686236e+01
GL_51 0 NS_51 NS_52 0 1.6372677698710228e-01
GL_52 0 NS_52 NS_51 0 -1.6372677698710228e-01
GS_51_3 0 NS_51 NA_3 0 6.0286980150450964e-01
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 1.3805021583364081e+01
RS_54 NS_54 0 1.3805021583364081e+01
GL_53 0 NS_53 NS_54 0 1.3053652152390091e-01
GL_54 0 NS_54 NS_53 0 -1.3053652152390091e-01
GS_53_3 0 NS_53 NA_3 0 6.0286980150450964e-01
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 1.7453012154519879e+01
RS_56 NS_56 0 1.7453012154519879e+01
GL_55 0 NS_55 NS_56 0 8.4170507635427994e-02
GL_56 0 NS_56 NS_55 0 -8.4170507635427994e-02
GS_55_3 0 NS_55 NA_3 0 6.0286980150450964e-01
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 1.7836078439168801e+01
RS_58 NS_58 0 1.7836078439168805e+01
GL_57 0 NS_57 NS_58 0 5.3586142573527437e-02
GL_58 0 NS_58 NS_57 0 -5.3586142573527437e-02
GS_57_3 0 NS_57 NA_3 0 6.0286980150450964e-01
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 1.9366404748437819e+01
RS_60 NS_60 0 1.9366404748437819e+01
GL_59 0 NS_59 NS_60 0 2.0213646406074141e-02
GL_60 0 NS_60 NS_59 0 -2.0213646406074141e-02
GS_59_3 0 NS_59 NA_3 0 6.0286980150450964e-01
*
* Real pole n. 61
CS_61 NS_61 0 9.9999999999999998e-13
RS_61 NS_61 0 6.8759459879260660e+01
GS_61_4 0 NS_61 NA_4 0 6.0286980150450964e-01
*
* Real pole n. 62
CS_62 NS_62 0 9.9999999999999998e-13
RS_62 NS_62 0 2.4827714035206478e+02
GS_62_4 0 NS_62 NA_4 0 6.0286980150450964e-01
*
* Real pole n. 63
CS_63 NS_63 0 9.9999999999999998e-13
RS_63 NS_63 0 5.8935503054175797e+03
GS_63_4 0 NS_63 NA_4 0 6.0286980150450964e-01
*
* Real pole n. 64
CS_64 NS_64 0 9.9999999999999998e-13
RS_64 NS_64 0 1.2841015484081297e+03
GS_64_4 0 NS_64 NA_4 0 6.0286980150450964e-01
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 2.8319423052259118e+01
RS_66 NS_66 0 2.8319423052259115e+01
GL_65 0 NS_65 NS_66 0 3.0726343572183612e-01
GL_66 0 NS_66 NS_65 0 -3.0726343572183612e-01
GS_65_4 0 NS_65 NA_4 0 6.0286980150450964e-01
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 1.8367949753848961e+01
RS_68 NS_68 0 1.8367949753848965e+01
GL_67 0 NS_67 NS_68 0 2.4584800021674161e-01
GL_68 0 NS_68 NS_67 0 -2.4584800021674161e-01
GS_67_4 0 NS_67 NA_4 0 6.0286980150450964e-01
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 1.4690910804179261e+01
RS_70 NS_70 0 1.4690910804179261e+01
GL_69 0 NS_69 NS_70 0 2.1320637363820186e-01
GL_70 0 NS_70 NS_69 0 -2.1320637363820186e-01
GS_69_4 0 NS_69 NA_4 0 6.0286980150450964e-01
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 1.6315799932686236e+01
RS_72 NS_72 0 1.6315799932686236e+01
GL_71 0 NS_71 NS_72 0 1.6372677698710228e-01
GL_72 0 NS_72 NS_71 0 -1.6372677698710228e-01
GS_71_4 0 NS_71 NA_4 0 6.0286980150450964e-01
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 1.3805021583364081e+01
RS_74 NS_74 0 1.3805021583364081e+01
GL_73 0 NS_73 NS_74 0 1.3053652152390091e-01
GL_74 0 NS_74 NS_73 0 -1.3053652152390091e-01
GS_73_4 0 NS_73 NA_4 0 6.0286980150450964e-01
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 1.7453012154519879e+01
RS_76 NS_76 0 1.7453012154519879e+01
GL_75 0 NS_75 NS_76 0 8.4170507635427994e-02
GL_76 0 NS_76 NS_75 0 -8.4170507635427994e-02
GS_75_4 0 NS_75 NA_4 0 6.0286980150450964e-01
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 1.7836078439168801e+01
RS_78 NS_78 0 1.7836078439168805e+01
GL_77 0 NS_77 NS_78 0 5.3586142573527437e-02
GL_78 0 NS_78 NS_77 0 -5.3586142573527437e-02
GS_77_4 0 NS_77 NA_4 0 6.0286980150450964e-01
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 1.9366404748437819e+01
RS_80 NS_80 0 1.9366404748437819e+01
GL_79 0 NS_79 NS_80 0 2.0213646406074141e-02
GL_80 0 NS_80 NS_79 0 -2.0213646406074141e-02
GS_79_4 0 NS_79 NA_4 0 6.0286980150450964e-01
*
* Real pole n. 81
CS_81 NS_81 0 9.9999999999999998e-13
RS_81 NS_81 0 6.8759459879260660e+01
GS_81_5 0 NS_81 NA_5 0 6.0286980150450964e-01
*
* Real pole n. 82
CS_82 NS_82 0 9.9999999999999998e-13
RS_82 NS_82 0 2.4827714035206478e+02
GS_82_5 0 NS_82 NA_5 0 6.0286980150450964e-01
*
* Real pole n. 83
CS_83 NS_83 0 9.9999999999999998e-13
RS_83 NS_83 0 5.8935503054175797e+03
GS_83_5 0 NS_83 NA_5 0 6.0286980150450964e-01
*
* Real pole n. 84
CS_84 NS_84 0 9.9999999999999998e-13
RS_84 NS_84 0 1.2841015484081297e+03
GS_84_5 0 NS_84 NA_5 0 6.0286980150450964e-01
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 2.8319423052259118e+01
RS_86 NS_86 0 2.8319423052259115e+01
GL_85 0 NS_85 NS_86 0 3.0726343572183612e-01
GL_86 0 NS_86 NS_85 0 -3.0726343572183612e-01
GS_85_5 0 NS_85 NA_5 0 6.0286980150450964e-01
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 1.8367949753848961e+01
RS_88 NS_88 0 1.8367949753848965e+01
GL_87 0 NS_87 NS_88 0 2.4584800021674161e-01
GL_88 0 NS_88 NS_87 0 -2.4584800021674161e-01
GS_87_5 0 NS_87 NA_5 0 6.0286980150450964e-01
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 1.4690910804179261e+01
RS_90 NS_90 0 1.4690910804179261e+01
GL_89 0 NS_89 NS_90 0 2.1320637363820186e-01
GL_90 0 NS_90 NS_89 0 -2.1320637363820186e-01
GS_89_5 0 NS_89 NA_5 0 6.0286980150450964e-01
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 1.6315799932686236e+01
RS_92 NS_92 0 1.6315799932686236e+01
GL_91 0 NS_91 NS_92 0 1.6372677698710228e-01
GL_92 0 NS_92 NS_91 0 -1.6372677698710228e-01
GS_91_5 0 NS_91 NA_5 0 6.0286980150450964e-01
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 1.3805021583364081e+01
RS_94 NS_94 0 1.3805021583364081e+01
GL_93 0 NS_93 NS_94 0 1.3053652152390091e-01
GL_94 0 NS_94 NS_93 0 -1.3053652152390091e-01
GS_93_5 0 NS_93 NA_5 0 6.0286980150450964e-01
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 1.7453012154519879e+01
RS_96 NS_96 0 1.7453012154519879e+01
GL_95 0 NS_95 NS_96 0 8.4170507635427994e-02
GL_96 0 NS_96 NS_95 0 -8.4170507635427994e-02
GS_95_5 0 NS_95 NA_5 0 6.0286980150450964e-01
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 1.7836078439168801e+01
RS_98 NS_98 0 1.7836078439168805e+01
GL_97 0 NS_97 NS_98 0 5.3586142573527437e-02
GL_98 0 NS_98 NS_97 0 -5.3586142573527437e-02
GS_97_5 0 NS_97 NA_5 0 6.0286980150450964e-01
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 1.9366404748437819e+01
RS_100 NS_100 0 1.9366404748437819e+01
GL_99 0 NS_99 NS_100 0 2.0213646406074141e-02
GL_100 0 NS_100 NS_99 0 -2.0213646406074141e-02
GS_99_5 0 NS_99 NA_5 0 6.0286980150450964e-01
*
* Real pole n. 101
CS_101 NS_101 0 9.9999999999999998e-13
RS_101 NS_101 0 6.8759459879260660e+01
GS_101_6 0 NS_101 NA_6 0 6.0286980150450964e-01
*
* Real pole n. 102
CS_102 NS_102 0 9.9999999999999998e-13
RS_102 NS_102 0 2.4827714035206478e+02
GS_102_6 0 NS_102 NA_6 0 6.0286980150450964e-01
*
* Real pole n. 103
CS_103 NS_103 0 9.9999999999999998e-13
RS_103 NS_103 0 5.8935503054175797e+03
GS_103_6 0 NS_103 NA_6 0 6.0286980150450964e-01
*
* Real pole n. 104
CS_104 NS_104 0 9.9999999999999998e-13
RS_104 NS_104 0 1.2841015484081297e+03
GS_104_6 0 NS_104 NA_6 0 6.0286980150450964e-01
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 2.8319423052259118e+01
RS_106 NS_106 0 2.8319423052259115e+01
GL_105 0 NS_105 NS_106 0 3.0726343572183612e-01
GL_106 0 NS_106 NS_105 0 -3.0726343572183612e-01
GS_105_6 0 NS_105 NA_6 0 6.0286980150450964e-01
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 1.8367949753848961e+01
RS_108 NS_108 0 1.8367949753848965e+01
GL_107 0 NS_107 NS_108 0 2.4584800021674161e-01
GL_108 0 NS_108 NS_107 0 -2.4584800021674161e-01
GS_107_6 0 NS_107 NA_6 0 6.0286980150450964e-01
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 1.4690910804179261e+01
RS_110 NS_110 0 1.4690910804179261e+01
GL_109 0 NS_109 NS_110 0 2.1320637363820186e-01
GL_110 0 NS_110 NS_109 0 -2.1320637363820186e-01
GS_109_6 0 NS_109 NA_6 0 6.0286980150450964e-01
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 1.6315799932686236e+01
RS_112 NS_112 0 1.6315799932686236e+01
GL_111 0 NS_111 NS_112 0 1.6372677698710228e-01
GL_112 0 NS_112 NS_111 0 -1.6372677698710228e-01
GS_111_6 0 NS_111 NA_6 0 6.0286980150450964e-01
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 1.3805021583364081e+01
RS_114 NS_114 0 1.3805021583364081e+01
GL_113 0 NS_113 NS_114 0 1.3053652152390091e-01
GL_114 0 NS_114 NS_113 0 -1.3053652152390091e-01
GS_113_6 0 NS_113 NA_6 0 6.0286980150450964e-01
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 1.7453012154519879e+01
RS_116 NS_116 0 1.7453012154519879e+01
GL_115 0 NS_115 NS_116 0 8.4170507635427994e-02
GL_116 0 NS_116 NS_115 0 -8.4170507635427994e-02
GS_115_6 0 NS_115 NA_6 0 6.0286980150450964e-01
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 1.7836078439168801e+01
RS_118 NS_118 0 1.7836078439168805e+01
GL_117 0 NS_117 NS_118 0 5.3586142573527437e-02
GL_118 0 NS_118 NS_117 0 -5.3586142573527437e-02
GS_117_6 0 NS_117 NA_6 0 6.0286980150450964e-01
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 1.9366404748437819e+01
RS_120 NS_120 0 1.9366404748437819e+01
GL_119 0 NS_119 NS_120 0 2.0213646406074141e-02
GL_120 0 NS_120 NS_119 0 -2.0213646406074141e-02
GS_119_6 0 NS_119 NA_6 0 6.0286980150450964e-01
*
* Real pole n. 121
CS_121 NS_121 0 9.9999999999999998e-13
RS_121 NS_121 0 6.8759459879260660e+01
GS_121_7 0 NS_121 NA_7 0 6.0286980150450964e-01
*
* Real pole n. 122
CS_122 NS_122 0 9.9999999999999998e-13
RS_122 NS_122 0 2.4827714035206478e+02
GS_122_7 0 NS_122 NA_7 0 6.0286980150450964e-01
*
* Real pole n. 123
CS_123 NS_123 0 9.9999999999999998e-13
RS_123 NS_123 0 5.8935503054175797e+03
GS_123_7 0 NS_123 NA_7 0 6.0286980150450964e-01
*
* Real pole n. 124
CS_124 NS_124 0 9.9999999999999998e-13
RS_124 NS_124 0 1.2841015484081297e+03
GS_124_7 0 NS_124 NA_7 0 6.0286980150450964e-01
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 2.8319423052259118e+01
RS_126 NS_126 0 2.8319423052259115e+01
GL_125 0 NS_125 NS_126 0 3.0726343572183612e-01
GL_126 0 NS_126 NS_125 0 -3.0726343572183612e-01
GS_125_7 0 NS_125 NA_7 0 6.0286980150450964e-01
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 1.8367949753848961e+01
RS_128 NS_128 0 1.8367949753848965e+01
GL_127 0 NS_127 NS_128 0 2.4584800021674161e-01
GL_128 0 NS_128 NS_127 0 -2.4584800021674161e-01
GS_127_7 0 NS_127 NA_7 0 6.0286980150450964e-01
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 1.4690910804179261e+01
RS_130 NS_130 0 1.4690910804179261e+01
GL_129 0 NS_129 NS_130 0 2.1320637363820186e-01
GL_130 0 NS_130 NS_129 0 -2.1320637363820186e-01
GS_129_7 0 NS_129 NA_7 0 6.0286980150450964e-01
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 1.6315799932686236e+01
RS_132 NS_132 0 1.6315799932686236e+01
GL_131 0 NS_131 NS_132 0 1.6372677698710228e-01
GL_132 0 NS_132 NS_131 0 -1.6372677698710228e-01
GS_131_7 0 NS_131 NA_7 0 6.0286980150450964e-01
*
* Complex pair n. 133/134
CS_133 NS_133 0 9.9999999999999998e-13
CS_134 NS_134 0 9.9999999999999998e-13
RS_133 NS_133 0 1.3805021583364081e+01
RS_134 NS_134 0 1.3805021583364081e+01
GL_133 0 NS_133 NS_134 0 1.3053652152390091e-01
GL_134 0 NS_134 NS_133 0 -1.3053652152390091e-01
GS_133_7 0 NS_133 NA_7 0 6.0286980150450964e-01
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 1.7453012154519879e+01
RS_136 NS_136 0 1.7453012154519879e+01
GL_135 0 NS_135 NS_136 0 8.4170507635427994e-02
GL_136 0 NS_136 NS_135 0 -8.4170507635427994e-02
GS_135_7 0 NS_135 NA_7 0 6.0286980150450964e-01
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 1.7836078439168801e+01
RS_138 NS_138 0 1.7836078439168805e+01
GL_137 0 NS_137 NS_138 0 5.3586142573527437e-02
GL_138 0 NS_138 NS_137 0 -5.3586142573527437e-02
GS_137_7 0 NS_137 NA_7 0 6.0286980150450964e-01
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 1.9366404748437819e+01
RS_140 NS_140 0 1.9366404748437819e+01
GL_139 0 NS_139 NS_140 0 2.0213646406074141e-02
GL_140 0 NS_140 NS_139 0 -2.0213646406074141e-02
GS_139_7 0 NS_139 NA_7 0 6.0286980150450964e-01
*
* Real pole n. 141
CS_141 NS_141 0 9.9999999999999998e-13
RS_141 NS_141 0 6.8759459879260660e+01
GS_141_8 0 NS_141 NA_8 0 6.0286980150450964e-01
*
* Real pole n. 142
CS_142 NS_142 0 9.9999999999999998e-13
RS_142 NS_142 0 2.4827714035206478e+02
GS_142_8 0 NS_142 NA_8 0 6.0286980150450964e-01
*
* Real pole n. 143
CS_143 NS_143 0 9.9999999999999998e-13
RS_143 NS_143 0 5.8935503054175797e+03
GS_143_8 0 NS_143 NA_8 0 6.0286980150450964e-01
*
* Real pole n. 144
CS_144 NS_144 0 9.9999999999999998e-13
RS_144 NS_144 0 1.2841015484081297e+03
GS_144_8 0 NS_144 NA_8 0 6.0286980150450964e-01
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 2.8319423052259118e+01
RS_146 NS_146 0 2.8319423052259115e+01
GL_145 0 NS_145 NS_146 0 3.0726343572183612e-01
GL_146 0 NS_146 NS_145 0 -3.0726343572183612e-01
GS_145_8 0 NS_145 NA_8 0 6.0286980150450964e-01
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 1.8367949753848961e+01
RS_148 NS_148 0 1.8367949753848965e+01
GL_147 0 NS_147 NS_148 0 2.4584800021674161e-01
GL_148 0 NS_148 NS_147 0 -2.4584800021674161e-01
GS_147_8 0 NS_147 NA_8 0 6.0286980150450964e-01
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 1.4690910804179261e+01
RS_150 NS_150 0 1.4690910804179261e+01
GL_149 0 NS_149 NS_150 0 2.1320637363820186e-01
GL_150 0 NS_150 NS_149 0 -2.1320637363820186e-01
GS_149_8 0 NS_149 NA_8 0 6.0286980150450964e-01
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 1.6315799932686236e+01
RS_152 NS_152 0 1.6315799932686236e+01
GL_151 0 NS_151 NS_152 0 1.6372677698710228e-01
GL_152 0 NS_152 NS_151 0 -1.6372677698710228e-01
GS_151_8 0 NS_151 NA_8 0 6.0286980150450964e-01
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 1.3805021583364081e+01
RS_154 NS_154 0 1.3805021583364081e+01
GL_153 0 NS_153 NS_154 0 1.3053652152390091e-01
GL_154 0 NS_154 NS_153 0 -1.3053652152390091e-01
GS_153_8 0 NS_153 NA_8 0 6.0286980150450964e-01
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 1.7453012154519879e+01
RS_156 NS_156 0 1.7453012154519879e+01
GL_155 0 NS_155 NS_156 0 8.4170507635427994e-02
GL_156 0 NS_156 NS_155 0 -8.4170507635427994e-02
GS_155_8 0 NS_155 NA_8 0 6.0286980150450964e-01
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 1.7836078439168801e+01
RS_158 NS_158 0 1.7836078439168805e+01
GL_157 0 NS_157 NS_158 0 5.3586142573527437e-02
GL_158 0 NS_158 NS_157 0 -5.3586142573527437e-02
GS_157_8 0 NS_157 NA_8 0 6.0286980150450964e-01
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 1.9366404748437819e+01
RS_160 NS_160 0 1.9366404748437819e+01
GL_159 0 NS_159 NS_160 0 2.0213646406074141e-02
GL_160 0 NS_160 NS_159 0 -2.0213646406074141e-02
GS_159_8 0 NS_159 NA_8 0 6.0286980150450964e-01
*
* Real pole n. 161
CS_161 NS_161 0 9.9999999999999998e-13
RS_161 NS_161 0 6.8759459879260660e+01
GS_161_9 0 NS_161 NA_9 0 6.0286980150450964e-01
*
* Real pole n. 162
CS_162 NS_162 0 9.9999999999999998e-13
RS_162 NS_162 0 2.4827714035206478e+02
GS_162_9 0 NS_162 NA_9 0 6.0286980150450964e-01
*
* Real pole n. 163
CS_163 NS_163 0 9.9999999999999998e-13
RS_163 NS_163 0 5.8935503054175797e+03
GS_163_9 0 NS_163 NA_9 0 6.0286980150450964e-01
*
* Real pole n. 164
CS_164 NS_164 0 9.9999999999999998e-13
RS_164 NS_164 0 1.2841015484081297e+03
GS_164_9 0 NS_164 NA_9 0 6.0286980150450964e-01
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 2.8319423052259118e+01
RS_166 NS_166 0 2.8319423052259115e+01
GL_165 0 NS_165 NS_166 0 3.0726343572183612e-01
GL_166 0 NS_166 NS_165 0 -3.0726343572183612e-01
GS_165_9 0 NS_165 NA_9 0 6.0286980150450964e-01
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 1.8367949753848961e+01
RS_168 NS_168 0 1.8367949753848965e+01
GL_167 0 NS_167 NS_168 0 2.4584800021674161e-01
GL_168 0 NS_168 NS_167 0 -2.4584800021674161e-01
GS_167_9 0 NS_167 NA_9 0 6.0286980150450964e-01
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 1.4690910804179261e+01
RS_170 NS_170 0 1.4690910804179261e+01
GL_169 0 NS_169 NS_170 0 2.1320637363820186e-01
GL_170 0 NS_170 NS_169 0 -2.1320637363820186e-01
GS_169_9 0 NS_169 NA_9 0 6.0286980150450964e-01
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 1.6315799932686236e+01
RS_172 NS_172 0 1.6315799932686236e+01
GL_171 0 NS_171 NS_172 0 1.6372677698710228e-01
GL_172 0 NS_172 NS_171 0 -1.6372677698710228e-01
GS_171_9 0 NS_171 NA_9 0 6.0286980150450964e-01
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 1.3805021583364081e+01
RS_174 NS_174 0 1.3805021583364081e+01
GL_173 0 NS_173 NS_174 0 1.3053652152390091e-01
GL_174 0 NS_174 NS_173 0 -1.3053652152390091e-01
GS_173_9 0 NS_173 NA_9 0 6.0286980150450964e-01
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 1.7453012154519879e+01
RS_176 NS_176 0 1.7453012154519879e+01
GL_175 0 NS_175 NS_176 0 8.4170507635427994e-02
GL_176 0 NS_176 NS_175 0 -8.4170507635427994e-02
GS_175_9 0 NS_175 NA_9 0 6.0286980150450964e-01
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 1.7836078439168801e+01
RS_178 NS_178 0 1.7836078439168805e+01
GL_177 0 NS_177 NS_178 0 5.3586142573527437e-02
GL_178 0 NS_178 NS_177 0 -5.3586142573527437e-02
GS_177_9 0 NS_177 NA_9 0 6.0286980150450964e-01
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 1.9366404748437819e+01
RS_180 NS_180 0 1.9366404748437819e+01
GL_179 0 NS_179 NS_180 0 2.0213646406074141e-02
GL_180 0 NS_180 NS_179 0 -2.0213646406074141e-02
GS_179_9 0 NS_179 NA_9 0 6.0286980150450964e-01
*
* Real pole n. 181
CS_181 NS_181 0 9.9999999999999998e-13
RS_181 NS_181 0 6.8759459879260660e+01
GS_181_10 0 NS_181 NA_10 0 6.0286980150450964e-01
*
* Real pole n. 182
CS_182 NS_182 0 9.9999999999999998e-13
RS_182 NS_182 0 2.4827714035206478e+02
GS_182_10 0 NS_182 NA_10 0 6.0286980150450964e-01
*
* Real pole n. 183
CS_183 NS_183 0 9.9999999999999998e-13
RS_183 NS_183 0 5.8935503054175797e+03
GS_183_10 0 NS_183 NA_10 0 6.0286980150450964e-01
*
* Real pole n. 184
CS_184 NS_184 0 9.9999999999999998e-13
RS_184 NS_184 0 1.2841015484081297e+03
GS_184_10 0 NS_184 NA_10 0 6.0286980150450964e-01
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 2.8319423052259118e+01
RS_186 NS_186 0 2.8319423052259115e+01
GL_185 0 NS_185 NS_186 0 3.0726343572183612e-01
GL_186 0 NS_186 NS_185 0 -3.0726343572183612e-01
GS_185_10 0 NS_185 NA_10 0 6.0286980150450964e-01
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 1.8367949753848961e+01
RS_188 NS_188 0 1.8367949753848965e+01
GL_187 0 NS_187 NS_188 0 2.4584800021674161e-01
GL_188 0 NS_188 NS_187 0 -2.4584800021674161e-01
GS_187_10 0 NS_187 NA_10 0 6.0286980150450964e-01
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 1.4690910804179261e+01
RS_190 NS_190 0 1.4690910804179261e+01
GL_189 0 NS_189 NS_190 0 2.1320637363820186e-01
GL_190 0 NS_190 NS_189 0 -2.1320637363820186e-01
GS_189_10 0 NS_189 NA_10 0 6.0286980150450964e-01
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 1.6315799932686236e+01
RS_192 NS_192 0 1.6315799932686236e+01
GL_191 0 NS_191 NS_192 0 1.6372677698710228e-01
GL_192 0 NS_192 NS_191 0 -1.6372677698710228e-01
GS_191_10 0 NS_191 NA_10 0 6.0286980150450964e-01
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 1.3805021583364081e+01
RS_194 NS_194 0 1.3805021583364081e+01
GL_193 0 NS_193 NS_194 0 1.3053652152390091e-01
GL_194 0 NS_194 NS_193 0 -1.3053652152390091e-01
GS_193_10 0 NS_193 NA_10 0 6.0286980150450964e-01
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 1.7453012154519879e+01
RS_196 NS_196 0 1.7453012154519879e+01
GL_195 0 NS_195 NS_196 0 8.4170507635427994e-02
GL_196 0 NS_196 NS_195 0 -8.4170507635427994e-02
GS_195_10 0 NS_195 NA_10 0 6.0286980150450964e-01
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 1.7836078439168801e+01
RS_198 NS_198 0 1.7836078439168805e+01
GL_197 0 NS_197 NS_198 0 5.3586142573527437e-02
GL_198 0 NS_198 NS_197 0 -5.3586142573527437e-02
GS_197_10 0 NS_197 NA_10 0 6.0286980150450964e-01
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 1.9366404748437819e+01
RS_200 NS_200 0 1.9366404748437819e+01
GL_199 0 NS_199 NS_200 0 2.0213646406074141e-02
GL_200 0 NS_200 NS_199 0 -2.0213646406074141e-02
GS_199_10 0 NS_199 NA_10 0 6.0286980150450964e-01
*
* Real pole n. 201
CS_201 NS_201 0 9.9999999999999998e-13
RS_201 NS_201 0 6.8759459879260660e+01
GS_201_11 0 NS_201 NA_11 0 6.0286980150450964e-01
*
* Real pole n. 202
CS_202 NS_202 0 9.9999999999999998e-13
RS_202 NS_202 0 2.4827714035206478e+02
GS_202_11 0 NS_202 NA_11 0 6.0286980150450964e-01
*
* Real pole n. 203
CS_203 NS_203 0 9.9999999999999998e-13
RS_203 NS_203 0 5.8935503054175797e+03
GS_203_11 0 NS_203 NA_11 0 6.0286980150450964e-01
*
* Real pole n. 204
CS_204 NS_204 0 9.9999999999999998e-13
RS_204 NS_204 0 1.2841015484081297e+03
GS_204_11 0 NS_204 NA_11 0 6.0286980150450964e-01
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 2.8319423052259118e+01
RS_206 NS_206 0 2.8319423052259115e+01
GL_205 0 NS_205 NS_206 0 3.0726343572183612e-01
GL_206 0 NS_206 NS_205 0 -3.0726343572183612e-01
GS_205_11 0 NS_205 NA_11 0 6.0286980150450964e-01
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 1.8367949753848961e+01
RS_208 NS_208 0 1.8367949753848965e+01
GL_207 0 NS_207 NS_208 0 2.4584800021674161e-01
GL_208 0 NS_208 NS_207 0 -2.4584800021674161e-01
GS_207_11 0 NS_207 NA_11 0 6.0286980150450964e-01
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 1.4690910804179261e+01
RS_210 NS_210 0 1.4690910804179261e+01
GL_209 0 NS_209 NS_210 0 2.1320637363820186e-01
GL_210 0 NS_210 NS_209 0 -2.1320637363820186e-01
GS_209_11 0 NS_209 NA_11 0 6.0286980150450964e-01
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 1.6315799932686236e+01
RS_212 NS_212 0 1.6315799932686236e+01
GL_211 0 NS_211 NS_212 0 1.6372677698710228e-01
GL_212 0 NS_212 NS_211 0 -1.6372677698710228e-01
GS_211_11 0 NS_211 NA_11 0 6.0286980150450964e-01
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 1.3805021583364081e+01
RS_214 NS_214 0 1.3805021583364081e+01
GL_213 0 NS_213 NS_214 0 1.3053652152390091e-01
GL_214 0 NS_214 NS_213 0 -1.3053652152390091e-01
GS_213_11 0 NS_213 NA_11 0 6.0286980150450964e-01
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 1.7453012154519879e+01
RS_216 NS_216 0 1.7453012154519879e+01
GL_215 0 NS_215 NS_216 0 8.4170507635427994e-02
GL_216 0 NS_216 NS_215 0 -8.4170507635427994e-02
GS_215_11 0 NS_215 NA_11 0 6.0286980150450964e-01
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 1.7836078439168801e+01
RS_218 NS_218 0 1.7836078439168805e+01
GL_217 0 NS_217 NS_218 0 5.3586142573527437e-02
GL_218 0 NS_218 NS_217 0 -5.3586142573527437e-02
GS_217_11 0 NS_217 NA_11 0 6.0286980150450964e-01
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 1.9366404748437819e+01
RS_220 NS_220 0 1.9366404748437819e+01
GL_219 0 NS_219 NS_220 0 2.0213646406074141e-02
GL_220 0 NS_220 NS_219 0 -2.0213646406074141e-02
GS_219_11 0 NS_219 NA_11 0 6.0286980150450964e-01
*
* Real pole n. 221
CS_221 NS_221 0 9.9999999999999998e-13
RS_221 NS_221 0 6.8759459879260660e+01
GS_221_12 0 NS_221 NA_12 0 6.0286980150450964e-01
*
* Real pole n. 222
CS_222 NS_222 0 9.9999999999999998e-13
RS_222 NS_222 0 2.4827714035206478e+02
GS_222_12 0 NS_222 NA_12 0 6.0286980150450964e-01
*
* Real pole n. 223
CS_223 NS_223 0 9.9999999999999998e-13
RS_223 NS_223 0 5.8935503054175797e+03
GS_223_12 0 NS_223 NA_12 0 6.0286980150450964e-01
*
* Real pole n. 224
CS_224 NS_224 0 9.9999999999999998e-13
RS_224 NS_224 0 1.2841015484081297e+03
GS_224_12 0 NS_224 NA_12 0 6.0286980150450964e-01
*
* Complex pair n. 225/226
CS_225 NS_225 0 9.9999999999999998e-13
CS_226 NS_226 0 9.9999999999999998e-13
RS_225 NS_225 0 2.8319423052259118e+01
RS_226 NS_226 0 2.8319423052259115e+01
GL_225 0 NS_225 NS_226 0 3.0726343572183612e-01
GL_226 0 NS_226 NS_225 0 -3.0726343572183612e-01
GS_225_12 0 NS_225 NA_12 0 6.0286980150450964e-01
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 1.8367949753848961e+01
RS_228 NS_228 0 1.8367949753848965e+01
GL_227 0 NS_227 NS_228 0 2.4584800021674161e-01
GL_228 0 NS_228 NS_227 0 -2.4584800021674161e-01
GS_227_12 0 NS_227 NA_12 0 6.0286980150450964e-01
*
* Complex pair n. 229/230
CS_229 NS_229 0 9.9999999999999998e-13
CS_230 NS_230 0 9.9999999999999998e-13
RS_229 NS_229 0 1.4690910804179261e+01
RS_230 NS_230 0 1.4690910804179261e+01
GL_229 0 NS_229 NS_230 0 2.1320637363820186e-01
GL_230 0 NS_230 NS_229 0 -2.1320637363820186e-01
GS_229_12 0 NS_229 NA_12 0 6.0286980150450964e-01
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 1.6315799932686236e+01
RS_232 NS_232 0 1.6315799932686236e+01
GL_231 0 NS_231 NS_232 0 1.6372677698710228e-01
GL_232 0 NS_232 NS_231 0 -1.6372677698710228e-01
GS_231_12 0 NS_231 NA_12 0 6.0286980150450964e-01
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 1.3805021583364081e+01
RS_234 NS_234 0 1.3805021583364081e+01
GL_233 0 NS_233 NS_234 0 1.3053652152390091e-01
GL_234 0 NS_234 NS_233 0 -1.3053652152390091e-01
GS_233_12 0 NS_233 NA_12 0 6.0286980150450964e-01
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 1.7453012154519879e+01
RS_236 NS_236 0 1.7453012154519879e+01
GL_235 0 NS_235 NS_236 0 8.4170507635427994e-02
GL_236 0 NS_236 NS_235 0 -8.4170507635427994e-02
GS_235_12 0 NS_235 NA_12 0 6.0286980150450964e-01
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 1.7836078439168801e+01
RS_238 NS_238 0 1.7836078439168805e+01
GL_237 0 NS_237 NS_238 0 5.3586142573527437e-02
GL_238 0 NS_238 NS_237 0 -5.3586142573527437e-02
GS_237_12 0 NS_237 NA_12 0 6.0286980150450964e-01
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 1.9366404748437819e+01
RS_240 NS_240 0 1.9366404748437819e+01
GL_239 0 NS_239 NS_240 0 2.0213646406074141e-02
GL_240 0 NS_240 NS_239 0 -2.0213646406074141e-02
GS_239_12 0 NS_239 NA_12 0 6.0286980150450964e-01
*
******************************


.ends
*******************
* End of subcircuit
*******************
