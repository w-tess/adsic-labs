**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [8 2 26] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_8_Module_wire_1mm_highloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 5.9934852708580545e-02
GC_1_2 b_1 NI_1 NS_2 0 -6.4654666394797083e-02
GC_1_3 b_1 NI_1 NS_3 0 -1.0233466126531187e-08
GC_1_4 b_1 NI_1 NS_4 0 -8.1983893351230079e-06
GC_1_5 b_1 NI_1 NS_5 0 -1.8758516813947932e-03
GC_1_6 b_1 NI_1 NS_6 0 -2.8706548412248973e-03
GC_1_7 b_1 NI_1 NS_7 0 -5.0998746470950910e-03
GC_1_8 b_1 NI_1 NS_8 0 1.9265479434409979e-03
GC_1_9 b_1 NI_1 NS_9 0 2.3837856116197599e-03
GC_1_10 b_1 NI_1 NS_10 0 -1.2477161950727601e-03
GC_1_11 b_1 NI_1 NS_11 0 -1.0661875966280447e-02
GC_1_12 b_1 NI_1 NS_12 0 1.1356529007343014e-03
GC_1_13 b_1 NI_1 NS_13 0 5.9634237015429538e-04
GC_1_14 b_1 NI_1 NS_14 0 1.7470517300509183e-03
GC_1_15 b_1 NI_1 NS_15 0 -9.6080888142928628e-04
GC_1_16 b_1 NI_1 NS_16 0 2.2969430138115262e-03
GC_1_17 b_1 NI_1 NS_17 0 5.3288097254274849e-04
GC_1_18 b_1 NI_1 NS_18 0 -5.8517879729081288e-03
GC_1_19 b_1 NI_1 NS_19 0 -8.5170547035245733e-03
GC_1_20 b_1 NI_1 NS_20 0 6.9045156927713706e-03
GC_1_21 b_1 NI_1 NS_21 0 2.5028306563983052e-03
GC_1_22 b_1 NI_1 NS_22 0 -3.6531650313559589e-03
GC_1_23 b_1 NI_1 NS_23 0 -2.5960265715554063e-03
GC_1_24 b_1 NI_1 NS_24 0 -5.3416983383630114e-04
GC_1_25 b_1 NI_1 NS_25 0 5.5354219558516306e-02
GC_1_26 b_1 NI_1 NS_26 0 1.8152608436065765e-03
GC_1_27 b_1 NI_1 NS_27 0 -5.0037226484896564e-02
GC_1_28 b_1 NI_1 NS_28 0 1.1076316952712911e-01
GC_1_29 b_1 NI_1 NS_29 0 1.1664253666469057e-08
GC_1_30 b_1 NI_1 NS_30 0 1.9861991793363391e-05
GC_1_31 b_1 NI_1 NS_31 0 -1.5739399321699425e-02
GC_1_32 b_1 NI_1 NS_32 0 2.4245664459279226e-02
GC_1_33 b_1 NI_1 NS_33 0 -7.8711120417003372e-03
GC_1_34 b_1 NI_1 NS_34 0 -1.4518767529591159e-02
GC_1_35 b_1 NI_1 NS_35 0 2.0325307732110536e-02
GC_1_36 b_1 NI_1 NS_36 0 6.6761255262385074e-03
GC_1_37 b_1 NI_1 NS_37 0 8.0658958356082562e-03
GC_1_38 b_1 NI_1 NS_38 0 4.4188585472529199e-02
GC_1_39 b_1 NI_1 NS_39 0 -1.1822666597684557e-02
GC_1_40 b_1 NI_1 NS_40 0 -3.1939241141848000e-03
GC_1_41 b_1 NI_1 NS_41 0 -5.1132719171693864e-03
GC_1_42 b_1 NI_1 NS_42 0 -4.0785569663554719e-03
GC_1_43 b_1 NI_1 NS_43 0 2.6802328466686398e-02
GC_1_44 b_1 NI_1 NS_44 0 1.2877213175474251e-04
GC_1_45 b_1 NI_1 NS_45 0 3.4101237119214825e-02
GC_1_46 b_1 NI_1 NS_46 0 3.1057523598419075e-02
GC_1_47 b_1 NI_1 NS_47 0 -1.5591733834292548e-02
GC_1_48 b_1 NI_1 NS_48 0 8.2163404205307707e-03
GC_1_49 b_1 NI_1 NS_49 0 -1.0700819399029685e-03
GC_1_50 b_1 NI_1 NS_50 0 -6.8532030435006627e-03
GC_1_51 b_1 NI_1 NS_51 0 -6.9887930908103357e-02
GC_1_52 b_1 NI_1 NS_52 0 1.6945028597021093e-03
GC_1_53 b_1 NI_1 NS_53 0 -7.4986630406882046e-03
GC_1_54 b_1 NI_1 NS_54 0 5.4463679169777113e-03
GC_1_55 b_1 NI_1 NS_55 0 -8.2819008038075067e-10
GC_1_56 b_1 NI_1 NS_56 0 -1.6858207847886790e-06
GC_1_57 b_1 NI_1 NS_57 0 2.5534451679427156e-04
GC_1_58 b_1 NI_1 NS_58 0 2.6645209554603607e-03
GC_1_59 b_1 NI_1 NS_59 0 4.5291717763011304e-03
GC_1_60 b_1 NI_1 NS_60 0 -2.7565535280063124e-03
GC_1_61 b_1 NI_1 NS_61 0 -5.4227002238950751e-03
GC_1_62 b_1 NI_1 NS_62 0 4.2041125753595278e-04
GC_1_63 b_1 NI_1 NS_63 0 8.8584598590663761e-03
GC_1_64 b_1 NI_1 NS_64 0 -6.2093760062330880e-04
GC_1_65 b_1 NI_1 NS_65 0 -2.8260892311363865e-03
GC_1_66 b_1 NI_1 NS_66 0 -2.3963222379300739e-03
GC_1_67 b_1 NI_1 NS_67 0 4.3105191748288669e-05
GC_1_68 b_1 NI_1 NS_68 0 -2.1139049360767801e-03
GC_1_69 b_1 NI_1 NS_69 0 -3.5070335195684062e-03
GC_1_70 b_1 NI_1 NS_70 0 5.5496239602017506e-03
GC_1_71 b_1 NI_1 NS_71 0 5.0984928002371400e-03
GC_1_72 b_1 NI_1 NS_72 0 -7.7604182478625263e-03
GC_1_73 b_1 NI_1 NS_73 0 -5.0389112787701555e-03
GC_1_74 b_1 NI_1 NS_74 0 3.0962138594566643e-03
GC_1_75 b_1 NI_1 NS_75 0 2.2446237576854038e-03
GC_1_76 b_1 NI_1 NS_76 0 -1.6873402428930846e-03
GC_1_77 b_1 NI_1 NS_77 0 -5.9469780546735291e-03
GC_1_78 b_1 NI_1 NS_78 0 3.8164552896847643e-03
GC_1_79 b_1 NI_1 NS_79 0 -1.3745899584277240e-03
GC_1_80 b_1 NI_1 NS_80 0 2.3328611511893287e-03
GC_1_81 b_1 NI_1 NS_81 0 7.5881727199374062e-10
GC_1_82 b_1 NI_1 NS_82 0 6.0065849244273874e-07
GC_1_83 b_1 NI_1 NS_83 0 -1.9596182586423825e-04
GC_1_84 b_1 NI_1 NS_84 0 -4.5534379655177878e-04
GC_1_85 b_1 NI_1 NS_85 0 -1.0665912540998624e-03
GC_1_86 b_1 NI_1 NS_86 0 -9.2132098612694681e-04
GC_1_87 b_1 NI_1 NS_87 0 -2.3173781109475668e-03
GC_1_88 b_1 NI_1 NS_88 0 3.1222785727115347e-04
GC_1_89 b_1 NI_1 NS_89 0 -3.4635653562912024e-04
GC_1_90 b_1 NI_1 NS_90 0 4.1981806371535566e-03
GC_1_91 b_1 NI_1 NS_91 0 9.7829065528359294e-04
GC_1_92 b_1 NI_1 NS_92 0 4.4367094388938669e-04
GC_1_93 b_1 NI_1 NS_93 0 -3.7329437083758268e-04
GC_1_94 b_1 NI_1 NS_94 0 7.9842631251566182e-05
GC_1_95 b_1 NI_1 NS_95 0 -3.1453545432697785e-04
GC_1_96 b_1 NI_1 NS_96 0 3.3540627908027420e-03
GC_1_97 b_1 NI_1 NS_97 0 5.2329373467686702e-03
GC_1_98 b_1 NI_1 NS_98 0 8.1284762372159727e-04
GC_1_99 b_1 NI_1 NS_99 0 1.3427520051352494e-03
GC_1_100 b_1 NI_1 NS_100 0 -1.9440147232562732e-03
GC_1_101 b_1 NI_1 NS_101 0 -8.8256310685517678e-04
GC_1_102 b_1 NI_1 NS_102 0 -6.3689546500520075e-04
GC_1_103 b_1 NI_1 NS_103 0 -1.4735533079394830e-03
GC_1_104 b_1 NI_1 NS_104 0 2.5664393804470035e-03
GC_1_105 b_1 NI_1 NS_105 0 3.9579046841301961e-04
GC_1_106 b_1 NI_1 NS_106 0 -2.0177620426844035e-03
GC_1_107 b_1 NI_1 NS_107 0 4.0760489900537490e-10
GC_1_108 b_1 NI_1 NS_108 0 -2.7072352122339902e-08
GC_1_109 b_1 NI_1 NS_109 0 1.8516035442806561e-05
GC_1_110 b_1 NI_1 NS_110 0 4.3377996232983926e-05
GC_1_111 b_1 NI_1 NS_111 0 8.1709677252975028e-05
GC_1_112 b_1 NI_1 NS_112 0 -3.0786352460080713e-05
GC_1_113 b_1 NI_1 NS_113 0 -1.3938884275204685e-05
GC_1_114 b_1 NI_1 NS_114 0 1.3650823884046396e-05
GC_1_115 b_1 NI_1 NS_115 0 1.9708922258612012e-04
GC_1_116 b_1 NI_1 NS_116 0 -9.8902008669821720e-05
GC_1_117 b_1 NI_1 NS_117 0 2.6744128272535009e-05
GC_1_118 b_1 NI_1 NS_118 0 -9.8059736628299107e-05
GC_1_119 b_1 NI_1 NS_119 0 -1.7490356617592001e-05
GC_1_120 b_1 NI_1 NS_120 0 -9.8091727031117634e-05
GC_1_121 b_1 NI_1 NS_121 0 9.8222350089192871e-06
GC_1_122 b_1 NI_1 NS_122 0 -9.7469478884276077e-05
GC_1_123 b_1 NI_1 NS_123 0 -9.8112201637410326e-05
GC_1_124 b_1 NI_1 NS_124 0 -3.1491541481183021e-04
GC_1_125 b_1 NI_1 NS_125 0 -1.3398287914741599e-04
GC_1_126 b_1 NI_1 NS_126 0 -1.1516245581740061e-04
GC_1_127 b_1 NI_1 NS_127 0 -1.9658470553434173e-05
GC_1_128 b_1 NI_1 NS_128 0 -1.9129802535379712e-04
GC_1_129 b_1 NI_1 NS_129 0 1.5212419498496677e-03
GC_1_130 b_1 NI_1 NS_130 0 -1.0185248679477031e-04
GC_1_131 b_1 NI_1 NS_131 0 1.5161330790076802e-04
GC_1_132 b_1 NI_1 NS_132 0 1.2758700896356437e-05
GC_1_133 b_1 NI_1 NS_133 0 -4.2742748849413949e-10
GC_1_134 b_1 NI_1 NS_134 0 4.5130525445575852e-08
GC_1_135 b_1 NI_1 NS_135 0 5.1582436663319681e-06
GC_1_136 b_1 NI_1 NS_136 0 7.5618140313775661e-05
GC_1_137 b_1 NI_1 NS_137 0 1.5335293772442113e-04
GC_1_138 b_1 NI_1 NS_138 0 1.3548425749522168e-04
GC_1_139 b_1 NI_1 NS_139 0 3.4656235527258671e-04
GC_1_140 b_1 NI_1 NS_140 0 -2.4743470012727381e-05
GC_1_141 b_1 NI_1 NS_141 0 5.1564520132888965e-05
GC_1_142 b_1 NI_1 NS_142 0 -5.8538770169051736e-04
GC_1_143 b_1 NI_1 NS_143 0 -1.4593695877479379e-04
GC_1_144 b_1 NI_1 NS_144 0 -6.8387289077554816e-05
GC_1_145 b_1 NI_1 NS_145 0 5.1712590847580669e-05
GC_1_146 b_1 NI_1 NS_146 0 -1.0508142888271244e-05
GC_1_147 b_1 NI_1 NS_147 0 4.7728655399018796e-05
GC_1_148 b_1 NI_1 NS_148 0 -4.5313210255697417e-04
GC_1_149 b_1 NI_1 NS_149 0 -7.0919247467915241e-04
GC_1_150 b_1 NI_1 NS_150 0 -8.3324118916299798e-05
GC_1_151 b_1 NI_1 NS_151 0 -1.7472496307247920e-04
GC_1_152 b_1 NI_1 NS_152 0 2.5870543259387221e-04
GC_1_153 b_1 NI_1 NS_153 0 1.0249916233569625e-04
GC_1_154 b_1 NI_1 NS_154 0 7.9809616708275628e-05
GC_1_155 b_1 NI_1 NS_155 0 -8.6720212128168909e-05
GC_1_156 b_1 NI_1 NS_156 0 -3.2996574262481629e-04
GC_1_157 b_1 NI_1 NS_157 0 -1.4356179722763130e-04
GC_1_158 b_1 NI_1 NS_158 0 6.6680320165499586e-04
GC_1_159 b_1 NI_1 NS_159 0 1.2440048262609677e-10
GC_1_160 b_1 NI_1 NS_160 0 -1.1384117274677266e-08
GC_1_161 b_1 NI_1 NS_161 0 -4.0172023090946738e-06
GC_1_162 b_1 NI_1 NS_162 0 -3.9916826629699495e-06
GC_1_163 b_1 NI_1 NS_163 0 -9.5853548007179893e-06
GC_1_164 b_1 NI_1 NS_164 0 -3.6874511784250466e-06
GC_1_165 b_1 NI_1 NS_165 0 -1.8731365441771954e-05
GC_1_166 b_1 NI_1 NS_166 0 -1.5342447691446096e-06
GC_1_167 b_1 NI_1 NS_167 0 -2.9271382837994811e-05
GC_1_168 b_1 NI_1 NS_168 0 2.7762771224331745e-05
GC_1_169 b_1 NI_1 NS_169 0 -2.1467904870280413e-05
GC_1_170 b_1 NI_1 NS_170 0 2.3556682983001287e-05
GC_1_171 b_1 NI_1 NS_171 0 6.1042869269607898e-06
GC_1_172 b_1 NI_1 NS_172 0 2.3439073137350275e-05
GC_1_173 b_1 NI_1 NS_173 0 -1.5895569095232862e-05
GC_1_174 b_1 NI_1 NS_174 0 5.5646866024925880e-05
GC_1_175 b_1 NI_1 NS_175 0 5.4417167331589520e-05
GC_1_176 b_1 NI_1 NS_176 0 6.5745678093507060e-05
GC_1_177 b_1 NI_1 NS_177 0 2.2593743191363518e-05
GC_1_178 b_1 NI_1 NS_178 0 4.5701641257726147e-05
GC_1_179 b_1 NI_1 NS_179 0 1.4942119515018684e-05
GC_1_180 b_1 NI_1 NS_180 0 4.9676076844950538e-05
GC_1_181 b_1 NI_1 NS_181 0 -5.1914710084349205e-04
GC_1_182 b_1 NI_1 NS_182 0 2.3890391099276964e-05
GC_1_183 b_1 NI_1 NS_183 0 -1.6380544611059055e-05
GC_1_184 b_1 NI_1 NS_184 0 -2.5702748792450663e-04
GC_1_185 b_1 NI_1 NS_185 0 -1.0826082679566479e-10
GC_1_186 b_1 NI_1 NS_186 0 4.7604531738260291e-09
GC_1_187 b_1 NI_1 NS_187 0 5.0802163161341772e-06
GC_1_188 b_1 NI_1 NS_188 0 9.6641027485829651e-06
GC_1_189 b_1 NI_1 NS_189 0 1.6473271665657563e-05
GC_1_190 b_1 NI_1 NS_190 0 1.3380149178603419e-05
GC_1_191 b_1 NI_1 NS_191 0 3.8420504254042955e-05
GC_1_192 b_1 NI_1 NS_192 0 -3.4928781919300877e-06
GC_1_193 b_1 NI_1 NS_193 0 1.4578073279133500e-05
GC_1_194 b_1 NI_1 NS_194 0 -6.2742694775200605e-05
GC_1_195 b_1 NI_1 NS_195 0 -1.1726885495882127e-05
GC_1_196 b_1 NI_1 NS_196 0 -9.0423434813204269e-06
GC_1_197 b_1 NI_1 NS_197 0 4.7447311751861810e-06
GC_1_198 b_1 NI_1 NS_198 0 -3.4993438124508949e-06
GC_1_199 b_1 NI_1 NS_199 0 9.7146746779431202e-06
GC_1_200 b_1 NI_1 NS_200 0 -5.0075302312417671e-05
GC_1_201 b_1 NI_1 NS_201 0 -6.6281364862631262e-05
GC_1_202 b_1 NI_1 NS_202 0 -2.1644694838285235e-05
GC_1_203 b_1 NI_1 NS_203 0 -1.6781843250420172e-05
GC_1_204 b_1 NI_1 NS_204 0 1.9314782077212255e-05
GC_1_205 b_1 NI_1 NS_205 0 1.6170796069631956e-05
GC_1_206 b_1 NI_1 NS_206 0 -1.3552352443299523e-06
GC_1_207 b_1 NI_1 NS_207 0 2.1848252754323478e-04
GC_1_208 b_1 NI_1 NS_208 0 7.6250188103439023e-06
GC_1_209 b_1 NI_1 NS_209 0 -2.7914673538223890e-05
GC_1_210 b_1 NI_1 NS_210 0 4.2480930955795539e-05
GC_1_211 b_1 NI_1 NS_211 0 3.6704873052262727e-11
GC_1_212 b_1 NI_1 NS_212 0 -2.7830065314644110e-10
GC_1_213 b_1 NI_1 NS_213 0 8.4367570954064381e-07
GC_1_214 b_1 NI_1 NS_214 0 4.8587722126687397e-07
GC_1_215 b_1 NI_1 NS_215 0 4.0290826542445129e-07
GC_1_216 b_1 NI_1 NS_216 0 -7.5371184311782107e-07
GC_1_217 b_1 NI_1 NS_217 0 -4.7578260464272994e-07
GC_1_218 b_1 NI_1 NS_218 0 9.9272452909558531e-07
GC_1_219 b_1 NI_1 NS_219 0 1.4092607134040200e-06
GC_1_220 b_1 NI_1 NS_220 0 1.8306206305212611e-07
GC_1_221 b_1 NI_1 NS_221 0 -4.2142650679951912e-07
GC_1_222 b_1 NI_1 NS_222 0 9.6875599445416464e-07
GC_1_223 b_1 NI_1 NS_223 0 5.7216895828136375e-07
GC_1_224 b_1 NI_1 NS_224 0 3.8282399404816205e-07
GC_1_225 b_1 NI_1 NS_225 0 5.5915977596157146e-07
GC_1_226 b_1 NI_1 NS_226 0 3.2458444072138624e-06
GC_1_227 b_1 NI_1 NS_227 0 4.0017169902102109e-06
GC_1_228 b_1 NI_1 NS_228 0 7.8432543068450710e-07
GC_1_229 b_1 NI_1 NS_229 0 9.0407613617344216e-07
GC_1_230 b_1 NI_1 NS_230 0 2.3922783613283715e-06
GC_1_231 b_1 NI_1 NS_231 0 1.1489417122555005e-06
GC_1_232 b_1 NI_1 NS_232 0 2.6151368145148415e-06
GC_1_233 b_1 NI_1 NS_233 0 -3.3615793333449168e-05
GC_1_234 b_1 NI_1 NS_234 0 4.1019974553364572e-07
GC_1_235 b_1 NI_1 NS_235 0 -2.4824765795583510e-05
GC_1_236 b_1 NI_1 NS_236 0 2.0783343812725676e-05
GC_1_237 b_1 NI_1 NS_237 0 -3.5006743958516238e-11
GC_1_238 b_1 NI_1 NS_238 0 -2.7089686914325185e-10
GC_1_239 b_1 NI_1 NS_239 0 1.6165286014681214e-06
GC_1_240 b_1 NI_1 NS_240 0 1.4394623648791514e-06
GC_1_241 b_1 NI_1 NS_241 0 2.5877681245395076e-07
GC_1_242 b_1 NI_1 NS_242 0 3.7182417152775981e-07
GC_1_243 b_1 NI_1 NS_243 0 1.7412280237372345e-06
GC_1_244 b_1 NI_1 NS_244 0 -2.0422220147307598e-07
GC_1_245 b_1 NI_1 NS_245 0 3.3659170384598686e-06
GC_1_246 b_1 NI_1 NS_246 0 -1.0270818601283743e-06
GC_1_247 b_1 NI_1 NS_247 0 4.2248035198067469e-07
GC_1_248 b_1 NI_1 NS_248 0 5.0189508004702002e-08
GC_1_249 b_1 NI_1 NS_249 0 2.5404315377544153e-07
GC_1_250 b_1 NI_1 NS_250 0 -2.9664617281188202e-07
GC_1_251 b_1 NI_1 NS_251 0 1.0839712693567370e-06
GC_1_252 b_1 NI_1 NS_252 0 -1.0041649501647894e-06
GC_1_253 b_1 NI_1 NS_253 0 1.6346566786296686e-06
GC_1_254 b_1 NI_1 NS_254 0 -1.2123161348136140e-06
GC_1_255 b_1 NI_1 NS_255 0 -5.8140746474907077e-08
GC_1_256 b_1 NI_1 NS_256 0 1.3019229587589354e-06
GC_1_257 b_1 NI_1 NS_257 0 3.3326943794327367e-07
GC_1_258 b_1 NI_1 NS_258 0 6.8673196801439136e-07
GC_1_259 b_1 NI_1 NS_259 0 -1.6980527964401524e-05
GC_1_260 b_1 NI_1 NS_260 0 -1.3435378273755001e-06
GC_1_261 b_1 NI_1 NS_261 0 -3.5487274396073843e-05
GC_1_262 b_1 NI_1 NS_262 0 4.3755692754004142e-05
GC_1_263 b_1 NI_1 NS_263 0 3.2703454565006975e-11
GC_1_264 b_1 NI_1 NS_264 0 -2.6824524670367912e-10
GC_1_265 b_1 NI_1 NS_265 0 1.0320796335245109e-06
GC_1_266 b_1 NI_1 NS_266 0 1.0605761593753714e-06
GC_1_267 b_1 NI_1 NS_267 0 1.7241338653784269e-06
GC_1_268 b_1 NI_1 NS_268 0 2.5964966358778387e-07
GC_1_269 b_1 NI_1 NS_269 0 1.0932111870167575e-06
GC_1_270 b_1 NI_1 NS_270 0 4.6059834254557620e-07
GC_1_271 b_1 NI_1 NS_271 0 2.9262620374096485e-06
GC_1_272 b_1 NI_1 NS_272 0 -4.3423253763669686e-07
GC_1_273 b_1 NI_1 NS_273 0 1.0132358677584838e-06
GC_1_274 b_1 NI_1 NS_274 0 5.3040535525338713e-09
GC_1_275 b_1 NI_1 NS_275 0 5.6285421835608502e-07
GC_1_276 b_1 NI_1 NS_276 0 -5.1625015573721805e-07
GC_1_277 b_1 NI_1 NS_277 0 1.6607430311026074e-06
GC_1_278 b_1 NI_1 NS_278 0 1.2910023897289594e-06
GC_1_279 b_1 NI_1 NS_279 0 2.8544590193673197e-06
GC_1_280 b_1 NI_1 NS_280 0 -1.2126692053098731e-06
GC_1_281 b_1 NI_1 NS_281 0 5.5986017256327180e-07
GC_1_282 b_1 NI_1 NS_282 0 1.1266010307485474e-06
GC_1_283 b_1 NI_1 NS_283 0 3.9045704721986212e-07
GC_1_284 b_1 NI_1 NS_284 0 1.5530727267952819e-06
GC_1_285 b_1 NI_1 NS_285 0 -3.6623114513638729e-05
GC_1_286 b_1 NI_1 NS_286 0 -3.7034576261482223e-06
GC_1_287 b_1 NI_1 NS_287 0 -1.1812994762128251e-05
GC_1_288 b_1 NI_1 NS_288 0 -5.5505898164968951e-06
GC_1_289 b_1 NI_1 NS_289 0 -3.0498030833888361e-11
GC_1_290 b_1 NI_1 NS_290 0 -1.3578566148752022e-10
GC_1_291 b_1 NI_1 NS_291 0 2.2976200171067841e-06
GC_1_292 b_1 NI_1 NS_292 0 1.7808637438308581e-06
GC_1_293 b_1 NI_1 NS_293 0 -6.4157924702450734e-07
GC_1_294 b_1 NI_1 NS_294 0 -3.8592712035544975e-07
GC_1_295 b_1 NI_1 NS_295 0 1.5505334447702363e-06
GC_1_296 b_1 NI_1 NS_296 0 -1.1518041682661032e-06
GC_1_297 b_1 NI_1 NS_297 0 1.8453794274492540e-06
GC_1_298 b_1 NI_1 NS_298 0 -4.3341838029909668e-07
GC_1_299 b_1 NI_1 NS_299 0 1.1932614477301316e-07
GC_1_300 b_1 NI_1 NS_300 0 -1.8767493446440110e-07
GC_1_301 b_1 NI_1 NS_301 0 5.5237203136157187e-08
GC_1_302 b_1 NI_1 NS_302 0 -3.1791031765603650e-07
GC_1_303 b_1 NI_1 NS_303 0 4.3573534421387249e-07
GC_1_304 b_1 NI_1 NS_304 0 -7.3740226441351977e-07
GC_1_305 b_1 NI_1 NS_305 0 9.1579267436966602e-07
GC_1_306 b_1 NI_1 NS_306 0 -1.3980117379597981e-06
GC_1_307 b_1 NI_1 NS_307 0 -1.8989909310324351e-07
GC_1_308 b_1 NI_1 NS_308 0 5.9848221669008170e-07
GC_1_309 b_1 NI_1 NS_309 0 3.5032407917798084e-07
GC_1_310 b_1 NI_1 NS_310 0 -1.4440495065055061e-08
GC_1_311 b_1 NI_1 NS_311 0 5.7887411022479193e-06
GC_1_312 b_1 NI_1 NS_312 0 2.3957892356863284e-06
GD_1_1 b_1 NI_1 NA_1 0 -2.9881630529505113e-02
GD_1_2 b_1 NI_1 NA_2 0 -2.0539317609763928e-02
GD_1_3 b_1 NI_1 NA_3 0 1.3427304153556941e-02
GD_1_4 b_1 NI_1 NA_4 0 -1.1219494574238587e-03
GD_1_5 b_1 NI_1 NA_5 0 1.6311756213701917e-04
GD_1_6 b_1 NI_1 NA_6 0 1.3323647169905203e-04
GD_1_7 b_1 NI_1 NA_7 0 7.4465326225461177e-07
GD_1_8 b_1 NI_1 NA_8 0 3.4878453060958149e-05
GD_1_9 b_1 NI_1 NA_9 0 8.9269178687395970e-06
GD_1_10 b_1 NI_1 NA_10 0 7.7381918748859573e-06
GD_1_11 b_1 NI_1 NA_11 0 1.1329729119207016e-05
GD_1_12 b_1 NI_1 NA_12 0 3.1921473820252031e-06
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 -5.0037719785017525e-02
GC_2_2 b_2 NI_2 NS_2 0 1.1076373767027689e-01
GC_2_3 b_2 NI_2 NS_3 0 1.1664279414513690e-08
GC_2_4 b_2 NI_2 NS_4 0 1.9861986912215787e-05
GC_2_5 b_2 NI_2 NS_5 0 -1.5739383571446577e-02
GC_2_6 b_2 NI_2 NS_6 0 2.4245657385051828e-02
GC_2_7 b_2 NI_2 NS_7 0 -7.8711093545999408e-03
GC_2_8 b_2 NI_2 NS_8 0 -1.4518741948540708e-02
GC_2_9 b_2 NI_2 NS_9 0 2.0325303696791499e-02
GC_2_10 b_2 NI_2 NS_10 0 6.6761488808325213e-03
GC_2_11 b_2 NI_2 NS_11 0 8.0659567308362500e-03
GC_2_12 b_2 NI_2 NS_12 0 4.4188588535655625e-02
GC_2_13 b_2 NI_2 NS_13 0 -1.1822644460416589e-02
GC_2_14 b_2 NI_2 NS_14 0 -3.1939196634110452e-03
GC_2_15 b_2 NI_2 NS_15 0 -5.1132613654034983e-03
GC_2_16 b_2 NI_2 NS_16 0 -4.0785578520759281e-03
GC_2_17 b_2 NI_2 NS_17 0 2.6802351255319507e-02
GC_2_18 b_2 NI_2 NS_18 0 1.2878838319268002e-04
GC_2_19 b_2 NI_2 NS_19 0 3.4101288351888165e-02
GC_2_20 b_2 NI_2 NS_20 0 3.1057522189457738e-02
GC_2_21 b_2 NI_2 NS_21 0 -1.5591715902611172e-02
GC_2_22 b_2 NI_2 NS_22 0 8.2163521308479762e-03
GC_2_23 b_2 NI_2 NS_23 0 -1.0700763171500364e-03
GC_2_24 b_2 NI_2 NS_24 0 -6.8531756839950242e-03
GC_2_25 b_2 NI_2 NS_25 0 -6.9888390242066653e-02
GC_2_26 b_2 NI_2 NS_26 0 1.6944830244588914e-03
GC_2_27 b_2 NI_2 NS_27 0 5.9934852708580469e-02
GC_2_28 b_2 NI_2 NS_28 0 -6.4654666394797000e-02
GC_2_29 b_2 NI_2 NS_29 0 -1.0233466126529798e-08
GC_2_30 b_2 NI_2 NS_30 0 -8.1983893351230147e-06
GC_2_31 b_2 NI_2 NS_31 0 -1.8758516813947932e-03
GC_2_32 b_2 NI_2 NS_32 0 -2.8706548412248995e-03
GC_2_33 b_2 NI_2 NS_33 0 -5.0998746470950927e-03
GC_2_34 b_2 NI_2 NS_34 0 1.9265479434409953e-03
GC_2_35 b_2 NI_2 NS_35 0 2.3837856116197516e-03
GC_2_36 b_2 NI_2 NS_36 0 -1.2477161950727610e-03
GC_2_37 b_2 NI_2 NS_37 0 -1.0661875966280447e-02
GC_2_38 b_2 NI_2 NS_38 0 1.1356529007343062e-03
GC_2_39 b_2 NI_2 NS_39 0 5.9634237015429321e-04
GC_2_40 b_2 NI_2 NS_40 0 1.7470517300509191e-03
GC_2_41 b_2 NI_2 NS_41 0 -9.6080888142928899e-04
GC_2_42 b_2 NI_2 NS_42 0 2.2969430138115280e-03
GC_2_43 b_2 NI_2 NS_43 0 5.3288097254274307e-04
GC_2_44 b_2 NI_2 NS_44 0 -5.8517879729081245e-03
GC_2_45 b_2 NI_2 NS_45 0 -8.5170547035245715e-03
GC_2_46 b_2 NI_2 NS_46 0 6.9045156927713819e-03
GC_2_47 b_2 NI_2 NS_47 0 2.5028306563983070e-03
GC_2_48 b_2 NI_2 NS_48 0 -3.6531650313559550e-03
GC_2_49 b_2 NI_2 NS_49 0 -2.5960265715554071e-03
GC_2_50 b_2 NI_2 NS_50 0 -5.3416983383629626e-04
GC_2_51 b_2 NI_2 NS_51 0 5.5354219558516236e-02
GC_2_52 b_2 NI_2 NS_52 0 1.8152608436065748e-03
GC_2_53 b_2 NI_2 NS_53 0 -1.3745704524008690e-03
GC_2_54 b_2 NI_2 NS_54 0 2.3328647324757524e-03
GC_2_55 b_2 NI_2 NS_55 0 7.5881762027234520e-10
GC_2_56 b_2 NI_2 NS_56 0 6.0065849899674574e-07
GC_2_57 b_2 NI_2 NS_57 0 -1.9596090223932992e-04
GC_2_58 b_2 NI_2 NS_58 0 -4.5533576207287493e-04
GC_2_59 b_2 NI_2 NS_59 0 -1.0665922628444703e-03
GC_2_60 b_2 NI_2 NS_60 0 -9.2132880615847245e-04
GC_2_61 b_2 NI_2 NS_61 0 -2.3173765228385978e-03
GC_2_62 b_2 NI_2 NS_62 0 3.1222083689818486e-04
GC_2_63 b_2 NI_2 NS_63 0 -3.4636422067155047e-04
GC_2_64 b_2 NI_2 NS_64 0 4.1981894755437257e-03
GC_2_65 b_2 NI_2 NS_65 0 9.7828934204943025e-04
GC_2_66 b_2 NI_2 NS_66 0 4.4367342765187139e-04
GC_2_67 b_2 NI_2 NS_67 0 -3.7329545536269503e-04
GC_2_68 b_2 NI_2 NS_68 0 7.9841425140933061e-05
GC_2_69 b_2 NI_2 NS_69 0 -3.1453904082015945e-04
GC_2_70 b_2 NI_2 NS_70 0 3.3540638103354359e-03
GC_2_71 b_2 NI_2 NS_71 0 5.2329406719678791e-03
GC_2_72 b_2 NI_2 NS_72 0 8.1285628475197616e-04
GC_2_73 b_2 NI_2 NS_73 0 1.3427545697935628e-03
GC_2_74 b_2 NI_2 NS_74 0 -1.9440140014151972e-03
GC_2_75 b_2 NI_2 NS_75 0 -8.8256221340532947e-04
GC_2_76 b_2 NI_2 NS_76 0 -6.3689647560772776e-04
GC_2_77 b_2 NI_2 NS_77 0 -1.4735563970516973e-03
GC_2_78 b_2 NI_2 NS_78 0 2.5664387109443892e-03
GC_2_79 b_2 NI_2 NS_79 0 -7.4975960757069681e-03
GC_2_80 b_2 NI_2 NS_80 0 5.4454235824727467e-03
GC_2_81 b_2 NI_2 NS_81 0 -8.2825467001905300e-10
GC_2_82 b_2 NI_2 NS_82 0 -1.6858108898331376e-06
GC_2_83 b_2 NI_2 NS_83 0 2.5528766609402405e-04
GC_2_84 b_2 NI_2 NS_84 0 2.6644769440055628e-03
GC_2_85 b_2 NI_2 NS_85 0 4.5291339501023018e-03
GC_2_86 b_2 NI_2 NS_86 0 -2.7565355677247054e-03
GC_2_87 b_2 NI_2 NS_87 0 -5.4227391907847484e-03
GC_2_88 b_2 NI_2 NS_88 0 4.2034577459685657e-04
GC_2_89 b_2 NI_2 NS_89 0 8.8583377785286174e-03
GC_2_90 b_2 NI_2 NS_90 0 -6.2088156242913570e-04
GC_2_91 b_2 NI_2 NS_91 0 -2.8261182324715926e-03
GC_2_92 b_2 NI_2 NS_92 0 -2.3963319295237846e-03
GC_2_93 b_2 NI_2 NS_93 0 4.3090589640461195e-05
GC_2_94 b_2 NI_2 NS_94 0 -2.1138834115335386e-03
GC_2_95 b_2 NI_2 NS_95 0 -3.5070931951752464e-03
GC_2_96 b_2 NI_2 NS_96 0 5.5495700728484393e-03
GC_2_97 b_2 NI_2 NS_97 0 5.0983693665808440e-03
GC_2_98 b_2 NI_2 NS_98 0 -7.7603757444736216e-03
GC_2_99 b_2 NI_2 NS_99 0 -5.0389557949857937e-03
GC_2_100 b_2 NI_2 NS_100 0 3.0962213485802763e-03
GC_2_101 b_2 NI_2 NS_101 0 2.2446186018856055e-03
GC_2_102 b_2 NI_2 NS_102 0 -1.6873571154541311e-03
GC_2_103 b_2 NI_2 NS_103 0 -5.9461873679980811e-03
GC_2_104 b_2 NI_2 NS_104 0 3.8165500824202197e-03
GC_2_105 b_2 NI_2 NS_105 0 1.5157434347576722e-04
GC_2_106 b_2 NI_2 NS_106 0 1.2809809140874620e-05
GC_2_107 b_2 NI_2 NS_107 0 -4.2742665395222229e-10
GC_2_108 b_2 NI_2 NS_108 0 4.5130301345949274e-08
GC_2_109 b_2 NI_2 NS_109 0 5.1596760519683039e-06
GC_2_110 b_2 NI_2 NS_110 0 7.5616107933734950e-05
GC_2_111 b_2 NI_2 NS_111 0 1.5335221836465564e-04
GC_2_112 b_2 NI_2 NS_112 0 1.3548710722301771e-04
GC_2_113 b_2 NI_2 NS_113 0 3.4656072079332009e-04
GC_2_114 b_2 NI_2 NS_114 0 -2.4741108271503300e-05
GC_2_115 b_2 NI_2 NS_115 0 5.1570183480894069e-05
GC_2_116 b_2 NI_2 NS_116 0 -5.8538715229608073e-04
GC_2_117 b_2 NI_2 NS_117 0 -1.4593519005951896e-04
GC_2_118 b_2 NI_2 NS_118 0 -6.8386950795887259e-05
GC_2_119 b_2 NI_2 NS_119 0 5.1713283732782018e-05
GC_2_120 b_2 NI_2 NS_120 0 -1.0507847617413628e-05
GC_2_121 b_2 NI_2 NS_121 0 4.7730213534758301e-05
GC_2_122 b_2 NI_2 NS_122 0 -4.5313042738881243e-04
GC_2_123 b_2 NI_2 NS_123 0 -7.0918794683506663e-04
GC_2_124 b_2 NI_2 NS_124 0 -8.3323698965071316e-05
GC_2_125 b_2 NI_2 NS_125 0 -1.7472346321385223e-04
GC_2_126 b_2 NI_2 NS_126 0 2.5870651860759923e-04
GC_2_127 b_2 NI_2 NS_127 0 1.0249954155007232e-04
GC_2_128 b_2 NI_2 NS_128 0 7.9812165568327902e-05
GC_2_129 b_2 NI_2 NS_129 0 -8.6761639444484198e-05
GC_2_130 b_2 NI_2 NS_130 0 -3.2996766262977670e-04
GC_2_131 b_2 NI_2 NS_131 0 3.9467687024090993e-04
GC_2_132 b_2 NI_2 NS_132 0 -2.0170416171404314e-03
GC_2_133 b_2 NI_2 NS_133 0 4.0764937719696678e-10
GC_2_134 b_2 NI_2 NS_134 0 -2.7091784441029882e-08
GC_2_135 b_2 NI_2 NS_135 0 1.8629832432831359e-05
GC_2_136 b_2 NI_2 NS_136 0 4.3391935934210435e-05
GC_2_137 b_2 NI_2 NS_137 0 8.1680057418210801e-05
GC_2_138 b_2 NI_2 NS_138 0 -3.0853931517876409e-05
GC_2_139 b_2 NI_2 NS_139 0 -1.3841629984959610e-05
GC_2_140 b_2 NI_2 NS_140 0 1.3779023028558621e-05
GC_2_141 b_2 NI_2 NS_141 0 1.9715185655923729e-04
GC_2_142 b_2 NI_2 NS_142 0 -9.9073456458437242e-05
GC_2_143 b_2 NI_2 NS_143 0 2.6774533893439978e-05
GC_2_144 b_2 NI_2 NS_144 0 -9.8009285484007937e-05
GC_2_145 b_2 NI_2 NS_145 0 -1.7495832621820412e-05
GC_2_146 b_2 NI_2 NS_146 0 -9.8105913661881053e-05
GC_2_147 b_2 NI_2 NS_147 0 9.9651051486111996e-06
GC_2_148 b_2 NI_2 NS_148 0 -9.7431746414185406e-05
GC_2_149 b_2 NI_2 NS_149 0 -9.8104245263925090e-05
GC_2_150 b_2 NI_2 NS_150 0 -3.1498379012690728e-04
GC_2_151 b_2 NI_2 NS_151 0 -1.3390325911973193e-04
GC_2_152 b_2 NI_2 NS_152 0 -1.1512948993797322e-04
GC_2_153 b_2 NI_2 NS_153 0 -1.9651413970535242e-05
GC_2_154 b_2 NI_2 NS_154 0 -1.9128949089750687e-04
GC_2_155 b_2 NI_2 NS_155 0 1.5206724221078630e-03
GC_2_156 b_2 NI_2 NS_156 0 -1.0185406213226167e-04
GC_2_157 b_2 NI_2 NS_157 0 -1.6167547132852096e-05
GC_2_158 b_2 NI_2 NS_158 0 -2.5713233982085400e-04
GC_2_159 b_2 NI_2 NS_159 0 -1.0826303175651568e-10
GC_2_160 b_2 NI_2 NS_160 0 4.7617827623041298e-09
GC_2_161 b_2 NI_2 NS_161 0 5.0889302852738434e-06
GC_2_162 b_2 NI_2 NS_162 0 9.7287696128188634e-06
GC_2_163 b_2 NI_2 NS_163 0 1.6466340399716960e-05
GC_2_164 b_2 NI_2 NS_164 0 1.3314056324544624e-05
GC_2_165 b_2 NI_2 NS_165 0 3.8436504831292203e-05
GC_2_166 b_2 NI_2 NS_166 0 -3.5538485728881405e-06
GC_2_167 b_2 NI_2 NS_167 0 1.4511380238905351e-05
GC_2_168 b_2 NI_2 NS_168 0 -6.2679408119752512e-05
GC_2_169 b_2 NI_2 NS_169 0 -1.1740220998157623e-05
GC_2_170 b_2 NI_2 NS_170 0 -9.0260278259952477e-06
GC_2_171 b_2 NI_2 NS_171 0 4.7333675123297289e-06
GC_2_172 b_2 NI_2 NS_172 0 -3.5102473048275405e-06
GC_2_173 b_2 NI_2 NS_173 0 9.6833327104846142e-06
GC_2_174 b_2 NI_2 NS_174 0 -5.0075247858060733e-05
GC_2_175 b_2 NI_2 NS_175 0 -6.6267409835535430e-05
GC_2_176 b_2 NI_2 NS_176 0 -2.1578366259689846e-05
GC_2_177 b_2 NI_2 NS_177 0 -1.6765733706235697e-05
GC_2_178 b_2 NI_2 NS_178 0 1.9317411422106590e-05
GC_2_179 b_2 NI_2 NS_179 0 1.6177485099280286e-05
GC_2_180 b_2 NI_2 NS_180 0 -1.3689171911959159e-06
GC_2_181 b_2 NI_2 NS_181 0 2.1856806026043459e-04
GC_2_182 b_2 NI_2 NS_182 0 7.6285008889322095e-06
GC_2_183 b_2 NI_2 NS_183 0 -1.4358277145971161e-04
GC_2_184 b_2 NI_2 NS_184 0 6.6681873057581730e-04
GC_2_185 b_2 NI_2 NS_185 0 1.2440178298572975e-10
GC_2_186 b_2 NI_2 NS_186 0 -1.1384667150893300e-08
GC_2_187 b_2 NI_2 NS_187 0 -4.0163430111585081e-06
GC_2_188 b_2 NI_2 NS_188 0 -3.9922643718637563e-06
GC_2_189 b_2 NI_2 NS_189 0 -9.5849406607737799e-06
GC_2_190 b_2 NI_2 NS_190 0 -3.6873690657765890e-06
GC_2_191 b_2 NI_2 NS_191 0 -1.8730175774520897e-05
GC_2_192 b_2 NI_2 NS_192 0 -1.5350584096156917e-06
GC_2_193 b_2 NI_2 NS_193 0 -2.9271138593072035e-05
GC_2_194 b_2 NI_2 NS_194 0 2.7762606583549018e-05
GC_2_195 b_2 NI_2 NS_195 0 -2.1466916807253203e-05
GC_2_196 b_2 NI_2 NS_196 0 2.3556306300507449e-05
GC_2_197 b_2 NI_2 NS_197 0 6.1046516509156917e-06
GC_2_198 b_2 NI_2 NS_198 0 2.3438810187248848e-05
GC_2_199 b_2 NI_2 NS_199 0 -1.5894478384880734e-05
GC_2_200 b_2 NI_2 NS_200 0 5.5645649557857500e-05
GC_2_201 b_2 NI_2 NS_201 0 5.4416753520409225e-05
GC_2_202 b_2 NI_2 NS_202 0 6.5745047910484297e-05
GC_2_203 b_2 NI_2 NS_203 0 2.2593814483453855e-05
GC_2_204 b_2 NI_2 NS_204 0 4.5702050087632227e-05
GC_2_205 b_2 NI_2 NS_205 0 1.4942180519755108e-05
GC_2_206 b_2 NI_2 NS_206 0 4.9676808354161423e-05
GC_2_207 b_2 NI_2 NS_207 0 -5.1915999362174147e-04
GC_2_208 b_2 NI_2 NS_208 0 2.3889064886626584e-05
GC_2_209 b_2 NI_2 NS_209 0 -2.4826036530227325e-05
GC_2_210 b_2 NI_2 NS_210 0 2.0783958272288957e-05
GC_2_211 b_2 NI_2 NS_211 0 -3.5006714723012686e-11
GC_2_212 b_2 NI_2 NS_212 0 -2.7090154647537828e-10
GC_2_213 b_2 NI_2 NS_213 0 1.6166640642600099e-06
GC_2_214 b_2 NI_2 NS_214 0 1.4393720392657486e-06
GC_2_215 b_2 NI_2 NS_215 0 2.5870846373965305e-07
GC_2_216 b_2 NI_2 NS_216 0 3.7190209921283601e-07
GC_2_217 b_2 NI_2 NS_217 0 1.7411259886259908e-06
GC_2_218 b_2 NI_2 NS_218 0 -2.0416400346592152e-07
GC_2_219 b_2 NI_2 NS_219 0 3.3661778535361783e-06
GC_2_220 b_2 NI_2 NS_220 0 -1.0270839900491294e-06
GC_2_221 b_2 NI_2 NS_221 0 4.2256026173139933e-07
GC_2_222 b_2 NI_2 NS_222 0 5.0171752915686385e-08
GC_2_223 b_2 NI_2 NS_223 0 2.5403826137322951e-07
GC_2_224 b_2 NI_2 NS_224 0 -2.9663364255119621e-07
GC_2_225 b_2 NI_2 NS_225 0 1.0840315432377508e-06
GC_2_226 b_2 NI_2 NS_226 0 -1.0041276345792633e-06
GC_2_227 b_2 NI_2 NS_227 0 1.6348101037127432e-06
GC_2_228 b_2 NI_2 NS_228 0 -1.2123855417853766e-06
GC_2_229 b_2 NI_2 NS_229 0 -5.8100920047221378e-08
GC_2_230 b_2 NI_2 NS_230 0 1.3019077527779525e-06
GC_2_231 b_2 NI_2 NS_231 0 3.3328558696613723e-07
GC_2_232 b_2 NI_2 NS_232 0 6.8675702847956561e-07
GC_2_233 b_2 NI_2 NS_233 0 -1.6981000880880379e-05
GC_2_234 b_2 NI_2 NS_234 0 -1.3435249282238657e-06
GC_2_235 b_2 NI_2 NS_235 0 -2.7825253256125678e-05
GC_2_236 b_2 NI_2 NS_236 0 4.2360480575986728e-05
GC_2_237 b_2 NI_2 NS_237 0 3.6705451978140027e-11
GC_2_238 b_2 NI_2 NS_238 0 -2.7773099246907627e-10
GC_2_239 b_2 NI_2 NS_239 0 8.4146527341151606e-07
GC_2_240 b_2 NI_2 NS_240 0 4.8946649089859325e-07
GC_2_241 b_2 NI_2 NS_241 0 4.0299542496338618e-07
GC_2_242 b_2 NI_2 NS_242 0 -7.5688550414603573e-07
GC_2_243 b_2 NI_2 NS_243 0 -4.8229317105046710e-07
GC_2_244 b_2 NI_2 NS_244 0 9.9668466938817942e-07
GC_2_245 b_2 NI_2 NS_245 0 1.4113530954863999e-06
GC_2_246 b_2 NI_2 NS_246 0 1.8134196361242915e-07
GC_2_247 b_2 NI_2 NS_247 0 -4.2582299037621908e-07
GC_2_248 b_2 NI_2 NS_248 0 9.6992937609970347e-07
GC_2_249 b_2 NI_2 NS_249 0 5.7117605753666229e-07
GC_2_250 b_2 NI_2 NS_250 0 3.8256426497921828e-07
GC_2_251 b_2 NI_2 NS_251 0 5.5721833197772435e-07
GC_2_252 b_2 NI_2 NS_252 0 3.2490416948925266e-06
GC_2_253 b_2 NI_2 NS_253 0 4.0010697371851770e-06
GC_2_254 b_2 NI_2 NS_254 0 7.7940025126073926e-07
GC_2_255 b_2 NI_2 NS_255 0 9.0180422205167500e-07
GC_2_256 b_2 NI_2 NS_256 0 2.3877079535690930e-06
GC_2_257 b_2 NI_2 NS_257 0 1.1488164942644996e-06
GC_2_258 b_2 NI_2 NS_258 0 2.6084903318736927e-06
GC_2_259 b_2 NI_2 NS_259 0 -3.3517704257428665e-05
GC_2_260 b_2 NI_2 NS_260 0 4.1416093417901734e-07
GC_2_261 b_2 NI_2 NS_261 0 -1.1797567943379813e-05
GC_2_262 b_2 NI_2 NS_262 0 -5.5691895589798676e-06
GC_2_263 b_2 NI_2 NS_263 0 -3.0498510320614440e-11
GC_2_264 b_2 NI_2 NS_264 0 -1.3564564778890608e-10
GC_2_265 b_2 NI_2 NS_265 0 2.2975254911130893e-06
GC_2_266 b_2 NI_2 NS_266 0 1.7812181868914601e-06
GC_2_267 b_2 NI_2 NS_267 0 -6.4111924354588978e-07
GC_2_268 b_2 NI_2 NS_268 0 -3.8629251411172964e-07
GC_2_269 b_2 NI_2 NS_269 0 1.5521516970849967e-06
GC_2_270 b_2 NI_2 NS_270 0 -1.1535837552488027e-06
GC_2_271 b_2 NI_2 NS_271 0 1.8422851262926460e-06
GC_2_272 b_2 NI_2 NS_272 0 -4.3467522868176573e-07
GC_2_273 b_2 NI_2 NS_273 0 1.1803393629659542e-07
GC_2_274 b_2 NI_2 NS_274 0 -1.8751676636145164e-07
GC_2_275 b_2 NI_2 NS_275 0 5.5244895483002028e-08
GC_2_276 b_2 NI_2 NS_276 0 -3.1825279856073647e-07
GC_2_277 b_2 NI_2 NS_277 0 4.3506150156330690e-07
GC_2_278 b_2 NI_2 NS_278 0 -7.3873650210580540e-07
GC_2_279 b_2 NI_2 NS_279 0 9.1283310865207233e-07
GC_2_280 b_2 NI_2 NS_280 0 -1.3978333964887706e-06
GC_2_281 b_2 NI_2 NS_281 0 -1.9067303241284792e-07
GC_2_282 b_2 NI_2 NS_282 0 5.9848021174789904e-07
GC_2_283 b_2 NI_2 NS_283 0 3.5017972574750206e-07
GC_2_284 b_2 NI_2 NS_284 0 -1.5154848590622499e-08
GC_2_285 b_2 NI_2 NS_285 0 5.8038864001412693e-06
GC_2_286 b_2 NI_2 NS_286 0 2.3966717895917926e-06
GC_2_287 b_2 NI_2 NS_287 0 -3.5487271757902390e-05
GC_2_288 b_2 NI_2 NS_288 0 4.3755698258612115e-05
GC_2_289 b_2 NI_2 NS_289 0 3.2703459322660947e-11
GC_2_290 b_2 NI_2 NS_290 0 -2.6824624542121541e-10
GC_2_291 b_2 NI_2 NS_291 0 1.0320798095662097e-06
GC_2_292 b_2 NI_2 NS_292 0 1.0605759667140500e-06
GC_2_293 b_2 NI_2 NS_293 0 1.7241328049422578e-06
GC_2_294 b_2 NI_2 NS_294 0 2.5964992032279362e-07
GC_2_295 b_2 NI_2 NS_295 0 1.0932120357998249e-06
GC_2_296 b_2 NI_2 NS_296 0 4.6059960874523228e-07
GC_2_297 b_2 NI_2 NS_297 0 2.9262620478441394e-06
GC_2_298 b_2 NI_2 NS_298 0 -4.3423347401779245e-07
GC_2_299 b_2 NI_2 NS_299 0 1.0132358749980138e-06
GC_2_300 b_2 NI_2 NS_300 0 5.3044812427702266e-09
GC_2_301 b_2 NI_2 NS_301 0 5.6285413814314435e-07
GC_2_302 b_2 NI_2 NS_302 0 -5.1625010337346877e-07
GC_2_303 b_2 NI_2 NS_303 0 1.6607435584903902e-06
GC_2_304 b_2 NI_2 NS_304 0 1.2910028386579395e-06
GC_2_305 b_2 NI_2 NS_305 0 2.8544592058570022e-06
GC_2_306 b_2 NI_2 NS_306 0 -1.2126697453387570e-06
GC_2_307 b_2 NI_2 NS_307 0 5.5986031676021257e-07
GC_2_308 b_2 NI_2 NS_308 0 1.1266008184679522e-06
GC_2_309 b_2 NI_2 NS_309 0 3.9045694302116883e-07
GC_2_310 b_2 NI_2 NS_310 0 1.5530721092318115e-06
GC_2_311 b_2 NI_2 NS_311 0 -3.6623120603906959e-05
GC_2_312 b_2 NI_2 NS_312 0 -3.7034616093951101e-06
GD_2_1 b_2 NI_2 NA_1 0 -2.0539192952172793e-02
GD_2_2 b_2 NI_2 NA_2 0 -2.9881630529505005e-02
GD_2_3 b_2 NI_2 NA_3 0 -1.1219611503046820e-03
GD_2_4 b_2 NI_2 NA_4 0 1.3427146547155416e-02
GD_2_5 b_2 NI_2 NA_5 0 1.3324649061085297e-04
GD_2_6 b_2 NI_2 NA_6 0 1.6315392054082708e-04
GD_2_7 b_2 NI_2 NA_7 0 3.4782104079854388e-05
GD_2_8 b_2 NI_2 NA_8 0 7.5813343018130616e-07
GD_2_9 b_2 NI_2 NA_9 0 7.7385921800857036e-06
GD_2_10 b_2 NI_2 NA_10 0 8.8774481950294364e-06
GD_2_11 b_2 NI_2 NA_11 0 3.1881942197431915e-06
GD_2_12 b_2 NI_2 NA_12 0 1.1329725045561610e-05
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 -7.4975960757069663e-03
GC_3_2 b_3 NI_3 NS_2 0 5.4454235824725073e-03
GC_3_3 b_3 NI_3 NS_3 0 -8.2825467001853611e-10
GC_3_4 b_3 NI_3 NS_4 0 -1.6858108898331999e-06
GC_3_5 b_3 NI_3 NS_5 0 2.5528766609402432e-04
GC_3_6 b_3 NI_3 NS_6 0 2.6644769440055662e-03
GC_3_7 b_3 NI_3 NS_7 0 4.5291339501023053e-03
GC_3_8 b_3 NI_3 NS_8 0 -2.7565355677247019e-03
GC_3_9 b_3 NI_3 NS_9 0 -5.4227391907847415e-03
GC_3_10 b_3 NI_3 NS_10 0 4.2034577459686053e-04
GC_3_11 b_3 NI_3 NS_11 0 8.8583377785286348e-03
GC_3_12 b_3 NI_3 NS_12 0 -6.2088156242914340e-04
GC_3_13 b_3 NI_3 NS_13 0 -2.8261182324715874e-03
GC_3_14 b_3 NI_3 NS_14 0 -2.3963319295237915e-03
GC_3_15 b_3 NI_3 NS_15 0 4.3090589640459914e-05
GC_3_16 b_3 NI_3 NS_16 0 -2.1138834115335446e-03
GC_3_17 b_3 NI_3 NS_17 0 -3.5070931951752412e-03
GC_3_18 b_3 NI_3 NS_18 0 5.5495700728484280e-03
GC_3_19 b_3 NI_3 NS_19 0 5.0983693665808362e-03
GC_3_20 b_3 NI_3 NS_20 0 -7.7603757444736380e-03
GC_3_21 b_3 NI_3 NS_21 0 -5.0389557949857937e-03
GC_3_22 b_3 NI_3 NS_22 0 3.0962213485802659e-03
GC_3_23 b_3 NI_3 NS_23 0 2.2446186018856081e-03
GC_3_24 b_3 NI_3 NS_24 0 -1.6873571154541421e-03
GC_3_25 b_3 NI_3 NS_25 0 -5.9461873679978799e-03
GC_3_26 b_3 NI_3 NS_26 0 3.8165500824202353e-03
GC_3_27 b_3 NI_3 NS_27 0 -1.3745899579498170e-03
GC_3_28 b_3 NI_3 NS_28 0 2.3328611430557451e-03
GC_3_29 b_3 NI_3 NS_29 0 7.5881727110688637e-10
GC_3_30 b_3 NI_3 NS_30 0 6.0065849286201200e-07
GC_3_31 b_3 NI_3 NS_31 0 -1.9596182595988700e-04
GC_3_32 b_3 NI_3 NS_32 0 -4.5534379655682807e-04
GC_3_33 b_3 NI_3 NS_33 0 -1.0665912541896300e-03
GC_3_34 b_3 NI_3 NS_34 0 -9.2132098607863736e-04
GC_3_35 b_3 NI_3 NS_35 0 -2.3173781110569524e-03
GC_3_36 b_3 NI_3 NS_36 0 3.1222785732386722e-04
GC_3_37 b_3 NI_3 NS_37 0 -3.4635653571128987e-04
GC_3_38 b_3 NI_3 NS_38 0 4.1981806373795191e-03
GC_3_39 b_3 NI_3 NS_39 0 9.7829065525191429e-04
GC_3_40 b_3 NI_3 NS_40 0 4.4367094401280929e-04
GC_3_41 b_3 NI_3 NS_41 0 -3.7329437078607571e-04
GC_3_42 b_3 NI_3 NS_42 0 7.9842631324595980e-05
GC_3_43 b_3 NI_3 NS_43 0 -3.1453545434071328e-04
GC_3_44 b_3 NI_3 NS_44 0 3.3540627909886562e-03
GC_3_45 b_3 NI_3 NS_45 0 5.2329373469934964e-03
GC_3_46 b_3 NI_3 NS_46 0 8.1284762392161468e-04
GC_3_47 b_3 NI_3 NS_47 0 1.3427520053122723e-03
GC_3_48 b_3 NI_3 NS_48 0 -1.9440147231157816e-03
GC_3_49 b_3 NI_3 NS_49 0 -8.8256310646948216e-04
GC_3_50 b_3 NI_3 NS_50 0 -6.3689546485460095e-04
GC_3_51 b_3 NI_3 NS_51 0 -1.4735533000609360e-03
GC_3_52 b_3 NI_3 NS_52 0 2.5664393832339765e-03
GC_3_53 b_3 NI_3 NS_53 0 5.9438136073012834e-02
GC_3_54 b_3 NI_3 NS_54 0 -6.3779997448680070e-02
GC_3_55 b_3 NI_3 NS_55 0 -1.0218715257316923e-08
GC_3_56 b_3 NI_3 NS_56 0 -8.2100868785480612e-06
GC_3_57 b_3 NI_3 NS_57 0 -1.8519166209792891e-03
GC_3_58 b_3 NI_3 NS_58 0 -2.8731340475971201e-03
GC_3_59 b_3 NI_3 NS_59 0 -5.1084756720848586e-03
GC_3_60 b_3 NI_3 NS_60 0 1.9400114889521790e-03
GC_3_61 b_3 NI_3 NS_61 0 2.4463666578743949e-03
GC_3_62 b_3 NI_3 NS_62 0 -1.2255434516112856e-03
GC_3_63 b_3 NI_3 NS_63 0 -1.0650799674863385e-02
GC_3_64 b_3 NI_3 NS_64 0 1.1045689712411105e-03
GC_3_65 b_3 NI_3 NS_65 0 6.4145744822000398e-04
GC_3_66 b_3 NI_3 NS_66 0 1.7543170152112596e-03
GC_3_67 b_3 NI_3 NS_67 0 -9.5624673213744670e-04
GC_3_68 b_3 NI_3 NS_68 0 2.2871421137470350e-03
GC_3_69 b_3 NI_3 NS_69 0 5.9413739439217756e-04
GC_3_70 b_3 NI_3 NS_70 0 -5.8937142081883862e-03
GC_3_71 b_3 NI_3 NS_71 0 -8.5380811876149439e-03
GC_3_72 b_3 NI_3 NS_72 0 6.8906920148834004e-03
GC_3_73 b_3 NI_3 NS_73 0 2.5187097649788420e-03
GC_3_74 b_3 NI_3 NS_74 0 -3.6778740922647824e-03
GC_3_75 b_3 NI_3 NS_75 0 -2.6381595052563205e-03
GC_3_76 b_3 NI_3 NS_76 0 -5.1433834238557251e-04
GC_3_77 b_3 NI_3 NS_77 0 5.4574972974246912e-02
GC_3_78 b_3 NI_3 NS_78 0 1.6205496302429696e-03
GC_3_79 b_3 NI_3 NS_79 0 -4.9957360006206875e-02
GC_3_80 b_3 NI_3 NS_80 0 1.0966284596734312e-01
GC_3_81 b_3 NI_3 NS_81 0 1.0579523109661094e-08
GC_3_82 b_3 NI_3 NS_82 0 1.9882063556629574e-05
GC_3_83 b_3 NI_3 NS_83 0 -1.5752602248633181e-02
GC_3_84 b_3 NI_3 NS_84 0 2.4251913232738787e-02
GC_3_85 b_3 NI_3 NS_85 0 -7.8021559516944297e-03
GC_3_86 b_3 NI_3 NS_86 0 -1.4485544701047265e-02
GC_3_87 b_3 NI_3 NS_87 0 2.0432729895326650e-02
GC_3_88 b_3 NI_3 NS_88 0 6.6858686342307263e-03
GC_3_89 b_3 NI_3 NS_89 0 8.0641705904882632e-03
GC_3_90 b_3 NI_3 NS_90 0 4.3992224131868873e-02
GC_3_91 b_3 NI_3 NS_91 0 -1.1854721044815861e-02
GC_3_92 b_3 NI_3 NS_92 0 -3.2297495410856954e-03
GC_3_93 b_3 NI_3 NS_93 0 -5.0941031615457776e-03
GC_3_94 b_3 NI_3 NS_94 0 -4.0920228885113069e-03
GC_3_95 b_3 NI_3 NS_95 0 2.6818340328436881e-02
GC_3_96 b_3 NI_3 NS_96 0 -1.0398369793334156e-05
GC_3_97 b_3 NI_3 NS_97 0 3.3876596522363425e-02
GC_3_98 b_3 NI_3 NS_98 0 3.0995863071548609e-02
GC_3_99 b_3 NI_3 NS_99 0 -1.5641050925009715e-02
GC_3_100 b_3 NI_3 NS_100 0 8.2858690252631435e-03
GC_3_101 b_3 NI_3 NS_101 0 -9.9915412322053505e-04
GC_3_102 b_3 NI_3 NS_102 0 -6.8608375351511845e-03
GC_3_103 b_3 NI_3 NS_103 0 -6.8944255118152636e-02
GC_3_104 b_3 NI_3 NS_104 0 1.7522185483934338e-03
GC_3_105 b_3 NI_3 NS_105 0 -1.2120664543369261e-03
GC_3_106 b_3 NI_3 NS_106 0 5.5288377915632095e-04
GC_3_107 b_3 NI_3 NS_107 0 3.0006679197599986e-10
GC_3_108 b_3 NI_3 NS_108 0 -5.7499735144104574e-07
GC_3_109 b_3 NI_3 NS_109 0 3.1147146205305917e-05
GC_3_110 b_3 NI_3 NS_110 0 6.3814449757213887e-04
GC_3_111 b_3 NI_3 NS_111 0 1.0887928372579334e-03
GC_3_112 b_3 NI_3 NS_112 0 -6.7568193551917897e-04
GC_3_113 b_3 NI_3 NS_113 0 -1.3741747924445843e-03
GC_3_114 b_3 NI_3 NS_114 0 7.5250725283126417e-05
GC_3_115 b_3 NI_3 NS_115 0 2.0942417593644582e-03
GC_3_116 b_3 NI_3 NS_116 0 -1.0656274011916027e-04
GC_3_117 b_3 NI_3 NS_117 0 -7.3383166357768531e-04
GC_3_118 b_3 NI_3 NS_118 0 -5.7289836294185904e-04
GC_3_119 b_3 NI_3 NS_119 0 5.7537690596903170e-06
GC_3_120 b_3 NI_3 NS_120 0 -4.8778998285053233e-04
GC_3_121 b_3 NI_3 NS_121 0 -9.0586722931610590e-04
GC_3_122 b_3 NI_3 NS_122 0 1.3910544906116581e-03
GC_3_123 b_3 NI_3 NS_123 0 1.2473495878830630e-03
GC_3_124 b_3 NI_3 NS_124 0 -1.8369134054800676e-03
GC_3_125 b_3 NI_3 NS_125 0 -1.2248408675950414e-03
GC_3_126 b_3 NI_3 NS_126 0 7.8178232634839835e-04
GC_3_127 b_3 NI_3 NS_127 0 5.7543582526925670e-04
GC_3_128 b_3 NI_3 NS_128 0 -4.1190529220703137e-04
GC_3_129 b_3 NI_3 NS_129 0 -7.3187183354730576e-04
GC_3_130 b_3 NI_3 NS_130 0 1.1403197329256207e-03
GC_3_131 b_3 NI_3 NS_131 0 -1.0992736620396356e-03
GC_3_132 b_3 NI_3 NS_132 0 1.9265919587895146e-03
GC_3_133 b_3 NI_3 NS_133 0 -9.9958187998483142e-11
GC_3_134 b_3 NI_3 NS_134 0 2.7260434669181933e-07
GC_3_135 b_3 NI_3 NS_135 0 5.8942674513287522e-05
GC_3_136 b_3 NI_3 NS_136 0 -8.7011292050877457e-05
GC_3_137 b_3 NI_3 NS_137 0 -2.6161328128995200e-04
GC_3_138 b_3 NI_3 NS_138 0 -1.7084760210281738e-04
GC_3_139 b_3 NI_3 NS_139 0 -5.2945252146459007e-04
GC_3_140 b_3 NI_3 NS_140 0 2.5205537383415256e-05
GC_3_141 b_3 NI_3 NS_141 0 4.2398994524010111e-05
GC_3_142 b_3 NI_3 NS_142 0 9.1577025606995311e-04
GC_3_143 b_3 NI_3 NS_143 0 2.4558174069285561e-04
GC_3_144 b_3 NI_3 NS_144 0 1.3074070458594299e-04
GC_3_145 b_3 NI_3 NS_145 0 -8.1504628124073653e-05
GC_3_146 b_3 NI_3 NS_146 0 2.6832874985938945e-05
GC_3_147 b_3 NI_3 NS_147 0 -7.0975044219698152e-05
GC_3_148 b_3 NI_3 NS_148 0 7.5355454199736336e-04
GC_3_149 b_3 NI_3 NS_149 0 1.2758459275053922e-03
GC_3_150 b_3 NI_3 NS_150 0 1.3806943393687501e-04
GC_3_151 b_3 NI_3 NS_151 0 3.2408622581356453e-04
GC_3_152 b_3 NI_3 NS_152 0 -4.2267378912753706e-04
GC_3_153 b_3 NI_3 NS_153 0 -2.4532879494754497e-04
GC_3_154 b_3 NI_3 NS_154 0 -1.0928772642395172e-04
GC_3_155 b_3 NI_3 NS_155 0 -1.5486299127683563e-03
GC_3_156 b_3 NI_3 NS_156 0 3.7254268501119085e-04
GC_3_157 b_3 NI_3 NS_157 0 3.8432217158260141e-04
GC_3_158 b_3 NI_3 NS_158 0 -2.0226219625256395e-03
GC_3_159 b_3 NI_3 NS_159 0 4.0280159777549734e-10
GC_3_160 b_3 NI_3 NS_160 0 -2.6940667068342456e-08
GC_3_161 b_3 NI_3 NS_161 0 1.8994438095025021e-05
GC_3_162 b_3 NI_3 NS_162 0 4.3663121534215328e-05
GC_3_163 b_3 NI_3 NS_163 0 8.2131171197734066e-05
GC_3_164 b_3 NI_3 NS_164 0 -3.0748892879030394e-05
GC_3_165 b_3 NI_3 NS_165 0 -1.3347310332522469e-05
GC_3_166 b_3 NI_3 NS_166 0 1.3987429634709880e-05
GC_3_167 b_3 NI_3 NS_167 0 1.9809683102856271e-04
GC_3_168 b_3 NI_3 NS_168 0 -9.9308113608500732e-05
GC_3_169 b_3 NI_3 NS_169 0 2.7246169269620235e-05
GC_3_170 b_3 NI_3 NS_170 0 -9.8014285668900401e-05
GC_3_171 b_3 NI_3 NS_171 0 -1.7287805152787286e-05
GC_3_172 b_3 NI_3 NS_172 0 -9.8335138648588066e-05
GC_3_173 b_3 NI_3 NS_173 0 1.0774117162266475e-05
GC_3_174 b_3 NI_3 NS_174 0 -9.7259054831402180e-05
GC_3_175 b_3 NI_3 NS_175 0 -9.7202756848590658e-05
GC_3_176 b_3 NI_3 NS_176 0 -3.1583836762545079e-04
GC_3_177 b_3 NI_3 NS_177 0 -1.3360484230555170e-04
GC_3_178 b_3 NI_3 NS_178 0 -1.1524848470247532e-04
GC_3_179 b_3 NI_3 NS_179 0 -1.9119749669929041e-05
GC_3_180 b_3 NI_3 NS_180 0 -1.9116379133716339e-04
GC_3_181 b_3 NI_3 NS_181 0 1.5264288676381046e-03
GC_3_182 b_3 NI_3 NS_182 0 -9.9582007608605257e-05
GC_3_183 b_3 NI_3 NS_183 0 1.2876808106926881e-04
GC_3_184 b_3 NI_3 NS_184 0 5.3480686938754187e-05
GC_3_185 b_3 NI_3 NS_185 0 -4.2223188231934821e-10
GC_3_186 b_3 NI_3 NS_186 0 4.4745808014121542e-08
GC_3_187 b_3 NI_3 NS_187 0 5.7032040322425014e-06
GC_3_188 b_3 NI_3 NS_188 0 7.6084092999094942e-05
GC_3_189 b_3 NI_3 NS_189 0 1.5379578601651994e-04
GC_3_190 b_3 NI_3 NS_190 0 1.3562047518786646e-04
GC_3_191 b_3 NI_3 NS_191 0 3.4705294744757421e-04
GC_3_192 b_3 NI_3 NS_192 0 -2.3958200864389601e-05
GC_3_193 b_3 NI_3 NS_193 0 5.3192882103688584e-05
GC_3_194 b_3 NI_3 NS_194 0 -5.8496672742671524e-04
GC_3_195 b_3 NI_3 NS_195 0 -1.4500295519276541e-04
GC_3_196 b_3 NI_3 NS_196 0 -6.8356343779096886e-05
GC_3_197 b_3 NI_3 NS_197 0 5.2203008415706122e-05
GC_3_198 b_3 NI_3 NS_198 0 -1.0716135874094718e-05
GC_3_199 b_3 NI_3 NS_199 0 4.8321262735931685e-05
GC_3_200 b_3 NI_3 NS_200 0 -4.5206125141611343e-04
GC_3_201 b_3 NI_3 NS_201 0 -7.0676813595342016e-04
GC_3_202 b_3 NI_3 NS_202 0 -8.3391004072922665e-05
GC_3_203 b_3 NI_3 NS_203 0 -1.7416244013703714e-04
GC_3_204 b_3 NI_3 NS_204 0 2.5967712440539683e-04
GC_3_205 b_3 NI_3 NS_205 0 1.0231320567971857e-04
GC_3_206 b_3 NI_3 NS_206 0 8.1092295578115954e-05
GC_3_207 b_3 NI_3 NS_207 0 -1.2122268443947334e-04
GC_3_208 b_3 NI_3 NS_208 0 -3.3414336225095429e-04
GC_3_209 b_3 NI_3 NS_209 0 -6.5847603818808798e-06
GC_3_210 b_3 NI_3 NS_210 0 9.9213319831600047e-05
GC_3_211 b_3 NI_3 NS_211 0 6.2415131154366316e-11
GC_3_212 b_3 NI_3 NS_212 0 -2.6617586479923546e-09
GC_3_213 b_3 NI_3 NS_213 0 -1.4903987536630648e-06
GC_3_214 b_3 NI_3 NS_214 0 -1.5556252129760585e-06
GC_3_215 b_3 NI_3 NS_215 0 -2.8329164324702218e-06
GC_3_216 b_3 NI_3 NS_216 0 -1.5878871543417275e-06
GC_3_217 b_3 NI_3 NS_217 0 -5.7178315259162902e-06
GC_3_218 b_3 NI_3 NS_218 0 -1.2614687092253027e-06
GC_3_219 b_3 NI_3 NS_219 0 -8.7595715862229738e-06
GC_3_220 b_3 NI_3 NS_220 0 6.4067722655862017e-06
GC_3_221 b_3 NI_3 NS_221 0 -6.4092262137874498e-06
GC_3_222 b_3 NI_3 NS_222 0 5.1019634023081062e-06
GC_3_223 b_3 NI_3 NS_223 0 8.4424842599446349e-07
GC_3_224 b_3 NI_3 NS_224 0 5.8470280648618639e-06
GC_3_225 b_3 NI_3 NS_225 0 -5.3961664926369774e-06
GC_3_226 b_3 NI_3 NS_226 0 1.2705485550367252e-05
GC_3_227 b_3 NI_3 NS_227 0 1.0828082278185205e-05
GC_3_228 b_3 NI_3 NS_228 0 1.5435688369863068e-05
GC_3_229 b_3 NI_3 NS_229 0 4.5989180010126433e-06
GC_3_230 b_3 NI_3 NS_230 0 1.0589226617051396e-05
GC_3_231 b_3 NI_3 NS_231 0 4.7903817671815576e-06
GC_3_232 b_3 NI_3 NS_232 0 9.9605559200955675e-06
GC_3_233 b_3 NI_3 NS_233 0 -7.2520428832457856e-05
GC_3_234 b_3 NI_3 NS_234 0 1.2870703152971838e-05
GC_3_235 b_3 NI_3 NS_235 0 -2.7806074816832438e-05
GC_3_236 b_3 NI_3 NS_236 0 -1.1427881551387101e-06
GC_3_237 b_3 NI_3 NS_237 0 -5.6802035694943189e-11
GC_3_238 b_3 NI_3 NS_238 0 1.0423995954566527e-09
GC_3_239 b_3 NI_3 NS_239 0 3.7494145118105939e-06
GC_3_240 b_3 NI_3 NS_240 0 4.4298205556197143e-06
GC_3_241 b_3 NI_3 NS_241 0 3.3687708038228649e-06
GC_3_242 b_3 NI_3 NS_242 0 3.3453251536813733e-06
GC_3_243 b_3 NI_3 NS_243 0 1.0419182671523847e-05
GC_3_244 b_3 NI_3 NS_244 0 -2.9807487198253946e-06
GC_3_245 b_3 NI_3 NS_245 0 6.6061140311962803e-06
GC_3_246 b_3 NI_3 NS_246 0 -1.4562633344443451e-05
GC_3_247 b_3 NI_3 NS_247 0 -3.0165739234952864e-06
GC_3_248 b_3 NI_3 NS_248 0 -1.0861344325599288e-06
GC_3_249 b_3 NI_3 NS_249 0 9.4457583805531733e-07
GC_3_250 b_3 NI_3 NS_250 0 -8.3627617094515229e-07
GC_3_251 b_3 NI_3 NS_251 0 2.9369381335583886e-06
GC_3_252 b_3 NI_3 NS_252 0 -1.2938430988979259e-05
GC_3_253 b_3 NI_3 NS_253 0 -1.3690770973809242e-05
GC_3_254 b_3 NI_3 NS_254 0 -3.7596288498825921e-06
GC_3_255 b_3 NI_3 NS_255 0 -3.5380576151247757e-06
GC_3_256 b_3 NI_3 NS_256 0 5.8960606241290375e-06
GC_3_257 b_3 NI_3 NS_257 0 2.7026888174348565e-06
GC_3_258 b_3 NI_3 NS_258 0 1.1370565085542508e-06
GC_3_259 b_3 NI_3 NS_259 0 1.7480838788589756e-07
GC_3_260 b_3 NI_3 NS_260 0 -5.8082580507293183e-06
GC_3_261 b_3 NI_3 NS_261 0 -2.7798142854524363e-05
GC_3_262 b_3 NI_3 NS_262 0 4.2303141145124232e-05
GC_3_263 b_3 NI_3 NS_263 0 3.6714333362034118e-11
GC_3_264 b_3 NI_3 NS_264 0 -2.7999033024791157e-10
GC_3_265 b_3 NI_3 NS_265 0 8.4060976767613601e-07
GC_3_266 b_3 NI_3 NS_266 0 4.8887836393644475e-07
GC_3_267 b_3 NI_3 NS_267 0 4.0308547667066406e-07
GC_3_268 b_3 NI_3 NS_268 0 -7.5631255084728013e-07
GC_3_269 b_3 NI_3 NS_269 0 -4.8232154876024897e-07
GC_3_270 b_3 NI_3 NS_270 0 9.9488195042252646e-07
GC_3_271 b_3 NI_3 NS_271 0 1.4097771957525017e-06
GC_3_272 b_3 NI_3 NS_272 0 1.8137231775667854e-07
GC_3_273 b_3 NI_3 NS_273 0 -4.2612467521537589e-07
GC_3_274 b_3 NI_3 NS_274 0 9.6865223929925907e-07
GC_3_275 b_3 NI_3 NS_275 0 5.7062319632246095e-07
GC_3_276 b_3 NI_3 NS_276 0 3.8250637939789425e-07
GC_3_277 b_3 NI_3 NS_277 0 5.5583613182565810e-07
GC_3_278 b_3 NI_3 NS_278 0 3.2468888653428789e-06
GC_3_279 b_3 NI_3 NS_279 0 3.9989909668582593e-06
GC_3_280 b_3 NI_3 NS_280 0 7.7857571826667737e-07
GC_3_281 b_3 NI_3 NS_281 0 9.0089336252147338e-07
GC_3_282 b_3 NI_3 NS_282 0 2.3851796036987364e-06
GC_3_283 b_3 NI_3 NS_283 0 1.1489768963654322e-06
GC_3_284 b_3 NI_3 NS_284 0 2.6054711378053921e-06
GC_3_285 b_3 NI_3 NS_285 0 -3.3471211483493070e-05
GC_3_286 b_3 NI_3 NS_286 0 4.1446803567796845e-07
GC_3_287 b_3 NI_3 NS_287 0 -2.4857670369630849e-05
GC_3_288 b_3 NI_3 NS_288 0 2.0849041530606262e-05
GC_3_289 b_3 NI_3 NS_289 0 -3.5016449158392393e-11
GC_3_290 b_3 NI_3 NS_290 0 -2.6866768637991908e-10
GC_3_291 b_3 NI_3 NS_291 0 1.6181042982806810e-06
GC_3_292 b_3 NI_3 NS_292 0 1.4408615991123771e-06
GC_3_293 b_3 NI_3 NS_293 0 2.6029538698761269e-07
GC_3_294 b_3 NI_3 NS_294 0 3.7175588318349607e-07
GC_3_295 b_3 NI_3 NS_295 0 1.7426638793692759e-06
GC_3_296 b_3 NI_3 NS_296 0 -2.0560494178861525e-07
GC_3_297 b_3 NI_3 NS_297 0 3.3661173232563902e-06
GC_3_298 b_3 NI_3 NS_298 0 -1.0275561886429571e-06
GC_3_299 b_3 NI_3 NS_299 0 4.2278218276759095e-07
GC_3_300 b_3 NI_3 NS_300 0 5.1394819117921561e-08
GC_3_301 b_3 NI_3 NS_301 0 2.5478031858720284e-07
GC_3_302 b_3 NI_3 NS_302 0 -2.9686672710056205e-07
GC_3_303 b_3 NI_3 NS_303 0 1.0838533163576374e-06
GC_3_304 b_3 NI_3 NS_304 0 -1.0037664897517268e-06
GC_3_305 b_3 NI_3 NS_305 0 1.6365250367165171e-06
GC_3_306 b_3 NI_3 NS_306 0 -1.2094852132953001e-06
GC_3_307 b_3 NI_3 NS_307 0 -5.6831722482021317e-08
GC_3_308 b_3 NI_3 NS_308 0 1.3046585281873994e-06
GC_3_309 b_3 NI_3 NS_309 0 3.3320737075395556e-07
GC_3_310 b_3 NI_3 NS_310 0 6.8983861517195726e-07
GC_3_311 b_3 NI_3 NS_311 0 -1.7034656755013925e-05
GC_3_312 b_3 NI_3 NS_312 0 -1.3465976239531934e-06
GD_3_1 b_3 NI_3 NA_1 0 1.3427146547155393e-02
GD_3_2 b_3 NI_3 NA_2 0 -1.1219494580257225e-03
GD_3_3 b_3 NI_3 NA_3 0 -2.9744124750322880e-02
GD_3_4 b_3 NI_3 NA_4 0 -2.0423328898149025e-02
GD_3_5 b_3 NI_3 NA_5 0 3.0059663067590475e-03
GD_3_6 b_3 NI_3 NA_6 0 -5.3669734924334352e-05
GD_3_7 b_3 NI_3 NA_7 0 1.6665991007296593e-04
GD_3_8 b_3 NI_3 NA_8 0 1.4002895124831384e-04
GD_3_9 b_3 NI_3 NA_9 0 -5.5170916907957148e-06
GD_3_10 b_3 NI_3 NA_10 0 1.2646759995208690e-05
GD_3_11 b_3 NI_3 NA_11 0 8.8710180443092484e-06
GD_3_12 b_3 NI_3 NA_12 0 7.7472950043768064e-06
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 -1.3745704524143981e-03
GC_4_2 b_4 NI_4 NS_2 0 2.3328647395210685e-03
GC_4_3 b_4 NI_4 NS_3 0 7.5881762047053013e-10
GC_4_4 b_4 NI_4 NS_4 0 6.0065849893445642e-07
GC_4_5 b_4 NI_4 NS_5 0 -1.9596090230233331e-04
GC_4_6 b_4 NI_4 NS_6 0 -4.5533576214058211e-04
GC_4_7 b_4 NI_4 NS_7 0 -1.0665922629642707e-03
GC_4_8 b_4 NI_4 NS_8 0 -9.2132880623234468e-04
GC_4_9 b_4 NI_4 NS_9 0 -2.3173765230588388e-03
GC_4_10 b_4 NI_4 NS_10 0 3.1222083675853138e-04
GC_4_11 b_4 NI_4 NS_11 0 -3.4636422129769717e-04
GC_4_12 b_4 NI_4 NS_12 0 4.1981894757741473e-03
GC_4_13 b_4 NI_4 NS_13 0 9.7828934157408783e-04
GC_4_14 b_4 NI_4 NS_14 0 4.4367342791590996e-04
GC_4_15 b_4 NI_4 NS_15 0 -3.7329545534134069e-04
GC_4_16 b_4 NI_4 NS_16 0 7.9841425643603002e-05
GC_4_17 b_4 NI_4 NS_17 0 -3.1453904086243552e-04
GC_4_18 b_4 NI_4 NS_18 0 3.3540638111544791e-03
GC_4_19 b_4 NI_4 NS_19 0 5.2329406726914860e-03
GC_4_20 b_4 NI_4 NS_20 0 8.1285628531144996e-04
GC_4_21 b_4 NI_4 NS_21 0 1.3427545700296971e-03
GC_4_22 b_4 NI_4 NS_22 0 -1.9440140011326480e-03
GC_4_23 b_4 NI_4 NS_23 0 -8.8256221336732320e-04
GC_4_24 b_4 NI_4 NS_24 0 -6.3689647527060485e-04
GC_4_25 b_4 NI_4 NS_25 0 -1.4735564028731604e-03
GC_4_26 b_4 NI_4 NS_26 0 2.5664387104945507e-03
GC_4_27 b_4 NI_4 NS_27 0 -7.4986630406880259e-03
GC_4_28 b_4 NI_4 NS_28 0 5.4463679169777183e-03
GC_4_29 b_4 NI_4 NS_29 0 -8.2819008038089098e-10
GC_4_30 b_4 NI_4 NS_30 0 -1.6858207847886993e-06
GC_4_31 b_4 NI_4 NS_31 0 2.5534451679426766e-04
GC_4_32 b_4 NI_4 NS_32 0 2.6645209554603528e-03
GC_4_33 b_4 NI_4 NS_33 0 4.5291717763011269e-03
GC_4_34 b_4 NI_4 NS_34 0 -2.7565535280063180e-03
GC_4_35 b_4 NI_4 NS_35 0 -5.4227002238950873e-03
GC_4_36 b_4 NI_4 NS_36 0 4.2041125753594248e-04
GC_4_37 b_4 NI_4 NS_37 0 8.8584598590663519e-03
GC_4_38 b_4 NI_4 NS_38 0 -6.2093760062331509e-04
GC_4_39 b_4 NI_4 NS_39 0 -2.8260892311364077e-03
GC_4_40 b_4 NI_4 NS_40 0 -2.3963222379300756e-03
GC_4_41 b_4 NI_4 NS_41 0 4.3105191748283411e-05
GC_4_42 b_4 NI_4 NS_42 0 -2.1139049360767706e-03
GC_4_43 b_4 NI_4 NS_43 0 -3.5070335195684262e-03
GC_4_44 b_4 NI_4 NS_44 0 5.5496239602017567e-03
GC_4_45 b_4 NI_4 NS_45 0 5.0984928002371357e-03
GC_4_46 b_4 NI_4 NS_46 0 -7.7604182478625047e-03
GC_4_47 b_4 NI_4 NS_47 0 -5.0389112787701624e-03
GC_4_48 b_4 NI_4 NS_48 0 3.0962138594566690e-03
GC_4_49 b_4 NI_4 NS_49 0 2.2446237576854008e-03
GC_4_50 b_4 NI_4 NS_50 0 -1.6873402428930829e-03
GC_4_51 b_4 NI_4 NS_51 0 -5.9469780546735429e-03
GC_4_52 b_4 NI_4 NS_52 0 3.8164552896847552e-03
GC_4_53 b_4 NI_4 NS_53 0 -4.9957171150348791e-02
GC_4_54 b_4 NI_4 NS_54 0 1.0966254766647213e-01
GC_4_55 b_4 NI_4 NS_55 0 1.0579502503450345e-08
GC_4_56 b_4 NI_4 NS_56 0 1.9882065471578493e-05
GC_4_57 b_4 NI_4 NS_57 0 -1.5752613716051411e-02
GC_4_58 b_4 NI_4 NS_58 0 2.4251933466342305e-02
GC_4_59 b_4 NI_4 NS_59 0 -7.8021463651088557e-03
GC_4_60 b_4 NI_4 NS_60 0 -1.4485562172606811e-02
GC_4_61 b_4 NI_4 NS_61 0 2.0432744143053690e-02
GC_4_62 b_4 NI_4 NS_62 0 6.6858548403368363e-03
GC_4_63 b_4 NI_4 NS_63 0 8.0641362852953528e-03
GC_4_64 b_4 NI_4 NS_64 0 4.3992228987664410e-02
GC_4_65 b_4 NI_4 NS_65 0 -1.1854727694379910e-02
GC_4_66 b_4 NI_4 NS_66 0 -3.2297456753758512e-03
GC_4_67 b_4 NI_4 NS_67 0 -5.0941014801587125e-03
GC_4_68 b_4 NI_4 NS_68 0 -4.0920275291115409e-03
GC_4_69 b_4 NI_4 NS_69 0 2.6818339765882254e-02
GC_4_70 b_4 NI_4 NS_70 0 -1.0406834673073906e-05
GC_4_71 b_4 NI_4 NS_71 0 3.3876575470817197e-02
GC_4_72 b_4 NI_4 NS_72 0 3.0995855490232507e-02
GC_4_73 b_4 NI_4 NS_73 0 -1.5641055958966428e-02
GC_4_74 b_4 NI_4 NS_74 0 8.2858614273286120e-03
GC_4_75 b_4 NI_4 NS_75 0 -9.9915425314631352e-04
GC_4_76 b_4 NI_4 NS_76 0 -6.8608537523428244e-03
GC_4_77 b_4 NI_4 NS_77 0 -6.8944011918482498e-02
GC_4_78 b_4 NI_4 NS_78 0 1.7522301711185649e-03
GC_4_79 b_4 NI_4 NS_79 0 5.9438136073012800e-02
GC_4_80 b_4 NI_4 NS_80 0 -6.3779997448680292e-02
GC_4_81 b_4 NI_4 NS_81 0 -1.0218715257320815e-08
GC_4_82 b_4 NI_4 NS_82 0 -8.2100868785479630e-06
GC_4_83 b_4 NI_4 NS_83 0 -1.8519166209792902e-03
GC_4_84 b_4 NI_4 NS_84 0 -2.8731340475971201e-03
GC_4_85 b_4 NI_4 NS_85 0 -5.1084756720848569e-03
GC_4_86 b_4 NI_4 NS_86 0 1.9400114889521767e-03
GC_4_87 b_4 NI_4 NS_87 0 2.4463666578743953e-03
GC_4_88 b_4 NI_4 NS_88 0 -1.2255434516112895e-03
GC_4_89 b_4 NI_4 NS_89 0 -1.0650799674863392e-02
GC_4_90 b_4 NI_4 NS_90 0 1.1045689712411066e-03
GC_4_91 b_4 NI_4 NS_91 0 6.4145744822000084e-04
GC_4_92 b_4 NI_4 NS_92 0 1.7543170152112600e-03
GC_4_93 b_4 NI_4 NS_93 0 -9.5624673213744714e-04
GC_4_94 b_4 NI_4 NS_94 0 2.2871421137470368e-03
GC_4_95 b_4 NI_4 NS_95 0 5.9413739439217919e-04
GC_4_96 b_4 NI_4 NS_96 0 -5.8937142081883801e-03
GC_4_97 b_4 NI_4 NS_97 0 -8.5380811876149317e-03
GC_4_98 b_4 NI_4 NS_98 0 6.8906920148833952e-03
GC_4_99 b_4 NI_4 NS_99 0 2.5187097649788455e-03
GC_4_100 b_4 NI_4 NS_100 0 -3.6778740922647898e-03
GC_4_101 b_4 NI_4 NS_101 0 -2.6381595052563131e-03
GC_4_102 b_4 NI_4 NS_102 0 -5.1433834238558021e-04
GC_4_103 b_4 NI_4 NS_103 0 5.4574972974247099e-02
GC_4_104 b_4 NI_4 NS_104 0 1.6205496302430103e-03
GC_4_105 b_4 NI_4 NS_105 0 -1.0993209339224840e-03
GC_4_106 b_4 NI_4 NS_106 0 1.9264488656125750e-03
GC_4_107 b_4 NI_4 NS_107 0 -9.9960441286759736e-11
GC_4_108 b_4 NI_4 NS_108 0 2.7260538805754594e-07
GC_4_109 b_4 NI_4 NS_109 0 5.8933463524565789e-05
GC_4_110 b_4 NI_4 NS_110 0 -8.7080058169892392e-05
GC_4_111 b_4 NI_4 NS_111 0 -2.6160836006586041e-04
GC_4_112 b_4 NI_4 NS_112 0 -1.7078573466833009e-04
GC_4_113 b_4 NI_4 NS_113 0 -5.2946919283830443e-04
GC_4_114 b_4 NI_4 NS_114 0 2.5259348619175401e-05
GC_4_115 b_4 NI_4 NS_115 0 4.2452468540268967e-05
GC_4_116 b_4 NI_4 NS_116 0 9.1569635473157530e-04
GC_4_117 b_4 NI_4 NS_117 0 2.4558828723111577e-04
GC_4_118 b_4 NI_4 NS_118 0 1.3071939791781717e-04
GC_4_119 b_4 NI_4 NS_119 0 -8.1498481443712531e-05
GC_4_120 b_4 NI_4 NS_120 0 2.6844114957338603e-05
GC_4_121 b_4 NI_4 NS_121 0 -7.0951258142956750e-05
GC_4_122 b_4 NI_4 NS_122 0 7.5354268404910062e-04
GC_4_123 b_4 NI_4 NS_123 0 1.2758086640151712e-03
GC_4_124 b_4 NI_4 NS_124 0 1.3799804233122792e-04
GC_4_125 b_4 NI_4 NS_125 0 3.2406021056442038e-04
GC_4_126 b_4 NI_4 NS_126 0 -4.2268318011576180e-04
GC_4_127 b_4 NI_4 NS_127 0 -2.4533855424971698e-04
GC_4_128 b_4 NI_4 NS_128 0 -1.0928505594099719e-04
GC_4_129 b_4 NI_4 NS_129 0 -1.5485139694443688e-03
GC_4_130 b_4 NI_4 NS_130 0 3.7255016766295186e-04
GC_4_131 b_4 NI_4 NS_131 0 -1.2121033466286288e-03
GC_4_132 b_4 NI_4 NS_132 0 5.5290802303188029e-04
GC_4_133 b_4 NI_4 NS_133 0 3.0006236193976750e-10
GC_4_134 b_4 NI_4 NS_134 0 -5.7499769591845096e-07
GC_4_135 b_4 NI_4 NS_135 0 3.1148052460973771e-05
GC_4_136 b_4 NI_4 NS_136 0 6.3814449314533533e-04
GC_4_137 b_4 NI_4 NS_137 0 1.0887951204821918e-03
GC_4_138 b_4 NI_4 NS_138 0 -6.7568288688358452e-04
GC_4_139 b_4 NI_4 NS_139 0 -1.3741759156993016e-03
GC_4_140 b_4 NI_4 NS_140 0 7.5249034282641339e-05
GC_4_141 b_4 NI_4 NS_141 0 2.0942445835718886e-03
GC_4_142 b_4 NI_4 NS_142 0 -1.0656098416821037e-04
GC_4_143 b_4 NI_4 NS_143 0 -7.3383076274294496e-04
GC_4_144 b_4 NI_4 NS_144 0 -5.7289970345373632e-04
GC_4_145 b_4 NI_4 NS_145 0 5.7546542128135375e-06
GC_4_146 b_4 NI_4 NS_146 0 -4.8779049432463406e-04
GC_4_147 b_4 NI_4 NS_147 0 -9.0586763068732450e-04
GC_4_148 b_4 NI_4 NS_148 0 1.3910529642514643e-03
GC_4_149 b_4 NI_4 NS_149 0 1.2473508898539992e-03
GC_4_150 b_4 NI_4 NS_150 0 -1.8369115743053250e-03
GC_4_151 b_4 NI_4 NS_151 0 -1.2248397785880110e-03
GC_4_152 b_4 NI_4 NS_152 0 7.8178305795523586e-04
GC_4_153 b_4 NI_4 NS_153 0 5.7543619705362106e-04
GC_4_154 b_4 NI_4 NS_154 0 -4.1190350944532602e-04
GC_4_155 b_4 NI_4 NS_155 0 -7.3189010619247399e-04
GC_4_156 b_4 NI_4 NS_156 0 1.1403220193143056e-03
GC_4_157 b_4 NI_4 NS_157 0 1.2876638751917045e-04
GC_4_158 b_4 NI_4 NS_158 0 5.3481972218915412e-05
GC_4_159 b_4 NI_4 NS_159 0 -4.2223195227664243e-10
GC_4_160 b_4 NI_4 NS_160 0 4.4745787412401936e-08
GC_4_161 b_4 NI_4 NS_161 0 5.7031009153498582e-06
GC_4_162 b_4 NI_4 NS_162 0 7.6084236064349057e-05
GC_4_163 b_4 NI_4 NS_163 0 1.5379601437865901e-04
GC_4_164 b_4 NI_4 NS_164 0 1.3562073377256556e-04
GC_4_165 b_4 NI_4 NS_165 0 3.4705326893460993e-04
GC_4_166 b_4 NI_4 NS_166 0 -2.3957912838638233e-05
GC_4_167 b_4 NI_4 NS_167 0 5.3193170814912721e-05
GC_4_168 b_4 NI_4 NS_168 0 -5.8496731938962123e-04
GC_4_169 b_4 NI_4 NS_169 0 -1.4500299471755077e-04
GC_4_170 b_4 NI_4 NS_170 0 -6.8356434737079663e-05
GC_4_171 b_4 NI_4 NS_171 0 5.2203095731019962e-05
GC_4_172 b_4 NI_4 NS_172 0 -1.0716015711468124e-05
GC_4_173 b_4 NI_4 NS_173 0 4.8321453309180503e-05
GC_4_174 b_4 NI_4 NS_174 0 -4.5206117137884777e-04
GC_4_175 b_4 NI_4 NS_175 0 -7.0676797156918921e-04
GC_4_176 b_4 NI_4 NS_176 0 -8.3391432965468425e-05
GC_4_177 b_4 NI_4 NS_177 0 -1.7416249565983339e-04
GC_4_178 b_4 NI_4 NS_178 0 2.5967704037050857e-04
GC_4_179 b_4 NI_4 NS_179 0 1.0231312799229876e-04
GC_4_180 b_4 NI_4 NS_180 0 8.1092285069053665e-05
GC_4_181 b_4 NI_4 NS_181 0 -1.2122385233829181e-04
GC_4_182 b_4 NI_4 NS_182 0 -3.3414360871326384e-04
GC_4_183 b_4 NI_4 NS_183 0 3.8540474142399674e-04
GC_4_184 b_4 NI_4 NS_184 0 -2.0233222536518063e-03
GC_4_185 b_4 NI_4 NS_185 0 4.0275552388057325e-10
GC_4_186 b_4 NI_4 NS_186 0 -2.6921603068563400e-08
GC_4_187 b_4 NI_4 NS_187 0 1.8880649696595821e-05
GC_4_188 b_4 NI_4 NS_188 0 4.3647508446278926e-05
GC_4_189 b_4 NI_4 NS_189 0 8.2161768404037707e-05
GC_4_190 b_4 NI_4 NS_190 0 -3.0679914494658285e-05
GC_4_191 b_4 NI_4 NS_191 0 -1.3443168508774842e-05
GC_4_192 b_4 NI_4 NS_192 0 1.3855590453880693e-05
GC_4_193 b_4 NI_4 NS_193 0 1.9803314084096464e-04
GC_4_194 b_4 NI_4 NS_194 0 -9.9134359268100394e-05
GC_4_195 b_4 NI_4 NS_195 0 2.7217482448308429e-05
GC_4_196 b_4 NI_4 NS_196 0 -9.8066136220361047e-05
GC_4_197 b_4 NI_4 NS_197 0 -1.7281658639674792e-05
GC_4_198 b_4 NI_4 NS_198 0 -9.8320967800103818e-05
GC_4_199 b_4 NI_4 NS_199 0 1.0631279048776298e-05
GC_4_200 b_4 NI_4 NS_200 0 -9.7299760656496535e-05
GC_4_201 b_4 NI_4 NS_201 0 -9.7211317437836814e-05
GC_4_202 b_4 NI_4 NS_202 0 -3.1576826254973230e-04
GC_4_203 b_4 NI_4 NS_203 0 -1.3368399231110078e-04
GC_4_204 b_4 NI_4 NS_204 0 -1.1528087978189936e-04
GC_4_205 b_4 NI_4 NS_205 0 -1.9126644286043095e-05
GC_4_206 b_4 NI_4 NS_206 0 -1.9117075076664015e-04
GC_4_207 b_4 NI_4 NS_207 0 1.5269827578651123e-03
GC_4_208 b_4 NI_4 NS_208 0 -9.9579655979461820e-05
GC_4_209 b_4 NI_4 NS_209 0 -2.7846432955870934e-05
GC_4_210 b_4 NI_4 NS_210 0 -1.1271728516093679e-06
GC_4_211 b_4 NI_4 NS_211 0 -5.6801599613188399e-11
GC_4_212 b_4 NI_4 NS_212 0 1.0421524662313318e-09
GC_4_213 b_4 NI_4 NS_213 0 3.7467179568558645e-06
GC_4_214 b_4 NI_4 NS_214 0 4.4128223052690662e-06
GC_4_215 b_4 NI_4 NS_215 0 3.3691630902850393e-06
GC_4_216 b_4 NI_4 NS_216 0 3.3616308858683882e-06
GC_4_217 b_4 NI_4 NS_217 0 1.0412999108337805e-05
GC_4_218 b_4 NI_4 NS_218 0 -2.9646621954399048e-06
GC_4_219 b_4 NI_4 NS_219 0 6.6233921179004571e-06
GC_4_220 b_4 NI_4 NS_220 0 -1.4577523668335172e-05
GC_4_221 b_4 NI_4 NS_221 0 -3.0131490707252050e-06
GC_4_222 b_4 NI_4 NS_222 0 -1.0905306776746729e-06
GC_4_223 b_4 NI_4 NS_223 0 9.4683076610660131e-07
GC_4_224 b_4 NI_4 NS_224 0 -8.3289932561304442e-07
GC_4_225 b_4 NI_4 NS_225 0 2.9441078002497657e-06
GC_4_226 b_4 NI_4 NS_226 0 -1.2938321176440312e-05
GC_4_227 b_4 NI_4 NS_227 0 -1.3694224642961080e-05
GC_4_228 b_4 NI_4 NS_228 0 -3.7760568196150076e-06
GC_4_229 b_4 NI_4 NS_229 0 -3.5424629858071511e-06
GC_4_230 b_4 NI_4 NS_230 0 5.8948709211703688e-06
GC_4_231 b_4 NI_4 NS_231 0 2.7008062272249341e-06
GC_4_232 b_4 NI_4 NS_232 0 1.1398779357831484e-06
GC_4_233 b_4 NI_4 NS_233 0 1.6185214306611624e-07
GC_4_234 b_4 NI_4 NS_234 0 -5.8089506098406671e-06
GC_4_235 b_4 NI_4 NS_235 0 -6.5847274316232357e-06
GC_4_236 b_4 NI_4 NS_236 0 9.9213278830947481e-05
GC_4_237 b_4 NI_4 NS_237 0 6.2415148832688892e-11
GC_4_238 b_4 NI_4 NS_238 0 -2.6617613128754473e-09
GC_4_239 b_4 NI_4 NS_239 0 -1.4903849485570984e-06
GC_4_240 b_4 NI_4 NS_240 0 -1.5556180071871688e-06
GC_4_241 b_4 NI_4 NS_241 0 -2.8329214595575688e-06
GC_4_242 b_4 NI_4 NS_242 0 -1.5879025458407536e-06
GC_4_243 b_4 NI_4 NS_243 0 -5.7178311398913939e-06
GC_4_244 b_4 NI_4 NS_244 0 -1.2614456170925704e-06
GC_4_245 b_4 NI_4 NS_245 0 -8.7595590080001223e-06
GC_4_246 b_4 NI_4 NS_246 0 6.4067485120221006e-06
GC_4_247 b_4 NI_4 NS_247 0 -6.4092312427770325e-06
GC_4_248 b_4 NI_4 NS_248 0 5.1019689501870078e-06
GC_4_249 b_4 NI_4 NS_249 0 8.4424484060106138e-07
GC_4_250 b_4 NI_4 NS_250 0 5.8470265130137457e-06
GC_4_251 b_4 NI_4 NS_251 0 -5.3961581623201367e-06
GC_4_252 b_4 NI_4 NS_252 0 1.2705497030195292e-05
GC_4_253 b_4 NI_4 NS_253 0 1.0828083287608439e-05
GC_4_254 b_4 NI_4 NS_254 0 1.5435675860371473e-05
GC_4_255 b_4 NI_4 NS_255 0 4.5989210084376476e-06
GC_4_256 b_4 NI_4 NS_256 0 1.0589226873889853e-05
GC_4_257 b_4 NI_4 NS_257 0 4.7903833024200509e-06
GC_4_258 b_4 NI_4 NS_258 0 9.9605484168792795e-06
GC_4_259 b_4 NI_4 NS_259 0 -7.2520399708693475e-05
GC_4_260 b_4 NI_4 NS_260 0 1.2870693321977114e-05
GC_4_261 b_4 NI_4 NS_261 0 -2.4858860148582116e-05
GC_4_262 b_4 NI_4 NS_262 0 2.0849541966624160e-05
GC_4_263 b_4 NI_4 NS_263 0 -3.5016417164848383e-11
GC_4_264 b_4 NI_4 NS_264 0 -2.6867101844036285e-10
GC_4_265 b_4 NI_4 NS_265 0 1.6182387100459861e-06
GC_4_266 b_4 NI_4 NS_266 0 1.4407743178202215e-06
GC_4_267 b_4 NI_4 NS_267 0 2.6022691975076801e-07
GC_4_268 b_4 NI_4 NS_268 0 3.7182517957361018e-07
GC_4_269 b_4 NI_4 NS_269 0 1.7425642394347806e-06
GC_4_270 b_4 NI_4 NS_270 0 -2.0555215435708460e-07
GC_4_271 b_4 NI_4 NS_271 0 3.3663628004412667e-06
GC_4_272 b_4 NI_4 NS_272 0 -1.0275575052314812e-06
GC_4_273 b_4 NI_4 NS_273 0 4.2285821666231169e-07
GC_4_274 b_4 NI_4 NS_274 0 5.1377028313063920e-08
GC_4_275 b_4 NI_4 NS_275 0 2.5477392734705698e-07
GC_4_276 b_4 NI_4 NS_276 0 -2.9685421799281024e-07
GC_4_277 b_4 NI_4 NS_277 0 1.0839096462961449e-06
GC_4_278 b_4 NI_4 NS_278 0 -1.0037312530528527e-06
GC_4_279 b_4 NI_4 NS_279 0 1.6366703576228641e-06
GC_4_280 b_4 NI_4 NS_280 0 -1.2095530647919578e-06
GC_4_281 b_4 NI_4 NS_281 0 -5.6794123695268620e-08
GC_4_282 b_4 NI_4 NS_282 0 1.3046417900450877e-06
GC_4_283 b_4 NI_4 NS_283 0 3.3322385508512826e-07
GC_4_284 b_4 NI_4 NS_284 0 6.8985930905650508e-07
GC_4_285 b_4 NI_4 NS_285 0 -1.7035034668298009e-05
GC_4_286 b_4 NI_4 NS_286 0 -1.3465760203921544e-06
GC_4_287 b_4 NI_4 NS_287 0 -2.7887633963388702e-05
GC_4_288 b_4 NI_4 NS_288 0 4.2423615486811728e-05
GC_4_289 b_4 NI_4 NS_289 0 3.6713791018910376e-11
GC_4_290 b_4 NI_4 NS_290 0 -2.8057040295841019e-10
GC_4_291 b_4 NI_4 NS_291 0 8.4282344685049989e-07
GC_4_292 b_4 NI_4 NS_292 0 4.8528865549570143e-07
GC_4_293 b_4 NI_4 NS_293 0 4.0300515655130835e-07
GC_4_294 b_4 NI_4 NS_294 0 -7.5313821654529246e-07
GC_4_295 b_4 NI_4 NS_295 0 -4.7580777485730920e-07
GC_4_296 b_4 NI_4 NS_296 0 9.9091369637113515e-07
GC_4_297 b_4 NI_4 NS_297 0 1.4076893751276455e-06
GC_4_298 b_4 NI_4 NS_298 0 1.8309231778812143e-07
GC_4_299 b_4 NI_4 NS_299 0 -4.2172399557456874e-07
GC_4_300 b_4 NI_4 NS_300 0 9.6747368032554851e-07
GC_4_301 b_4 NI_4 NS_301 0 5.7161783311229323e-07
GC_4_302 b_4 NI_4 NS_302 0 3.8276271834516744e-07
GC_4_303 b_4 NI_4 NS_303 0 5.5777862407850857e-07
GC_4_304 b_4 NI_4 NS_304 0 3.2436840808789862e-06
GC_4_305 b_4 NI_4 NS_305 0 3.9996423381050667e-06
GC_4_306 b_4 NI_4 NS_306 0 7.8349351928560944e-07
GC_4_307 b_4 NI_4 NS_307 0 9.0316508783260223e-07
GC_4_308 b_4 NI_4 NS_308 0 2.3897394850790474e-06
GC_4_309 b_4 NI_4 NS_309 0 1.1491003222692528e-06
GC_4_310 b_4 NI_4 NS_310 0 2.6121086810137782e-06
GC_4_311 b_4 NI_4 NS_311 0 -3.3569338745703027e-05
GC_4_312 b_4 NI_4 NS_312 0 4.1045995230193090e-07
GD_4_1 b_4 NI_4 NA_1 0 -1.1219611508926921e-03
GD_4_2 b_4 NI_4 NA_2 0 1.3427304153556871e-02
GD_4_3 b_4 NI_4 NA_3 0 -2.0423391285306812e-02
GD_4_4 b_4 NI_4 NA_4 0 -2.9744124750322714e-02
GD_4_5 b_4 NI_4 NA_5 0 -5.3604005821996413e-05
GD_4_6 b_4 NI_4 NA_6 0 3.0059891770120553e-03
GD_4_7 b_4 NI_4 NA_7 0 1.4002930277488501e-04
GD_4_8 b_4 NI_4 NA_8 0 1.6665145175970050e-04
GD_4_9 b_4 NI_4 NA_9 0 1.2667335689303253e-05
GD_4_10 b_4 NI_4 NA_10 0 -5.5171968108644407e-06
GD_4_11 b_4 NI_4 NA_11 0 7.7476748188097460e-06
GD_4_12 b_4 NI_4 NA_12 0 8.9205540572978247e-06
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 3.9467687032897691e-04
GC_5_2 b_5 NI_5 NS_2 0 -2.0170416171539402e-03
GC_5_3 b_5 NI_5 NS_3 0 4.0764937719759125e-10
GC_5_4 b_5 NI_5 NS_4 0 -2.7091784441528768e-08
GC_5_5 b_5 NI_5 NS_5 0 1.8629832432254174e-05
GC_5_6 b_5 NI_5 NS_6 0 4.3391935931797746e-05
GC_5_7 b_5 NI_5 NS_7 0 8.1680057416494116e-05
GC_5_8 b_5 NI_5 NS_8 0 -3.0853931520430810e-05
GC_5_9 b_5 NI_5 NS_9 0 -1.3841629986494910e-05
GC_5_10 b_5 NI_5 NS_10 0 1.3779023024987995e-05
GC_5_11 b_5 NI_5 NS_11 0 1.9715185655194513e-04
GC_5_12 b_5 NI_5 NS_12 0 -9.9073456462967906e-05
GC_5_13 b_5 NI_5 NS_13 0 2.6774533889887827e-05
GC_5_14 b_5 NI_5 NS_14 0 -9.8009285487182359e-05
GC_5_15 b_5 NI_5 NS_15 0 -1.7495832625523529e-05
GC_5_16 b_5 NI_5 NS_16 0 -9.8105913661928975e-05
GC_5_17 b_5 NI_5 NS_17 0 9.9651051412419351e-06
GC_5_18 b_5 NI_5 NS_18 0 -9.7431746421277498e-05
GC_5_19 b_5 NI_5 NS_19 0 -9.8104245280797065e-05
GC_5_20 b_5 NI_5 NS_20 0 -3.1498379012328783e-04
GC_5_21 b_5 NI_5 NS_21 0 -1.3390325912625319e-04
GC_5_22 b_5 NI_5 NS_22 0 -1.1512948993539613e-04
GC_5_23 b_5 NI_5 NS_23 0 -1.9651413973917018e-05
GC_5_24 b_5 NI_5 NS_24 0 -1.9128949089743555e-04
GC_5_25 b_5 NI_5 NS_25 0 1.5206724221139792e-03
GC_5_26 b_5 NI_5 NS_26 0 -1.0185406213861956e-04
GC_5_27 b_5 NI_5 NS_27 0 1.5161331202599761e-04
GC_5_28 b_5 NI_5 NS_28 0 1.2758695189803312e-05
GC_5_29 b_5 NI_5 NS_29 0 -4.2742748854259139e-10
GC_5_30 b_5 NI_5 NS_30 0 4.5130525477756281e-08
GC_5_31 b_5 NI_5 NS_31 0 5.1582437104964261e-06
GC_5_32 b_5 NI_5 NS_32 0 7.5618140244996246e-05
GC_5_33 b_5 NI_5 NS_33 0 1.5335293777481984e-04
GC_5_34 b_5 NI_5 NS_34 0 1.3548425737556116e-04
GC_5_35 b_5 NI_5 NS_35 0 3.4656235537696757e-04
GC_5_36 b_5 NI_5 NS_36 0 -2.4743470229438334e-05
GC_5_37 b_5 NI_5 NS_37 0 5.1564519903269019e-05
GC_5_38 b_5 NI_5 NS_38 0 -5.8538770221130715e-04
GC_5_39 b_5 NI_5 NS_39 0 -1.4593695891179642e-04
GC_5_40 b_5 NI_5 NS_40 0 -6.8387289374700059e-05
GC_5_41 b_5 NI_5 NS_41 0 5.1712590612903231e-05
GC_5_42 b_5 NI_5 NS_42 0 -1.0508142976454757e-05
GC_5_43 b_5 NI_5 NS_43 0 4.7728655042746513e-05
GC_5_44 b_5 NI_5 NS_44 0 -4.5313210307075508e-04
GC_5_45 b_5 NI_5 NS_45 0 -7.0919247553276863e-04
GC_5_46 b_5 NI_5 NS_46 0 -8.3324118971539533e-05
GC_5_47 b_5 NI_5 NS_47 0 -1.7472496339957695e-04
GC_5_48 b_5 NI_5 NS_48 0 2.5870543245382012e-04
GC_5_49 b_5 NI_5 NS_49 0 1.0249916219591510e-04
GC_5_50 b_5 NI_5 NS_50 0 7.9809616443885271e-05
GC_5_51 b_5 NI_5 NS_51 0 -8.6720207596101167e-05
GC_5_52 b_5 NI_5 NS_52 0 -3.2996574253456849e-04
GC_5_53 b_5 NI_5 NS_53 0 -1.2121033466290173e-03
GC_5_54 b_5 NI_5 NS_54 0 5.5290802303253114e-04
GC_5_55 b_5 NI_5 NS_55 0 3.0006236193993707e-10
GC_5_56 b_5 NI_5 NS_56 0 -5.7499769591846694e-07
GC_5_57 b_5 NI_5 NS_57 0 3.1148052460964067e-05
GC_5_58 b_5 NI_5 NS_58 0 6.3814449314533327e-04
GC_5_59 b_5 NI_5 NS_59 0 1.0887951204821729e-03
GC_5_60 b_5 NI_5 NS_60 0 -6.7568288688357617e-04
GC_5_61 b_5 NI_5 NS_61 0 -1.3741759156993393e-03
GC_5_62 b_5 NI_5 NS_62 0 7.5249034282667333e-05
GC_5_63 b_5 NI_5 NS_63 0 2.0942445835719211e-03
GC_5_64 b_5 NI_5 NS_64 0 -1.0656098416810272e-04
GC_5_65 b_5 NI_5 NS_65 0 -7.3383076274290138e-04
GC_5_66 b_5 NI_5 NS_66 0 -5.7289970345369772e-04
GC_5_67 b_5 NI_5 NS_67 0 5.7546542128465117e-06
GC_5_68 b_5 NI_5 NS_68 0 -4.8779049432464197e-04
GC_5_69 b_5 NI_5 NS_69 0 -9.0586763068728276e-04
GC_5_70 b_5 NI_5 NS_70 0 1.3910529642514966e-03
GC_5_71 b_5 NI_5 NS_71 0 1.2473508898540714e-03
GC_5_72 b_5 NI_5 NS_72 0 -1.8369115743053250e-03
GC_5_73 b_5 NI_5 NS_73 0 -1.2248397785879839e-03
GC_5_74 b_5 NI_5 NS_74 0 7.8178305795525017e-04
GC_5_75 b_5 NI_5 NS_75 0 5.7543619705362984e-04
GC_5_76 b_5 NI_5 NS_76 0 -4.1190350944529750e-04
GC_5_77 b_5 NI_5 NS_77 0 -7.3189010619300124e-04
GC_5_78 b_5 NI_5 NS_78 0 1.1403220193142794e-03
GC_5_79 b_5 NI_5 NS_79 0 -1.0992736657821672e-03
GC_5_80 b_5 NI_5 NS_80 0 1.9265919499781867e-03
GC_5_81 b_5 NI_5 NS_81 0 -9.9958119731328968e-11
GC_5_82 b_5 NI_5 NS_82 0 2.7260434700994913e-07
GC_5_83 b_5 NI_5 NS_83 0 5.8942674719951255e-05
GC_5_84 b_5 NI_5 NS_84 0 -8.7011292073306917e-05
GC_5_85 b_5 NI_5 NS_85 0 -2.6161328109190328e-04
GC_5_86 b_5 NI_5 NS_86 0 -1.7084760208701700e-04
GC_5_87 b_5 NI_5 NS_87 0 -5.2945252103955777e-04
GC_5_88 b_5 NI_5 NS_88 0 2.5205537233216399e-05
GC_5_89 b_5 NI_5 NS_89 0 4.2398994481917676e-05
GC_5_90 b_5 NI_5 NS_90 0 9.1577025531136059e-04
GC_5_91 b_5 NI_5 NS_91 0 2.4558174024738897e-04
GC_5_92 b_5 NI_5 NS_92 0 1.3074070442489565e-04
GC_5_93 b_5 NI_5 NS_93 0 -8.1504628241374299e-05
GC_5_94 b_5 NI_5 NS_94 0 2.6832875303487565e-05
GC_5_95 b_5 NI_5 NS_95 0 -7.0975044167335402e-05
GC_5_96 b_5 NI_5 NS_96 0 7.5355454260140784e-04
GC_5_97 b_5 NI_5 NS_97 0 1.2758459284037086e-03
GC_5_98 b_5 NI_5 NS_98 0 1.3806943399139474e-04
GC_5_99 b_5 NI_5 NS_99 0 3.2408622636345615e-04
GC_5_100 b_5 NI_5 NS_100 0 -4.2267378930148234e-04
GC_5_101 b_5 NI_5 NS_101 0 -2.4532879446818948e-04
GC_5_102 b_5 NI_5 NS_102 0 -1.0928772673865638e-04
GC_5_103 b_5 NI_5 NS_103 0 -1.5486299047001420e-03
GC_5_104 b_5 NI_5 NS_104 0 3.7254268685880970e-04
GC_5_105 b_5 NI_5 NS_105 0 5.9215489962724764e-02
GC_5_106 b_5 NI_5 NS_106 0 -6.3407636300857259e-02
GC_5_107 b_5 NI_5 NS_107 0 -1.0211750104087057e-08
GC_5_108 b_5 NI_5 NS_108 0 -8.2108571934109275e-06
GC_5_109 b_5 NI_5 NS_109 0 -1.8466567588426846e-03
GC_5_110 b_5 NI_5 NS_110 0 -2.8683123701404847e-03
GC_5_111 b_5 NI_5 NS_111 0 -5.1018049687674870e-03
GC_5_112 b_5 NI_5 NS_112 0 1.9432405042730510e-03
GC_5_113 b_5 NI_5 NS_113 0 2.4539731021212363e-03
GC_5_114 b_5 NI_5 NS_114 0 -1.2214745377999380e-03
GC_5_115 b_5 NI_5 NS_115 0 -1.0637008586728598e-02
GC_5_116 b_5 NI_5 NS_116 0 1.1057795139107671e-03
GC_5_117 b_5 NI_5 NS_117 0 6.4906104355947421e-04
GC_5_118 b_5 NI_5 NS_118 0 1.7568055400822653e-03
GC_5_119 b_5 NI_5 NS_119 0 -9.5190922325557995e-04
GC_5_120 b_5 NI_5 NS_120 0 2.2857457167483677e-03
GC_5_121 b_5 NI_5 NS_121 0 6.0496281193835977e-04
GC_5_122 b_5 NI_5 NS_122 0 -5.8869625838110801e-03
GC_5_123 b_5 NI_5 NS_123 0 -8.5212789070572975e-03
GC_5_124 b_5 NI_5 NS_124 0 6.8916057982835064e-03
GC_5_125 b_5 NI_5 NS_125 0 2.5250257717987518e-03
GC_5_126 b_5 NI_5 NS_126 0 -3.6699130634487071e-03
GC_5_127 b_5 NI_5 NS_127 0 -2.6398888960123277e-03
GC_5_128 b_5 NI_5 NS_128 0 -5.0014762094001321e-04
GC_5_129 b_5 NI_5 NS_129 0 5.4262590367559010e-02
GC_5_130 b_5 NI_5 NS_130 0 1.5891713896911003e-03
GC_5_131 b_5 NI_5 NS_131 0 -4.9912563744016029e-02
GC_5_132 b_5 NI_5 NS_132 0 1.0946196122956110e-01
GC_5_133 b_5 NI_5 NS_133 0 1.0782684477160389e-08
GC_5_134 b_5 NI_5 NS_134 0 1.9879857699720465e-05
GC_5_135 b_5 NI_5 NS_135 0 -1.5753192442280312e-02
GC_5_136 b_5 NI_5 NS_136 0 2.4251006398907114e-02
GC_5_137 b_5 NI_5 NS_137 0 -7.8027687570088209e-03
GC_5_138 b_5 NI_5 NS_138 0 -1.4488573082192722e-02
GC_5_139 b_5 NI_5 NS_139 0 2.0433212269113828e-02
GC_5_140 b_5 NI_5 NS_140 0 6.6873577305288567e-03
GC_5_141 b_5 NI_5 NS_141 0 8.0583335496318461e-03
GC_5_142 b_5 NI_5 NS_142 0 4.3992668860862172e-02
GC_5_143 b_5 NI_5 NS_143 0 -1.1853720034492695e-02
GC_5_144 b_5 NI_5 NS_144 0 -3.2338870078374906e-03
GC_5_145 b_5 NI_5 NS_145 0 -5.0942080903603965e-03
GC_5_146 b_5 NI_5 NS_146 0 -4.0938825194097219e-03
GC_5_147 b_5 NI_5 NS_147 0 2.6816834479478937e-02
GC_5_148 b_5 NI_5 NS_148 0 -8.8216820012392885e-06
GC_5_149 b_5 NI_5 NS_149 0 3.3872764837874686e-02
GC_5_150 b_5 NI_5 NS_150 0 3.0990203991718819e-02
GC_5_151 b_5 NI_5 NS_151 0 -1.5640925585210644e-02
GC_5_152 b_5 NI_5 NS_152 0 8.2834129277136442e-03
GC_5_153 b_5 NI_5 NS_153 0 -9.9439840955380479e-04
GC_5_154 b_5 NI_5 NS_154 0 -6.8670016975417294e-03
GC_5_155 b_5 NI_5 NS_155 0 -6.8769710450590035e-02
GC_5_156 b_5 NI_5 NS_156 0 1.7777698504401580e-03
GC_5_157 b_5 NI_5 NS_157 0 -7.6472780163478818e-03
GC_5_158 b_5 NI_5 NS_158 0 5.8567235176520110e-03
GC_5_159 b_5 NI_5 NS_159 0 -8.4251215129149537e-10
GC_5_160 b_5 NI_5 NS_160 0 -1.6876108882019738e-06
GC_5_161 b_5 NI_5 NS_161 0 2.5405881226810866e-04
GC_5_162 b_5 NI_5 NS_162 0 2.6638827778355592e-03
GC_5_163 b_5 NI_5 NS_163 0 4.5287651405927585e-03
GC_5_164 b_5 NI_5 NS_164 0 -2.7517441800721785e-03
GC_5_165 b_5 NI_5 NS_165 0 -5.4237649933211261e-03
GC_5_166 b_5 NI_5 NS_166 0 4.1627734726820920e-04
GC_5_167 b_5 NI_5 NS_167 0 8.8489949678563252e-03
GC_5_168 b_5 NI_5 NS_168 0 -6.0329856067813743e-04
GC_5_169 b_5 NI_5 NS_169 0 -2.8273784151117949e-03
GC_5_170 b_5 NI_5 NS_170 0 -2.3878794998851579e-03
GC_5_171 b_5 NI_5 NS_171 0 4.8268255975313299e-05
GC_5_172 b_5 NI_5 NS_172 0 -2.1045587677131824e-03
GC_5_173 b_5 NI_5 NS_173 0 -3.5071477919363559e-03
GC_5_174 b_5 NI_5 NS_174 0 5.5654796014008856e-03
GC_5_175 b_5 NI_5 NS_175 0 5.1183014482111908e-03
GC_5_176 b_5 NI_5 NS_176 0 -7.7286276105334980e-03
GC_5_177 b_5 NI_5 NS_177 0 -5.0253323951217335e-03
GC_5_178 b_5 NI_5 NS_178 0 3.1189362088843097e-03
GC_5_179 b_5 NI_5 NS_179 0 2.2497873906578364e-03
GC_5_180 b_5 NI_5 NS_180 0 -1.6595376233848728e-03
GC_5_181 b_5 NI_5 NS_181 0 -6.2720699667936303e-03
GC_5_182 b_5 NI_5 NS_182 0 3.8172623940376182e-03
GC_5_183 b_5 NI_5 NS_183 0 -1.3159048032284912e-03
GC_5_184 b_5 NI_5 NS_184 0 2.1722207299458012e-03
GC_5_185 b_5 NI_5 NS_185 0 7.7247492039753620e-10
GC_5_186 b_5 NI_5 NS_186 0 6.0126661879104851e-07
GC_5_187 b_5 NI_5 NS_187 0 -1.9612989217871986e-04
GC_5_188 b_5 NI_5 NS_188 0 -4.5795047464408249e-04
GC_5_189 b_5 NI_5 NS_189 0 -1.0663204084601916e-03
GC_5_190 b_5 NI_5 NS_190 0 -9.2689119069791698e-04
GC_5_191 b_5 NI_5 NS_191 0 -2.3216409846091679e-03
GC_5_192 b_5 NI_5 NS_192 0 3.0885303422369126e-04
GC_5_193 b_5 NI_5 NS_193 0 -3.5739848773951814e-04
GC_5_194 b_5 NI_5 NS_194 0 4.2021104394642092e-03
GC_5_195 b_5 NI_5 NS_195 0 9.8001058276248553e-04
GC_5_196 b_5 NI_5 NS_196 0 4.4275210728321793e-04
GC_5_197 b_5 NI_5 NS_197 0 -3.7449348107852808e-04
GC_5_198 b_5 NI_5 NS_198 0 7.7738857288901415e-05
GC_5_199 b_5 NI_5 NS_199 0 -3.1870783947904243e-04
GC_5_200 b_5 NI_5 NS_200 0 3.3550914906553134e-03
GC_5_201 b_5 NI_5 NS_201 0 5.2311011365012887e-03
GC_5_202 b_5 NI_5 NS_202 0 8.1047424476673980e-04
GC_5_203 b_5 NI_5 NS_203 0 1.3422336715926666e-03
GC_5_204 b_5 NI_5 NS_204 0 -1.9491672036624989e-03
GC_5_205 b_5 NI_5 NS_205 0 -8.8183379038938290e-04
GC_5_206 b_5 NI_5 NS_206 0 -6.4378730917925961e-04
GC_5_207 b_5 NI_5 NS_207 0 -1.3370800512422171e-03
GC_5_208 b_5 NI_5 NS_208 0 2.5847967361392467e-03
GC_5_209 b_5 NI_5 NS_209 0 3.8620814434733104e-04
GC_5_210 b_5 NI_5 NS_210 0 -2.0252878232734435e-03
GC_5_211 b_5 NI_5 NS_211 0 4.0260186355572215e-10
GC_5_212 b_5 NI_5 NS_212 0 -2.6893743813703713e-08
GC_5_213 b_5 NI_5 NS_213 0 1.8850642765433500e-05
GC_5_214 b_5 NI_5 NS_214 0 4.3631168231041981e-05
GC_5_215 b_5 NI_5 NS_215 0 8.2151685450270037e-05
GC_5_216 b_5 NI_5 NS_216 0 -3.0666300331728400e-05
GC_5_217 b_5 NI_5 NS_217 0 -1.3460177778958137e-05
GC_5_218 b_5 NI_5 NS_218 0 1.3808944579456746e-05
GC_5_219 b_5 NI_5 NS_219 0 1.9797123512973691e-04
GC_5_220 b_5 NI_5 NS_220 0 -9.9099563142820659e-05
GC_5_221 b_5 NI_5 NS_221 0 2.7210975527597455e-05
GC_5_222 b_5 NI_5 NS_222 0 -9.8085102442501985e-05
GC_5_223 b_5 NI_5 NS_223 0 -1.7289683397512035e-05
GC_5_224 b_5 NI_5 NS_224 0 -9.8313648943239212e-05
GC_5_225 b_5 NI_5 NS_225 0 1.0597728096093220e-05
GC_5_226 b_5 NI_5 NS_226 0 -9.7356896215138907e-05
GC_5_227 b_5 NI_5 NS_227 0 -9.7278143303828479e-05
GC_5_228 b_5 NI_5 NS_228 0 -3.1575652856578629e-04
GC_5_229 b_5 NI_5 NS_229 0 -1.3369272192936260e-04
GC_5_230 b_5 NI_5 NS_230 0 -1.1532242258339623e-04
GC_5_231 b_5 NI_5 NS_231 0 -1.9101665678708535e-05
GC_5_232 b_5 NI_5 NS_232 0 -1.9122446465119085e-04
GC_5_233 b_5 NI_5 NS_233 0 1.5286795436102152e-03
GC_5_234 b_5 NI_5 NS_234 0 -9.9338068026158684e-05
GC_5_235 b_5 NI_5 NS_235 0 1.2824482306885644e-04
GC_5_236 b_5 NI_5 NS_236 0 5.5586348136646450e-05
GC_5_237 b_5 NI_5 NS_237 0 -4.2209249755030364e-10
GC_5_238 b_5 NI_5 NS_238 0 4.4721732704204236e-08
GC_5_239 b_5 NI_5 NS_239 0 5.7604319562637968e-06
GC_5_240 b_5 NI_5 NS_240 0 7.6123947814389395e-05
GC_5_241 b_5 NI_5 NS_241 0 1.5376806714730313e-04
GC_5_242 b_5 NI_5 NS_242 0 1.3563431510885953e-04
GC_5_243 b_5 NI_5 NS_243 0 3.4707304590821884e-04
GC_5_244 b_5 NI_5 NS_244 0 -2.4008687633251271e-05
GC_5_245 b_5 NI_5 NS_245 0 5.3250621399498880e-05
GC_5_246 b_5 NI_5 NS_246 0 -5.8494565304011788e-04
GC_5_247 b_5 NI_5 NS_247 0 -1.4501223029903096e-04
GC_5_248 b_5 NI_5 NS_248 0 -6.8322989841542716e-05
GC_5_249 b_5 NI_5 NS_249 0 5.2206224592302893e-05
GC_5_250 b_5 NI_5 NS_250 0 -1.0707672343166772e-05
GC_5_251 b_5 NI_5 NS_251 0 4.8324650363863878e-05
GC_5_252 b_5 NI_5 NS_252 0 -4.5206767776138299e-04
GC_5_253 b_5 NI_5 NS_253 0 -7.0671503590279106e-04
GC_5_254 b_5 NI_5 NS_254 0 -8.3345688590489284e-05
GC_5_255 b_5 NI_5 NS_255 0 -1.7415344927532828e-04
GC_5_256 b_5 NI_5 NS_256 0 2.5972212781021347e-04
GC_5_257 b_5 NI_5 NS_257 0 1.0227107636011362e-04
GC_5_258 b_5 NI_5 NS_258 0 8.1142078855284841e-05
GC_5_259 b_5 NI_5 NS_259 0 -1.2306561458993906e-04
GC_5_260 b_5 NI_5 NS_260 0 -3.3447033409318027e-04
GC_5_261 b_5 NI_5 NS_261 0 -1.4271473645287945e-04
GC_5_262 b_5 NI_5 NS_262 0 6.6398827996723593e-04
GC_5_263 b_5 NI_5 NS_263 0 1.2463229585532024e-10
GC_5_264 b_5 NI_5 NS_264 0 -1.1464989794897443e-08
GC_5_265 b_5 NI_5 NS_265 0 -4.0098324486847746e-06
GC_5_266 b_5 NI_5 NS_266 0 -3.9985351622961009e-06
GC_5_267 b_5 NI_5 NS_267 0 -9.6089759356155400e-06
GC_5_268 b_5 NI_5 NS_268 0 -3.7333276638023070e-06
GC_5_269 b_5 NI_5 NS_269 0 -1.8752441301156251e-05
GC_5_270 b_5 NI_5 NS_270 0 -1.5170146370238504e-06
GC_5_271 b_5 NI_5 NS_271 0 -2.9293434693476312e-05
GC_5_272 b_5 NI_5 NS_272 0 2.7695969803338952e-05
GC_5_273 b_5 NI_5 NS_273 0 -2.1495343541213936e-05
GC_5_274 b_5 NI_5 NS_274 0 2.3548508581561971e-05
GC_5_275 b_5 NI_5 NS_275 0 6.0794688673387181e-06
GC_5_276 b_5 NI_5 NS_276 0 2.3428414745216090e-05
GC_5_277 b_5 NI_5 NS_277 0 -1.5898351460727427e-05
GC_5_278 b_5 NI_5 NS_278 0 5.5619624334109508e-05
GC_5_279 b_5 NI_5 NS_279 0 5.4333376425170029e-05
GC_5_280 b_5 NI_5 NS_280 0 6.5658593039493951e-05
GC_5_281 b_5 NI_5 NS_281 0 2.2574648483868615e-05
GC_5_282 b_5 NI_5 NS_282 0 4.5652058038796665e-05
GC_5_283 b_5 NI_5 NS_283 0 1.4988655919955863e-05
GC_5_284 b_5 NI_5 NS_284 0 4.9568130607333322e-05
GC_5_285 b_5 NI_5 NS_285 0 -5.1674629761129553e-04
GC_5_286 b_5 NI_5 NS_286 0 2.4176486422227245e-05
GC_5_287 b_5 NI_5 NS_287 0 -1.7525454302717305e-05
GC_5_288 b_5 NI_5 NS_288 0 -2.5351705720961186e-04
GC_5_289 b_5 NI_5 NS_289 0 -1.0840951270630802e-10
GC_5_290 b_5 NI_5 NS_290 0 4.8101624129240496e-09
GC_5_291 b_5 NI_5 NS_291 0 5.0649840488125913e-06
GC_5_292 b_5 NI_5 NS_292 0 9.6682506636548561e-06
GC_5_293 b_5 NI_5 NS_293 0 1.6493793564062969e-05
GC_5_294 b_5 NI_5 NS_294 0 1.3404317820306904e-05
GC_5_295 b_5 NI_5 NS_295 0 3.8423175084940796e-05
GC_5_296 b_5 NI_5 NS_296 0 -3.4230206775914035e-06
GC_5_297 b_5 NI_5 NS_297 0 1.4655240385743540e-05
GC_5_298 b_5 NI_5 NS_298 0 -6.2678549799526448e-05
GC_5_299 b_5 NI_5 NS_299 0 -1.1682861386834360e-05
GC_5_300 b_5 NI_5 NS_300 0 -9.0308616475710930e-06
GC_5_301 b_5 NI_5 NS_301 0 4.7729739212910418e-06
GC_5_302 b_5 NI_5 NS_302 0 -3.5003845247526719e-06
GC_5_303 b_5 NI_5 NS_303 0 9.7656286939428857e-06
GC_5_304 b_5 NI_5 NS_304 0 -4.9987526921034184e-05
GC_5_305 b_5 NI_5 NS_305 0 -6.6158996259598052e-05
GC_5_306 b_5 NI_5 NS_306 0 -2.1604507498575765e-05
GC_5_307 b_5 NI_5 NS_307 0 -1.6750712796528477e-05
GC_5_308 b_5 NI_5 NS_308 0 1.9351803528070888e-05
GC_5_309 b_5 NI_5 NS_309 0 1.6103498710328603e-05
GC_5_310 b_5 NI_5 NS_310 0 -1.2511215110176941e-06
GC_5_311 b_5 NI_5 NS_311 0 2.1545969180508743e-04
GC_5_312 b_5 NI_5 NS_312 0 7.2320056652959500e-06
GD_5_1 b_5 NI_5 NA_1 0 1.6315392052185300e-04
GD_5_2 b_5 NI_5 NA_2 0 1.3323647119903653e-04
GD_5_3 b_5 NI_5 NA_3 0 3.0059891770121056e-03
GD_5_4 b_5 NI_5 NA_4 0 -5.3669732937386012e-05
GD_5_5 b_5 NI_5 NA_5 0 -2.9682552450643926e-02
GD_5_6 b_5 NI_5 NA_6 0 -2.0430178913138922e-02
GD_5_7 b_5 NI_5 NA_7 0 1.3447778880549956e-02
GD_5_8 b_5 NI_5 NA_8 0 -1.1284130958466509e-03
GD_5_9 b_5 NI_5 NA_9 0 1.6640052713515682e-04
GD_5_10 b_5 NI_5 NA_10 0 1.4009478178153364e-04
GD_5_11 b_5 NI_5 NA_11 0 5.6434017117627705e-07
GD_5_12 b_5 NI_5 NA_12 0 3.5144870028929442e-05
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 1.5157434031294110e-04
GC_6_2 b_6 NI_6 NS_2 0 1.2809807721790264e-05
GC_6_3 b_6 NI_6 NS_3 0 -4.2742665402475290e-10
GC_6_4 b_6 NI_6 NS_4 0 4.5130301353889023e-08
GC_6_5 b_6 NI_6 NS_5 0 5.1596762151418862e-06
GC_6_6 b_6 NI_6 NS_6 0 7.5616107998997050e-05
GC_6_7 b_6 NI_6 NS_7 0 1.5335221855013498e-04
GC_6_8 b_6 NI_6 NS_8 0 1.3548710716536545e-04
GC_6_9 b_6 NI_6 NS_9 0 3.4656072090659049e-04
GC_6_10 b_6 NI_6 NS_10 0 -2.4741108396141590e-05
GC_6_11 b_6 NI_6 NS_11 0 5.1570183439346215e-05
GC_6_12 b_6 NI_6 NS_12 0 -5.8538715235579642e-04
GC_6_13 b_6 NI_6 NS_13 0 -1.4593519007921206e-04
GC_6_14 b_6 NI_6 NS_14 0 -6.8386950673637745e-05
GC_6_15 b_6 NI_6 NS_15 0 5.1713283850788880e-05
GC_6_16 b_6 NI_6 NS_16 0 -1.0507847524648707e-05
GC_6_17 b_6 NI_6 NS_17 0 4.7730213934262387e-05
GC_6_18 b_6 NI_6 NS_18 0 -4.5313042713358164e-04
GC_6_19 b_6 NI_6 NS_19 0 -7.0918794637193948e-04
GC_6_20 b_6 NI_6 NS_20 0 -8.3323699330682910e-05
GC_6_21 b_6 NI_6 NS_21 0 -1.7472346305612188e-04
GC_6_22 b_6 NI_6 NS_22 0 2.5870651847223789e-04
GC_6_23 b_6 NI_6 NS_23 0 1.0249954168076233e-04
GC_6_24 b_6 NI_6 NS_24 0 7.9812165480014363e-05
GC_6_25 b_6 NI_6 NS_25 0 -8.6761638088865090e-05
GC_6_26 b_6 NI_6 NS_26 0 -3.2996766228861161e-04
GC_6_27 b_6 NI_6 NS_27 0 3.9579047094818012e-04
GC_6_28 b_6 NI_6 NS_28 0 -2.0177620441232521e-03
GC_6_29 b_6 NI_6 NS_29 0 4.0760489902501630e-10
GC_6_30 b_6 NI_6 NS_30 0 -2.7072352132898621e-08
GC_6_31 b_6 NI_6 NS_31 0 1.8516035402822967e-05
GC_6_32 b_6 NI_6 NS_32 0 4.3377996176531647e-05
GC_6_33 b_6 NI_6 NS_33 0 8.1709677196281161e-05
GC_6_34 b_6 NI_6 NS_34 0 -3.0786352502017423e-05
GC_6_35 b_6 NI_6 NS_35 0 -1.3938884324080366e-05
GC_6_36 b_6 NI_6 NS_36 0 1.3650823813618939e-05
GC_6_37 b_6 NI_6 NS_37 0 1.9708922241116954e-04
GC_6_38 b_6 NI_6 NS_38 0 -9.8902008739698563e-05
GC_6_39 b_6 NI_6 NS_39 0 2.6744128190183247e-05
GC_6_40 b_6 NI_6 NS_40 0 -9.8059736673188479e-05
GC_6_41 b_6 NI_6 NS_41 0 -1.7490356676107947e-05
GC_6_42 b_6 NI_6 NS_42 0 -9.8091727016159534e-05
GC_6_43 b_6 NI_6 NS_43 0 9.8222349470372809e-06
GC_6_44 b_6 NI_6 NS_44 0 -9.7469479017807406e-05
GC_6_45 b_6 NI_6 NS_45 0 -9.8112201951225381e-05
GC_6_46 b_6 NI_6 NS_46 0 -3.1491541495352963e-04
GC_6_47 b_6 NI_6 NS_47 0 -1.3398287937104307e-04
GC_6_48 b_6 NI_6 NS_48 0 -1.1516245593084510e-04
GC_6_49 b_6 NI_6 NS_49 0 -1.9658470699634692e-05
GC_6_50 b_6 NI_6 NS_50 0 -1.9129802544966940e-04
GC_6_51 b_6 NI_6 NS_51 0 1.5212419508357064e-03
GC_6_52 b_6 NI_6 NS_52 0 -1.0185248702054264e-04
GC_6_53 b_6 NI_6 NS_53 0 -1.0993209279456827e-03
GC_6_54 b_6 NI_6 NS_54 0 1.9264488602822526e-03
GC_6_55 b_6 NI_6 NS_55 0 -9.9960372328513066e-11
GC_6_56 b_6 NI_6 NS_56 0 2.7260538808841335e-07
GC_6_57 b_6 NI_6 NS_57 0 5.8933463610379077e-05
GC_6_58 b_6 NI_6 NS_58 0 -8.7080058339564096e-05
GC_6_59 b_6 NI_6 NS_59 0 -2.6160836006459346e-04
GC_6_60 b_6 NI_6 NS_60 0 -1.7078573490407188e-04
GC_6_61 b_6 NI_6 NS_61 0 -5.2946919279402149e-04
GC_6_62 b_6 NI_6 NS_62 0 2.5259348307462496e-05
GC_6_63 b_6 NI_6 NS_63 0 4.2452468201349448e-05
GC_6_64 b_6 NI_6 NS_64 0 9.1569635414498745e-04
GC_6_65 b_6 NI_6 NS_65 0 2.4558828711875773e-04
GC_6_66 b_6 NI_6 NS_66 0 1.3071939753188204e-04
GC_6_67 b_6 NI_6 NS_67 0 -8.1498481741995373e-05
GC_6_68 b_6 NI_6 NS_68 0 2.6844114795914232e-05
GC_6_69 b_6 NI_6 NS_69 0 -7.0951258499657083e-05
GC_6_70 b_6 NI_6 NS_70 0 7.5354268323844429e-04
GC_6_71 b_6 NI_6 NS_71 0 1.2758086626034595e-03
GC_6_72 b_6 NI_6 NS_72 0 1.3799804198716902e-04
GC_6_73 b_6 NI_6 NS_73 0 3.2406020988702441e-04
GC_6_74 b_6 NI_6 NS_74 0 -4.2268318030886021e-04
GC_6_75 b_6 NI_6 NS_75 0 -2.4533855461694498e-04
GC_6_76 b_6 NI_6 NS_76 0 -1.0928505623243643e-04
GC_6_77 b_6 NI_6 NS_77 0 -1.5485139655560373e-03
GC_6_78 b_6 NI_6 NS_78 0 3.7255016722565881e-04
GC_6_79 b_6 NI_6 NS_79 0 -1.2120664070484606e-03
GC_6_80 b_6 NI_6 NS_80 0 5.5288358058765304e-04
GC_6_81 b_6 NI_6 NS_81 0 3.0006673123479246e-10
GC_6_82 b_6 NI_6 NS_82 0 -5.7499733148222036e-07
GC_6_83 b_6 NI_6 NS_83 0 3.1147145751544431e-05
GC_6_84 b_6 NI_6 NS_84 0 6.3814449665242719e-04
GC_6_85 b_6 NI_6 NS_85 0 1.0887928365402900e-03
GC_6_86 b_6 NI_6 NS_86 0 -6.7568193631959350e-04
GC_6_87 b_6 NI_6 NS_87 0 -1.3741747929434428e-03
GC_6_88 b_6 NI_6 NS_88 0 7.5250724066521814e-05
GC_6_89 b_6 NI_6 NS_89 0 2.0942417570502013e-03
GC_6_90 b_6 NI_6 NS_90 0 -1.0656274188195585e-04
GC_6_91 b_6 NI_6 NS_91 0 -7.3383166448999797e-04
GC_6_92 b_6 NI_6 NS_92 0 -5.7289836410679242e-04
GC_6_93 b_6 NI_6 NS_93 0 5.7537680211187741e-06
GC_6_94 b_6 NI_6 NS_94 0 -4.8778998313019778e-04
GC_6_95 b_6 NI_6 NS_95 0 -9.0586723004564104e-04
GC_6_96 b_6 NI_6 NS_96 0 1.3910544878334402e-03
GC_6_97 b_6 NI_6 NS_97 0 1.2473495838130019e-03
GC_6_98 b_6 NI_6 NS_98 0 -1.8369134090307835e-03
GC_6_99 b_6 NI_6 NS_99 0 -1.2248408683873033e-03
GC_6_100 b_6 NI_6 NS_100 0 7.8178232261206571e-04
GC_6_101 b_6 NI_6 NS_101 0 5.7543582813650448e-04
GC_6_102 b_6 NI_6 NS_102 0 -4.1190529759865287e-04
GC_6_103 b_6 NI_6 NS_103 0 -7.3187165943608531e-04
GC_6_104 b_6 NI_6 NS_104 0 1.1403197669149487e-03
GC_6_105 b_6 NI_6 NS_105 0 -4.9912546863792144e-02
GC_6_106 b_6 NI_6 NS_106 0 1.0946193887043948e-01
GC_6_107 b_6 NI_6 NS_107 0 1.0782683154866814e-08
GC_6_108 b_6 NI_6 NS_108 0 1.9879858069175796e-05
GC_6_109 b_6 NI_6 NS_109 0 -1.5753191826808798e-02
GC_6_110 b_6 NI_6 NS_110 0 2.4251006273635318e-02
GC_6_111 b_6 NI_6 NS_111 0 -7.8027682414024430e-03
GC_6_112 b_6 NI_6 NS_112 0 -1.4488574680566796e-02
GC_6_113 b_6 NI_6 NS_113 0 2.0433212336492396e-02
GC_6_114 b_6 NI_6 NS_114 0 6.6873557365669392e-03
GC_6_115 b_6 NI_6 NS_115 0 8.0583305635608064e-03
GC_6_116 b_6 NI_6 NS_116 0 4.3992667030562600e-02
GC_6_117 b_6 NI_6 NS_117 0 -1.1853721549012219e-02
GC_6_118 b_6 NI_6 NS_118 0 -3.2338876291069085e-03
GC_6_119 b_6 NI_6 NS_119 0 -5.0942089297391965e-03
GC_6_120 b_6 NI_6 NS_120 0 -4.0938822611839634e-03
GC_6_121 b_6 NI_6 NS_121 0 2.6816832856513109e-02
GC_6_122 b_6 NI_6 NS_122 0 -8.8227355233235298e-06
GC_6_123 b_6 NI_6 NS_123 0 3.3872762160008819e-02
GC_6_124 b_6 NI_6 NS_124 0 3.0990204682648199e-02
GC_6_125 b_6 NI_6 NS_125 0 -1.5640926444160309e-02
GC_6_126 b_6 NI_6 NS_126 0 8.2834126754453025e-03
GC_6_127 b_6 NI_6 NS_127 0 -9.9439865912615043e-04
GC_6_128 b_6 NI_6 NS_128 0 -6.8670025706375889e-03
GC_6_129 b_6 NI_6 NS_129 0 -6.8769692222333353e-02
GC_6_130 b_6 NI_6 NS_130 0 1.7777710403328218e-03
GC_6_131 b_6 NI_6 NS_131 0 5.9215489962724771e-02
GC_6_132 b_6 NI_6 NS_132 0 -6.3407636300857301e-02
GC_6_133 b_6 NI_6 NS_133 0 -1.0211750104088715e-08
GC_6_134 b_6 NI_6 NS_134 0 -8.2108571934109800e-06
GC_6_135 b_6 NI_6 NS_135 0 -1.8466567588426841e-03
GC_6_136 b_6 NI_6 NS_136 0 -2.8683123701404843e-03
GC_6_137 b_6 NI_6 NS_137 0 -5.1018049687674861e-03
GC_6_138 b_6 NI_6 NS_138 0 1.9432405042730508e-03
GC_6_139 b_6 NI_6 NS_139 0 2.4539731021212346e-03
GC_6_140 b_6 NI_6 NS_140 0 -1.2214745377999367e-03
GC_6_141 b_6 NI_6 NS_141 0 -1.0637008586728593e-02
GC_6_142 b_6 NI_6 NS_142 0 1.1057795139107721e-03
GC_6_143 b_6 NI_6 NS_143 0 6.4906104355947475e-04
GC_6_144 b_6 NI_6 NS_144 0 1.7568055400822690e-03
GC_6_145 b_6 NI_6 NS_145 0 -9.5190922325557442e-04
GC_6_146 b_6 NI_6 NS_146 0 2.2857457167483656e-03
GC_6_147 b_6 NI_6 NS_147 0 6.0496281193836714e-04
GC_6_148 b_6 NI_6 NS_148 0 -5.8869625838110810e-03
GC_6_149 b_6 NI_6 NS_149 0 -8.5212789070572906e-03
GC_6_150 b_6 NI_6 NS_150 0 6.8916057982835047e-03
GC_6_151 b_6 NI_6 NS_151 0 2.5250257717987557e-03
GC_6_152 b_6 NI_6 NS_152 0 -3.6699130634487106e-03
GC_6_153 b_6 NI_6 NS_153 0 -2.6398888960123251e-03
GC_6_154 b_6 NI_6 NS_154 0 -5.0014762094001668e-04
GC_6_155 b_6 NI_6 NS_155 0 5.4262590367559024e-02
GC_6_156 b_6 NI_6 NS_156 0 1.5891713896910914e-03
GC_6_157 b_6 NI_6 NS_157 0 -1.3158639643578573e-03
GC_6_158 b_6 NI_6 NS_158 0 2.1722220842503208e-03
GC_6_159 b_6 NI_6 NS_159 0 7.7247550756717771e-10
GC_6_160 b_6 NI_6 NS_160 0 6.0126670905628429e-07
GC_6_161 b_6 NI_6 NS_161 0 -1.9612813500747295e-04
GC_6_162 b_6 NI_6 NS_162 0 -4.5793429396958778e-04
GC_6_163 b_6 NI_6 NS_163 0 -1.0663224132107358e-03
GC_6_164 b_6 NI_6 NS_164 0 -9.2690698893680096e-04
GC_6_165 b_6 NI_6 NS_165 0 -2.3216377405190108e-03
GC_6_166 b_6 NI_6 NS_166 0 3.0883884497085666e-04
GC_6_167 b_6 NI_6 NS_167 0 -3.5741414742638411e-04
GC_6_168 b_6 NI_6 NS_168 0 4.2021284042135735e-03
GC_6_169 b_6 NI_6 NS_169 0 9.8000801436476576e-04
GC_6_170 b_6 NI_6 NS_170 0 4.4275717495589531e-04
GC_6_171 b_6 NI_6 NS_171 0 -3.7449557410897978e-04
GC_6_172 b_6 NI_6 NS_172 0 7.7736282895278250e-05
GC_6_173 b_6 NI_6 NS_173 0 -3.1871488331706966e-04
GC_6_174 b_6 NI_6 NS_174 0 3.3550933326881435e-03
GC_6_175 b_6 NI_6 NS_175 0 5.2311075295818328e-03
GC_6_176 b_6 NI_6 NS_176 0 8.1049137193250442e-04
GC_6_177 b_6 NI_6 NS_177 0 1.3422387448348693e-03
GC_6_178 b_6 NI_6 NS_178 0 -1.9491659262996321e-03
GC_6_179 b_6 NI_6 NS_179 0 -8.8183193801034054e-04
GC_6_180 b_6 NI_6 NS_180 0 -6.4378956060342162e-04
GC_6_181 b_6 NI_6 NS_181 0 -1.3370813001153188e-03
GC_6_182 b_6 NI_6 NS_182 0 2.5847959779491843e-03
GC_6_183 b_6 NI_6 NS_183 0 -7.6472777598518048e-03
GC_6_184 b_6 NI_6 NS_184 0 5.8567239269299055e-03
GC_6_185 b_6 NI_6 NS_185 0 -8.4251219674268920e-10
GC_6_186 b_6 NI_6 NS_186 0 -1.6876108431264379e-06
GC_6_187 b_6 NI_6 NS_187 0 2.5405881628339015e-04
GC_6_188 b_6 NI_6 NS_188 0 2.6638827817409977e-03
GC_6_189 b_6 NI_6 NS_189 0 4.5287651879800618e-03
GC_6_190 b_6 NI_6 NS_190 0 -2.7517441758933424e-03
GC_6_191 b_6 NI_6 NS_191 0 -5.4237649446824462e-03
GC_6_192 b_6 NI_6 NS_192 0 4.1627728340774036e-04
GC_6_193 b_6 NI_6 NS_193 0 8.8489949382731820e-03
GC_6_194 b_6 NI_6 NS_194 0 -6.0329864409836671e-04
GC_6_195 b_6 NI_6 NS_195 0 -2.8273784113507332e-03
GC_6_196 b_6 NI_6 NS_196 0 -2.3878795498347913e-03
GC_6_197 b_6 NI_6 NS_197 0 4.8268229086503788e-05
GC_6_198 b_6 NI_6 NS_198 0 -2.1045587978107171e-03
GC_6_199 b_6 NI_6 NS_199 0 -3.5071478368893872e-03
GC_6_200 b_6 NI_6 NS_200 0 5.5654795023737701e-03
GC_6_201 b_6 NI_6 NS_201 0 5.1183013216546521e-03
GC_6_202 b_6 NI_6 NS_202 0 -7.7286276384112562e-03
GC_6_203 b_6 NI_6 NS_203 0 -5.0253324617630614e-03
GC_6_204 b_6 NI_6 NS_204 0 3.1189361712689627e-03
GC_6_205 b_6 NI_6 NS_205 0 2.2497873076311827e-03
GC_6_206 b_6 NI_6 NS_206 0 -1.6595376517622323e-03
GC_6_207 b_6 NI_6 NS_207 0 -6.2720704311510275e-03
GC_6_208 b_6 NI_6 NS_208 0 3.8172621860017913e-03
GC_6_209 b_6 NI_6 NS_209 0 1.2824311394141427e-04
GC_6_210 b_6 NI_6 NS_210 0 5.5587841082956335e-05
GC_6_211 b_6 NI_6 NS_211 0 -4.2209257114574173e-10
GC_6_212 b_6 NI_6 NS_212 0 4.4721715132282386e-08
GC_6_213 b_6 NI_6 NS_213 0 5.7603063039913100e-06
GC_6_214 b_6 NI_6 NS_214 0 7.6124133486296376e-05
GC_6_215 b_6 NI_6 NS_215 0 1.5376831906569748e-04
GC_6_216 b_6 NI_6 NS_216 0 1.3563455001290006e-04
GC_6_217 b_6 NI_6 NS_217 0 3.4707338916729582e-04
GC_6_218 b_6 NI_6 NS_218 0 -2.4008417429795056e-05
GC_6_219 b_6 NI_6 NS_219 0 5.3250879351751137e-05
GC_6_220 b_6 NI_6 NS_220 0 -5.8494622635987044e-04
GC_6_221 b_6 NI_6 NS_221 0 -1.4501227652516174e-04
GC_6_222 b_6 NI_6 NS_222 0 -6.8323073059257215e-05
GC_6_223 b_6 NI_6 NS_223 0 5.2206312738218990e-05
GC_6_224 b_6 NI_6 NS_224 0 -1.0707557948624030e-05
GC_6_225 b_6 NI_6 NS_225 0 4.8324829232930010e-05
GC_6_226 b_6 NI_6 NS_226 0 -4.5206759624715929e-04
GC_6_227 b_6 NI_6 NS_227 0 -7.0671486047070217e-04
GC_6_228 b_6 NI_6 NS_228 0 -8.3346071387218265e-05
GC_6_229 b_6 NI_6 NS_229 0 -1.7415349044114033e-04
GC_6_230 b_6 NI_6 NS_230 0 2.5972205185926042e-04
GC_6_231 b_6 NI_6 NS_231 0 1.0227100313805719e-04
GC_6_232 b_6 NI_6 NS_232 0 8.1142071246262094e-05
GC_6_233 b_6 NI_6 NS_233 0 -1.2306695903762502e-04
GC_6_234 b_6 NI_6 NS_234 0 -3.3447060399634156e-04
GC_6_235 b_6 NI_6 NS_235 0 3.8512279777697876e-04
GC_6_236 b_6 NI_6 NS_236 0 -2.0245853368198903e-03
GC_6_237 b_6 NI_6 NS_237 0 4.0264790320202008e-10
GC_6_238 b_6 NI_6 NS_238 0 -2.6912814438385387e-08
GC_6_239 b_6 NI_6 NS_239 0 1.8964557414198234e-05
GC_6_240 b_6 NI_6 NS_240 0 4.3646769281857876e-05
GC_6_241 b_6 NI_6 NS_241 0 8.2121180927012544e-05
GC_6_242 b_6 NI_6 NS_242 0 -3.0735340110135757e-05
GC_6_243 b_6 NI_6 NS_243 0 -1.3364254676164405e-05
GC_6_244 b_6 NI_6 NS_244 0 1.3940739760461222e-05
GC_6_245 b_6 NI_6 NS_245 0 1.9803504369048517e-04
GC_6_246 b_6 NI_6 NS_246 0 -9.9273347596798251e-05
GC_6_247 b_6 NI_6 NS_247 0 2.7239745476864380e-05
GC_6_248 b_6 NI_6 NS_248 0 -9.8033292470488815e-05
GC_6_249 b_6 NI_6 NS_249 0 -1.7295797825711810e-05
GC_6_250 b_6 NI_6 NS_250 0 -9.8327848341321517e-05
GC_6_251 b_6 NI_6 NS_251 0 1.0740655651299258e-05
GC_6_252 b_6 NI_6 NS_252 0 -9.7316253665893603e-05
GC_6_253 b_6 NI_6 NS_253 0 -9.7269565161823217e-05
GC_6_254 b_6 NI_6 NS_254 0 -3.1582661462218090e-04
GC_6_255 b_6 NI_6 NS_255 0 -1.3361352247895879e-04
GC_6_256 b_6 NI_6 NS_256 0 -1.1528990621764768e-04
GC_6_257 b_6 NI_6 NS_257 0 -1.9094748617127504e-05
GC_6_258 b_6 NI_6 NS_258 0 -1.9121733296413720e-04
GC_6_259 b_6 NI_6 NS_259 0 1.5281239975381150e-03
GC_6_260 b_6 NI_6 NS_260 0 -9.9340182694242365e-05
GC_6_261 b_6 NI_6 NS_261 0 -1.7314431751576996e-05
GC_6_262 b_6 NI_6 NS_262 0 -2.5362085792600988e-04
GC_6_263 b_6 NI_6 NS_263 0 -1.0841168062052938e-10
GC_6_264 b_6 NI_6 NS_264 0 4.8114852621272048e-09
GC_6_265 b_6 NI_6 NS_265 0 5.0737559788472487e-06
GC_6_266 b_6 NI_6 NS_266 0 9.7330064481711001e-06
GC_6_267 b_6 NI_6 NS_267 0 1.6486990394528898e-05
GC_6_268 b_6 NI_6 NS_268 0 1.3338260819662094e-05
GC_6_269 b_6 NI_6 NS_269 0 3.8439306943016742e-05
GC_6_270 b_6 NI_6 NS_270 0 -3.4839413254294801e-06
GC_6_271 b_6 NI_6 NS_271 0 1.4588787649207907e-05
GC_6_272 b_6 NI_6 NS_272 0 -6.2615390995567719e-05
GC_6_273 b_6 NI_6 NS_273 0 -1.1696091761869410e-05
GC_6_274 b_6 NI_6 NS_274 0 -9.0145924823973183e-06
GC_6_275 b_6 NI_6 NS_275 0 4.7616308790345091e-06
GC_6_276 b_6 NI_6 NS_276 0 -3.5113517564930895e-06
GC_6_277 b_6 NI_6 NS_277 0 9.7343948044611219e-06
GC_6_278 b_6 NI_6 NS_278 0 -4.9987537153408024e-05
GC_6_279 b_6 NI_6 NS_279 0 -6.6144971472922298e-05
GC_6_280 b_6 NI_6 NS_280 0 -2.1538293524517717e-05
GC_6_281 b_6 NI_6 NS_281 0 -1.6734573111957356e-05
GC_6_282 b_6 NI_6 NS_282 0 1.9354403787013914e-05
GC_6_283 b_6 NI_6 NS_283 0 1.6110181987210749e-05
GC_6_284 b_6 NI_6 NS_284 0 -1.2647831865924396e-06
GC_6_285 b_6 NI_6 NS_285 0 2.1554434729260661e-04
GC_6_286 b_6 NI_6 NS_286 0 7.2353968812132916e-06
GC_6_287 b_6 NI_6 NS_287 0 -1.4269275397553645e-04
GC_6_288 b_6 NI_6 NS_288 0 6.6397302122472976e-04
GC_6_289 b_6 NI_6 NS_289 0 1.2463082438824942e-10
GC_6_290 b_6 NI_6 NS_290 0 -1.1464438557577187e-08
GC_6_291 b_6 NI_6 NS_291 0 -4.0106801564010904e-06
GC_6_292 b_6 NI_6 NS_292 0 -3.9979564403153309e-06
GC_6_293 b_6 NI_6 NS_293 0 -9.6094390300754869e-06
GC_6_294 b_6 NI_6 NS_294 0 -3.7334837008931137e-06
GC_6_295 b_6 NI_6 NS_295 0 -1.8753686054914598e-05
GC_6_296 b_6 NI_6 NS_296 0 -1.5161594207862936e-06
GC_6_297 b_6 NI_6 NS_297 0 -2.9293756257726810e-05
GC_6_298 b_6 NI_6 NS_298 0 2.7696087662670570e-05
GC_6_299 b_6 NI_6 NS_299 0 -2.1496390417925533e-05
GC_6_300 b_6 NI_6 NS_300 0 2.3548923295515979e-05
GC_6_301 b_6 NI_6 NS_301 0 6.0790762442166064e-06
GC_6_302 b_6 NI_6 NS_302 0 2.3428696215242751e-05
GC_6_303 b_6 NI_6 NS_303 0 -1.5899459151453798e-05
GC_6_304 b_6 NI_6 NS_304 0 5.5620861786215712e-05
GC_6_305 b_6 NI_6 NS_305 0 5.4333653054705104e-05
GC_6_306 b_6 NI_6 NS_306 0 6.5659238849733980e-05
GC_6_307 b_6 NI_6 NS_307 0 2.2574534151218602e-05
GC_6_308 b_6 NI_6 NS_308 0 4.5651720352407810e-05
GC_6_309 b_6 NI_6 NS_309 0 1.4988559502574870e-05
GC_6_310 b_6 NI_6 NS_310 0 4.9567425854880780e-05
GC_6_311 b_6 NI_6 NS_311 0 -5.1673363762118330e-04
GC_6_312 b_6 NI_6 NS_312 0 2.4177847931116264e-05
GD_6_1 b_6 NI_6 NA_1 0 1.3324649184630303e-04
GD_6_2 b_6 NI_6 NA_2 0 1.6311756150690884e-04
GD_6_3 b_6 NI_6 NA_3 0 -5.3604006295013688e-05
GD_6_4 b_6 NI_6 NA_4 0 3.0059662968141233e-03
GD_6_5 b_6 NI_6 NA_5 0 -2.0430180464526975e-02
GD_6_6 b_6 NI_6 NA_6 0 -2.9682552450643988e-02
GD_6_7 b_6 NI_6 NA_7 0 -1.1284369305508274e-03
GD_6_8 b_6 NI_6 NA_8 0 1.3447779025221051e-02
GD_6_9 b_6 NI_6 NA_9 0 1.4009512861829632e-04
GD_6_10 b_6 NI_6 NA_10 0 1.6641036580786558e-04
GD_6_11 b_6 NI_6 NA_11 0 3.5049212710817529e-05
GD_6_12 b_6 NI_6 NA_12 0 5.5021198772757272e-07
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 -1.4358277110201553e-04
GC_7_2 b_7 NI_7 NS_2 0 6.6681872828090781e-04
GC_7_3 b_7 NI_7 NS_3 0 1.2440178283328307e-10
GC_7_4 b_7 NI_7 NS_4 0 -1.1384667119624718e-08
GC_7_5 b_7 NI_7 NS_5 0 -4.0163430042962893e-06
GC_7_6 b_7 NI_7 NS_6 0 -3.9922643762725221e-06
GC_7_7 b_7 NI_7 NS_7 0 -9.5849406527026045e-06
GC_7_8 b_7 NI_7 NS_8 0 -3.6873690727635584e-06
GC_7_9 b_7 NI_7 NS_9 0 -1.8730175754591587e-05
GC_7_10 b_7 NI_7 NS_10 0 -1.5350584180591134e-06
GC_7_11 b_7 NI_7 NS_11 0 -2.9271138580354818e-05
GC_7_12 b_7 NI_7 NS_12 0 2.7762606522213624e-05
GC_7_13 b_7 NI_7 NS_13 0 -2.1466916807246698e-05
GC_7_14 b_7 NI_7 NS_14 0 2.3556306258608005e-05
GC_7_15 b_7 NI_7 NS_15 0 6.1046516259146977e-06
GC_7_16 b_7 NI_7 NS_16 0 2.3438810170057101e-05
GC_7_17 b_7 NI_7 NS_17 0 -1.5894478397270282e-05
GC_7_18 b_7 NI_7 NS_18 0 5.5645649505206454e-05
GC_7_19 b_7 NI_7 NS_19 0 5.4416753461782856e-05
GC_7_20 b_7 NI_7 NS_20 0 6.5745047860699590e-05
GC_7_21 b_7 NI_7 NS_21 0 2.2593814480823682e-05
GC_7_22 b_7 NI_7 NS_22 0 4.5702050038966620e-05
GC_7_23 b_7 NI_7 NS_23 0 1.4942180562961764e-05
GC_7_24 b_7 NI_7 NS_24 0 4.9676808271689084e-05
GC_7_25 b_7 NI_7 NS_25 0 -5.1915999164438666e-04
GC_7_26 b_7 NI_7 NS_26 0 2.3889065164902189e-05
GC_7_27 b_7 NI_7 NS_27 0 -1.6380544945699784e-05
GC_7_28 b_7 NI_7 NS_28 0 -2.5702749152125138e-04
GC_7_29 b_7 NI_7 NS_29 0 -1.0826082725884329e-10
GC_7_30 b_7 NI_7 NS_30 0 4.7604533602204582e-09
GC_7_31 b_7 NI_7 NS_31 0 5.0802163689597004e-06
GC_7_32 b_7 NI_7 NS_32 0 9.6641027957594155e-06
GC_7_33 b_7 NI_7 NS_33 0 1.6473271735193750e-05
GC_7_34 b_7 NI_7 NS_34 0 1.3380149159107653e-05
GC_7_35 b_7 NI_7 NS_35 0 3.8420504286303967e-05
GC_7_36 b_7 NI_7 NS_36 0 -3.4928781790882534e-06
GC_7_37 b_7 NI_7 NS_37 0 1.4578073426117889e-05
GC_7_38 b_7 NI_7 NS_38 0 -6.2742694805009862e-05
GC_7_39 b_7 NI_7 NS_39 0 -1.1726885375707036e-05
GC_7_40 b_7 NI_7 NS_40 0 -9.0423435090529887e-06
GC_7_41 b_7 NI_7 NS_41 0 4.7447311947537729e-06
GC_7_42 b_7 NI_7 NS_42 0 -3.4993439195339796e-06
GC_7_43 b_7 NI_7 NS_43 0 9.7146747727948895e-06
GC_7_44 b_7 NI_7 NS_44 0 -5.0075302455725603e-05
GC_7_45 b_7 NI_7 NS_45 0 -6.6281364920266528e-05
GC_7_46 b_7 NI_7 NS_46 0 -2.1644695060868092e-05
GC_7_47 b_7 NI_7 NS_47 0 -1.6781843254161608e-05
GC_7_48 b_7 NI_7 NS_48 0 1.9314781944041681e-05
GC_7_49 b_7 NI_7 NS_49 0 1.6170796120583617e-05
GC_7_50 b_7 NI_7 NS_50 0 -1.3552353883624818e-06
GC_7_51 b_7 NI_7 NS_51 0 2.1848253065247930e-04
GC_7_52 b_7 NI_7 NS_52 0 7.6250192927573152e-06
GC_7_53 b_7 NI_7 NS_53 0 3.8540474143316329e-04
GC_7_54 b_7 NI_7 NS_54 0 -2.0233222528372365e-03
GC_7_55 b_7 NI_7 NS_55 0 4.0275552422384426e-10
GC_7_56 b_7 NI_7 NS_56 0 -2.6921602856865795e-08
GC_7_57 b_7 NI_7 NS_57 0 1.8880649690223802e-05
GC_7_58 b_7 NI_7 NS_58 0 4.3647508444377784e-05
GC_7_59 b_7 NI_7 NS_59 0 8.2161768395391953e-05
GC_7_60 b_7 NI_7 NS_60 0 -3.0679914495366656e-05
GC_7_61 b_7 NI_7 NS_61 0 -1.3443168522730596e-05
GC_7_62 b_7 NI_7 NS_62 0 1.3855590452207539e-05
GC_7_63 b_7 NI_7 NS_63 0 1.9803314081816973e-04
GC_7_64 b_7 NI_7 NS_64 0 -9.9134359246950225e-05
GC_7_65 b_7 NI_7 NS_65 0 2.7217482437235157e-05
GC_7_66 b_7 NI_7 NS_66 0 -9.8066136207506773e-05
GC_7_67 b_7 NI_7 NS_67 0 -1.7281658638423555e-05
GC_7_68 b_7 NI_7 NS_68 0 -9.8320967788343626e-05
GC_7_69 b_7 NI_7 NS_69 0 1.0631279030577422e-05
GC_7_70 b_7 NI_7 NS_70 0 -9.7299760636741179e-05
GC_7_71 b_7 NI_7 NS_71 0 -9.7211317435389282e-05
GC_7_72 b_7 NI_7 NS_72 0 -3.1576826249880754e-04
GC_7_73 b_7 NI_7 NS_73 0 -1.3368399231572116e-04
GC_7_74 b_7 NI_7 NS_74 0 -1.1528087974328368e-04
GC_7_75 b_7 NI_7 NS_75 0 -1.9126644302841283e-05
GC_7_76 b_7 NI_7 NS_76 0 -1.9117075071604158e-04
GC_7_77 b_7 NI_7 NS_77 0 1.5269827571986040e-03
GC_7_78 b_7 NI_7 NS_78 0 -9.9579655959236259e-05
GC_7_79 b_7 NI_7 NS_79 0 1.2876808315160588e-04
GC_7_80 b_7 NI_7 NS_80 0 5.3480700736054919e-05
GC_7_81 b_7 NI_7 NS_81 0 -4.2223190660913456e-10
GC_7_82 b_7 NI_7 NS_82 0 4.4745807335896226e-08
GC_7_83 b_7 NI_7 NS_83 0 5.7032040621346380e-06
GC_7_84 b_7 NI_7 NS_84 0 7.6084092926938915e-05
GC_7_85 b_7 NI_7 NS_85 0 1.5379578602551733e-04
GC_7_86 b_7 NI_7 NS_86 0 1.3562047509033882e-04
GC_7_87 b_7 NI_7 NS_87 0 3.4705294757742590e-04
GC_7_88 b_7 NI_7 NS_88 0 -2.3958201025522658e-05
GC_7_89 b_7 NI_7 NS_89 0 5.3192881825739770e-05
GC_7_90 b_7 NI_7 NS_90 0 -5.8496672809420789e-04
GC_7_91 b_7 NI_7 NS_91 0 -1.4500295560809971e-04
GC_7_92 b_7 NI_7 NS_92 0 -6.8356344218469084e-05
GC_7_93 b_7 NI_7 NS_93 0 5.2203007970130633e-05
GC_7_94 b_7 NI_7 NS_94 0 -1.0716135752307108e-05
GC_7_95 b_7 NI_7 NS_95 0 4.8321261798390794e-05
GC_7_96 b_7 NI_7 NS_96 0 -4.5206125148872174e-04
GC_7_97 b_7 NI_7 NS_97 0 -7.0676813662949687e-04
GC_7_98 b_7 NI_7 NS_98 0 -8.3391003003821572e-05
GC_7_99 b_7 NI_7 NS_99 0 -1.7416244046720319e-04
GC_7_100 b_7 NI_7 NS_100 0 2.5967712502026366e-04
GC_7_101 b_7 NI_7 NS_101 0 1.0231320530265359e-04
GC_7_102 b_7 NI_7 NS_102 0 8.1092296256021304e-05
GC_7_103 b_7 NI_7 NS_103 0 -1.2122269645667476e-04
GC_7_104 b_7 NI_7 NS_104 0 -3.3414336407553010e-04
GC_7_105 b_7 NI_7 NS_105 0 -7.6472777598514631e-03
GC_7_106 b_7 NI_7 NS_106 0 5.8567239269293383e-03
GC_7_107 b_7 NI_7 NS_107 0 -8.4251219674278836e-10
GC_7_108 b_7 NI_7 NS_108 0 -1.6876108431264057e-06
GC_7_109 b_7 NI_7 NS_109 0 2.5405881628338413e-04
GC_7_110 b_7 NI_7 NS_110 0 2.6638827817409877e-03
GC_7_111 b_7 NI_7 NS_111 0 4.5287651879800470e-03
GC_7_112 b_7 NI_7 NS_112 0 -2.7517441758933493e-03
GC_7_113 b_7 NI_7 NS_113 0 -5.4237649446824566e-03
GC_7_114 b_7 NI_7 NS_114 0 4.1627728340773191e-04
GC_7_115 b_7 NI_7 NS_115 0 8.8489949382731525e-03
GC_7_116 b_7 NI_7 NS_116 0 -6.0329864409836812e-04
GC_7_117 b_7 NI_7 NS_117 0 -2.8273784113507440e-03
GC_7_118 b_7 NI_7 NS_118 0 -2.3878795498347921e-03
GC_7_119 b_7 NI_7 NS_119 0 4.8268229086495656e-05
GC_7_120 b_7 NI_7 NS_120 0 -2.1045587978107141e-03
GC_7_121 b_7 NI_7 NS_121 0 -3.5071478368894019e-03
GC_7_122 b_7 NI_7 NS_122 0 5.5654795023737640e-03
GC_7_123 b_7 NI_7 NS_123 0 5.1183013216546227e-03
GC_7_124 b_7 NI_7 NS_124 0 -7.7286276384112571e-03
GC_7_125 b_7 NI_7 NS_125 0 -5.0253324617630735e-03
GC_7_126 b_7 NI_7 NS_126 0 3.1189361712689527e-03
GC_7_127 b_7 NI_7 NS_127 0 2.2497873076311849e-03
GC_7_128 b_7 NI_7 NS_128 0 -1.6595376517622511e-03
GC_7_129 b_7 NI_7 NS_129 0 -6.2720704311505461e-03
GC_7_130 b_7 NI_7 NS_130 0 3.8172621860018572e-03
GC_7_131 b_7 NI_7 NS_131 0 -1.3159048032284910e-03
GC_7_132 b_7 NI_7 NS_132 0 2.1722207299458012e-03
GC_7_133 b_7 NI_7 NS_133 0 7.7247492039753692e-10
GC_7_134 b_7 NI_7 NS_134 0 6.0126661879104851e-07
GC_7_135 b_7 NI_7 NS_135 0 -1.9612989217871986e-04
GC_7_136 b_7 NI_7 NS_136 0 -4.5795047464408260e-04
GC_7_137 b_7 NI_7 NS_137 0 -1.0663204084601916e-03
GC_7_138 b_7 NI_7 NS_138 0 -9.2689119069791698e-04
GC_7_139 b_7 NI_7 NS_139 0 -2.3216409846091679e-03
GC_7_140 b_7 NI_7 NS_140 0 3.0885303422369126e-04
GC_7_141 b_7 NI_7 NS_141 0 -3.5739848773951814e-04
GC_7_142 b_7 NI_7 NS_142 0 4.2021104394642092e-03
GC_7_143 b_7 NI_7 NS_143 0 9.8001058276248553e-04
GC_7_144 b_7 NI_7 NS_144 0 4.4275210728321793e-04
GC_7_145 b_7 NI_7 NS_145 0 -3.7449348107852808e-04
GC_7_146 b_7 NI_7 NS_146 0 7.7738857288901415e-05
GC_7_147 b_7 NI_7 NS_147 0 -3.1870783947904243e-04
GC_7_148 b_7 NI_7 NS_148 0 3.3550914906553134e-03
GC_7_149 b_7 NI_7 NS_149 0 5.2311011365012887e-03
GC_7_150 b_7 NI_7 NS_150 0 8.1047424476673980e-04
GC_7_151 b_7 NI_7 NS_151 0 1.3422336715926666e-03
GC_7_152 b_7 NI_7 NS_152 0 -1.9491672036624989e-03
GC_7_153 b_7 NI_7 NS_153 0 -8.8183379038938290e-04
GC_7_154 b_7 NI_7 NS_154 0 -6.4378730917925961e-04
GC_7_155 b_7 NI_7 NS_155 0 -1.3370800512422169e-03
GC_7_156 b_7 NI_7 NS_156 0 2.5847967361392467e-03
GC_7_157 b_7 NI_7 NS_157 0 5.9215545716411133e-02
GC_7_158 b_7 NI_7 NS_158 0 -6.3409888186437544e-02
GC_7_159 b_7 NI_7 NS_159 0 -1.0212118891351630e-08
GC_7_160 b_7 NI_7 NS_160 0 -8.2107767580865346e-06
GC_7_161 b_7 NI_7 NS_161 0 -1.8466559761794066e-03
GC_7_162 b_7 NI_7 NS_162 0 -2.8683128459668209e-03
GC_7_163 b_7 NI_7 NS_163 0 -5.1018024122670607e-03
GC_7_164 b_7 NI_7 NS_164 0 1.9432400523765054e-03
GC_7_165 b_7 NI_7 NS_165 0 2.4539734551011333e-03
GC_7_166 b_7 NI_7 NS_166 0 -1.2214794358196928e-03
GC_7_167 b_7 NI_7 NS_167 0 -1.0637006231012392e-02
GC_7_168 b_7 NI_7 NS_168 0 1.1057812879340645e-03
GC_7_169 b_7 NI_7 NS_169 0 6.4906461332207822e-04
GC_7_170 b_7 NI_7 NS_170 0 1.7568004895305227e-03
GC_7_171 b_7 NI_7 NS_171 0 -9.5190817421228621e-04
GC_7_172 b_7 NI_7 NS_172 0 2.2857441665880100e-03
GC_7_173 b_7 NI_7 NS_173 0 6.0496815202646325e-04
GC_7_174 b_7 NI_7 NS_174 0 -5.8869707909627797e-03
GC_7_175 b_7 NI_7 NS_175 0 -8.5212747052947971e-03
GC_7_176 b_7 NI_7 NS_176 0 6.8915948240748457e-03
GC_7_177 b_7 NI_7 NS_177 0 2.5250460717155931e-03
GC_7_178 b_7 NI_7 NS_178 0 -3.6699197998128364e-03
GC_7_179 b_7 NI_7 NS_179 0 -2.6398225470247033e-03
GC_7_180 b_7 NI_7 NS_180 0 -5.0015549797038320e-04
GC_7_181 b_7 NI_7 NS_181 0 5.4264680611438965e-02
GC_7_182 b_7 NI_7 NS_182 0 1.5897801271940819e-03
GC_7_183 b_7 NI_7 NS_183 0 -4.9912650990698186e-02
GC_7_184 b_7 NI_7 NS_184 0 1.0945976773453428e-01
GC_7_185 b_7 NI_7 NS_185 0 1.0779369496324964e-08
GC_7_186 b_7 NI_7 NS_186 0 1.9879994952018852e-05
GC_7_187 b_7 NI_7 NS_187 0 -1.5753182069471884e-02
GC_7_188 b_7 NI_7 NS_188 0 2.4251007673335396e-02
GC_7_189 b_7 NI_7 NS_189 0 -7.8027599945105254e-03
GC_7_190 b_7 NI_7 NS_190 0 -1.4488578218151228e-02
GC_7_191 b_7 NI_7 NS_191 0 2.0433220556028926e-02
GC_7_192 b_7 NI_7 NS_192 0 6.6873493377433641e-03
GC_7_193 b_7 NI_7 NS_193 0 8.0583355117086041e-03
GC_7_194 b_7 NI_7 NS_194 0 4.3992655741508326e-02
GC_7_195 b_7 NI_7 NS_195 0 -1.1853719755617198e-02
GC_7_196 b_7 NI_7 NS_196 0 -3.2338872784580873e-03
GC_7_197 b_7 NI_7 NS_197 0 -5.0942056376577860e-03
GC_7_198 b_7 NI_7 NS_198 0 -4.0938844441229492e-03
GC_7_199 b_7 NI_7 NS_199 0 2.6816844875280930e-02
GC_7_200 b_7 NI_7 NS_200 0 -8.8235822316711230e-06
GC_7_201 b_7 NI_7 NS_201 0 3.3872779953340620e-02
GC_7_202 b_7 NI_7 NS_202 0 3.0990188914985870e-02
GC_7_203 b_7 NI_7 NS_203 0 -1.5640908425233500e-02
GC_7_204 b_7 NI_7 NS_204 0 8.2834064567377588e-03
GC_7_205 b_7 NI_7 NS_205 0 -9.9433631433919786e-04
GC_7_206 b_7 NI_7 NS_206 0 -6.8669924362394982e-03
GC_7_207 b_7 NI_7 NS_207 0 -6.8767643625414099e-02
GC_7_208 b_7 NI_7 NS_208 0 1.7784390956096098e-03
GC_7_209 b_7 NI_7 NS_209 0 -1.2147766850268246e-03
GC_7_210 b_7 NI_7 NS_210 0 5.5868900861232636e-04
GC_7_211 b_7 NI_7 NS_211 0 3.0016424142646743e-10
GC_7_212 b_7 NI_7 NS_212 0 -5.7498731518362927e-07
GC_7_213 b_7 NI_7 NS_213 0 3.1227428524697041e-05
GC_7_214 b_7 NI_7 NS_214 0 6.3819814794441646e-04
GC_7_215 b_7 NI_7 NS_215 0 1.0888451722027603e-03
GC_7_216 b_7 NI_7 NS_216 0 -6.7567693431046358e-04
GC_7_217 b_7 NI_7 NS_217 0 -1.3740906963273965e-03
GC_7_218 b_7 NI_7 NS_218 0 7.5344570739183713e-05
GC_7_219 b_7 NI_7 NS_219 0 2.0944073047581401e-03
GC_7_220 b_7 NI_7 NS_220 0 -1.0659929526179310e-04
GC_7_221 b_7 NI_7 NS_221 0 -7.3376592626040816e-04
GC_7_222 b_7 NI_7 NS_222 0 -5.7284925311756765e-04
GC_7_223 b_7 NI_7 NS_223 0 5.7948715350829092e-06
GC_7_224 b_7 NI_7 NS_224 0 -4.8780379405073725e-04
GC_7_225 b_7 NI_7 NS_225 0 -9.0574312811513588e-04
GC_7_226 b_7 NI_7 NS_226 0 1.3911734445568227e-03
GC_7_227 b_7 NI_7 NS_227 0 1.2475487313830730e-03
GC_7_228 b_7 NI_7 NS_228 0 -1.8368924176892596e-03
GC_7_229 b_7 NI_7 NS_229 0 -1.2247766870124926e-03
GC_7_230 b_7 NI_7 NS_230 0 7.8190148089467987e-04
GC_7_231 b_7 NI_7 NS_231 0 5.7537113204741063e-04
GC_7_232 b_7 NI_7 NS_232 0 -4.1171102837814216e-04
GC_7_233 b_7 NI_7 NS_233 0 -7.3681762282656383e-04
GC_7_234 b_7 NI_7 NS_234 0 1.1397080052426328e-03
GC_7_235 b_7 NI_7 NS_235 0 -1.0982578765505117e-03
GC_7_236 b_7 NI_7 NS_236 0 1.9217212903037911e-03
GC_7_237 b_7 NI_7 NS_237 0 -1.0011976176653372e-10
GC_7_238 b_7 NI_7 NS_238 0 2.7261063218283314e-07
GC_7_239 b_7 NI_7 NS_239 0 5.8926676878478605e-05
GC_7_240 b_7 NI_7 NS_240 0 -8.7036768569161762e-05
GC_7_241 b_7 NI_7 NS_241 0 -2.6162990224484853e-04
GC_7_242 b_7 NI_7 NS_242 0 -1.7088135146712871e-04
GC_7_243 b_7 NI_7 NS_243 0 -5.2946161901550937e-04
GC_7_244 b_7 NI_7 NS_244 0 2.5218972936618971e-05
GC_7_245 b_7 NI_7 NS_245 0 4.2319761081346728e-05
GC_7_246 b_7 NI_7 NS_246 0 9.1574023628012346e-04
GC_7_247 b_7 NI_7 NS_247 0 2.4557870487389925e-04
GC_7_248 b_7 NI_7 NS_248 0 1.3068614065450641e-04
GC_7_249 b_7 NI_7 NS_249 0 -8.1516797593017833e-05
GC_7_250 b_7 NI_7 NS_250 0 2.6822493933045613e-05
GC_7_251 b_7 NI_7 NS_251 0 -7.1002100061892375e-05
GC_7_252 b_7 NI_7 NS_252 0 7.5354698037330924e-04
GC_7_253 b_7 NI_7 NS_253 0 1.2757768788860769e-03
GC_7_254 b_7 NI_7 NS_254 0 1.3796385185575147e-04
GC_7_255 b_7 NI_7 NS_255 0 3.2408105528303991e-04
GC_7_256 b_7 NI_7 NS_256 0 -4.2273775452169270e-04
GC_7_257 b_7 NI_7 NS_257 0 -2.4521740115315046e-04
GC_7_258 b_7 NI_7 NS_258 0 -1.0940951196285528e-04
GC_7_259 b_7 NI_7 NS_259 0 -1.5443533403494019e-03
GC_7_260 b_7 NI_7 NS_260 0 3.7327962330254127e-04
GC_7_261 b_7 NI_7 NS_261 0 3.9420725835198340e-04
GC_7_262 b_7 NI_7 NS_262 0 -2.0158041651288311e-03
GC_7_263 b_7 NI_7 NS_263 0 4.0775106436988400e-10
GC_7_264 b_7 NI_7 NS_264 0 -2.7128610086892232e-08
GC_7_265 b_7 NI_7 NS_265 0 1.8621476136846073e-05
GC_7_266 b_7 NI_7 NS_266 0 4.3392278918428386e-05
GC_7_267 b_7 NI_7 NS_267 0 8.1698018720038678e-05
GC_7_268 b_7 NI_7 NS_268 0 -3.0805112125441941e-05
GC_7_269 b_7 NI_7 NS_269 0 -1.3803874603529112e-05
GC_7_270 b_7 NI_7 NS_270 0 1.3744897747533755e-05
GC_7_271 b_7 NI_7 NS_271 0 1.9714653708874499e-04
GC_7_272 b_7 NI_7 NS_272 0 -9.9016356832570059e-05
GC_7_273 b_7 NI_7 NS_273 0 2.6817244362375208e-05
GC_7_274 b_7 NI_7 NS_274 0 -9.8015267835985706e-05
GC_7_275 b_7 NI_7 NS_275 0 -1.7477954192465305e-05
GC_7_276 b_7 NI_7 NS_276 0 -9.8100283084745585e-05
GC_7_277 b_7 NI_7 NS_277 0 9.9799348357493491e-06
GC_7_278 b_7 NI_7 NS_278 0 -9.7467350242713135e-05
GC_7_279 b_7 NI_7 NS_279 0 -9.8080466018231379e-05
GC_7_280 b_7 NI_7 NS_280 0 -3.1492223593655228e-04
GC_7_281 b_7 NI_7 NS_281 0 -1.3387635388897618e-04
GC_7_282 b_7 NI_7 NS_282 0 -1.1513419566297736e-04
GC_7_283 b_7 NI_7 NS_283 0 -1.9677621069679770e-05
GC_7_284 b_7 NI_7 NS_284 0 -1.9124507653991624e-04
GC_7_285 b_7 NI_7 NS_285 0 1.5196010033117551e-03
GC_7_286 b_7 NI_7 NS_286 0 -1.0206151654094538e-04
GC_7_287 b_7 NI_7 NS_287 0 1.5107002052955974e-04
GC_7_288 b_7 NI_7 NS_288 0 1.2317849256770206e-05
GC_7_289 b_7 NI_7 NS_289 0 -4.2760172502667801e-10
GC_7_290 b_7 NI_7 NS_290 0 4.5173474046794331e-08
GC_7_291 b_7 NI_7 NS_291 0 5.2778162143966404e-06
GC_7_292 b_7 NI_7 NS_292 0 7.5702684489769553e-05
GC_7_293 b_7 NI_7 NS_293 0 1.5331514859052856e-04
GC_7_294 b_7 NI_7 NS_294 0 1.3549625503205613e-04
GC_7_295 b_7 NI_7 NS_295 0 3.4661306293453785e-04
GC_7_296 b_7 NI_7 NS_296 0 -2.4832170563755508e-05
GC_7_297 b_7 NI_7 NS_297 0 5.1685677294125370e-05
GC_7_298 b_7 NI_7 NS_298 0 -5.8541630005264609e-04
GC_7_299 b_7 NI_7 NS_299 0 -1.4594533283728448e-04
GC_7_300 b_7 NI_7 NS_300 0 -6.8352176568999343e-05
GC_7_301 b_7 NI_7 NS_301 0 5.1710238290031612e-05
GC_7_302 b_7 NI_7 NS_302 0 -1.0508038789129435e-05
GC_7_303 b_7 NI_7 NS_303 0 4.7742078682248066e-05
GC_7_304 b_7 NI_7 NS_304 0 -4.5319513899674493e-04
GC_7_305 b_7 NI_7 NS_305 0 -7.0912994675149813e-04
GC_7_306 b_7 NI_7 NS_306 0 -8.3358421138813598e-05
GC_7_307 b_7 NI_7 NS_307 0 -1.7471253501016203e-04
GC_7_308 b_7 NI_7 NS_308 0 2.5874041175590317e-04
GC_7_309 b_7 NI_7 NS_309 0 1.0252651123468313e-04
GC_7_310 b_7 NI_7 NS_310 0 7.9813427780555760e-05
GC_7_311 b_7 NI_7 NS_311 0 -8.6272404746300850e-05
GC_7_312 b_7 NI_7 NS_312 0 -3.2981071536103824e-04
GD_7_1 b_7 NI_7 NA_1 0 7.5813342782774465e-07
GD_7_2 b_7 NI_7 NA_2 0 3.4878453258523752e-05
GD_7_3 b_7 NI_7 NA_3 0 1.6665145170272858e-04
GD_7_4 b_7 NI_7 NA_4 0 1.4002895097130997e-04
GD_7_5 b_7 NI_7 NA_5 0 1.3447779025220976e-02
GD_7_6 b_7 NI_7 NA_6 0 -1.1284130958466509e-03
GD_7_7 b_7 NI_7 NA_7 0 -2.9682548536956586e-02
GD_7_8 b_7 NI_7 NA_8 0 -2.0430107712356163e-02
GD_7_9 b_7 NI_7 NA_9 0 3.0067237936815421e-03
GD_7_10 b_7 NI_7 NA_10 0 -5.3852870598373075e-05
GD_7_11 b_7 NI_7 NA_11 0 1.6323049487556560e-04
GD_7_12 b_7 NI_7 NA_12 0 1.3331433768776040e-04
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 -1.6167546346001212e-05
GC_8_2 b_8 NI_8 NS_2 0 -2.5713233941492626e-04
GC_8_3 b_8 NI_8 NS_3 0 -1.0826303208586181e-10
GC_8_4 b_8 NI_8 NS_4 0 4.7617827419555280e-09
GC_8_5 b_8 NI_8 NS_5 0 5.0889302443760544e-06
GC_8_6 b_8 NI_8 NS_6 0 9.7287695765667816e-06
GC_8_7 b_8 NI_8 NS_7 0 1.6466340319762671e-05
GC_8_8 b_8 NI_8 NS_8 0 1.3314056333776607e-05
GC_8_9 b_8 NI_8 NS_9 0 3.8436504779952025e-05
GC_8_10 b_8 NI_8 NS_10 0 -3.5538485196520503e-06
GC_8_11 b_8 NI_8 NS_11 0 1.4511380251945124e-05
GC_8_12 b_8 NI_8 NS_12 0 -6.2679408067528377e-05
GC_8_13 b_8 NI_8 NS_13 0 -1.1740220998701557e-05
GC_8_14 b_8 NI_8 NS_14 0 -9.0260278370894769e-06
GC_8_15 b_8 NI_8 NS_15 0 4.7333674940266429e-06
GC_8_16 b_8 NI_8 NS_16 0 -3.5102473065850996e-06
GC_8_17 b_8 NI_8 NS_17 0 9.6833326691443547e-06
GC_8_18 b_8 NI_8 NS_18 0 -5.0075247857790665e-05
GC_8_19 b_8 NI_8 NS_19 0 -6.6267409859366994e-05
GC_8_20 b_8 NI_8 NS_20 0 -2.1578366250738504e-05
GC_8_21 b_8 NI_8 NS_21 0 -1.6765733735519055e-05
GC_8_22 b_8 NI_8 NS_22 0 1.9317411380766195e-05
GC_8_23 b_8 NI_8 NS_23 0 1.6177485038959895e-05
GC_8_24 b_8 NI_8 NS_24 0 -1.3689172287323076e-06
GC_8_25 b_8 NI_8 NS_25 0 2.1856805979095537e-04
GC_8_26 b_8 NI_8 NS_26 0 7.6285006144600530e-06
GC_8_27 b_8 NI_8 NS_27 0 -1.4356179702673877e-04
GC_8_28 b_8 NI_8 NS_28 0 6.6680320097223906e-04
GC_8_29 b_8 NI_8 NS_29 0 1.2440048255517016e-10
GC_8_30 b_8 NI_8 NS_30 0 -1.1384117251325469e-08
GC_8_31 b_8 NI_8 NS_31 0 -4.0172023088898646e-06
GC_8_32 b_8 NI_8 NS_32 0 -3.9916826661073943e-06
GC_8_33 b_8 NI_8 NS_33 0 -9.5853548017728028e-06
GC_8_34 b_8 NI_8 NS_34 0 -3.6874511816323813e-06
GC_8_35 b_8 NI_8 NS_35 0 -1.8731365440536228e-05
GC_8_36 b_8 NI_8 NS_36 0 -1.5342447717560008e-06
GC_8_37 b_8 NI_8 NS_37 0 -2.9271382836074807e-05
GC_8_38 b_8 NI_8 NS_38 0 2.7762771212752415e-05
GC_8_39 b_8 NI_8 NS_39 0 -2.1467904866000576e-05
GC_8_40 b_8 NI_8 NS_40 0 2.3556682973693485e-05
GC_8_41 b_8 NI_8 NS_41 0 6.1042869238306745e-06
GC_8_42 b_8 NI_8 NS_42 0 2.3439073128338383e-05
GC_8_43 b_8 NI_8 NS_43 0 -1.5895569090154768e-05
GC_8_44 b_8 NI_8 NS_44 0 5.5646865993752913e-05
GC_8_45 b_8 NI_8 NS_45 0 5.4417167291327347e-05
GC_8_46 b_8 NI_8 NS_46 0 6.5745678060251544e-05
GC_8_47 b_8 NI_8 NS_47 0 2.2593743178577830e-05
GC_8_48 b_8 NI_8 NS_48 0 4.5701641236649271e-05
GC_8_49 b_8 NI_8 NS_49 0 1.4942119515944652e-05
GC_8_50 b_8 NI_8 NS_50 0 4.9676076813549103e-05
GC_8_51 b_8 NI_8 NS_51 0 -5.1914710027336564e-04
GC_8_52 b_8 NI_8 NS_52 0 2.3890391155129313e-05
GC_8_53 b_8 NI_8 NS_53 0 1.2876638926023485e-04
GC_8_54 b_8 NI_8 NS_54 0 5.3481976805741583e-05
GC_8_55 b_8 NI_8 NS_55 0 -4.2223195079865327e-10
GC_8_56 b_8 NI_8 NS_56 0 4.4745786293387590e-08
GC_8_57 b_8 NI_8 NS_57 0 5.7031009502788389e-06
GC_8_58 b_8 NI_8 NS_58 0 7.6084235980778767e-05
GC_8_59 b_8 NI_8 NS_59 0 1.5379601437128689e-04
GC_8_60 b_8 NI_8 NS_60 0 1.3562073366501511e-04
GC_8_61 b_8 NI_8 NS_61 0 3.4705326895678723e-04
GC_8_62 b_8 NI_8 NS_62 0 -2.3957913000097628e-05
GC_8_63 b_8 NI_8 NS_63 0 5.3193170542316967e-05
GC_8_64 b_8 NI_8 NS_64 0 -5.8496731973744359e-04
GC_8_65 b_8 NI_8 NS_65 0 -1.4500299497281926e-04
GC_8_66 b_8 NI_8 NS_66 0 -6.8356434967202509e-05
GC_8_67 b_8 NI_8 NS_67 0 5.2203095453777032e-05
GC_8_68 b_8 NI_8 NS_68 0 -1.0716015634691465e-05
GC_8_69 b_8 NI_8 NS_69 0 4.8321452738715421e-05
GC_8_70 b_8 NI_8 NS_70 0 -4.5206117130000063e-04
GC_8_71 b_8 NI_8 NS_71 0 -7.0676797170387553e-04
GC_8_72 b_8 NI_8 NS_72 0 -8.3391432372071402e-05
GC_8_73 b_8 NI_8 NS_73 0 -1.7416249563174339e-04
GC_8_74 b_8 NI_8 NS_74 0 2.5967704049033492e-04
GC_8_75 b_8 NI_8 NS_75 0 1.0231312789714045e-04
GC_8_76 b_8 NI_8 NS_76 0 8.1092285045744335e-05
GC_8_77 b_8 NI_8 NS_77 0 -1.2122385674743239e-04
GC_8_78 b_8 NI_8 NS_78 0 -3.3414361046165216e-04
GC_8_79 b_8 NI_8 NS_79 0 3.8432217036462398e-04
GC_8_80 b_8 NI_8 NS_80 0 -2.0226219634084256e-03
GC_8_81 b_8 NI_8 NS_81 0 4.0280159499782288e-10
GC_8_82 b_8 NI_8 NS_82 0 -2.6940666819761023e-08
GC_8_83 b_8 NI_8 NS_83 0 1.8994438107017242e-05
GC_8_84 b_8 NI_8 NS_84 0 4.3663121558033101e-05
GC_8_85 b_8 NI_8 NS_85 0 8.2131171215708309e-05
GC_8_86 b_8 NI_8 NS_86 0 -3.0748892858536859e-05
GC_8_87 b_8 NI_8 NS_87 0 -1.3347310322054155e-05
GC_8_88 b_8 NI_8 NS_88 0 1.3987429665906454e-05
GC_8_89 b_8 NI_8 NS_89 0 1.9809683108304720e-04
GC_8_90 b_8 NI_8 NS_90 0 -9.9308113555127085e-05
GC_8_91 b_8 NI_8 NS_91 0 2.7246169287065153e-05
GC_8_92 b_8 NI_8 NS_92 0 -9.8014285630353652e-05
GC_8_93 b_8 NI_8 NS_93 0 -1.7287805123024855e-05
GC_8_94 b_8 NI_8 NS_94 0 -9.8335138630231494e-05
GC_8_95 b_8 NI_8 NS_95 0 1.0774117184646937e-05
GC_8_96 b_8 NI_8 NS_96 0 -9.7259054709234157e-05
GC_8_97 b_8 NI_8 NS_97 0 -9.7202756623346288e-05
GC_8_98 b_8 NI_8 NS_98 0 -3.1583836751997445e-04
GC_8_99 b_8 NI_8 NS_99 0 -1.3360484216877401e-04
GC_8_100 b_8 NI_8 NS_100 0 -1.1524848463245590e-04
GC_8_101 b_8 NI_8 NS_101 0 -1.9119749525387771e-05
GC_8_102 b_8 NI_8 NS_102 0 -1.9116379125838048e-04
GC_8_103 b_8 NI_8 NS_103 0 1.5264288686948335e-03
GC_8_104 b_8 NI_8 NS_104 0 -9.9582006932615597e-05
GC_8_105 b_8 NI_8 NS_105 0 -1.3158639644326115e-03
GC_8_106 b_8 NI_8 NS_106 0 2.1722220845998936e-03
GC_8_107 b_8 NI_8 NS_107 0 7.7247550757486874e-10
GC_8_108 b_8 NI_8 NS_108 0 6.0126670905295524e-07
GC_8_109 b_8 NI_8 NS_109 0 -1.9612813500728332e-04
GC_8_110 b_8 NI_8 NS_110 0 -4.5793429396826885e-04
GC_8_111 b_8 NI_8 NS_111 0 -1.0663224132102577e-03
GC_8_112 b_8 NI_8 NS_112 0 -9.2690698893546002e-04
GC_8_113 b_8 NI_8 NS_113 0 -2.3216377405192307e-03
GC_8_114 b_8 NI_8 NS_114 0 3.0883884497287772e-04
GC_8_115 b_8 NI_8 NS_115 0 -3.5741414742391684e-04
GC_8_116 b_8 NI_8 NS_116 0 4.2021284042181133e-03
GC_8_117 b_8 NI_8 NS_117 0 9.8000801436571748e-04
GC_8_118 b_8 NI_8 NS_118 0 4.4275717495873094e-04
GC_8_119 b_8 NI_8 NS_119 0 -3.7449557410707489e-04
GC_8_120 b_8 NI_8 NS_120 0 7.7736282896408463e-05
GC_8_121 b_8 NI_8 NS_121 0 -3.1871488331666010e-04
GC_8_122 b_8 NI_8 NS_122 0 3.3550933326939670e-03
GC_8_123 b_8 NI_8 NS_123 0 5.2311075295889799e-03
GC_8_124 b_8 NI_8 NS_124 0 8.1049137194075152e-04
GC_8_125 b_8 NI_8 NS_125 0 1.3422387448358958e-03
GC_8_126 b_8 NI_8 NS_126 0 -1.9491659262917194e-03
GC_8_127 b_8 NI_8 NS_127 0 -8.8183193801590184e-04
GC_8_128 b_8 NI_8 NS_128 0 -6.4378956059178596e-04
GC_8_129 b_8 NI_8 NS_129 0 -1.3370813004176705e-03
GC_8_130 b_8 NI_8 NS_130 0 2.5847959779031621e-03
GC_8_131 b_8 NI_8 NS_131 0 -7.6472780163477803e-03
GC_8_132 b_8 NI_8 NS_132 0 5.8567235176520483e-03
GC_8_133 b_8 NI_8 NS_133 0 -8.4251215129073530e-10
GC_8_134 b_8 NI_8 NS_134 0 -1.6876108882020200e-06
GC_8_135 b_8 NI_8 NS_135 0 2.5405881226811040e-04
GC_8_136 b_8 NI_8 NS_136 0 2.6638827778355570e-03
GC_8_137 b_8 NI_8 NS_137 0 4.5287651405927628e-03
GC_8_138 b_8 NI_8 NS_138 0 -2.7517441800721867e-03
GC_8_139 b_8 NI_8 NS_139 0 -5.4237649933211269e-03
GC_8_140 b_8 NI_8 NS_140 0 4.1627734726819797e-04
GC_8_141 b_8 NI_8 NS_141 0 8.8489949678563148e-03
GC_8_142 b_8 NI_8 NS_142 0 -6.0329856067815304e-04
GC_8_143 b_8 NI_8 NS_143 0 -2.8273784151118023e-03
GC_8_144 b_8 NI_8 NS_144 0 -2.3878794998851700e-03
GC_8_145 b_8 NI_8 NS_145 0 4.8268255975300471e-05
GC_8_146 b_8 NI_8 NS_146 0 -2.1045587677131837e-03
GC_8_147 b_8 NI_8 NS_147 0 -3.5071477919363728e-03
GC_8_148 b_8 NI_8 NS_148 0 5.5654796014008743e-03
GC_8_149 b_8 NI_8 NS_149 0 5.1183014482111613e-03
GC_8_150 b_8 NI_8 NS_150 0 -7.7286276105334884e-03
GC_8_151 b_8 NI_8 NS_151 0 -5.0253323951217474e-03
GC_8_152 b_8 NI_8 NS_152 0 3.1189362088843114e-03
GC_8_153 b_8 NI_8 NS_153 0 2.2497873906578260e-03
GC_8_154 b_8 NI_8 NS_154 0 -1.6595376233848702e-03
GC_8_155 b_8 NI_8 NS_155 0 -6.2720699667936728e-03
GC_8_156 b_8 NI_8 NS_156 0 3.8172623940375913e-03
GC_8_157 b_8 NI_8 NS_157 0 -4.9912615939729947e-02
GC_8_158 b_8 NI_8 NS_158 0 1.0945969476384075e-01
GC_8_159 b_8 NI_8 NS_159 0 1.0779367068884287e-08
GC_8_160 b_8 NI_8 NS_160 0 1.9879995593761137e-05
GC_8_161 b_8 NI_8 NS_161 0 -1.5753182422540347e-02
GC_8_162 b_8 NI_8 NS_162 0 2.4251006314715374e-02
GC_8_163 b_8 NI_8 NS_163 0 -7.8027610944894727e-03
GC_8_164 b_8 NI_8 NS_164 0 -1.4488579407464010e-02
GC_8_165 b_8 NI_8 NS_165 0 2.0433219688962192e-02
GC_8_166 b_8 NI_8 NS_166 0 6.6873482868715188e-03
GC_8_167 b_8 NI_8 NS_167 0 8.0583333712676633e-03
GC_8_168 b_8 NI_8 NS_168 0 4.3992655391015323e-02
GC_8_169 b_8 NI_8 NS_169 0 -1.1853720040041734e-02
GC_8_170 b_8 NI_8 NS_170 0 -3.2338883181902201e-03
GC_8_171 b_8 NI_8 NS_171 0 -5.0942066676139897e-03
GC_8_172 b_8 NI_8 NS_172 0 -4.0938851571480422e-03
GC_8_173 b_8 NI_8 NS_173 0 2.6816843409736439e-02
GC_8_174 b_8 NI_8 NS_174 0 -8.8262891987884688e-06
GC_8_175 b_8 NI_8 NS_175 0 3.3872775525771386e-02
GC_8_176 b_8 NI_8 NS_176 0 3.0990187487154479e-02
GC_8_177 b_8 NI_8 NS_177 0 -1.5640909823766754e-02
GC_8_178 b_8 NI_8 NS_178 0 8.2834043849423899e-03
GC_8_179 b_8 NI_8 NS_179 0 -9.9433627412317681e-04
GC_8_180 b_8 NI_8 NS_180 0 -6.8669959580531332e-03
GC_8_181 b_8 NI_8 NS_181 0 -6.8767583485058223e-02
GC_8_182 b_8 NI_8 NS_182 0 1.7784432136259277e-03
GC_8_183 b_8 NI_8 NS_183 0 5.9215545716411196e-02
GC_8_184 b_8 NI_8 NS_184 0 -6.3409888186437655e-02
GC_8_185 b_8 NI_8 NS_185 0 -1.0212118891352486e-08
GC_8_186 b_8 NI_8 NS_186 0 -8.2107767580865820e-06
GC_8_187 b_8 NI_8 NS_187 0 -1.8466559761794066e-03
GC_8_188 b_8 NI_8 NS_188 0 -2.8683128459668257e-03
GC_8_189 b_8 NI_8 NS_189 0 -5.1018024122670624e-03
GC_8_190 b_8 NI_8 NS_190 0 1.9432400523765022e-03
GC_8_191 b_8 NI_8 NS_191 0 2.4539734551011225e-03
GC_8_192 b_8 NI_8 NS_192 0 -1.2214794358196969e-03
GC_8_193 b_8 NI_8 NS_193 0 -1.0637006231012398e-02
GC_8_194 b_8 NI_8 NS_194 0 1.1057812879340678e-03
GC_8_195 b_8 NI_8 NS_195 0 6.4906461332207095e-04
GC_8_196 b_8 NI_8 NS_196 0 1.7568004895305255e-03
GC_8_197 b_8 NI_8 NS_197 0 -9.5190817421228469e-04
GC_8_198 b_8 NI_8 NS_198 0 2.2857441665880131e-03
GC_8_199 b_8 NI_8 NS_199 0 6.0496815202646130e-04
GC_8_200 b_8 NI_8 NS_200 0 -5.8869707909627797e-03
GC_8_201 b_8 NI_8 NS_201 0 -8.5212747052948023e-03
GC_8_202 b_8 NI_8 NS_202 0 6.8915948240748474e-03
GC_8_203 b_8 NI_8 NS_203 0 2.5250460717155926e-03
GC_8_204 b_8 NI_8 NS_204 0 -3.6699197998128394e-03
GC_8_205 b_8 NI_8 NS_205 0 -2.6398225470247029e-03
GC_8_206 b_8 NI_8 NS_206 0 -5.0015549797038776e-04
GC_8_207 b_8 NI_8 NS_207 0 5.4264680611439062e-02
GC_8_208 b_8 NI_8 NS_208 0 1.5897801271940947e-03
GC_8_209 b_8 NI_8 NS_209 0 -1.0983047198724612e-03
GC_8_210 b_8 NI_8 NS_210 0 1.9215778567149241e-03
GC_8_211 b_8 NI_8 NS_211 0 -1.0012200778960880e-10
GC_8_212 b_8 NI_8 NS_212 0 2.7261165841861971e-07
GC_8_213 b_8 NI_8 NS_213 0 5.8917471588614681e-05
GC_8_214 b_8 NI_8 NS_214 0 -8.7105571411952260e-05
GC_8_215 b_8 NI_8 NS_215 0 -2.6162502003455255e-04
GC_8_216 b_8 NI_8 NS_216 0 -1.7081949714302621e-04
GC_8_217 b_8 NI_8 NS_217 0 -5.2947831462674545e-04
GC_8_218 b_8 NI_8 NS_218 0 2.5272764143830444e-05
GC_8_219 b_8 NI_8 NS_219 0 4.2373178823795556e-05
GC_8_220 b_8 NI_8 NS_220 0 9.1566637871523927e-04
GC_8_221 b_8 NI_8 NS_221 0 2.4558524419294547e-04
GC_8_222 b_8 NI_8 NS_222 0 1.3066484492986829e-04
GC_8_223 b_8 NI_8 NS_223 0 -8.1510649632403763e-05
GC_8_224 b_8 NI_8 NS_224 0 2.6833724058776324e-05
GC_8_225 b_8 NI_8 NS_225 0 -7.0978323293623491e-05
GC_8_226 b_8 NI_8 NS_226 0 7.5353511020353223e-04
GC_8_227 b_8 NI_8 NS_227 0 1.2757395607046178e-03
GC_8_228 b_8 NI_8 NS_228 0 1.3789245542054302e-04
GC_8_229 b_8 NI_8 NS_229 0 3.2405502316563240e-04
GC_8_230 b_8 NI_8 NS_230 0 -4.2274714571759582e-04
GC_8_231 b_8 NI_8 NS_231 0 -2.4522716599664329e-04
GC_8_232 b_8 NI_8 NS_232 0 -1.0940685519728147e-04
GC_8_233 b_8 NI_8 NS_233 0 -1.5442371277728636e-03
GC_8_234 b_8 NI_8 NS_234 0 3.7328710229100366e-04
GC_8_235 b_8 NI_8 NS_235 0 -1.2147410732494101e-03
GC_8_236 b_8 NI_8 NS_236 0 5.5866870161100281e-04
GC_8_237 b_8 NI_8 NS_237 0 3.0016891516189231e-10
GC_8_238 b_8 NI_8 NS_238 0 -5.7498703536090579e-07
GC_8_239 b_8 NI_8 NS_239 0 3.1226506345418348e-05
GC_8_240 b_8 NI_8 NS_240 0 6.3819819137128555e-04
GC_8_241 b_8 NI_8 NS_241 0 1.0888429695922648e-03
GC_8_242 b_8 NI_8 NS_242 0 -6.7567588582472524e-04
GC_8_243 b_8 NI_8 NS_243 0 -1.3740894625347596e-03
GC_8_244 b_8 NI_8 NS_244 0 7.5346247359486755e-05
GC_8_245 b_8 NI_8 NS_245 0 2.0944046447536643e-03
GC_8_246 b_8 NI_8 NS_246 0 -1.0660111672496194e-04
GC_8_247 b_8 NI_8 NS_247 0 -7.3376676690411959e-04
GC_8_248 b_8 NI_8 NS_248 0 -5.7284806421391634e-04
GC_8_249 b_8 NI_8 NS_249 0 5.7939154522137194e-06
GC_8_250 b_8 NI_8 NS_250 0 -4.8780333068000593e-04
GC_8_251 b_8 NI_8 NS_251 0 -9.0574288576900064e-04
GC_8_252 b_8 NI_8 NS_252 0 1.3911749225337592e-03
GC_8_253 b_8 NI_8 NS_253 0 1.2475474352374131e-03
GC_8_254 b_8 NI_8 NS_254 0 -1.8368940342357038e-03
GC_8_255 b_8 NI_8 NS_255 0 -1.2247777879912086e-03
GC_8_256 b_8 NI_8 NS_256 0 7.8190085781550513e-04
GC_8_257 b_8 NI_8 NS_257 0 5.7537071758387195e-04
GC_8_258 b_8 NI_8 NS_258 0 -4.1171263888531884e-04
GC_8_259 b_8 NI_8 NS_259 0 -7.3680273455707754e-04
GC_8_260 b_8 NI_8 NS_260 0 1.1397051971127291e-03
GC_8_261 b_8 NI_8 NS_261 0 1.5103108357690696e-04
GC_8_262 b_8 NI_8 NS_262 0 1.2368461311741488e-05
GC_8_263 b_8 NI_8 NS_263 0 -4.2760090215683310e-10
GC_8_264 b_8 NI_8 NS_264 0 4.5173254185240784e-08
GC_8_265 b_8 NI_8 NS_265 0 5.2792762435066730e-06
GC_8_266 b_8 NI_8 NS_266 0 7.5700598064378969e-05
GC_8_267 b_8 NI_8 NS_267 0 1.5331439972273000e-04
GC_8_268 b_8 NI_8 NS_268 0 1.3549913111244533e-04
GC_8_269 b_8 NI_8 NS_269 0 3.4661139668886321e-04
GC_8_270 b_8 NI_8 NS_270 0 -2.4829789413242371e-05
GC_8_271 b_8 NI_8 NS_271 0 5.1691377674675405e-05
GC_8_272 b_8 NI_8 NS_272 0 -5.8541576760627123e-04
GC_8_273 b_8 NI_8 NS_273 0 -1.4594355466272620e-04
GC_8_274 b_8 NI_8 NS_274 0 -6.8351846251356869e-05
GC_8_275 b_8 NI_8 NS_275 0 5.1710930944460901e-05
GC_8_276 b_8 NI_8 NS_276 0 -1.0507735904095151e-05
GC_8_277 b_8 NI_8 NS_277 0 4.7743656745994047e-05
GC_8_278 b_8 NI_8 NS_278 0 -4.5319346338904779e-04
GC_8_279 b_8 NI_8 NS_279 0 -7.0912542376299096e-04
GC_8_280 b_8 NI_8 NS_280 0 -8.3358066986932938e-05
GC_8_281 b_8 NI_8 NS_281 0 -1.7471104938664121e-04
GC_8_282 b_8 NI_8 NS_282 0 2.5874147755709982e-04
GC_8_283 b_8 NI_8 NS_283 0 1.0252688935255387e-04
GC_8_284 b_8 NI_8 NS_284 0 7.9815961575267362e-05
GC_8_285 b_8 NI_8 NS_285 0 -8.6313407181137954e-05
GC_8_286 b_8 NI_8 NS_286 0 -3.2981257549434312e-04
GC_8_287 b_8 NI_8 NS_287 0 3.9532339352367192e-04
GC_8_288 b_8 NI_8 NS_288 0 -2.0165266085578133e-03
GC_8_289 b_8 NI_8 NS_289 0 4.0770693374240989e-10
GC_8_290 b_8 NI_8 NS_290 0 -2.7109177959273493e-08
GC_8_291 b_8 NI_8 NS_291 0 1.8507561981177049e-05
GC_8_292 b_8 NI_8 NS_292 0 4.3378359690435352e-05
GC_8_293 b_8 NI_8 NS_293 0 8.1727560238208755e-05
GC_8_294 b_8 NI_8 NS_294 0 -3.0737467716388291e-05
GC_8_295 b_8 NI_8 NS_295 0 -1.3901175957216243e-05
GC_8_296 b_8 NI_8 NS_296 0 1.3616746976200068e-05
GC_8_297 b_8 NI_8 NS_297 0 1.9708381335272452e-04
GC_8_298 b_8 NI_8 NS_298 0 -9.8844897497924765e-05
GC_8_299 b_8 NI_8 NS_299 0 2.6786766085916242e-05
GC_8_300 b_8 NI_8 NS_300 0 -9.8065688745305313e-05
GC_8_301 b_8 NI_8 NS_301 0 -1.7472511380316244e-05
GC_8_302 b_8 NI_8 NS_302 0 -9.8086077282896847e-05
GC_8_303 b_8 NI_8 NS_303 0 9.8369786541569102e-06
GC_8_304 b_8 NI_8 NS_304 0 -9.7505027330488942e-05
GC_8_305 b_8 NI_8 NS_305 0 -9.8088434170964616e-05
GC_8_306 b_8 NI_8 NS_306 0 -3.1485388161739674e-04
GC_8_307 b_8 NI_8 NS_307 0 -1.3395601705570241e-04
GC_8_308 b_8 NI_8 NS_308 0 -1.1516728148377077e-04
GC_8_309 b_8 NI_8 NS_309 0 -1.9684699152375215e-05
GC_8_310 b_8 NI_8 NS_310 0 -1.9125377951374921e-04
GC_8_311 b_8 NI_8 NS_311 0 1.5201720367583221e-03
GC_8_312 b_8 NI_8 NS_312 0 -1.0206019962982020e-04
GD_8_1 b_8 NI_8 NA_1 0 3.4782103774728116e-05
GD_8_2 b_8 NI_8 NA_2 0 7.4465323313469096e-07
GD_8_3 b_8 NI_8 NA_3 0 1.4002930261906244e-04
GD_8_4 b_8 NI_8 NA_4 0 1.6665991033260245e-04
GD_8_5 b_8 NI_8 NA_5 0 -1.1284369305385969e-03
GD_8_6 b_8 NI_8 NA_6 0 1.3447778880549989e-02
GD_8_7 b_8 NI_8 NA_7 0 -2.0430112943460196e-02
GD_8_8 b_8 NI_8 NA_8 0 -2.9682548536956510e-02
GD_8_9 b_8 NI_8 NA_9 0 -5.3787250140997398e-05
GD_8_10 b_8 NI_8 NA_10 0 3.0067015982982387e-03
GD_8_11 b_8 NI_8 NA_11 0 1.3332437404675219e-04
GD_8_12 b_8 NI_8 NA_12 0 1.6319284778228848e-04
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 -2.7825253317720535e-05
GC_9_2 b_9 NI_9 NS_2 0 4.2360480970062478e-05
GC_9_3 b_9 NI_9 NS_3 0 3.6705452149573874e-11
GC_9_4 b_9 NI_9 NS_4 0 -2.7773099347400120e-10
GC_9_5 b_9 NI_9 NS_5 0 8.4146527350424023e-07
GC_9_6 b_9 NI_9 NS_6 0 4.8946649218755071e-07
GC_9_7 b_9 NI_9 NS_7 0 4.0299542583822256e-07
GC_9_8 b_9 NI_9 NS_8 0 -7.5688550334365094e-07
GC_9_9 b_9 NI_9 NS_9 0 -4.8229317115985230e-07
GC_9_10 b_9 NI_9 NS_10 0 9.9668466970067931e-07
GC_9_11 b_9 NI_9 NS_11 0 1.4113530950785409e-06
GC_9_12 b_9 NI_9 NS_12 0 1.8134196639004098e-07
GC_9_13 b_9 NI_9 NS_13 0 -4.2582299094129303e-07
GC_9_14 b_9 NI_9 NS_14 0 9.6992937776628908e-07
GC_9_15 b_9 NI_9 NS_15 0 5.7117605787853569e-07
GC_9_16 b_9 NI_9 NS_16 0 3.8256426642473781e-07
GC_9_17 b_9 NI_9 NS_17 0 5.5721832766273417e-07
GC_9_18 b_9 NI_9 NS_18 0 3.2490416989827340e-06
GC_9_19 b_9 NI_9 NS_19 0 4.0010697382329025e-06
GC_9_20 b_9 NI_9 NS_20 0 7.7940026603567249e-07
GC_9_21 b_9 NI_9 NS_21 0 9.0180422010192130e-07
GC_9_22 b_9 NI_9 NS_22 0 2.3877079675032606e-06
GC_9_23 b_9 NI_9 NS_23 0 1.1488164887782043e-06
GC_9_24 b_9 NI_9 NS_24 0 2.6084903508666871e-06
GC_9_25 b_9 NI_9 NS_25 0 -3.3517704592232139e-05
GC_9_26 b_9 NI_9 NS_26 0 4.1416089652152652e-07
GC_9_27 b_9 NI_9 NS_27 0 -2.4824765179544829e-05
GC_9_28 b_9 NI_9 NS_28 0 2.0783343909777786e-05
GC_9_29 b_9 NI_9 NS_29 0 -3.5006742735123628e-11
GC_9_30 b_9 NI_9 NS_30 0 -2.7089689726622501e-10
GC_9_31 b_9 NI_9 NS_31 0 1.6165286210569925e-06
GC_9_32 b_9 NI_9 NS_32 0 1.4394623452483613e-06
GC_9_33 b_9 NI_9 NS_33 0 2.5877682590230377e-07
GC_9_34 b_9 NI_9 NS_34 0 3.7182413012778879e-07
GC_9_35 b_9 NI_9 NS_35 0 1.7412280379383222e-06
GC_9_36 b_9 NI_9 NS_36 0 -2.0422228138728400e-07
GC_9_37 b_9 NI_9 NS_37 0 3.3659168890189227e-06
GC_9_38 b_9 NI_9 NS_38 0 -1.0270819605054827e-06
GC_9_39 b_9 NI_9 NS_39 0 4.2248026054265377e-07
GC_9_40 b_9 NI_9 NS_40 0 5.0189528753038571e-08
GC_9_41 b_9 NI_9 NS_41 0 2.5404315542185467e-07
GC_9_42 b_9 NI_9 NS_42 0 -2.9664613625610492e-07
GC_9_43 b_9 NI_9 NS_43 0 1.0839712532254712e-06
GC_9_44 b_9 NI_9 NS_44 0 -1.0041649823866649e-06
GC_9_45 b_9 NI_9 NS_45 0 1.6346565800343606e-06
GC_9_46 b_9 NI_9 NS_46 0 -1.2123161557508548e-06
GC_9_47 b_9 NI_9 NS_47 0 -5.8140804426424332e-08
GC_9_48 b_9 NI_9 NS_48 0 1.3019229353536975e-06
GC_9_49 b_9 NI_9 NS_49 0 3.3326938358625586e-07
GC_9_50 b_9 NI_9 NS_50 0 6.8673194077664838e-07
GC_9_51 b_9 NI_9 NS_51 0 -1.6980528151601013e-05
GC_9_52 b_9 NI_9 NS_52 0 -1.3435380259202514e-06
GC_9_53 b_9 NI_9 NS_53 0 -6.5847272516456971e-06
GC_9_54 b_9 NI_9 NS_54 0 9.9213280311678722e-05
GC_9_55 b_9 NI_9 NS_55 0 6.2415148636732235e-11
GC_9_56 b_9 NI_9 NS_56 0 -2.6617611451689750e-09
GC_9_57 b_9 NI_9 NS_57 0 -1.4903849639240146e-06
GC_9_58 b_9 NI_9 NS_58 0 -1.5556180129947433e-06
GC_9_59 b_9 NI_9 NS_59 0 -2.8329214769700996e-06
GC_9_60 b_9 NI_9 NS_60 0 -1.5879025450239912e-06
GC_9_61 b_9 NI_9 NS_61 0 -5.7178311624726976e-06
GC_9_62 b_9 NI_9 NS_62 0 -1.2614456191399888e-06
GC_9_63 b_9 NI_9 NS_63 0 -8.7595590444695392e-06
GC_9_64 b_9 NI_9 NS_64 0 6.4067485413983382e-06
GC_9_65 b_9 NI_9 NS_65 0 -6.4092312594614174e-06
GC_9_66 b_9 NI_9 NS_66 0 5.1019689659470569e-06
GC_9_67 b_9 NI_9 NS_67 0 8.4424483951109653e-07
GC_9_68 b_9 NI_9 NS_68 0 5.8470265283187179e-06
GC_9_69 b_9 NI_9 NS_69 0 -5.3961581876285884e-06
GC_9_70 b_9 NI_9 NS_70 0 1.2705497053305607e-05
GC_9_71 b_9 NI_9 NS_71 0 1.0828083282777947e-05
GC_9_72 b_9 NI_9 NS_72 0 1.5435675911834708e-05
GC_9_73 b_9 NI_9 NS_73 0 4.5989209896435773e-06
GC_9_74 b_9 NI_9 NS_74 0 1.0589226905583486e-05
GC_9_75 b_9 NI_9 NS_75 0 4.7903832595351659e-06
GC_9_76 b_9 NI_9 NS_76 0 9.9605484615789344e-06
GC_9_77 b_9 NI_9 NS_77 0 -7.2520401022305129e-05
GC_9_78 b_9 NI_9 NS_78 0 1.2870693080633802e-05
GC_9_79 b_9 NI_9 NS_79 0 -2.7806073643109790e-05
GC_9_80 b_9 NI_9 NS_80 0 -1.1427843456095774e-06
GC_9_81 b_9 NI_9 NS_81 0 -5.6802035487823329e-11
GC_9_82 b_9 NI_9 NS_82 0 1.0423995783348966e-09
GC_9_83 b_9 NI_9 NS_83 0 3.7494144587854289e-06
GC_9_84 b_9 NI_9 NS_84 0 4.4298204415077601e-06
GC_9_85 b_9 NI_9 NS_85 0 3.3687706566898657e-06
GC_9_86 b_9 NI_9 NS_86 0 3.3453251196240462e-06
GC_9_87 b_9 NI_9 NS_87 0 1.0419182530001227e-05
GC_9_88 b_9 NI_9 NS_88 0 -2.9807487347751072e-06
GC_9_89 b_9 NI_9 NS_89 0 6.6061138309756580e-06
GC_9_90 b_9 NI_9 NS_90 0 -1.4562633198855352e-05
GC_9_91 b_9 NI_9 NS_91 0 -3.0165739893926087e-06
GC_9_92 b_9 NI_9 NS_92 0 -1.0861343721468929e-06
GC_9_93 b_9 NI_9 NS_93 0 9.4457582140669989e-07
GC_9_94 b_9 NI_9 NS_94 0 -8.3627612097326185e-07
GC_9_95 b_9 NI_9 NS_95 0 2.9369379841157936e-06
GC_9_96 b_9 NI_9 NS_96 0 -1.2938430937170143e-05
GC_9_97 b_9 NI_9 NS_97 0 -1.3690771053465228e-05
GC_9_98 b_9 NI_9 NS_98 0 -3.7596286181055994e-06
GC_9_99 b_9 NI_9 NS_99 0 -3.5380576875046690e-06
GC_9_100 b_9 NI_9 NS_100 0 5.8960607497122954e-06
GC_9_101 b_9 NI_9 NS_101 0 2.7026886968700820e-06
GC_9_102 b_9 NI_9 NS_102 0 1.1370566590409766e-06
GC_9_103 b_9 NI_9 NS_103 0 1.7480503162410350e-07
GC_9_104 b_9 NI_9 NS_104 0 -5.8082586159609685e-06
GC_9_105 b_9 NI_9 NS_105 0 3.8512279775502383e-04
GC_9_106 b_9 NI_9 NS_106 0 -2.0245853373034727e-03
GC_9_107 b_9 NI_9 NS_107 0 4.0264790318012384e-10
GC_9_108 b_9 NI_9 NS_108 0 -2.6912814427789660e-08
GC_9_109 b_9 NI_9 NS_109 0 1.8964557408948703e-05
GC_9_110 b_9 NI_9 NS_110 0 4.3646769283366990e-05
GC_9_111 b_9 NI_9 NS_111 0 8.2121180923165130e-05
GC_9_112 b_9 NI_9 NS_112 0 -3.0735340105735475e-05
GC_9_113 b_9 NI_9 NS_113 0 -1.3364254681332558e-05
GC_9_114 b_9 NI_9 NS_114 0 1.3940739764703039e-05
GC_9_115 b_9 NI_9 NS_115 0 1.9803504368590054e-04
GC_9_116 b_9 NI_9 NS_116 0 -9.9273347580171970e-05
GC_9_117 b_9 NI_9 NS_117 0 2.7239745475352741e-05
GC_9_118 b_9 NI_9 NS_118 0 -9.8033292455776056e-05
GC_9_119 b_9 NI_9 NS_119 0 -1.7295797815720240e-05
GC_9_120 b_9 NI_9 NS_120 0 -9.8327848335149669e-05
GC_9_121 b_9 NI_9 NS_121 0 1.0740655661349599e-05
GC_9_122 b_9 NI_9 NS_122 0 -9.7316253649717496e-05
GC_9_123 b_9 NI_9 NS_123 0 -9.7269565132599537e-05
GC_9_124 b_9 NI_9 NS_124 0 -3.1582661461632692e-04
GC_9_125 b_9 NI_9 NS_125 0 -1.3361352245252648e-04
GC_9_126 b_9 NI_9 NS_126 0 -1.1528990621692888e-04
GC_9_127 b_9 NI_9 NS_127 0 -1.9094748588045034e-05
GC_9_128 b_9 NI_9 NS_128 0 -1.9121733297875447e-04
GC_9_129 b_9 NI_9 NS_129 0 1.5281239979811731e-03
GC_9_130 b_9 NI_9 NS_130 0 -9.9340182592612153e-05
GC_9_131 b_9 NI_9 NS_131 0 1.2824482784304245e-04
GC_9_132 b_9 NI_9 NS_132 0 5.5586338990865712e-05
GC_9_133 b_9 NI_9 NS_133 0 -4.2209249767122762e-10
GC_9_134 b_9 NI_9 NS_134 0 4.4721732783179159e-08
GC_9_135 b_9 NI_9 NS_135 0 5.7604319127083250e-06
GC_9_136 b_9 NI_9 NS_136 0 7.6123947643920057e-05
GC_9_137 b_9 NI_9 NS_137 0 1.5376806698385386e-04
GC_9_138 b_9 NI_9 NS_138 0 1.3563431492034887e-04
GC_9_139 b_9 NI_9 NS_139 0 3.4707304563695406e-04
GC_9_140 b_9 NI_9 NS_140 0 -2.4008687850771267e-05
GC_9_141 b_9 NI_9 NS_141 0 5.3250620887962043e-05
GC_9_142 b_9 NI_9 NS_142 0 -5.8494565294516193e-04
GC_9_143 b_9 NI_9 NS_143 0 -1.4501223050704506e-04
GC_9_144 b_9 NI_9 NS_144 0 -6.8322989817517514e-05
GC_9_145 b_9 NI_9 NS_145 0 5.2206224525304681e-05
GC_9_146 b_9 NI_9 NS_146 0 -1.0707672238993501e-05
GC_9_147 b_9 NI_9 NS_147 0 4.8324650209925473e-05
GC_9_148 b_9 NI_9 NS_148 0 -4.5206767781065136e-04
GC_9_149 b_9 NI_9 NS_149 0 -7.0671503615724691e-04
GC_9_150 b_9 NI_9 NS_150 0 -8.3345688649039102e-05
GC_9_151 b_9 NI_9 NS_151 0 -1.7415344933027540e-04
GC_9_152 b_9 NI_9 NS_152 0 2.5972212759007549e-04
GC_9_153 b_9 NI_9 NS_153 0 1.0227107644378453e-04
GC_9_154 b_9 NI_9 NS_154 0 8.1142078434611728e-05
GC_9_155 b_9 NI_9 NS_155 0 -1.2306560694197455e-04
GC_9_156 b_9 NI_9 NS_156 0 -3.3447033340213729e-04
GC_9_157 b_9 NI_9 NS_157 0 -1.2147410755369739e-03
GC_9_158 b_9 NI_9 NS_158 0 5.5866869281773082e-04
GC_9_159 b_9 NI_9 NS_159 0 3.0016891468441797e-10
GC_9_160 b_9 NI_9 NS_160 0 -5.7498703510631130e-07
GC_9_161 b_9 NI_9 NS_161 0 3.1226506211848767e-05
GC_9_162 b_9 NI_9 NS_162 0 6.3819819143119054e-04
GC_9_163 b_9 NI_9 NS_163 0 1.0888429694894662e-03
GC_9_164 b_9 NI_9 NS_164 0 -6.7567588567620733e-04
GC_9_165 b_9 NI_9 NS_165 0 -1.3740894626869833e-03
GC_9_166 b_9 NI_9 NS_166 0 7.5346247553915308e-05
GC_9_167 b_9 NI_9 NS_167 0 2.0944046448194338e-03
GC_9_168 b_9 NI_9 NS_168 0 -1.0660111617937601e-04
GC_9_169 b_9 NI_9 NS_169 0 -7.3376676685907316e-04
GC_9_170 b_9 NI_9 NS_170 0 -5.7284806389186634e-04
GC_9_171 b_9 NI_9 NS_171 0 5.7939156526512609e-06
GC_9_172 b_9 NI_9 NS_172 0 -4.8780333053988282e-04
GC_9_173 b_9 NI_9 NS_173 0 -9.0574288561763995e-04
GC_9_174 b_9 NI_9 NS_174 0 1.3911749231120402e-03
GC_9_175 b_9 NI_9 NS_175 0 1.2475474362186815e-03
GC_9_176 b_9 NI_9 NS_176 0 -1.8368940338072354e-03
GC_9_177 b_9 NI_9 NS_177 0 -1.2247777872286469e-03
GC_9_178 b_9 NI_9 NS_178 0 7.8190085804032388e-04
GC_9_179 b_9 NI_9 NS_179 0 5.7537071841502882e-04
GC_9_180 b_9 NI_9 NS_180 0 -4.1171263898725265e-04
GC_9_181 b_9 NI_9 NS_181 0 -7.3680272603912178e-04
GC_9_182 b_9 NI_9 NS_182 0 1.1397051997029657e-03
GC_9_183 b_9 NI_9 NS_183 0 -1.0982578697247168e-03
GC_9_184 b_9 NI_9 NS_184 0 1.9217212486725844e-03
GC_9_185 b_9 NI_9 NS_185 0 -1.0011977933921596e-10
GC_9_186 b_9 NI_9 NS_186 0 2.7261063438915587e-07
GC_9_187 b_9 NI_9 NS_187 0 5.8926677126540295e-05
GC_9_188 b_9 NI_9 NS_188 0 -8.7036768548511085e-05
GC_9_189 b_9 NI_9 NS_189 0 -2.6162990191140703e-04
GC_9_190 b_9 NI_9 NS_190 0 -1.7088135161437857e-04
GC_9_191 b_9 NI_9 NS_191 0 -5.2946161843356147e-04
GC_9_192 b_9 NI_9 NS_192 0 2.5218972718356703e-05
GC_9_193 b_9 NI_9 NS_193 0 4.2319761513302712e-05
GC_9_194 b_9 NI_9 NS_194 0 9.1574023472713786e-04
GC_9_195 b_9 NI_9 NS_195 0 2.4557870477003003e-04
GC_9_196 b_9 NI_9 NS_196 0 1.3068613957945420e-04
GC_9_197 b_9 NI_9 NS_197 0 -8.1516798159253395e-05
GC_9_198 b_9 NI_9 NS_198 0 2.6822493678379699e-05
GC_9_199 b_9 NI_9 NS_199 0 -7.1002100108367934e-05
GC_9_200 b_9 NI_9 NS_200 0 7.5354697931167755e-04
GC_9_201 b_9 NI_9 NS_201 0 1.2757768777081097e-03
GC_9_202 b_9 NI_9 NS_202 0 1.3796385031185674e-04
GC_9_203 b_9 NI_9 NS_203 0 3.2408105494257153e-04
GC_9_204 b_9 NI_9 NS_204 0 -4.2273775586633601e-04
GC_9_205 b_9 NI_9 NS_205 0 -2.4521740082313347e-04
GC_9_206 b_9 NI_9 NS_206 0 -1.0940951370403582e-04
GC_9_207 b_9 NI_9 NS_207 0 -1.5443533049606063e-03
GC_9_208 b_9 NI_9 NS_208 0 3.7327962780640410e-04
GC_9_209 b_9 NI_9 NS_209 0 5.9438174500982210e-02
GC_9_210 b_9 NI_9 NS_210 0 -6.3780044320492071e-02
GC_9_211 b_9 NI_9 NS_211 0 -1.0218717795266404e-08
GC_9_212 b_9 NI_9 NS_212 0 -8.2100850940507151e-06
GC_9_213 b_9 NI_9 NS_213 0 -1.8519170180632131e-03
GC_9_214 b_9 NI_9 NS_214 0 -2.8731348100675467e-03
GC_9_215 b_9 NI_9 NS_215 0 -5.1084750342265655e-03
GC_9_216 b_9 NI_9 NS_216 0 1.9400105759025915e-03
GC_9_217 b_9 NI_9 NS_217 0 2.4463645136159331e-03
GC_9_218 b_9 NI_9 NS_218 0 -1.2255485306284367e-03
GC_9_219 b_9 NI_9 NS_219 0 -1.0650803114645691e-02
GC_9_220 b_9 NI_9 NS_220 0 1.1045727226969598e-03
GC_9_221 b_9 NI_9 NS_221 0 6.4145724032083854e-04
GC_9_222 b_9 NI_9 NS_222 0 1.7543134321693213e-03
GC_9_223 b_9 NI_9 NS_223 0 -9.5624731274385102e-04
GC_9_224 b_9 NI_9 NS_224 0 2.2871429574059395e-03
GC_9_225 b_9 NI_9 NS_225 0 5.9413402762514920e-04
GC_9_226 b_9 NI_9 NS_226 0 -5.8937211153621966e-03
GC_9_227 b_9 NI_9 NS_227 0 -8.5380903516811425e-03
GC_9_228 b_9 NI_9 NS_228 0 6.8906956142890646e-03
GC_9_229 b_9 NI_9 NS_229 0 2.5187079356760200e-03
GC_9_230 b_9 NI_9 NS_230 0 -3.6778727026020087e-03
GC_9_231 b_9 NI_9 NS_231 0 -2.6381597244180210e-03
GC_9_232 b_9 NI_9 NS_232 0 -5.1433843996302752e-04
GC_9_233 b_9 NI_9 NS_233 0 5.4575014107666929e-02
GC_9_234 b_9 NI_9 NS_234 0 1.6205591348719189e-03
GC_9_235 b_9 NI_9 NS_235 0 -4.9957335227356889e-02
GC_9_236 b_9 NI_9 NS_236 0 1.0966288254923440e-01
GC_9_237 b_9 NI_9 NS_237 0 1.0580850978741676e-08
GC_9_238 b_9 NI_9 NS_238 0 1.9882058041269511e-05
GC_9_239 b_9 NI_9 NS_239 0 -1.5752600624722560e-02
GC_9_240 b_9 NI_9 NS_240 0 2.4251911151477595e-02
GC_9_241 b_9 NI_9 NS_241 0 -7.8021574088024560e-03
GC_9_242 b_9 NI_9 NS_242 0 -1.4485548315517844e-02
GC_9_243 b_9 NI_9 NS_243 0 2.0432726147173751e-02
GC_9_244 b_9 NI_9 NS_244 0 6.6858618356341335e-03
GC_9_245 b_9 NI_9 NS_245 0 8.0641598453024040e-03
GC_9_246 b_9 NI_9 NS_246 0 4.3992228789321138e-02
GC_9_247 b_9 NI_9 NS_247 0 -1.1854720828864383e-02
GC_9_248 b_9 NI_9 NS_248 0 -3.2297431212269445e-03
GC_9_249 b_9 NI_9 NS_249 0 -5.0941020364672447e-03
GC_9_250 b_9 NI_9 NS_250 0 -4.0920246487202950e-03
GC_9_251 b_9 NI_9 NS_251 0 2.6818336758005375e-02
GC_9_252 b_9 NI_9 NS_252 0 -1.0400387337788498e-05
GC_9_253 b_9 NI_9 NS_253 0 3.3876594811035950e-02
GC_9_254 b_9 NI_9 NS_254 0 3.0995868422760524e-02
GC_9_255 b_9 NI_9 NS_255 0 -1.5641050364042747e-02
GC_9_256 b_9 NI_9 NS_256 0 8.2858690226329350e-03
GC_9_257 b_9 NI_9 NS_257 0 -9.9915577813659536e-04
GC_9_258 b_9 NI_9 NS_258 0 -6.8608391491022606e-03
GC_9_259 b_9 NI_9 NS_259 0 -6.8944292129345330e-02
GC_9_260 b_9 NI_9 NS_260 0 1.7522024121739486e-03
GC_9_261 b_9 NI_9 NS_261 0 -7.4976050247960438e-03
GC_9_262 b_9 NI_9 NS_262 0 5.4454474121713127e-03
GC_9_263 b_9 NI_9 NS_263 0 -8.2825504284356087e-10
GC_9_264 b_9 NI_9 NS_264 0 -1.6858110465050761e-06
GC_9_265 b_9 NI_9 NS_265 0 2.5528979621843376e-04
GC_9_266 b_9 NI_9 NS_266 0 2.6644770986489616e-03
GC_9_267 b_9 NI_9 NS_267 0 4.5291311737956433e-03
GC_9_268 b_9 NI_9 NS_268 0 -2.7565392768417228e-03
GC_9_269 b_9 NI_9 NS_269 0 -5.4227402040446125e-03
GC_9_270 b_9 NI_9 NS_270 0 4.2035093949704911e-04
GC_9_271 b_9 NI_9 NS_271 0 8.8583384359765191e-03
GC_9_272 b_9 NI_9 NS_272 0 -6.2088505594412493e-04
GC_9_273 b_9 NI_9 NS_273 0 -2.8261194604404182e-03
GC_9_274 b_9 NI_9 NS_274 0 -2.3963291279584442e-03
GC_9_275 b_9 NI_9 NS_275 0 4.3090299723284219e-05
GC_9_276 b_9 NI_9 NS_276 0 -2.1138831481322898e-03
GC_9_277 b_9 NI_9 NS_277 0 -3.5070906803346636e-03
GC_9_278 b_9 NI_9 NS_278 0 5.5495734927849313e-03
GC_9_279 b_9 NI_9 NS_279 0 5.0983691843059587e-03
GC_9_280 b_9 NI_9 NS_280 0 -7.7603767194391717e-03
GC_9_281 b_9 NI_9 NS_281 0 -5.0389546366635257e-03
GC_9_282 b_9 NI_9 NS_282 0 3.0962239743942493e-03
GC_9_283 b_9 NI_9 NS_283 0 2.2446188648831845e-03
GC_9_284 b_9 NI_9 NS_284 0 -1.6873558985848465e-03
GC_9_285 b_9 NI_9 NS_285 0 -5.9462060208454338e-03
GC_9_286 b_9 NI_9 NS_286 0 3.8165511269497212e-03
GC_9_287 b_9 NI_9 NS_287 0 -1.3746089080371303e-03
GC_9_288 b_9 NI_9 NS_288 0 2.3328708467421004e-03
GC_9_289 b_9 NI_9 NS_289 0 7.5881858999508210e-10
GC_9_290 b_9 NI_9 NS_290 0 6.0065829866922035e-07
GC_9_291 b_9 NI_9 NS_291 0 -1.9596140498731016e-04
GC_9_292 b_9 NI_9 NS_292 0 -4.5534341782619192e-04
GC_9_293 b_9 NI_9 NS_293 0 -1.0665939101090565e-03
GC_9_294 b_9 NI_9 NS_294 0 -9.2131959233472335e-04
GC_9_295 b_9 NI_9 NS_295 0 -2.3173790648370524e-03
GC_9_296 b_9 NI_9 NS_296 0 3.1223076785602495e-04
GC_9_297 b_9 NI_9 NS_297 0 -3.4634935108651368e-04
GC_9_298 b_9 NI_9 NS_298 0 4.1981837629813772e-03
GC_9_299 b_9 NI_9 NS_299 0 9.7829186500863943e-04
GC_9_300 b_9 NI_9 NS_300 0 4.4367013036742011e-04
GC_9_301 b_9 NI_9 NS_301 0 -3.7329483155213274e-04
GC_9_302 b_9 NI_9 NS_302 0 7.9843243359172943e-05
GC_9_303 b_9 NI_9 NS_303 0 -3.1453282997478016e-04
GC_9_304 b_9 NI_9 NS_304 0 3.3540654670163005e-03
GC_9_305 b_9 NI_9 NS_305 0 5.2329434371575180e-03
GC_9_306 b_9 NI_9 NS_306 0 8.1284473435285843e-04
GC_9_307 b_9 NI_9 NS_307 0 1.3427527634437227e-03
GC_9_308 b_9 NI_9 NS_308 0 -1.9440163306120872e-03
GC_9_309 b_9 NI_9 NS_309 0 -8.8256362515712393e-04
GC_9_310 b_9 NI_9 NS_310 0 -6.3689550758349700e-04
GC_9_311 b_9 NI_9 NS_311 0 -1.4735606988318204e-03
GC_9_312 b_9 NI_9 NS_312 0 2.5664403223774547e-03
GD_9_1 b_9 NI_9 NA_1 0 8.8774482025347023e-06
GD_9_2 b_9 NI_9 NA_2 0 7.7381918374771894e-06
GD_9_3 b_9 NI_9 NA_3 0 -5.5171969360454257e-06
GD_9_4 b_9 NI_9 NA_4 0 1.2646759611220681e-05
GD_9_5 b_9 NI_9 NA_5 0 1.6641036578223781e-04
GD_9_6 b_9 NI_9 NA_6 0 1.4009478068831448e-04
GD_9_7 b_9 NI_9 NA_7 0 3.0067015979806768e-03
GD_9_8 b_9 NI_9 NA_8 0 -5.3852870516734467e-05
GD_9_9 b_9 NI_9 NA_9 0 -2.9744132406365524e-02
GD_9_10 b_9 NI_9 NA_10 0 -2.0423329308840246e-02
GD_9_11 b_9 NI_9 NA_11 0 1.3427147738053148e-02
GD_9_12 b_9 NI_9 NA_12 0 -1.1219485718105334e-03
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 -2.4826037075934336e-05
GC_10_2 b_10 NI_10 NS_2 0 2.0783954904167742e-05
GC_10_3 b_10 NI_10 NS_3 0 -3.5006716145202000e-11
GC_10_4 b_10 NI_10 NS_4 0 -2.7090146222543380e-10
GC_10_5 b_10 NI_10 NS_5 0 1.6166640647054870e-06
GC_10_6 b_10 NI_10 NS_6 0 1.4393720474517962e-06
GC_10_7 b_10 NI_10 NS_7 0 2.5870845097806143e-07
GC_10_8 b_10 NI_10 NS_8 0 3.7190211864472098e-07
GC_10_9 b_10 NI_10 NS_9 0 1.7411259490500930e-06
GC_10_10 b_10 NI_10 NS_10 0 -2.0416395007247797e-07
GC_10_11 b_10 NI_10 NS_11 0 3.3661779716103820e-06
GC_10_12 b_10 NI_10 NS_12 0 -1.0270838020369747e-06
GC_10_13 b_10 NI_10 NS_13 0 4.2256042203256025e-07
GC_10_14 b_10 NI_10 NS_14 0 5.0171846016213856e-08
GC_10_15 b_10 NI_10 NS_15 0 2.5403837189028662e-07
GC_10_16 b_10 NI_10 NS_16 0 -2.9663372563991967e-07
GC_10_17 b_10 NI_10 NS_17 0 1.0840317650617250e-06
GC_10_18 b_10 NI_10 NS_18 0 -1.0041276965004177e-06
GC_10_19 b_10 NI_10 NS_19 0 1.6348101783968348e-06
GC_10_20 b_10 NI_10 NS_20 0 -1.2123858302711978e-06
GC_10_21 b_10 NI_10 NS_21 0 -5.8100883767638879e-08
GC_10_22 b_10 NI_10 NS_22 0 1.3019076199981360e-06
GC_10_23 b_10 NI_10 NS_23 0 3.3328567064268641e-07
GC_10_24 b_10 NI_10 NS_24 0 6.8675688990575883e-07
GC_10_25 b_10 NI_10 NS_25 0 -1.6980997934209409e-05
GC_10_26 b_10 NI_10 NS_26 0 -1.3435244436664302e-06
GC_10_27 b_10 NI_10 NS_27 0 -2.7914673503538703e-05
GC_10_28 b_10 NI_10 NS_28 0 4.2480930506973719e-05
GC_10_29 b_10 NI_10 NS_29 0 3.6704872886122803e-11
GC_10_30 b_10 NI_10 NS_30 0 -2.7830063985858140e-10
GC_10_31 b_10 NI_10 NS_31 0 8.4367571393639816e-07
GC_10_32 b_10 NI_10 NS_32 0 4.8587722432010174e-07
GC_10_33 b_10 NI_10 NS_33 0 4.0290827303665512e-07
GC_10_34 b_10 NI_10 NS_34 0 -7.5371184182549380e-07
GC_10_35 b_10 NI_10 NS_35 0 -4.7578259270368927e-07
GC_10_36 b_10 NI_10 NS_36 0 9.9272453165939375e-07
GC_10_37 b_10 NI_10 NS_37 0 1.4092607393600989e-06
GC_10_38 b_10 NI_10 NS_38 0 1.8306204235572403e-07
GC_10_39 b_10 NI_10 NS_39 0 -4.2142649185272873e-07
GC_10_40 b_10 NI_10 NS_40 0 9.6875597104670624e-07
GC_10_41 b_10 NI_10 NS_41 0 5.7216894530404513e-07
GC_10_42 b_10 NI_10 NS_42 0 3.8282397747621660e-07
GC_10_43 b_10 NI_10 NS_43 0 5.5915977172539907e-07
GC_10_44 b_10 NI_10 NS_44 0 3.2458443800314024e-06
GC_10_45 b_10 NI_10 NS_45 0 4.0017169622802075e-06
GC_10_46 b_10 NI_10 NS_46 0 7.8432540845401400e-07
GC_10_47 b_10 NI_10 NS_47 0 9.0407612707941629e-07
GC_10_48 b_10 NI_10 NS_48 0 2.3922783460478133e-06
GC_10_49 b_10 NI_10 NS_49 0 1.1489417131207028e-06
GC_10_50 b_10 NI_10 NS_50 0 2.6151367956788612e-06
GC_10_51 b_10 NI_10 NS_51 0 -3.3615792955377090e-05
GC_10_52 b_10 NI_10 NS_52 0 4.1019978778532906e-07
GC_10_53 b_10 NI_10 NS_53 0 -2.7846429771757052e-05
GC_10_54 b_10 NI_10 NS_54 0 -1.1271766206249247e-06
GC_10_55 b_10 NI_10 NS_55 0 -5.6801602037097494e-11
GC_10_56 b_10 NI_10 NS_56 0 1.0421525253437477e-09
GC_10_57 b_10 NI_10 NS_57 0 3.7467178472331476e-06
GC_10_58 b_10 NI_10 NS_58 0 4.4128221556255503e-06
GC_10_59 b_10 NI_10 NS_59 0 3.3691629041667820e-06
GC_10_60 b_10 NI_10 NS_60 0 3.3616308532012670e-06
GC_10_61 b_10 NI_10 NS_61 0 1.0412998947686062e-05
GC_10_62 b_10 NI_10 NS_62 0 -2.9646622272336261e-06
GC_10_63 b_10 NI_10 NS_63 0 6.6233918688102596e-06
GC_10_64 b_10 NI_10 NS_64 0 -1.4577523588194197e-05
GC_10_65 b_10 NI_10 NS_65 0 -3.0131491718583588e-06
GC_10_66 b_10 NI_10 NS_66 0 -1.0905306749877885e-06
GC_10_67 b_10 NI_10 NS_67 0 9.4683070721502279e-07
GC_10_68 b_10 NI_10 NS_68 0 -8.3289928909491212e-07
GC_10_69 b_10 NI_10 NS_69 0 2.9441076171736370e-06
GC_10_70 b_10 NI_10 NS_70 0 -1.2938321250661405e-05
GC_10_71 b_10 NI_10 NS_71 0 -1.3694224907280689e-05
GC_10_72 b_10 NI_10 NS_72 0 -3.7760567192249914e-06
GC_10_73 b_10 NI_10 NS_73 0 -3.5424630949320633e-06
GC_10_74 b_10 NI_10 NS_74 0 5.8948709086331775e-06
GC_10_75 b_10 NI_10 NS_75 0 2.7008062273237545e-06
GC_10_76 b_10 NI_10 NS_76 0 1.1398778705268446e-06
GC_10_77 b_10 NI_10 NS_77 0 1.6185539141399628e-07
GC_10_78 b_10 NI_10 NS_78 0 -5.8089500386629109e-06
GC_10_79 b_10 NI_10 NS_79 0 -6.5847609936882730e-06
GC_10_80 b_10 NI_10 NS_80 0 9.9213322487484064e-05
GC_10_81 b_10 NI_10 NS_81 0 6.2415130812325453e-11
GC_10_82 b_10 NI_10 NS_82 0 -2.6617588604870679e-09
GC_10_83 b_10 NI_10 NS_83 0 -1.4903987545883219e-06
GC_10_84 b_10 NI_10 NS_84 0 -1.5556252031771703e-06
GC_10_85 b_10 NI_10 NS_85 0 -2.8329164322282960e-06
GC_10_86 b_10 NI_10 NS_86 0 -1.5878871419688042e-06
GC_10_87 b_10 NI_10 NS_87 0 -5.7178315325385344e-06
GC_10_88 b_10 NI_10 NS_88 0 -1.2614686893842145e-06
GC_10_89 b_10 NI_10 NS_89 0 -8.7595715638538128e-06
GC_10_90 b_10 NI_10 NS_90 0 6.4067723149840816e-06
GC_10_91 b_10 NI_10 NS_91 0 -6.4092262017494328e-06
GC_10_92 b_10 NI_10 NS_92 0 5.1019634314827991e-06
GC_10_93 b_10 NI_10 NS_93 0 8.4424844664790300e-07
GC_10_94 b_10 NI_10 NS_94 0 5.8470280732011489e-06
GC_10_95 b_10 NI_10 NS_95 0 -5.3961664823685020e-06
GC_10_96 b_10 NI_10 NS_96 0 1.2705485600613561e-05
GC_10_97 b_10 NI_10 NS_97 0 1.0828082346797669e-05
GC_10_98 b_10 NI_10 NS_98 0 1.5435688432917414e-05
GC_10_99 b_10 NI_10 NS_99 0 4.5989180199088617e-06
GC_10_100 b_10 NI_10 NS_100 0 1.0589226678132116e-05
GC_10_101 b_10 NI_10 NS_101 0 4.7903817381849534e-06
GC_10_102 b_10 NI_10 NS_102 0 9.9605560025077804e-06
GC_10_103 b_10 NI_10 NS_103 0 -7.2520431138663606e-05
GC_10_104 b_10 NI_10 NS_104 0 1.2870702746351485e-05
GC_10_105 b_10 NI_10 NS_105 0 1.2824310917558922e-04
GC_10_106 b_10 NI_10 NS_106 0 5.5587852479288083e-05
GC_10_107 b_10 NI_10 NS_107 0 -4.2209257118022369e-10
GC_10_108 b_10 NI_10 NS_108 0 4.4721715130756648e-08
GC_10_109 b_10 NI_10 NS_109 0 5.7603062221437970e-06
GC_10_110 b_10 NI_10 NS_110 0 7.6124133529409987e-05
GC_10_111 b_10 NI_10 NS_111 0 1.5376831893820862e-04
GC_10_112 b_10 NI_10 NS_112 0 1.3563455013548839e-04
GC_10_113 b_10 NI_10 NS_113 0 3.4707338886461872e-04
GC_10_114 b_10 NI_10 NS_114 0 -2.4008417156469861e-05
GC_10_115 b_10 NI_10 NS_115 0 5.3250879683860037e-05
GC_10_116 b_10 NI_10 NS_116 0 -5.8494622534182997e-04
GC_10_117 b_10 NI_10 NS_117 0 -1.4501227604991833e-04
GC_10_118 b_10 NI_10 NS_118 0 -6.8323072577714580e-05
GC_10_119 b_10 NI_10 NS_119 0 5.2206313148536705e-05
GC_10_120 b_10 NI_10 NS_120 0 -1.0707558084672238e-05
GC_10_121 b_10 NI_10 NS_121 0 4.8324829654605725e-05
GC_10_122 b_10 NI_10 NS_122 0 -4.5206759616783396e-04
GC_10_123 b_10 NI_10 NS_123 0 -7.0671486017394205e-04
GC_10_124 b_10 NI_10 NS_124 0 -8.3346071169656592e-05
GC_10_125 b_10 NI_10 NS_125 0 -1.7415349030986850e-04
GC_10_126 b_10 NI_10 NS_126 0 2.5972205241186233e-04
GC_10_127 b_10 NI_10 NS_127 0 1.0227100322312986e-04
GC_10_128 b_10 NI_10 NS_128 0 8.1142072008156833e-05
GC_10_129 b_10 NI_10 NS_129 0 -1.2306696817145812e-04
GC_10_130 b_10 NI_10 NS_130 0 -3.3447060411824920e-04
GC_10_131 b_10 NI_10 NS_131 0 3.8620814640400852e-04
GC_10_132 b_10 NI_10 NS_132 0 -2.0252878404763111e-03
GC_10_133 b_10 NI_10 NS_133 0 4.0260186039709338e-10
GC_10_134 b_10 NI_10 NS_134 0 -2.6893743210117818e-08
GC_10_135 b_10 NI_10 NS_135 0 1.8850642810153096e-05
GC_10_136 b_10 NI_10 NS_136 0 4.3631168195547953e-05
GC_10_137 b_10 NI_10 NS_137 0 8.2151685482455066e-05
GC_10_138 b_10 NI_10 NS_138 0 -3.0666300397258061e-05
GC_10_139 b_10 NI_10 NS_139 0 -1.3460177720490712e-05
GC_10_140 b_10 NI_10 NS_140 0 1.3808944495887105e-05
GC_10_141 b_10 NI_10 NS_141 0 1.9797123510814914e-04
GC_10_142 b_10 NI_10 NS_142 0 -9.9099563376684382e-05
GC_10_143 b_10 NI_10 NS_143 0 2.7210975526635565e-05
GC_10_144 b_10 NI_10 NS_144 0 -9.8085102577170452e-05
GC_10_145 b_10 NI_10 NS_145 0 -1.7289683466273591e-05
GC_10_146 b_10 NI_10 NS_146 0 -9.8313649014516235e-05
GC_10_147 b_10 NI_10 NS_147 0 1.0597728133220182e-05
GC_10_148 b_10 NI_10 NS_148 0 -9.7356896454588819e-05
GC_10_149 b_10 NI_10 NS_149 0 -9.7278143526596152e-05
GC_10_150 b_10 NI_10 NS_150 0 -3.1575652896329248e-04
GC_10_151 b_10 NI_10 NS_151 0 -1.3369272192560155e-04
GC_10_152 b_10 NI_10 NS_152 0 -1.1532242291810430e-04
GC_10_153 b_10 NI_10 NS_153 0 -1.9101665375565842e-05
GC_10_154 b_10 NI_10 NS_154 0 -1.9122446510101687e-04
GC_10_155 b_10 NI_10 NS_155 0 1.5286795588133895e-03
GC_10_156 b_10 NI_10 NS_156 0 -9.9338064924617159e-05
GC_10_157 b_10 NI_10 NS_157 0 -1.0983047129905286e-03
GC_10_158 b_10 NI_10 NS_158 0 1.9215778666370293e-03
GC_10_159 b_10 NI_10 NS_159 0 -1.0012200748424698e-10
GC_10_160 b_10 NI_10 NS_160 0 2.7261165828906014e-07
GC_10_161 b_10 NI_10 NS_161 0 5.8917471633448603e-05
GC_10_162 b_10 NI_10 NS_162 0 -8.7105571923830832e-05
GC_10_163 b_10 NI_10 NS_163 0 -2.6162502034395929e-04
GC_10_164 b_10 NI_10 NS_164 0 -1.7081949783936766e-04
GC_10_165 b_10 NI_10 NS_165 0 -5.2947831522617730e-04
GC_10_166 b_10 NI_10 NS_166 0 2.5272762972283214e-05
GC_10_167 b_10 NI_10 NS_167 0 4.2373175763682535e-05
GC_10_168 b_10 NI_10 NS_168 0 9.1566637864842553e-04
GC_10_169 b_10 NI_10 NS_169 0 2.4558524257576648e-04
GC_10_170 b_10 NI_10 NS_170 0 1.3066484562038755e-04
GC_10_171 b_10 NI_10 NS_171 0 -8.1510649852482004e-05
GC_10_172 b_10 NI_10 NS_172 0 2.6833725231839720e-05
GC_10_173 b_10 NI_10 NS_173 0 -7.0978324456389365e-05
GC_10_174 b_10 NI_10 NS_174 0 7.5353511188094142e-04
GC_10_175 b_10 NI_10 NS_175 0 1.2757395617001297e-03
GC_10_176 b_10 NI_10 NS_176 0 1.3789245743877046e-04
GC_10_177 b_10 NI_10 NS_177 0 3.2405502347661894e-04
GC_10_178 b_10 NI_10 NS_178 0 -4.2274714510477109e-04
GC_10_179 b_10 NI_10 NS_179 0 -2.4522716600903496e-04
GC_10_180 b_10 NI_10 NS_180 0 -1.0940685466369367e-04
GC_10_181 b_10 NI_10 NS_181 0 -1.5442371361053505e-03
GC_10_182 b_10 NI_10 NS_182 0 3.7328710149219521e-04
GC_10_183 b_10 NI_10 NS_183 0 -1.2147766846229674e-03
GC_10_184 b_10 NI_10 NS_184 0 5.5868900144230571e-04
GC_10_185 b_10 NI_10 NS_185 0 3.0016424138339034e-10
GC_10_186 b_10 NI_10 NS_186 0 -5.7498731504946888e-07
GC_10_187 b_10 NI_10 NS_187 0 3.1227428539180193e-05
GC_10_188 b_10 NI_10 NS_188 0 6.3819814794280902e-04
GC_10_189 b_10 NI_10 NS_189 0 1.0888451722179020e-03
GC_10_190 b_10 NI_10 NS_190 0 -6.7567693432021598e-04
GC_10_191 b_10 NI_10 NS_191 0 -1.3740906963046222e-03
GC_10_192 b_10 NI_10 NS_192 0 7.5344570729055232e-05
GC_10_193 b_10 NI_10 NS_193 0 2.0944073047835798e-03
GC_10_194 b_10 NI_10 NS_194 0 -1.0659929531357928e-04
GC_10_195 b_10 NI_10 NS_195 0 -7.3376592624205240e-04
GC_10_196 b_10 NI_10 NS_196 0 -5.7284925314569771e-04
GC_10_197 b_10 NI_10 NS_197 0 5.7948715315435287e-06
GC_10_198 b_10 NI_10 NS_198 0 -4.8780379407593579e-04
GC_10_199 b_10 NI_10 NS_199 0 -9.0574312806516804e-04
GC_10_200 b_10 NI_10 NS_200 0 1.3911734445058621e-03
GC_10_201 b_10 NI_10 NS_201 0 1.2475487313940486e-03
GC_10_202 b_10 NI_10 NS_202 0 -1.8368924178396675e-03
GC_10_203 b_10 NI_10 NS_203 0 -1.2247766869372780e-03
GC_10_204 b_10 NI_10 NS_204 0 7.8190148077005321e-04
GC_10_205 b_10 NI_10 NS_205 0 5.7537113226200775e-04
GC_10_206 b_10 NI_10 NS_206 0 -4.1171102859299336e-04
GC_10_207 b_10 NI_10 NS_207 0 -7.3681761651263149e-04
GC_10_208 b_10 NI_10 NS_208 0 1.1397080063322229e-03
GC_10_209 b_10 NI_10 NS_209 0 -4.9957157009269768e-02
GC_10_210 b_10 NI_10 NS_210 0 1.0966274658728527e-01
GC_10_211 b_10 NI_10 NS_211 0 1.0580846965555003e-08
GC_10_212 b_10 NI_10 NS_212 0 1.9882056793241710e-05
GC_10_213 b_10 NI_10 NS_213 0 -1.5752613758823357e-02
GC_10_214 b_10 NI_10 NS_214 0 2.4251930397095497e-02
GC_10_215 b_10 NI_10 NS_215 0 -7.8021495503761990e-03
GC_10_216 b_10 NI_10 NS_216 0 -1.4485564272828677e-02
GC_10_217 b_10 NI_10 NS_217 0 2.0432739291833445e-02
GC_10_218 b_10 NI_10 NS_218 0 6.6858498285347579e-03
GC_10_219 b_10 NI_10 NS_219 0 8.0641272309114817e-03
GC_10_220 b_10 NI_10 NS_220 0 4.3992236373296592e-02
GC_10_221 b_10 NI_10 NS_221 0 -1.1854727393366951e-02
GC_10_222 b_10 NI_10 NS_222 0 -3.2297409055207257e-03
GC_10_223 b_10 NI_10 NS_223 0 -5.0941021446472522e-03
GC_10_224 b_10 NI_10 NS_224 0 -4.0920283263967076e-03
GC_10_225 b_10 NI_10 NS_225 0 2.6818332759259156e-02
GC_10_226 b_10 NI_10 NS_226 0 -1.0405901739955536e-05
GC_10_227 b_10 NI_10 NS_227 0 3.3876574607631861e-02
GC_10_228 b_10 NI_10 NS_228 0 3.0995868061728403e-02
GC_10_229 b_10 NI_10 NS_229 0 -1.5641056192866147e-02
GC_10_230 b_10 NI_10 NS_230 0 8.2858669010746760e-03
GC_10_231 b_10 NI_10 NS_231 0 -9.9915869430774692e-04
GC_10_232 b_10 NI_10 NS_232 0 -6.8608480926139722e-03
GC_10_233 b_10 NI_10 NS_233 0 -6.8944187882407859e-02
GC_10_234 b_10 NI_10 NS_234 0 1.7521962529281172e-03
GC_10_235 b_10 NI_10 NS_235 0 5.9438174500982294e-02
GC_10_236 b_10 NI_10 NS_236 0 -6.3780044320491919e-02
GC_10_237 b_10 NI_10 NS_237 0 -1.0218717795266189e-08
GC_10_238 b_10 NI_10 NS_238 0 -8.2100850940506508e-06
GC_10_239 b_10 NI_10 NS_239 0 -1.8519170180632102e-03
GC_10_240 b_10 NI_10 NS_240 0 -2.8731348100675467e-03
GC_10_241 b_10 NI_10 NS_241 0 -5.1084750342265655e-03
GC_10_242 b_10 NI_10 NS_242 0 1.9400105759025902e-03
GC_10_243 b_10 NI_10 NS_243 0 2.4463645136159331e-03
GC_10_244 b_10 NI_10 NS_244 0 -1.2255485306284385e-03
GC_10_245 b_10 NI_10 NS_245 0 -1.0650803114645694e-02
GC_10_246 b_10 NI_10 NS_246 0 1.1045727226969614e-03
GC_10_247 b_10 NI_10 NS_247 0 6.4145724032083822e-04
GC_10_248 b_10 NI_10 NS_248 0 1.7543134321693218e-03
GC_10_249 b_10 NI_10 NS_249 0 -9.5624731274385135e-04
GC_10_250 b_10 NI_10 NS_250 0 2.2871429574059425e-03
GC_10_251 b_10 NI_10 NS_251 0 5.9413402762514670e-04
GC_10_252 b_10 NI_10 NS_252 0 -5.8937211153621931e-03
GC_10_253 b_10 NI_10 NS_253 0 -8.5380903516811390e-03
GC_10_254 b_10 NI_10 NS_254 0 6.8906956142890724e-03
GC_10_255 b_10 NI_10 NS_255 0 2.5187079356760234e-03
GC_10_256 b_10 NI_10 NS_256 0 -3.6778727026020031e-03
GC_10_257 b_10 NI_10 NS_257 0 -2.6381597244180223e-03
GC_10_258 b_10 NI_10 NS_258 0 -5.1433843996302091e-04
GC_10_259 b_10 NI_10 NS_259 0 5.4575014107666804e-02
GC_10_260 b_10 NI_10 NS_260 0 1.6205591348719070e-03
GC_10_261 b_10 NI_10 NS_261 0 -1.3745905451381098e-03
GC_10_262 b_10 NI_10 NS_262 0 2.3328751956352952e-03
GC_10_263 b_10 NI_10 NS_263 0 7.5881886160042663e-10
GC_10_264 b_10 NI_10 NS_264 0 6.0065828798477989e-07
GC_10_265 b_10 NI_10 NS_265 0 -1.9596046860603485e-04
GC_10_266 b_10 NI_10 NS_266 0 -4.5533533220927275e-04
GC_10_267 b_10 NI_10 NS_267 0 -1.0665948721612427e-03
GC_10_268 b_10 NI_10 NS_268 0 -9.2132735416159783e-04
GC_10_269 b_10 NI_10 NS_269 0 -2.3173774124387470e-03
GC_10_270 b_10 NI_10 NS_270 0 3.1222384568039511e-04
GC_10_271 b_10 NI_10 NS_271 0 -3.4635675297816325e-04
GC_10_272 b_10 NI_10 NS_272 0 4.1981926069968182e-03
GC_10_273 b_10 NI_10 NS_273 0 9.7829070586936224e-04
GC_10_274 b_10 NI_10 NS_274 0 4.4367255478046770e-04
GC_10_275 b_10 NI_10 NS_275 0 -3.7329590593141105e-04
GC_10_276 b_10 NI_10 NS_276 0 7.9841939005989728e-05
GC_10_277 b_10 NI_10 NS_277 0 -3.1453628485497969e-04
GC_10_278 b_10 NI_10 NS_278 0 3.3540664095542553e-03
GC_10_279 b_10 NI_10 NS_279 0 5.2329467711993158e-03
GC_10_280 b_10 NI_10 NS_280 0 8.1285316902855796e-04
GC_10_281 b_10 NI_10 NS_281 0 1.3427552736417615e-03
GC_10_282 b_10 NI_10 NS_282 0 -1.9440156821573179e-03
GC_10_283 b_10 NI_10 NS_283 0 -8.8256278729533140e-04
GC_10_284 b_10 NI_10 NS_284 0 -6.3689652085268560e-04
GC_10_285 b_10 NI_10 NS_285 0 -1.4735645022307153e-03
GC_10_286 b_10 NI_10 NS_286 0 2.5664394616210116e-03
GC_10_287 b_10 NI_10 NS_287 0 -7.4986728019016870e-03
GC_10_288 b_10 NI_10 NS_288 0 5.4463736044302220e-03
GC_10_289 b_10 NI_10 NS_289 0 -8.2819008874232171e-10
GC_10_290 b_10 NI_10 NS_290 0 -1.6858209024942455e-06
GC_10_291 b_10 NI_10 NS_291 0 2.5534683118825325e-04
GC_10_292 b_10 NI_10 NS_292 0 2.6645211981117570e-03
GC_10_293 b_10 NI_10 NS_293 0 4.5291691759910642e-03
GC_10_294 b_10 NI_10 NS_294 0 -2.7565572830191920e-03
GC_10_295 b_10 NI_10 NS_295 0 -5.4227010287392187e-03
GC_10_296 b_10 NI_10 NS_296 0 4.2041651361554062e-04
GC_10_297 b_10 NI_10 NS_297 0 8.8584610087896268e-03
GC_10_298 b_10 NI_10 NS_298 0 -6.2094131486168324e-04
GC_10_299 b_10 NI_10 NS_299 0 -2.8260900937832020e-03
GC_10_300 b_10 NI_10 NS_300 0 -2.3963195077242277e-03
GC_10_301 b_10 NI_10 NS_301 0 4.3105060396030606e-05
GC_10_302 b_10 NI_10 NS_302 0 -2.1139049464674025e-03
GC_10_303 b_10 NI_10 NS_303 0 -3.5070302768425671e-03
GC_10_304 b_10 NI_10 NS_304 0 5.5496268167169226e-03
GC_10_305 b_10 NI_10 NS_305 0 5.0984923970970753e-03
GC_10_306 b_10 NI_10 NS_306 0 -7.7604205411807804e-03
GC_10_307 b_10 NI_10 NS_307 0 -5.0389100498201347e-03
GC_10_308 b_10 NI_10 NS_308 0 3.0962157420722351e-03
GC_10_309 b_10 NI_10 NS_309 0 2.2446243261625932e-03
GC_10_310 b_10 NI_10 NS_310 0 -1.6873400590580396e-03
GC_10_311 b_10 NI_10 NS_311 0 -5.9469814837945093e-03
GC_10_312 b_10 NI_10 NS_312 0 3.8164576042803576e-03
GD_10_1 b_10 NI_10 NA_1 0 7.7385923302773625e-06
GD_10_2 b_10 NI_10 NA_2 0 8.9269178903577362e-06
GD_10_3 b_10 NI_10 NA_3 0 1.2667334859890936e-05
GD_10_4 b_10 NI_10 NA_4 0 -5.5170915967900383e-06
GD_10_5 b_10 NI_10 NA_5 0 1.4009512909082065e-04
GD_10_6 b_10 NI_10 NA_6 0 1.6640052708753871e-04
GD_10_7 b_10 NI_10 NA_7 0 -5.3787251821943267e-05
GD_10_8 b_10 NI_10 NA_8 0 3.0067237937127594e-03
GD_10_9 b_10 NI_10 NA_9 0 -2.0423393897813610e-02
GD_10_10 b_10 NI_10 NA_10 0 -2.9744132406365822e-02
GD_10_11 b_10 NI_10 NA_11 0 -1.1219599193645952e-03
GD_10_12 b_10 NI_10 NA_12 0 1.3427306305630196e-02
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 -3.5487272118791538e-05
GC_11_2 b_11 NI_11 NS_2 0 4.3755697548911845e-05
GC_11_3 b_11 NI_11 NS_3 0 3.2703458169589655e-11
GC_11_4 b_11 NI_11 NS_4 0 -2.6824612755362823e-10
GC_11_5 b_11 NI_11 NS_5 0 1.0320798086996838e-06
GC_11_6 b_11 NI_11 NS_6 0 1.0605759765109829e-06
GC_11_7 b_11 NI_11 NS_7 0 1.7241328069064181e-06
GC_11_8 b_11 NI_11 NS_8 0 2.5964993302961068e-07
GC_11_9 b_11 NI_11 NS_9 0 1.0932120348244174e-06
GC_11_10 b_11 NI_11 NS_10 0 4.6059962957482023e-07
GC_11_11 b_11 NI_11 NS_11 0 2.9262620813076854e-06
GC_11_12 b_11 NI_11 NS_12 0 -4.3423343455232166e-07
GC_11_13 b_11 NI_11 NS_13 0 1.0132358973283233e-06
GC_11_14 b_11 NI_11 NS_14 0 5.3045095197681734e-09
GC_11_15 b_11 NI_11 NS_15 0 5.6285416852712747e-07
GC_11_16 b_11 NI_11 NS_16 0 -5.1625010430550455e-07
GC_11_17 b_11 NI_11 NS_17 0 1.6607436160140879e-06
GC_11_18 b_11 NI_11 NS_18 0 1.2910028624499153e-06
GC_11_19 b_11 NI_11 NS_19 0 2.8544592743976204e-06
GC_11_20 b_11 NI_11 NS_20 0 -1.2126697849448984e-06
GC_11_21 b_11 NI_11 NS_21 0 5.5986035005755069e-07
GC_11_22 b_11 NI_11 NS_22 0 1.1266008068719638e-06
GC_11_23 b_11 NI_11 NS_23 0 3.9045698306902999e-07
GC_11_24 b_11 NI_11 NS_24 0 1.5530721039942667e-06
GC_11_25 b_11 NI_11 NS_25 0 -3.6623119920681246e-05
GC_11_26 b_11 NI_11 NS_26 0 -3.7034613793420238e-06
GC_11_27 b_11 NI_11 NS_27 0 -1.1812995353083849e-05
GC_11_28 b_11 NI_11 NS_28 0 -5.5505897429587533e-06
GC_11_29 b_11 NI_11 NS_29 0 -3.0498032305890395e-11
GC_11_30 b_11 NI_11 NS_30 0 -1.3578568612893242e-10
GC_11_31 b_11 NI_11 NS_31 0 2.2976201026816278e-06
GC_11_32 b_11 NI_11 NS_32 0 1.7808637747388546e-06
GC_11_33 b_11 NI_11 NS_33 0 -6.4157914550578336e-07
GC_11_34 b_11 NI_11 NS_34 0 -3.8592716755342714e-07
GC_11_35 b_11 NI_11 NS_35 0 1.5505335309380986e-06
GC_11_36 b_11 NI_11 NS_36 0 -1.1518042436362913e-06
GC_11_37 b_11 NI_11 NS_37 0 1.8453794300833869e-06
GC_11_38 b_11 NI_11 NS_38 0 -4.3341854551171949e-07
GC_11_39 b_11 NI_11 NS_39 0 1.1932615206241478e-07
GC_11_40 b_11 NI_11 NS_40 0 -1.8767499590490944e-07
GC_11_41 b_11 NI_11 NS_41 0 5.5237171778032610e-08
GC_11_42 b_11 NI_11 NS_42 0 -3.1791035723000316e-07
GC_11_43 b_11 NI_11 NS_43 0 4.3573530828375422e-07
GC_11_44 b_11 NI_11 NS_44 0 -7.3740235922405811e-07
GC_11_45 b_11 NI_11 NS_45 0 9.1579257701023676e-07
GC_11_46 b_11 NI_11 NS_46 0 -1.3980117412017951e-06
GC_11_47 b_11 NI_11 NS_47 0 -1.8989911287167984e-07
GC_11_48 b_11 NI_11 NS_48 0 5.9848222640797466e-07
GC_11_49 b_11 NI_11 NS_49 0 3.5032407144180114e-07
GC_11_50 b_11 NI_11 NS_50 0 -1.4440491770217840e-08
GC_11_51 b_11 NI_11 NS_51 0 5.7887410294409160e-06
GC_11_52 b_11 NI_11 NS_52 0 2.3957892099664491e-06
GC_11_53 b_11 NI_11 NS_53 0 -2.7887634369773307e-05
GC_11_54 b_11 NI_11 NS_54 0 4.2423618403911843e-05
GC_11_55 b_11 NI_11 NS_55 0 3.6713789341458320e-11
GC_11_56 b_11 NI_11 NS_56 0 -2.8057047226726072e-10
GC_11_57 b_11 NI_11 NS_57 0 8.4282344369351079e-07
GC_11_58 b_11 NI_11 NS_58 0 4.8528865757814962e-07
GC_11_59 b_11 NI_11 NS_59 0 4.0300514981681646e-07
GC_11_60 b_11 NI_11 NS_60 0 -7.5313821367140634e-07
GC_11_61 b_11 NI_11 NS_61 0 -4.7580779673088141e-07
GC_11_62 b_11 NI_11 NS_62 0 9.9091370053516267e-07
GC_11_63 b_11 NI_11 NS_63 0 1.4076893618144319e-06
GC_11_64 b_11 NI_11 NS_64 0 1.8309238647855173e-07
GC_11_65 b_11 NI_11 NS_65 0 -4.2172397997824648e-07
GC_11_66 b_11 NI_11 NS_66 0 9.6747371775648502e-07
GC_11_67 b_11 NI_11 NS_67 0 5.7161785158921943e-07
GC_11_68 b_11 NI_11 NS_68 0 3.8276272405044288e-07
GC_11_69 b_11 NI_11 NS_69 0 5.5777862401169323e-07
GC_11_70 b_11 NI_11 NS_70 0 3.2436841224742264e-06
GC_11_71 b_11 NI_11 NS_71 0 3.9996423812253922e-06
GC_11_72 b_11 NI_11 NS_72 0 7.8349358484028772e-07
GC_11_73 b_11 NI_11 NS_73 0 9.0316508682121874e-07
GC_11_74 b_11 NI_11 NS_74 0 2.3897395456446958e-06
GC_11_75 b_11 NI_11 NS_75 0 1.1491002713746738e-06
GC_11_76 b_11 NI_11 NS_76 0 2.6121087675904197e-06
GC_11_77 b_11 NI_11 NS_77 0 -3.3569341302838053e-05
GC_11_78 b_11 NI_11 NS_78 0 4.1045948020516811e-07
GC_11_79 b_11 NI_11 NS_79 0 -2.4857671230368115e-05
GC_11_80 b_11 NI_11 NS_80 0 2.0849043296820922e-05
GC_11_81 b_11 NI_11 NS_81 0 -3.5016448676964662e-11
GC_11_82 b_11 NI_11 NS_82 0 -2.6866770601366137e-10
GC_11_83 b_11 NI_11 NS_83 0 1.6181043321283270e-06
GC_11_84 b_11 NI_11 NS_84 0 1.4408616037561001e-06
GC_11_85 b_11 NI_11 NS_85 0 2.6029540698287562e-07
GC_11_86 b_11 NI_11 NS_86 0 3.7175586398012264e-07
GC_11_87 b_11 NI_11 NS_87 0 1.7426638823205763e-06
GC_11_88 b_11 NI_11 NS_88 0 -2.0560495061497625e-07
GC_11_89 b_11 NI_11 NS_89 0 3.3661173197982537e-06
GC_11_90 b_11 NI_11 NS_90 0 -1.0275561830523912e-06
GC_11_91 b_11 NI_11 NS_91 0 4.2278216623601885e-07
GC_11_92 b_11 NI_11 NS_92 0 5.1394840273672097e-08
GC_11_93 b_11 NI_11 NS_93 0 2.5478033210834520e-07
GC_11_94 b_11 NI_11 NS_94 0 -2.9686669741970702e-07
GC_11_95 b_11 NI_11 NS_95 0 1.0838533425271015e-06
GC_11_96 b_11 NI_11 NS_96 0 -1.0037664201181465e-06
GC_11_97 b_11 NI_11 NS_97 0 1.6365251103874489e-06
GC_11_98 b_11 NI_11 NS_98 0 -1.2094851648296976e-06
GC_11_99 b_11 NI_11 NS_99 0 -5.6831706249236157e-08
GC_11_100 b_11 NI_11 NS_100 0 1.3046586127802238e-06
GC_11_101 b_11 NI_11 NS_101 0 3.3320738282436543e-07
GC_11_102 b_11 NI_11 NS_102 0 6.8983872815124084e-07
GC_11_103 b_11 NI_11 NS_103 0 -1.7034658179480959e-05
GC_11_104 b_11 NI_11 NS_104 0 -1.3465976607043752e-06
GC_11_105 b_11 NI_11 NS_105 0 -1.4269275345295108e-04
GC_11_106 b_11 NI_11 NS_106 0 6.6397301983326317e-04
GC_11_107 b_11 NI_11 NS_107 0 1.2463080421614215e-10
GC_11_108 b_11 NI_11 NS_108 0 -1.1464438668294725e-08
GC_11_109 b_11 NI_11 NS_109 0 -4.0106801629813447e-06
GC_11_110 b_11 NI_11 NS_110 0 -3.9979564519983141e-06
GC_11_111 b_11 NI_11 NS_111 0 -9.6094390415244721e-06
GC_11_112 b_11 NI_11 NS_112 0 -3.7334837100273836e-06
GC_11_113 b_11 NI_11 NS_113 0 -1.8753686067535531e-05
GC_11_114 b_11 NI_11 NS_114 0 -1.5161594332193001e-06
GC_11_115 b_11 NI_11 NS_115 0 -2.9293756288006828e-05
GC_11_116 b_11 NI_11 NS_116 0 2.7696087664219725e-05
GC_11_117 b_11 NI_11 NS_117 0 -2.1496390418427844e-05
GC_11_118 b_11 NI_11 NS_118 0 2.3548923302955025e-05
GC_11_119 b_11 NI_11 NS_119 0 6.0790762495934513e-06
GC_11_120 b_11 NI_11 NS_120 0 2.3428696209196983e-05
GC_11_121 b_11 NI_11 NS_121 0 -1.5899459126598287e-05
GC_11_122 b_11 NI_11 NS_122 0 5.5620861755864306e-05
GC_11_123 b_11 NI_11 NS_123 0 5.4333653022300063e-05
GC_11_124 b_11 NI_11 NS_124 0 6.5659238760355199e-05
GC_11_125 b_11 NI_11 NS_125 0 2.2574534132986993e-05
GC_11_126 b_11 NI_11 NS_126 0 4.5651720279058430e-05
GC_11_127 b_11 NI_11 NS_127 0 1.4988559504347248e-05
GC_11_128 b_11 NI_11 NS_128 0 4.9567425758152815e-05
GC_11_129 b_11 NI_11 NS_129 0 -5.1673363651487066e-04
GC_11_130 b_11 NI_11 NS_130 0 2.4177847896412243e-05
GC_11_131 b_11 NI_11 NS_131 0 -1.7525452095133627e-05
GC_11_132 b_11 NI_11 NS_132 0 -2.5351705939687986e-04
GC_11_133 b_11 NI_11 NS_133 0 -1.0840951116474921e-10
GC_11_134 b_11 NI_11 NS_134 0 4.8101624044058115e-09
GC_11_135 b_11 NI_11 NS_135 0 5.0649840232325952e-06
GC_11_136 b_11 NI_11 NS_136 0 9.6682506236630324e-06
GC_11_137 b_11 NI_11 NS_137 0 1.6493793536150346e-05
GC_11_138 b_11 NI_11 NS_138 0 1.3404317775622513e-05
GC_11_139 b_11 NI_11 NS_139 0 3.8423175046213176e-05
GC_11_140 b_11 NI_11 NS_140 0 -3.4230207504710022e-06
GC_11_141 b_11 NI_11 NS_141 0 1.4655240253047387e-05
GC_11_142 b_11 NI_11 NS_142 0 -6.2678549867060642e-05
GC_11_143 b_11 NI_11 NS_143 0 -1.1682861416242784e-05
GC_11_144 b_11 NI_11 NS_144 0 -9.0308617023093165e-06
GC_11_145 b_11 NI_11 NS_145 0 4.7729738618559334e-06
GC_11_146 b_11 NI_11 NS_146 0 -3.5003845606341421e-06
GC_11_147 b_11 NI_11 NS_147 0 9.7656285918642550e-06
GC_11_148 b_11 NI_11 NS_148 0 -4.9987527104862736e-05
GC_11_149 b_11 NI_11 NS_149 0 -6.6158996585859449e-05
GC_11_150 b_11 NI_11 NS_150 0 -2.1604507570584313e-05
GC_11_151 b_11 NI_11 NS_151 0 -1.6750712944858810e-05
GC_11_152 b_11 NI_11 NS_152 0 1.9351803436505492e-05
GC_11_153 b_11 NI_11 NS_153 0 1.6103498621857804e-05
GC_11_154 b_11 NI_11 NS_154 0 -1.2511216447052201e-06
GC_11_155 b_11 NI_11 NS_155 0 2.1545969347177502e-04
GC_11_156 b_11 NI_11 NS_156 0 7.2320055730428795e-06
GC_11_157 b_11 NI_11 NS_157 0 3.9532339171836548e-04
GC_11_158 b_11 NI_11 NS_158 0 -2.0165265755622960e-03
GC_11_159 b_11 NI_11 NS_159 0 4.0770678058206364e-10
GC_11_160 b_11 NI_11 NS_160 0 -2.7109182572589901e-08
GC_11_161 b_11 NI_11 NS_161 0 1.8507561832485304e-05
GC_11_162 b_11 NI_11 NS_162 0 4.3378359708821096e-05
GC_11_163 b_11 NI_11 NS_163 0 8.1727560098113734e-05
GC_11_164 b_11 NI_11 NS_164 0 -3.0737467612997545e-05
GC_11_165 b_11 NI_11 NS_165 0 -1.3901176150742021e-05
GC_11_166 b_11 NI_11 NS_166 0 1.3616747093684171e-05
GC_11_167 b_11 NI_11 NS_167 0 1.9708381321716263e-04
GC_11_168 b_11 NI_11 NS_168 0 -9.8844897031513527e-05
GC_11_169 b_11 NI_11 NS_169 0 2.6786766006532836e-05
GC_11_170 b_11 NI_11 NS_170 0 -9.8065688494444213e-05
GC_11_171 b_11 NI_11 NS_171 0 -1.7472511297423367e-05
GC_11_172 b_11 NI_11 NS_172 0 -9.8086077113027670e-05
GC_11_173 b_11 NI_11 NS_173 0 9.8369784629573268e-06
GC_11_174 b_11 NI_11 NS_174 0 -9.7505026915439613e-05
GC_11_175 b_11 NI_11 NS_175 0 -9.8088433941717791e-05
GC_11_176 b_11 NI_11 NS_176 0 -3.1485388079871741e-04
GC_11_177 b_11 NI_11 NS_177 0 -1.3395601718407184e-04
GC_11_178 b_11 NI_11 NS_178 0 -1.1516728085802833e-04
GC_11_179 b_11 NI_11 NS_179 0 -1.9684699850390934e-05
GC_11_180 b_11 NI_11 NS_180 0 -1.9125377866070095e-04
GC_11_181 b_11 NI_11 NS_181 0 1.5201720074701211e-03
GC_11_182 b_11 NI_11 NS_182 0 -1.0206020577446964e-04
GC_11_183 b_11 NI_11 NS_183 0 1.5107002763036428e-04
GC_11_184 b_11 NI_11 NS_184 0 1.2317844495784135e-05
GC_11_185 b_11 NI_11 NS_185 0 -4.2760172506881040e-10
GC_11_186 b_11 NI_11 NS_186 0 4.5173474093349532e-08
GC_11_187 b_11 NI_11 NS_187 0 5.2778161262714664e-06
GC_11_188 b_11 NI_11 NS_188 0 7.5702684104743287e-05
GC_11_189 b_11 NI_11 NS_189 0 1.5331514819327995e-04
GC_11_190 b_11 NI_11 NS_190 0 1.3549625473952627e-04
GC_11_191 b_11 NI_11 NS_191 0 3.4661306248518983e-04
GC_11_192 b_11 NI_11 NS_192 0 -2.4832170881305117e-05
GC_11_193 b_11 NI_11 NS_193 0 5.1685676330989786e-05
GC_11_194 b_11 NI_11 NS_194 0 -5.8541629982868733e-04
GC_11_195 b_11 NI_11 NS_195 0 -1.4594533316179058e-04
GC_11_196 b_11 NI_11 NS_196 0 -6.8352176427198845e-05
GC_11_197 b_11 NI_11 NS_197 0 5.1710238203805061e-05
GC_11_198 b_11 NI_11 NS_198 0 -1.0508038636386444e-05
GC_11_199 b_11 NI_11 NS_199 0 4.7742078299037750e-05
GC_11_200 b_11 NI_11 NS_200 0 -4.5319513908694253e-04
GC_11_201 b_11 NI_11 NS_201 0 -7.0912994732521000e-04
GC_11_202 b_11 NI_11 NS_202 0 -8.3358420923229659e-05
GC_11_203 b_11 NI_11 NS_203 0 -1.7471253528139483e-04
GC_11_204 b_11 NI_11 NS_204 0 2.5874041171093784e-04
GC_11_205 b_11 NI_11 NS_205 0 1.0252651110903021e-04
GC_11_206 b_11 NI_11 NS_206 0 7.9813427600584772e-05
GC_11_207 b_11 NI_11 NS_207 0 -8.6272400965968385e-05
GC_11_208 b_11 NI_11 NS_208 0 -3.2981071525530701e-04
GC_11_209 b_11 NI_11 NS_209 0 -7.4986728019017443e-03
GC_11_210 b_11 NI_11 NS_210 0 5.4463736044302576e-03
GC_11_211 b_11 NI_11 NS_211 0 -8.2819008874237703e-10
GC_11_212 b_11 NI_11 NS_212 0 -1.6858209024942493e-06
GC_11_213 b_11 NI_11 NS_213 0 2.5534683118825260e-04
GC_11_214 b_11 NI_11 NS_214 0 2.6645211981117609e-03
GC_11_215 b_11 NI_11 NS_215 0 4.5291691759910668e-03
GC_11_216 b_11 NI_11 NS_216 0 -2.7565572830191860e-03
GC_11_217 b_11 NI_11 NS_217 0 -5.4227010287392092e-03
GC_11_218 b_11 NI_11 NS_218 0 4.2041651361554870e-04
GC_11_219 b_11 NI_11 NS_219 0 8.8584610087896476e-03
GC_11_220 b_11 NI_11 NS_220 0 -6.2094131486169094e-04
GC_11_221 b_11 NI_11 NS_221 0 -2.8260900937831881e-03
GC_11_222 b_11 NI_11 NS_222 0 -2.3963195077242390e-03
GC_11_223 b_11 NI_11 NS_223 0 4.3105060396027231e-05
GC_11_224 b_11 NI_11 NS_224 0 -2.1139049464674129e-03
GC_11_225 b_11 NI_11 NS_225 0 -3.5070302768425658e-03
GC_11_226 b_11 NI_11 NS_226 0 5.5496268167169053e-03
GC_11_227 b_11 NI_11 NS_227 0 5.0984923970970562e-03
GC_11_228 b_11 NI_11 NS_228 0 -7.7604205411807899e-03
GC_11_229 b_11 NI_11 NS_229 0 -5.0389100498201408e-03
GC_11_230 b_11 NI_11 NS_230 0 3.0962157420722364e-03
GC_11_231 b_11 NI_11 NS_231 0 2.2446243261625906e-03
GC_11_232 b_11 NI_11 NS_232 0 -1.6873400590580387e-03
GC_11_233 b_11 NI_11 NS_233 0 -5.9469814837945431e-03
GC_11_234 b_11 NI_11 NS_234 0 3.8164576042803455e-03
GC_11_235 b_11 NI_11 NS_235 0 -1.3746089080371303e-03
GC_11_236 b_11 NI_11 NS_236 0 2.3328708467421004e-03
GC_11_237 b_11 NI_11 NS_237 0 7.5881858999508427e-10
GC_11_238 b_11 NI_11 NS_238 0 6.0065829866922035e-07
GC_11_239 b_11 NI_11 NS_239 0 -1.9596140498731016e-04
GC_11_240 b_11 NI_11 NS_240 0 -4.5534341782619192e-04
GC_11_241 b_11 NI_11 NS_241 0 -1.0665939101090565e-03
GC_11_242 b_11 NI_11 NS_242 0 -9.2131959233472335e-04
GC_11_243 b_11 NI_11 NS_243 0 -2.3173790648370524e-03
GC_11_244 b_11 NI_11 NS_244 0 3.1223076785602495e-04
GC_11_245 b_11 NI_11 NS_245 0 -3.4634935108651368e-04
GC_11_246 b_11 NI_11 NS_246 0 4.1981837629813772e-03
GC_11_247 b_11 NI_11 NS_247 0 9.7829186500863943e-04
GC_11_248 b_11 NI_11 NS_248 0 4.4367013036742011e-04
GC_11_249 b_11 NI_11 NS_249 0 -3.7329483155213274e-04
GC_11_250 b_11 NI_11 NS_250 0 7.9843243359172943e-05
GC_11_251 b_11 NI_11 NS_251 0 -3.1453282997478016e-04
GC_11_252 b_11 NI_11 NS_252 0 3.3540654670163005e-03
GC_11_253 b_11 NI_11 NS_253 0 5.2329434371575180e-03
GC_11_254 b_11 NI_11 NS_254 0 8.1284473435285843e-04
GC_11_255 b_11 NI_11 NS_255 0 1.3427527634437227e-03
GC_11_256 b_11 NI_11 NS_256 0 -1.9440163306120872e-03
GC_11_257 b_11 NI_11 NS_257 0 -8.8256362515712393e-04
GC_11_258 b_11 NI_11 NS_258 0 -6.3689550758349700e-04
GC_11_259 b_11 NI_11 NS_259 0 -1.4735606988318206e-03
GC_11_260 b_11 NI_11 NS_260 0 2.5664403223774547e-03
GC_11_261 b_11 NI_11 NS_261 0 5.9934872176725558e-02
GC_11_262 b_11 NI_11 NS_262 0 -6.4654688880769473e-02
GC_11_263 b_11 NI_11 NS_263 0 -1.0233459242464464e-08
GC_11_264 b_11 NI_11 NS_264 0 -8.1983890893134588e-06
GC_11_265 b_11 NI_11 NS_265 0 -1.8758509241864956e-03
GC_11_266 b_11 NI_11 NS_266 0 -2.8706552577083470e-03
GC_11_267 b_11 NI_11 NS_267 0 -5.0998749713799460e-03
GC_11_268 b_11 NI_11 NS_268 0 1.9265463411645828e-03
GC_11_269 b_11 NI_11 NS_269 0 2.3837857309807384e-03
GC_11_270 b_11 NI_11 NS_270 0 -1.2477164560036559e-03
GC_11_271 b_11 NI_11 NS_271 0 -1.0661877419294493e-02
GC_11_272 b_11 NI_11 NS_272 0 1.1356494290803651e-03
GC_11_273 b_11 NI_11 NS_273 0 5.9634084239520643e-04
GC_11_274 b_11 NI_11 NS_274 0 1.7470507596459629e-03
GC_11_275 b_11 NI_11 NS_275 0 -9.6081025971570064e-04
GC_11_276 b_11 NI_11 NS_276 0 2.2969430900836450e-03
GC_11_277 b_11 NI_11 NS_277 0 5.3287960886574850e-04
GC_11_278 b_11 NI_11 NS_278 0 -5.8517889776854163e-03
GC_11_279 b_11 NI_11 NS_279 0 -8.5170581773715542e-03
GC_11_280 b_11 NI_11 NS_280 0 6.9045152310177500e-03
GC_11_281 b_11 NI_11 NS_281 0 2.5028293539788135e-03
GC_11_282 b_11 NI_11 NS_282 0 -3.6531654157300575e-03
GC_11_283 b_11 NI_11 NS_283 0 -2.5960272420183991e-03
GC_11_284 b_11 NI_11 NS_284 0 -5.3417109205793978e-04
GC_11_285 b_11 NI_11 NS_285 0 5.5354237091426325e-02
GC_11_286 b_11 NI_11 NS_286 0 1.8152607095886688e-03
GC_11_287 b_11 NI_11 NS_287 0 -5.0037327829396315e-02
GC_11_288 b_11 NI_11 NS_288 0 1.1076328461393392e-01
GC_11_289 b_11 NI_11 NS_289 0 1.1665773251622735e-08
GC_11_290 b_11 NI_11 NS_290 0 1.9861986579842647e-05
GC_11_291 b_11 NI_11 NS_291 0 -1.5739397893329860e-02
GC_11_292 b_11 NI_11 NS_292 0 2.4245668900486857e-02
GC_11_293 b_11 NI_11 NS_293 0 -7.8711079956238321e-03
GC_11_294 b_11 NI_11 NS_294 0 -1.4518764823294446e-02
GC_11_295 b_11 NI_11 NS_295 0 2.0325311073735711e-02
GC_11_296 b_11 NI_11 NS_296 0 6.6761281774983137e-03
GC_11_297 b_11 NI_11 NS_297 0 8.0659041034618819e-03
GC_11_298 b_11 NI_11 NS_298 0 4.4188587774245537e-02
GC_11_299 b_11 NI_11 NS_299 0 -1.1822662229691951e-02
GC_11_300 b_11 NI_11 NS_300 0 -3.1939218945757123e-03
GC_11_301 b_11 NI_11 NS_301 0 -5.1132688764593797e-03
GC_11_302 b_11 NI_11 NS_302 0 -4.0785583363014471e-03
GC_11_303 b_11 NI_11 NS_303 0 2.6802333498360361e-02
GC_11_304 b_11 NI_11 NS_304 0 1.2877611304160569e-04
GC_11_305 b_11 NI_11 NS_305 0 3.4101248503789233e-02
GC_11_306 b_11 NI_11 NS_306 0 3.1057524260687835e-02
GC_11_307 b_11 NI_11 NS_307 0 -1.5591728455634200e-02
GC_11_308 b_11 NI_11 NS_308 0 8.2163429262317560e-03
GC_11_309 b_11 NI_11 NS_309 0 -1.0700800155233480e-03
GC_11_310 b_11 NI_11 NS_310 0 -6.8531986409254573e-03
GC_11_311 b_11 NI_11 NS_311 0 -6.9888024605155433e-02
GC_11_312 b_11 NI_11 NS_312 0 1.6944964169878815e-03
GD_11_1 b_11 NI_11 NA_1 0 1.1329725107923389e-05
GD_11_2 b_11 NI_11 NA_2 0 3.1921477912352178e-06
GD_11_3 b_11 NI_11 NA_3 0 8.9205540932762657e-06
GD_11_4 b_11 NI_11 NA_4 0 7.7472952676729611e-06
GD_11_5 b_11 NI_11 NA_5 0 5.5021187994817243e-07
GD_11_6 b_11 NI_11 NA_6 0 3.5144869535856608e-05
GD_11_7 b_11 NI_11 NA_7 0 1.6319284715978337e-04
GD_11_8 b_11 NI_11 NA_8 0 1.3331433614870728e-04
GD_11_9 b_11 NI_11 NA_9 0 1.3427306305630242e-02
GD_11_10 b_11 NI_11 NA_10 0 -1.1219485718105334e-03
GD_11_11 b_11 NI_11 NA_11 0 -2.9881632654782862e-02
GD_11_12 b_11 NI_11 NA_12 0 -2.0539297881308625e-02
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -1.1797570252669703e-05
GC_12_2 b_12 NI_12 NS_2 0 -5.5691853433838269e-06
GC_12_3 b_12 NI_12 NS_3 0 -3.0498513015992871e-11
GC_12_4 b_12 NI_12 NS_4 0 -1.3564556114991476e-10
GC_12_5 b_12 NI_12 NS_5 0 2.2975255125355737e-06
GC_12_6 b_12 NI_12 NS_6 0 1.7812182265993157e-06
GC_12_7 b_12 NI_12 NS_7 0 -6.4111922510698784e-07
GC_12_8 b_12 NI_12 NS_8 0 -3.8629249152882822e-07
GC_12_9 b_12 NI_12 NS_9 0 1.5521516806902440e-06
GC_12_10 b_12 NI_12 NS_10 0 -1.1535837110341623e-06
GC_12_11 b_12 NI_12 NS_11 0 1.8422851526251265e-06
GC_12_12 b_12 NI_12 NS_12 0 -4.3467506702939397e-07
GC_12_13 b_12 NI_12 NS_13 0 1.1803394576520930e-07
GC_12_14 b_12 NI_12 NS_14 0 -1.8751662639441011e-07
GC_12_15 b_12 NI_12 NS_15 0 5.5244992053347525e-08
GC_12_16 b_12 NI_12 NS_16 0 -3.1825272840054238e-07
GC_12_17 b_12 NI_12 NS_17 0 4.3506160587420214e-07
GC_12_18 b_12 NI_12 NS_18 0 -7.3873623929982073e-07
GC_12_19 b_12 NI_12 NS_19 0 9.1283351560315807e-07
GC_12_20 b_12 NI_12 NS_20 0 -1.3978332452319775e-06
GC_12_21 b_12 NI_12 NS_21 0 -1.9067286661987305e-07
GC_12_22 b_12 NI_12 NS_22 0 5.9848034657615100e-07
GC_12_23 b_12 NI_12 NS_23 0 3.5017977628176399e-07
GC_12_24 b_12 NI_12 NS_24 0 -1.5154643106458540e-08
GC_12_25 b_12 NI_12 NS_25 0 5.8038829913424421e-06
GC_12_26 b_12 NI_12 NS_26 0 2.3966716566912995e-06
GC_12_27 b_12 NI_12 NS_27 0 -3.5487274974771937e-05
GC_12_28 b_12 NI_12 NS_28 0 4.3755693920935175e-05
GC_12_29 b_12 NI_12 NS_29 0 3.2703454529600078e-11
GC_12_30 b_12 NI_12 NS_30 0 -2.6824524781632964e-10
GC_12_31 b_12 NI_12 NS_31 0 1.0320796327419903e-06
GC_12_32 b_12 NI_12 NS_32 0 1.0605761692636599e-06
GC_12_33 b_12 NI_12 NS_33 0 1.7241338669414169e-06
GC_12_34 b_12 NI_12 NS_34 0 2.5964967543165208e-07
GC_12_35 b_12 NI_12 NS_35 0 1.0932111829717883e-06
GC_12_36 b_12 NI_12 NS_36 0 4.6059835919624293e-07
GC_12_37 b_12 NI_12 NS_37 0 2.9262620517772246e-06
GC_12_38 b_12 NI_12 NS_38 0 -4.3423249646901929e-07
GC_12_39 b_12 NI_12 NS_39 0 1.0132358698160301e-06
GC_12_40 b_12 NI_12 NS_40 0 5.3040815337453892e-09
GC_12_41 b_12 NI_12 NS_41 0 5.6285423503848203e-07
GC_12_42 b_12 NI_12 NS_42 0 -5.1625013856882879e-07
GC_12_43 b_12 NI_12 NS_43 0 1.6607430423062694e-06
GC_12_44 b_12 NI_12 NS_44 0 1.2910024602005999e-06
GC_12_45 b_12 NI_12 NS_45 0 2.8544591178677821e-06
GC_12_46 b_12 NI_12 NS_46 0 -1.2126691420498421e-06
GC_12_47 b_12 NI_12 NS_47 0 5.5986021873745868e-07
GC_12_48 b_12 NI_12 NS_48 0 1.1266010851967697e-06
GC_12_49 b_12 NI_12 NS_49 0 3.9045706989159638e-07
GC_12_50 b_12 NI_12 NS_50 0 1.5530727911605897e-06
GC_12_51 b_12 NI_12 NS_51 0 -3.6623115448116268e-05
GC_12_52 b_12 NI_12 NS_52 0 -3.7034576498221664e-06
GC_12_53 b_12 NI_12 NS_53 0 -2.4858860783792326e-05
GC_12_54 b_12 NI_12 NS_54 0 2.0849540608071523e-05
GC_12_55 b_12 NI_12 NS_55 0 -3.5016416924174342e-11
GC_12_56 b_12 NI_12 NS_56 0 -2.6867107882395603e-10
GC_12_57 b_12 NI_12 NS_57 0 1.6182387216772835e-06
GC_12_58 b_12 NI_12 NS_58 0 1.4407743386463441e-06
GC_12_59 b_12 NI_12 NS_59 0 2.6022693911595453e-07
GC_12_60 b_12 NI_12 NS_60 0 3.7182518690874001e-07
GC_12_61 b_12 NI_12 NS_61 0 1.7425642445498522e-06
GC_12_62 b_12 NI_12 NS_62 0 -2.0555215158228333e-07
GC_12_63 b_12 NI_12 NS_63 0 3.3663628089467519e-06
GC_12_64 b_12 NI_12 NS_64 0 -1.0275574567843550e-06
GC_12_65 b_12 NI_12 NS_65 0 4.2285822679489970e-07
GC_12_66 b_12 NI_12 NS_66 0 5.1377087750729743e-08
GC_12_67 b_12 NI_12 NS_67 0 2.5477397766724403e-07
GC_12_68 b_12 NI_12 NS_68 0 -2.9685419630507140e-07
GC_12_69 b_12 NI_12 NS_69 0 1.0839097553855493e-06
GC_12_70 b_12 NI_12 NS_70 0 -1.0037311593885309e-06
GC_12_71 b_12 NI_12 NS_71 0 1.6366705546044817e-06
GC_12_72 b_12 NI_12 NS_72 0 -1.2095531562853831e-06
GC_12_73 b_12 NI_12 NS_73 0 -5.6794037365246510e-08
GC_12_74 b_12 NI_12 NS_74 0 1.3046417165856357e-06
GC_12_75 b_12 NI_12 NS_75 0 3.3322391731526925e-07
GC_12_76 b_12 NI_12 NS_76 0 6.8985923699759929e-07
GC_12_77 b_12 NI_12 NS_77 0 -1.7035033448717149e-05
GC_12_78 b_12 NI_12 NS_78 0 -1.3465757904357997e-06
GC_12_79 b_12 NI_12 NS_79 0 -2.7798142785676495e-05
GC_12_80 b_12 NI_12 NS_80 0 4.2303139645931034e-05
GC_12_81 b_12 NI_12 NS_81 0 3.6714333312259701e-11
GC_12_82 b_12 NI_12 NS_82 0 -2.7999033049334339e-10
GC_12_83 b_12 NI_12 NS_83 0 8.4060977623393487e-07
GC_12_84 b_12 NI_12 NS_84 0 4.8887836706243212e-07
GC_12_85 b_12 NI_12 NS_85 0 4.0308548777246327e-07
GC_12_86 b_12 NI_12 NS_86 0 -7.5631255150269464e-07
GC_12_87 b_12 NI_12 NS_87 0 -4.8232153491443750e-07
GC_12_88 b_12 NI_12 NS_88 0 9.9488195182904415e-07
GC_12_89 b_12 NI_12 NS_89 0 1.4097772266015355e-06
GC_12_90 b_12 NI_12 NS_90 0 1.8137230284899505e-07
GC_12_91 b_12 NI_12 NS_91 0 -4.2612465129644331e-07
GC_12_92 b_12 NI_12 NS_92 0 9.6865223307110882e-07
GC_12_93 b_12 NI_12 NS_93 0 5.7062320849582725e-07
GC_12_94 b_12 NI_12 NS_94 0 3.8250636042150613e-07
GC_12_95 b_12 NI_12 NS_95 0 5.5583619722727032e-07
GC_12_96 b_12 NI_12 NS_96 0 3.2468888222682127e-06
GC_12_97 b_12 NI_12 NS_97 0 3.9989909454333139e-06
GC_12_98 b_12 NI_12 NS_98 0 7.7857558612711763e-07
GC_12_99 b_12 NI_12 NS_99 0 9.0089335274510423e-07
GC_12_100 b_12 NI_12 NS_100 0 2.3851795247572355e-06
GC_12_101 b_12 NI_12 NS_101 0 1.1489769064503067e-06
GC_12_102 b_12 NI_12 NS_102 0 2.6054710429043479e-06
GC_12_103 b_12 NI_12 NS_103 0 -3.3471210253637544e-05
GC_12_104 b_12 NI_12 NS_104 0 4.1446808705433656e-07
GC_12_105 b_12 NI_12 NS_105 0 -1.7314430851867561e-05
GC_12_106 b_12 NI_12 NS_106 0 -2.5362085271826056e-04
GC_12_107 b_12 NI_12 NS_107 0 -1.0841168075004451e-10
GC_12_108 b_12 NI_12 NS_108 0 4.8114849797877035e-09
GC_12_109 b_12 NI_12 NS_109 0 5.0737559379129060e-06
GC_12_110 b_12 NI_12 NS_110 0 9.7330063808582592e-06
GC_12_111 b_12 NI_12 NS_111 0 1.6486990290205782e-05
GC_12_112 b_12 NI_12 NS_112 0 1.3338260786005966e-05
GC_12_113 b_12 NI_12 NS_113 0 3.8439306823446135e-05
GC_12_114 b_12 NI_12 NS_114 0 -3.4839413371776869e-06
GC_12_115 b_12 NI_12 NS_115 0 1.4588787507649230e-05
GC_12_116 b_12 NI_12 NS_116 0 -6.2615390869304421e-05
GC_12_117 b_12 NI_12 NS_117 0 -1.1696091813055320e-05
GC_12_118 b_12 NI_12 NS_118 0 -9.0145924369200109e-06
GC_12_119 b_12 NI_12 NS_119 0 4.7616308776375468e-06
GC_12_120 b_12 NI_12 NS_120 0 -3.5113517123472294e-06
GC_12_121 b_12 NI_12 NS_121 0 9.7343947116579984e-06
GC_12_122 b_12 NI_12 NS_122 0 -4.9987537154976831e-05
GC_12_123 b_12 NI_12 NS_123 0 -6.6144971614622060e-05
GC_12_124 b_12 NI_12 NS_124 0 -2.1538293350384389e-05
GC_12_125 b_12 NI_12 NS_125 0 -1.6734573206362417e-05
GC_12_126 b_12 NI_12 NS_126 0 1.9354403919175079e-05
GC_12_127 b_12 NI_12 NS_127 0 1.6110181829437117e-05
GC_12_128 b_12 NI_12 NS_128 0 -1.2647830462061793e-06
GC_12_129 b_12 NI_12 NS_129 0 2.1554434261218265e-04
GC_12_130 b_12 NI_12 NS_130 0 7.2353958549903964e-06
GC_12_131 b_12 NI_12 NS_131 0 -1.4271473596395669e-04
GC_12_132 b_12 NI_12 NS_132 0 6.6398827876130138e-04
GC_12_133 b_12 NI_12 NS_133 0 1.2463229555689493e-10
GC_12_134 b_12 NI_12 NS_134 0 -1.1464989740430575e-08
GC_12_135 b_12 NI_12 NS_135 0 -4.0098324462559567e-06
GC_12_136 b_12 NI_12 NS_136 0 -3.9985351751454620e-06
GC_12_137 b_12 NI_12 NS_137 0 -9.6089759389006607e-06
GC_12_138 b_12 NI_12 NS_138 0 -3.7333276799216413e-06
GC_12_139 b_12 NI_12 NS_139 0 -1.8752441300746589e-05
GC_12_140 b_12 NI_12 NS_140 0 -1.5170146602137774e-06
GC_12_141 b_12 NI_12 NS_141 0 -2.9293434729683400e-05
GC_12_142 b_12 NI_12 NS_142 0 2.7695969760869983e-05
GC_12_143 b_12 NI_12 NS_143 0 -2.1495343563124574e-05
GC_12_144 b_12 NI_12 NS_144 0 2.3548508556752217e-05
GC_12_145 b_12 NI_12 NS_145 0 6.0794688422185585e-06
GC_12_146 b_12 NI_12 NS_146 0 2.3428414745650035e-05
GC_12_147 b_12 NI_12 NS_147 0 -1.5898351493266746e-05
GC_12_148 b_12 NI_12 NS_148 0 5.5619624309295508e-05
GC_12_149 b_12 NI_12 NS_149 0 5.4333376373670778e-05
GC_12_150 b_12 NI_12 NS_150 0 6.5658593028113839e-05
GC_12_151 b_12 NI_12 NS_151 0 2.2574648470536394e-05
GC_12_152 b_12 NI_12 NS_152 0 4.5652058009623420e-05
GC_12_153 b_12 NI_12 NS_153 0 1.4988655931686414e-05
GC_12_154 b_12 NI_12 NS_154 0 4.9568130553067425e-05
GC_12_155 b_12 NI_12 NS_155 0 -5.1674629660697824e-04
GC_12_156 b_12 NI_12 NS_156 0 2.4176486500369352e-05
GC_12_157 b_12 NI_12 NS_157 0 1.5103108378874467e-04
GC_12_158 b_12 NI_12 NS_158 0 1.2368480906084946e-05
GC_12_159 b_12 NI_12 NS_159 0 -4.2760090181003391e-10
GC_12_160 b_12 NI_12 NS_160 0 4.5173253872570853e-08
GC_12_161 b_12 NI_12 NS_161 0 5.2792760994392944e-06
GC_12_162 b_12 NI_12 NS_162 0 7.5700598123346706e-05
GC_12_163 b_12 NI_12 NS_163 0 1.5331439973078275e-04
GC_12_164 b_12 NI_12 NS_164 0 1.3549913128115600e-04
GC_12_165 b_12 NI_12 NS_165 0 3.4661139678540741e-04
GC_12_166 b_12 NI_12 NS_166 0 -2.4829789413269622e-05
GC_12_167 b_12 NI_12 NS_167 0 5.1691377570406889e-05
GC_12_168 b_12 NI_12 NS_168 0 -5.8541576767621127e-04
GC_12_169 b_12 NI_12 NS_169 0 -1.4594355476029485e-04
GC_12_170 b_12 NI_12 NS_170 0 -6.8351846270686662e-05
GC_12_171 b_12 NI_12 NS_171 0 5.1710930868625107e-05
GC_12_172 b_12 NI_12 NS_172 0 -1.0507735863531382e-05
GC_12_173 b_12 NI_12 NS_173 0 4.7743656413783091e-05
GC_12_174 b_12 NI_12 NS_174 0 -4.5319346341065469e-04
GC_12_175 b_12 NI_12 NS_175 0 -7.0912542411346333e-04
GC_12_176 b_12 NI_12 NS_176 0 -8.3358066384554345e-05
GC_12_177 b_12 NI_12 NS_177 0 -1.7471104969526307e-04
GC_12_178 b_12 NI_12 NS_178 0 2.5874147803089042e-04
GC_12_179 b_12 NI_12 NS_179 0 1.0252688875223691e-04
GC_12_180 b_12 NI_12 NS_180 0 7.9815962274817711e-05
GC_12_181 b_12 NI_12 NS_181 0 -8.6313424366681266e-05
GC_12_182 b_12 NI_12 NS_182 0 -3.2981257827635147e-04
GC_12_183 b_12 NI_12 NS_183 0 3.9420726176487333e-04
GC_12_184 b_12 NI_12 NS_184 0 -2.0158041665361789e-03
GC_12_185 b_12 NI_12 NS_185 0 4.0775106433844452e-10
GC_12_186 b_12 NI_12 NS_186 0 -2.7128610073401757e-08
GC_12_187 b_12 NI_12 NS_187 0 1.8621476085839802e-05
GC_12_188 b_12 NI_12 NS_188 0 4.3392278802842948e-05
GC_12_189 b_12 NI_12 NS_189 0 8.1698018620902728e-05
GC_12_190 b_12 NI_12 NS_190 0 -3.0805112238808512e-05
GC_12_191 b_12 NI_12 NS_191 0 -1.3803874706525713e-05
GC_12_192 b_12 NI_12 NS_192 0 1.3744897547408532e-05
GC_12_193 b_12 NI_12 NS_193 0 1.9714653653355192e-04
GC_12_194 b_12 NI_12 NS_194 0 -9.9016357006212775e-05
GC_12_195 b_12 NI_12 NS_195 0 2.6817243944477409e-05
GC_12_196 b_12 NI_12 NS_196 0 -9.8015267852158181e-05
GC_12_197 b_12 NI_12 NS_197 0 -1.7477954309332206e-05
GC_12_198 b_12 NI_12 NS_198 0 -9.8100282824301223e-05
GC_12_199 b_12 NI_12 NS_199 0 9.9799345416017455e-06
GC_12_200 b_12 NI_12 NS_200 0 -9.7467350081518401e-05
GC_12_201 b_12 NI_12 NS_201 0 -9.8080466142243819e-05
GC_12_202 b_12 NI_12 NS_202 0 -3.1492223561225901e-04
GC_12_203 b_12 NI_12 NS_203 0 -1.3387635393416960e-04
GC_12_204 b_12 NI_12 NS_204 0 -1.1513419560661489e-04
GC_12_205 b_12 NI_12 NS_205 0 -1.9677621086664163e-05
GC_12_206 b_12 NI_12 NS_206 0 -1.9124507657278171e-04
GC_12_207 b_12 NI_12 NS_207 0 1.5196010044442139e-03
GC_12_208 b_12 NI_12 NS_208 0 -1.0206151647923588e-04
GC_12_209 b_12 NI_12 NS_209 0 -1.3745905451381098e-03
GC_12_210 b_12 NI_12 NS_210 0 2.3328751956352952e-03
GC_12_211 b_12 NI_12 NS_211 0 7.5881886160042663e-10
GC_12_212 b_12 NI_12 NS_212 0 6.0065828798477989e-07
GC_12_213 b_12 NI_12 NS_213 0 -1.9596046860603485e-04
GC_12_214 b_12 NI_12 NS_214 0 -4.5533533220927275e-04
GC_12_215 b_12 NI_12 NS_215 0 -1.0665948721612427e-03
GC_12_216 b_12 NI_12 NS_216 0 -9.2132735416159783e-04
GC_12_217 b_12 NI_12 NS_217 0 -2.3173774124387470e-03
GC_12_218 b_12 NI_12 NS_218 0 3.1222384568039511e-04
GC_12_219 b_12 NI_12 NS_219 0 -3.4635675297816325e-04
GC_12_220 b_12 NI_12 NS_220 0 4.1981926069968182e-03
GC_12_221 b_12 NI_12 NS_221 0 9.7829070586936224e-04
GC_12_222 b_12 NI_12 NS_222 0 4.4367255478046770e-04
GC_12_223 b_12 NI_12 NS_223 0 -3.7329590593141105e-04
GC_12_224 b_12 NI_12 NS_224 0 7.9841939005989728e-05
GC_12_225 b_12 NI_12 NS_225 0 -3.1453628485497969e-04
GC_12_226 b_12 NI_12 NS_226 0 3.3540664095542553e-03
GC_12_227 b_12 NI_12 NS_227 0 5.2329467711993158e-03
GC_12_228 b_12 NI_12 NS_228 0 8.1285316902855796e-04
GC_12_229 b_12 NI_12 NS_229 0 1.3427552736417615e-03
GC_12_230 b_12 NI_12 NS_230 0 -1.9440156821573179e-03
GC_12_231 b_12 NI_12 NS_231 0 -8.8256278729533140e-04
GC_12_232 b_12 NI_12 NS_232 0 -6.3689652085268560e-04
GC_12_233 b_12 NI_12 NS_233 0 -1.4735645022307155e-03
GC_12_234 b_12 NI_12 NS_234 0 2.5664394616210116e-03
GC_12_235 b_12 NI_12 NS_235 0 -7.4976050247960759e-03
GC_12_236 b_12 NI_12 NS_236 0 5.4454474121714159e-03
GC_12_237 b_12 NI_12 NS_237 0 -8.2825504284325460e-10
GC_12_238 b_12 NI_12 NS_238 0 -1.6858110465050547e-06
GC_12_239 b_12 NI_12 NS_239 0 2.5528979621843576e-04
GC_12_240 b_12 NI_12 NS_240 0 2.6644770986489607e-03
GC_12_241 b_12 NI_12 NS_241 0 4.5291311737956459e-03
GC_12_242 b_12 NI_12 NS_242 0 -2.7565392768417268e-03
GC_12_243 b_12 NI_12 NS_243 0 -5.4227402040446160e-03
GC_12_244 b_12 NI_12 NS_244 0 4.2035093949704299e-04
GC_12_245 b_12 NI_12 NS_245 0 8.8583384359765070e-03
GC_12_246 b_12 NI_12 NS_246 0 -6.2088505594412482e-04
GC_12_247 b_12 NI_12 NS_247 0 -2.8261194604404238e-03
GC_12_248 b_12 NI_12 NS_248 0 -2.3963291279584420e-03
GC_12_249 b_12 NI_12 NS_249 0 4.3090299723284856e-05
GC_12_250 b_12 NI_12 NS_250 0 -2.1138831481322842e-03
GC_12_251 b_12 NI_12 NS_251 0 -3.5070906803346654e-03
GC_12_252 b_12 NI_12 NS_252 0 5.5495734927849382e-03
GC_12_253 b_12 NI_12 NS_253 0 5.0983691843059648e-03
GC_12_254 b_12 NI_12 NS_254 0 -7.7603767194391613e-03
GC_12_255 b_12 NI_12 NS_255 0 -5.0389546366635214e-03
GC_12_256 b_12 NI_12 NS_256 0 3.0962239743942566e-03
GC_12_257 b_12 NI_12 NS_257 0 2.2446188648831871e-03
GC_12_258 b_12 NI_12 NS_258 0 -1.6873558985848404e-03
GC_12_259 b_12 NI_12 NS_259 0 -5.9462060208455196e-03
GC_12_260 b_12 NI_12 NS_260 0 3.8165511269497160e-03
GC_12_261 b_12 NI_12 NS_261 0 -5.0037766385717712e-02
GC_12_262 b_12 NI_12 NS_262 0 1.1076371941789569e-01
GC_12_263 b_12 NI_12 NS_263 0 1.1665793020626096e-08
GC_12_264 b_12 NI_12 NS_264 0 1.9861984027535971e-05
GC_12_265 b_12 NI_12 NS_265 0 -1.5739382493761923e-02
GC_12_266 b_12 NI_12 NS_266 0 2.4245660171461274e-02
GC_12_267 b_12 NI_12 NS_267 0 -7.8711063318772853e-03
GC_12_268 b_12 NI_12 NS_268 0 -1.4518740526456809e-02
GC_12_269 b_12 NI_12 NS_269 0 2.0325306008332569e-02
GC_12_270 b_12 NI_12 NS_270 0 6.6761496592268902e-03
GC_12_271 b_12 NI_12 NS_271 0 8.0659618563202855e-03
GC_12_272 b_12 NI_12 NS_272 0 4.4188589531114611e-02
GC_12_273 b_12 NI_12 NS_273 0 -1.1822640386574837e-02
GC_12_274 b_12 NI_12 NS_274 0 -3.1939187542997893e-03
GC_12_275 b_12 NI_12 NS_275 0 -5.1132594620222635e-03
GC_12_276 b_12 NI_12 NS_276 0 -4.0785602649854157e-03
GC_12_277 b_12 NI_12 NS_277 0 2.6802354868561164e-02
GC_12_278 b_12 NI_12 NS_278 0 1.2878766545135572e-04
GC_12_279 b_12 NI_12 NS_279 0 3.4101292925104797e-02
GC_12_280 b_12 NI_12 NS_280 0 3.1057519141005411e-02
GC_12_281 b_12 NI_12 NS_281 0 -1.5591712749512550e-02
GC_12_282 b_12 NI_12 NS_282 0 8.2163503952508883e-03
GC_12_283 b_12 NI_12 NS_283 0 -1.0700744194643440e-03
GC_12_284 b_12 NI_12 NS_284 0 -6.8531774377402722e-03
GC_12_285 b_12 NI_12 NS_285 0 -6.9888373032334125e-02
GC_12_286 b_12 NI_12 NS_286 0 1.6944864943063435e-03
GC_12_287 b_12 NI_12 NS_287 0 5.9934872176725572e-02
GC_12_288 b_12 NI_12 NS_288 0 -6.4654688880769556e-02
GC_12_289 b_12 NI_12 NS_289 0 -1.0233459242464641e-08
GC_12_290 b_12 NI_12 NS_290 0 -8.1983890893134673e-06
GC_12_291 b_12 NI_12 NS_291 0 -1.8758509241864954e-03
GC_12_292 b_12 NI_12 NS_292 0 -2.8706552577083492e-03
GC_12_293 b_12 NI_12 NS_293 0 -5.0998749713799460e-03
GC_12_294 b_12 NI_12 NS_294 0 1.9265463411645798e-03
GC_12_295 b_12 NI_12 NS_295 0 2.3837857309807380e-03
GC_12_296 b_12 NI_12 NS_296 0 -1.2477164560036581e-03
GC_12_297 b_12 NI_12 NS_297 0 -1.0661877419294493e-02
GC_12_298 b_12 NI_12 NS_298 0 1.1356494290803618e-03
GC_12_299 b_12 NI_12 NS_299 0 5.9634084239520687e-04
GC_12_300 b_12 NI_12 NS_300 0 1.7470507596459581e-03
GC_12_301 b_12 NI_12 NS_301 0 -9.6081025971570173e-04
GC_12_302 b_12 NI_12 NS_302 0 2.2969430900836411e-03
GC_12_303 b_12 NI_12 NS_303 0 5.3287960886574427e-04
GC_12_304 b_12 NI_12 NS_304 0 -5.8517889776854232e-03
GC_12_305 b_12 NI_12 NS_305 0 -8.5170581773715611e-03
GC_12_306 b_12 NI_12 NS_306 0 6.9045152310177466e-03
GC_12_307 b_12 NI_12 NS_307 0 2.5028293539788101e-03
GC_12_308 b_12 NI_12 NS_308 0 -3.6531654157300605e-03
GC_12_309 b_12 NI_12 NS_309 0 -2.5960272420184013e-03
GC_12_310 b_12 NI_12 NS_310 0 -5.3417109205794347e-04
GC_12_311 b_12 NI_12 NS_311 0 5.5354237091426381e-02
GC_12_312 b_12 NI_12 NS_312 0 1.8152607095886768e-03
GD_12_1 b_12 NI_12 NA_1 0 3.1881946227987220e-06
GD_12_2 b_12 NI_12 NA_2 0 1.1329729207406400e-05
GD_12_3 b_12 NI_12 NA_3 0 7.7476749672612469e-06
GD_12_4 b_12 NI_12 NA_4 0 8.8710180982852016e-06
GD_12_5 b_12 NI_12 NA_5 0 3.5049212387849538e-05
GD_12_6 b_12 NI_12 NA_6 0 5.6434010322872382e-07
GD_12_7 b_12 NI_12 NA_7 0 1.3332437336799685e-04
GD_12_8 b_12 NI_12 NA_8 0 1.6323049397341525e-04
GD_12_9 b_12 NI_12 NA_9 0 -1.1219599193645952e-03
GD_12_10 b_12 NI_12 NA_10 0 1.3427147738053138e-02
GD_12_11 b_12 NI_12 NA_11 0 -2.0539182651673933e-02
GD_12_12 b_12 NI_12 NA_12 0 -2.9881632654782862e-02
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 4.2343545449649795e+00
GS_1_1 0 NS_1 NA_1 0 6.6612210139581451e-01
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 3.2831077413326582e+01
GS_2_1 0 NS_2 NA_1 0 6.6612210139581451e-01
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 2.6080429374782270e+04
GS_3_1 0 NS_3 NA_1 0 6.6612210139581451e-01
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 3.7725017732018654e+02
GS_4_1 0 NS_4 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 3.3374995756891884e+01
RS_6 NS_6 0 3.3374995756891884e+01
GL_5 0 NS_5 NS_6 0 2.6701555989767023e-01
GL_6 0 NS_6 NS_5 0 -2.6701555989767023e-01
GS_5_1 0 NS_5 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 2.9295701153420790e+01
RS_8 NS_8 0 2.9295701153420794e+01
GL_7 0 NS_7 NS_8 0 2.3487955264476459e-01
GL_8 0 NS_8 NS_7 0 -2.3487955264476459e-01
GS_7_1 0 NS_7 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 2.8507729740122922e+01
RS_10 NS_10 0 2.8507729740122926e+01
GL_9 0 NS_9 NS_10 0 2.0394625738154515e-01
GL_10 0 NS_10 NS_9 0 -2.0394625738154515e-01
GS_9_1 0 NS_9 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 2.4864874006578756e+01
RS_12 NS_12 0 2.4864874006578756e+01
GL_11 0 NS_11 NS_12 0 1.7909712637378425e-01
GL_12 0 NS_12 NS_11 0 -1.7909712637378425e-01
GS_11_1 0 NS_11 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 3.3007896983248521e+01
RS_14 NS_14 0 3.3007896983248521e+01
GL_13 0 NS_13 NS_14 0 1.5156613511308689e-01
GL_14 0 NS_14 NS_13 0 -1.5156613511308689e-01
GS_13_1 0 NS_13 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 3.6604236705818273e+01
RS_16 NS_16 0 3.6604236705818266e+01
GL_15 0 NS_15 NS_16 0 1.3563092831954773e-01
GL_16 0 NS_16 NS_15 0 -1.3563092831954773e-01
GS_15_1 0 NS_15 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 2.9177663054419767e+01
RS_18 NS_18 0 2.9177663054419764e+01
GL_17 0 NS_17 NS_18 0 1.0672464725066795e-01
GL_18 0 NS_18 NS_17 0 -1.0672464725066795e-01
GS_17_1 0 NS_17 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 2.6438828877664562e+01
RS_20 NS_20 0 2.6438828877664562e+01
GL_19 0 NS_19 NS_20 0 8.4783325096234138e-02
GL_20 0 NS_20 NS_19 0 -8.4783325096234138e-02
GS_19_1 0 NS_19 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 3.2035193249046884e+01
RS_22 NS_22 0 3.2035193249046884e+01
GL_21 0 NS_21 NS_22 0 5.4984278123817384e-02
GL_22 0 NS_22 NS_21 0 -5.4984278123817384e-02
GS_21_1 0 NS_21 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 3.6868268229015122e+01
RS_24 NS_24 0 3.6868268229015115e+01
GL_23 0 NS_23 NS_24 0 3.0685149591018136e-02
GL_24 0 NS_24 NS_23 0 -3.0685149591018136e-02
GS_23_1 0 NS_23 NA_1 0 6.6612210139581451e-01
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 3.6553981154890621e+01
RS_26 NS_26 0 3.6553981154890629e+01
GL_25 0 NS_25 NS_26 0 3.8052754090332945e-03
GL_26 0 NS_26 NS_25 0 -3.8052754090332945e-03
GS_25_1 0 NS_25 NA_1 0 6.6612210139581451e-01
*
* Real pole n. 27
CS_27 NS_27 0 9.9999999999999998e-13
RS_27 NS_27 0 4.2343545449649795e+00
GS_27_2 0 NS_27 NA_2 0 6.6612210139581451e-01
*
* Real pole n. 28
CS_28 NS_28 0 9.9999999999999998e-13
RS_28 NS_28 0 3.2831077413326582e+01
GS_28_2 0 NS_28 NA_2 0 6.6612210139581451e-01
*
* Real pole n. 29
CS_29 NS_29 0 9.9999999999999998e-13
RS_29 NS_29 0 2.6080429374782270e+04
GS_29_2 0 NS_29 NA_2 0 6.6612210139581451e-01
*
* Real pole n. 30
CS_30 NS_30 0 9.9999999999999998e-13
RS_30 NS_30 0 3.7725017732018654e+02
GS_30_2 0 NS_30 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 3.3374995756891884e+01
RS_32 NS_32 0 3.3374995756891884e+01
GL_31 0 NS_31 NS_32 0 2.6701555989767023e-01
GL_32 0 NS_32 NS_31 0 -2.6701555989767023e-01
GS_31_2 0 NS_31 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 2.9295701153420790e+01
RS_34 NS_34 0 2.9295701153420794e+01
GL_33 0 NS_33 NS_34 0 2.3487955264476459e-01
GL_34 0 NS_34 NS_33 0 -2.3487955264476459e-01
GS_33_2 0 NS_33 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 2.8507729740122922e+01
RS_36 NS_36 0 2.8507729740122926e+01
GL_35 0 NS_35 NS_36 0 2.0394625738154515e-01
GL_36 0 NS_36 NS_35 0 -2.0394625738154515e-01
GS_35_2 0 NS_35 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 2.4864874006578756e+01
RS_38 NS_38 0 2.4864874006578756e+01
GL_37 0 NS_37 NS_38 0 1.7909712637378425e-01
GL_38 0 NS_38 NS_37 0 -1.7909712637378425e-01
GS_37_2 0 NS_37 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 3.3007896983248521e+01
RS_40 NS_40 0 3.3007896983248521e+01
GL_39 0 NS_39 NS_40 0 1.5156613511308689e-01
GL_40 0 NS_40 NS_39 0 -1.5156613511308689e-01
GS_39_2 0 NS_39 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 3.6604236705818273e+01
RS_42 NS_42 0 3.6604236705818266e+01
GL_41 0 NS_41 NS_42 0 1.3563092831954773e-01
GL_42 0 NS_42 NS_41 0 -1.3563092831954773e-01
GS_41_2 0 NS_41 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 2.9177663054419767e+01
RS_44 NS_44 0 2.9177663054419764e+01
GL_43 0 NS_43 NS_44 0 1.0672464725066795e-01
GL_44 0 NS_44 NS_43 0 -1.0672464725066795e-01
GS_43_2 0 NS_43 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 2.6438828877664562e+01
RS_46 NS_46 0 2.6438828877664562e+01
GL_45 0 NS_45 NS_46 0 8.4783325096234138e-02
GL_46 0 NS_46 NS_45 0 -8.4783325096234138e-02
GS_45_2 0 NS_45 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 3.2035193249046884e+01
RS_48 NS_48 0 3.2035193249046884e+01
GL_47 0 NS_47 NS_48 0 5.4984278123817384e-02
GL_48 0 NS_48 NS_47 0 -5.4984278123817384e-02
GS_47_2 0 NS_47 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 3.6868268229015122e+01
RS_50 NS_50 0 3.6868268229015115e+01
GL_49 0 NS_49 NS_50 0 3.0685149591018136e-02
GL_50 0 NS_50 NS_49 0 -3.0685149591018136e-02
GS_49_2 0 NS_49 NA_2 0 6.6612210139581451e-01
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 3.6553981154890621e+01
RS_52 NS_52 0 3.6553981154890629e+01
GL_51 0 NS_51 NS_52 0 3.8052754090332945e-03
GL_52 0 NS_52 NS_51 0 -3.8052754090332945e-03
GS_51_2 0 NS_51 NA_2 0 6.6612210139581451e-01
*
* Real pole n. 53
CS_53 NS_53 0 9.9999999999999998e-13
RS_53 NS_53 0 4.2343545449649795e+00
GS_53_3 0 NS_53 NA_3 0 6.6612210139581451e-01
*
* Real pole n. 54
CS_54 NS_54 0 9.9999999999999998e-13
RS_54 NS_54 0 3.2831077413326582e+01
GS_54_3 0 NS_54 NA_3 0 6.6612210139581451e-01
*
* Real pole n. 55
CS_55 NS_55 0 9.9999999999999998e-13
RS_55 NS_55 0 2.6080429374782270e+04
GS_55_3 0 NS_55 NA_3 0 6.6612210139581451e-01
*
* Real pole n. 56
CS_56 NS_56 0 9.9999999999999998e-13
RS_56 NS_56 0 3.7725017732018654e+02
GS_56_3 0 NS_56 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 3.3374995756891884e+01
RS_58 NS_58 0 3.3374995756891884e+01
GL_57 0 NS_57 NS_58 0 2.6701555989767023e-01
GL_58 0 NS_58 NS_57 0 -2.6701555989767023e-01
GS_57_3 0 NS_57 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 2.9295701153420790e+01
RS_60 NS_60 0 2.9295701153420794e+01
GL_59 0 NS_59 NS_60 0 2.3487955264476459e-01
GL_60 0 NS_60 NS_59 0 -2.3487955264476459e-01
GS_59_3 0 NS_59 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 2.8507729740122922e+01
RS_62 NS_62 0 2.8507729740122926e+01
GL_61 0 NS_61 NS_62 0 2.0394625738154515e-01
GL_62 0 NS_62 NS_61 0 -2.0394625738154515e-01
GS_61_3 0 NS_61 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 2.4864874006578756e+01
RS_64 NS_64 0 2.4864874006578756e+01
GL_63 0 NS_63 NS_64 0 1.7909712637378425e-01
GL_64 0 NS_64 NS_63 0 -1.7909712637378425e-01
GS_63_3 0 NS_63 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 3.3007896983248521e+01
RS_66 NS_66 0 3.3007896983248521e+01
GL_65 0 NS_65 NS_66 0 1.5156613511308689e-01
GL_66 0 NS_66 NS_65 0 -1.5156613511308689e-01
GS_65_3 0 NS_65 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 3.6604236705818273e+01
RS_68 NS_68 0 3.6604236705818266e+01
GL_67 0 NS_67 NS_68 0 1.3563092831954773e-01
GL_68 0 NS_68 NS_67 0 -1.3563092831954773e-01
GS_67_3 0 NS_67 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 2.9177663054419767e+01
RS_70 NS_70 0 2.9177663054419764e+01
GL_69 0 NS_69 NS_70 0 1.0672464725066795e-01
GL_70 0 NS_70 NS_69 0 -1.0672464725066795e-01
GS_69_3 0 NS_69 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 2.6438828877664562e+01
RS_72 NS_72 0 2.6438828877664562e+01
GL_71 0 NS_71 NS_72 0 8.4783325096234138e-02
GL_72 0 NS_72 NS_71 0 -8.4783325096234138e-02
GS_71_3 0 NS_71 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 3.2035193249046884e+01
RS_74 NS_74 0 3.2035193249046884e+01
GL_73 0 NS_73 NS_74 0 5.4984278123817384e-02
GL_74 0 NS_74 NS_73 0 -5.4984278123817384e-02
GS_73_3 0 NS_73 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 3.6868268229015122e+01
RS_76 NS_76 0 3.6868268229015115e+01
GL_75 0 NS_75 NS_76 0 3.0685149591018136e-02
GL_76 0 NS_76 NS_75 0 -3.0685149591018136e-02
GS_75_3 0 NS_75 NA_3 0 6.6612210139581451e-01
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 3.6553981154890621e+01
RS_78 NS_78 0 3.6553981154890629e+01
GL_77 0 NS_77 NS_78 0 3.8052754090332945e-03
GL_78 0 NS_78 NS_77 0 -3.8052754090332945e-03
GS_77_3 0 NS_77 NA_3 0 6.6612210139581451e-01
*
* Real pole n. 79
CS_79 NS_79 0 9.9999999999999998e-13
RS_79 NS_79 0 4.2343545449649795e+00
GS_79_4 0 NS_79 NA_4 0 6.6612210139581451e-01
*
* Real pole n. 80
CS_80 NS_80 0 9.9999999999999998e-13
RS_80 NS_80 0 3.2831077413326582e+01
GS_80_4 0 NS_80 NA_4 0 6.6612210139581451e-01
*
* Real pole n. 81
CS_81 NS_81 0 9.9999999999999998e-13
RS_81 NS_81 0 2.6080429374782270e+04
GS_81_4 0 NS_81 NA_4 0 6.6612210139581451e-01
*
* Real pole n. 82
CS_82 NS_82 0 9.9999999999999998e-13
RS_82 NS_82 0 3.7725017732018654e+02
GS_82_4 0 NS_82 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 3.3374995756891884e+01
RS_84 NS_84 0 3.3374995756891884e+01
GL_83 0 NS_83 NS_84 0 2.6701555989767023e-01
GL_84 0 NS_84 NS_83 0 -2.6701555989767023e-01
GS_83_4 0 NS_83 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 2.9295701153420790e+01
RS_86 NS_86 0 2.9295701153420794e+01
GL_85 0 NS_85 NS_86 0 2.3487955264476459e-01
GL_86 0 NS_86 NS_85 0 -2.3487955264476459e-01
GS_85_4 0 NS_85 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 2.8507729740122922e+01
RS_88 NS_88 0 2.8507729740122926e+01
GL_87 0 NS_87 NS_88 0 2.0394625738154515e-01
GL_88 0 NS_88 NS_87 0 -2.0394625738154515e-01
GS_87_4 0 NS_87 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 2.4864874006578756e+01
RS_90 NS_90 0 2.4864874006578756e+01
GL_89 0 NS_89 NS_90 0 1.7909712637378425e-01
GL_90 0 NS_90 NS_89 0 -1.7909712637378425e-01
GS_89_4 0 NS_89 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 3.3007896983248521e+01
RS_92 NS_92 0 3.3007896983248521e+01
GL_91 0 NS_91 NS_92 0 1.5156613511308689e-01
GL_92 0 NS_92 NS_91 0 -1.5156613511308689e-01
GS_91_4 0 NS_91 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 3.6604236705818273e+01
RS_94 NS_94 0 3.6604236705818266e+01
GL_93 0 NS_93 NS_94 0 1.3563092831954773e-01
GL_94 0 NS_94 NS_93 0 -1.3563092831954773e-01
GS_93_4 0 NS_93 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 2.9177663054419767e+01
RS_96 NS_96 0 2.9177663054419764e+01
GL_95 0 NS_95 NS_96 0 1.0672464725066795e-01
GL_96 0 NS_96 NS_95 0 -1.0672464725066795e-01
GS_95_4 0 NS_95 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 2.6438828877664562e+01
RS_98 NS_98 0 2.6438828877664562e+01
GL_97 0 NS_97 NS_98 0 8.4783325096234138e-02
GL_98 0 NS_98 NS_97 0 -8.4783325096234138e-02
GS_97_4 0 NS_97 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 3.2035193249046884e+01
RS_100 NS_100 0 3.2035193249046884e+01
GL_99 0 NS_99 NS_100 0 5.4984278123817384e-02
GL_100 0 NS_100 NS_99 0 -5.4984278123817384e-02
GS_99_4 0 NS_99 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 3.6868268229015122e+01
RS_102 NS_102 0 3.6868268229015115e+01
GL_101 0 NS_101 NS_102 0 3.0685149591018136e-02
GL_102 0 NS_102 NS_101 0 -3.0685149591018136e-02
GS_101_4 0 NS_101 NA_4 0 6.6612210139581451e-01
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 3.6553981154890621e+01
RS_104 NS_104 0 3.6553981154890629e+01
GL_103 0 NS_103 NS_104 0 3.8052754090332945e-03
GL_104 0 NS_104 NS_103 0 -3.8052754090332945e-03
GS_103_4 0 NS_103 NA_4 0 6.6612210139581451e-01
*
* Real pole n. 105
CS_105 NS_105 0 9.9999999999999998e-13
RS_105 NS_105 0 4.2343545449649795e+00
GS_105_5 0 NS_105 NA_5 0 6.6612210139581451e-01
*
* Real pole n. 106
CS_106 NS_106 0 9.9999999999999998e-13
RS_106 NS_106 0 3.2831077413326582e+01
GS_106_5 0 NS_106 NA_5 0 6.6612210139581451e-01
*
* Real pole n. 107
CS_107 NS_107 0 9.9999999999999998e-13
RS_107 NS_107 0 2.6080429374782270e+04
GS_107_5 0 NS_107 NA_5 0 6.6612210139581451e-01
*
* Real pole n. 108
CS_108 NS_108 0 9.9999999999999998e-13
RS_108 NS_108 0 3.7725017732018654e+02
GS_108_5 0 NS_108 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 3.3374995756891884e+01
RS_110 NS_110 0 3.3374995756891884e+01
GL_109 0 NS_109 NS_110 0 2.6701555989767023e-01
GL_110 0 NS_110 NS_109 0 -2.6701555989767023e-01
GS_109_5 0 NS_109 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 2.9295701153420790e+01
RS_112 NS_112 0 2.9295701153420794e+01
GL_111 0 NS_111 NS_112 0 2.3487955264476459e-01
GL_112 0 NS_112 NS_111 0 -2.3487955264476459e-01
GS_111_5 0 NS_111 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 2.8507729740122922e+01
RS_114 NS_114 0 2.8507729740122926e+01
GL_113 0 NS_113 NS_114 0 2.0394625738154515e-01
GL_114 0 NS_114 NS_113 0 -2.0394625738154515e-01
GS_113_5 0 NS_113 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 2.4864874006578756e+01
RS_116 NS_116 0 2.4864874006578756e+01
GL_115 0 NS_115 NS_116 0 1.7909712637378425e-01
GL_116 0 NS_116 NS_115 0 -1.7909712637378425e-01
GS_115_5 0 NS_115 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 3.3007896983248521e+01
RS_118 NS_118 0 3.3007896983248521e+01
GL_117 0 NS_117 NS_118 0 1.5156613511308689e-01
GL_118 0 NS_118 NS_117 0 -1.5156613511308689e-01
GS_117_5 0 NS_117 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 3.6604236705818273e+01
RS_120 NS_120 0 3.6604236705818266e+01
GL_119 0 NS_119 NS_120 0 1.3563092831954773e-01
GL_120 0 NS_120 NS_119 0 -1.3563092831954773e-01
GS_119_5 0 NS_119 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 2.9177663054419767e+01
RS_122 NS_122 0 2.9177663054419764e+01
GL_121 0 NS_121 NS_122 0 1.0672464725066795e-01
GL_122 0 NS_122 NS_121 0 -1.0672464725066795e-01
GS_121_5 0 NS_121 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 2.6438828877664562e+01
RS_124 NS_124 0 2.6438828877664562e+01
GL_123 0 NS_123 NS_124 0 8.4783325096234138e-02
GL_124 0 NS_124 NS_123 0 -8.4783325096234138e-02
GS_123_5 0 NS_123 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 3.2035193249046884e+01
RS_126 NS_126 0 3.2035193249046884e+01
GL_125 0 NS_125 NS_126 0 5.4984278123817384e-02
GL_126 0 NS_126 NS_125 0 -5.4984278123817384e-02
GS_125_5 0 NS_125 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 3.6868268229015122e+01
RS_128 NS_128 0 3.6868268229015115e+01
GL_127 0 NS_127 NS_128 0 3.0685149591018136e-02
GL_128 0 NS_128 NS_127 0 -3.0685149591018136e-02
GS_127_5 0 NS_127 NA_5 0 6.6612210139581451e-01
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 3.6553981154890621e+01
RS_130 NS_130 0 3.6553981154890629e+01
GL_129 0 NS_129 NS_130 0 3.8052754090332945e-03
GL_130 0 NS_130 NS_129 0 -3.8052754090332945e-03
GS_129_5 0 NS_129 NA_5 0 6.6612210139581451e-01
*
* Real pole n. 131
CS_131 NS_131 0 9.9999999999999998e-13
RS_131 NS_131 0 4.2343545449649795e+00
GS_131_6 0 NS_131 NA_6 0 6.6612210139581451e-01
*
* Real pole n. 132
CS_132 NS_132 0 9.9999999999999998e-13
RS_132 NS_132 0 3.2831077413326582e+01
GS_132_6 0 NS_132 NA_6 0 6.6612210139581451e-01
*
* Real pole n. 133
CS_133 NS_133 0 9.9999999999999998e-13
RS_133 NS_133 0 2.6080429374782270e+04
GS_133_6 0 NS_133 NA_6 0 6.6612210139581451e-01
*
* Real pole n. 134
CS_134 NS_134 0 9.9999999999999998e-13
RS_134 NS_134 0 3.7725017732018654e+02
GS_134_6 0 NS_134 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 3.3374995756891884e+01
RS_136 NS_136 0 3.3374995756891884e+01
GL_135 0 NS_135 NS_136 0 2.6701555989767023e-01
GL_136 0 NS_136 NS_135 0 -2.6701555989767023e-01
GS_135_6 0 NS_135 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 2.9295701153420790e+01
RS_138 NS_138 0 2.9295701153420794e+01
GL_137 0 NS_137 NS_138 0 2.3487955264476459e-01
GL_138 0 NS_138 NS_137 0 -2.3487955264476459e-01
GS_137_6 0 NS_137 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 2.8507729740122922e+01
RS_140 NS_140 0 2.8507729740122926e+01
GL_139 0 NS_139 NS_140 0 2.0394625738154515e-01
GL_140 0 NS_140 NS_139 0 -2.0394625738154515e-01
GS_139_6 0 NS_139 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 2.4864874006578756e+01
RS_142 NS_142 0 2.4864874006578756e+01
GL_141 0 NS_141 NS_142 0 1.7909712637378425e-01
GL_142 0 NS_142 NS_141 0 -1.7909712637378425e-01
GS_141_6 0 NS_141 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 3.3007896983248521e+01
RS_144 NS_144 0 3.3007896983248521e+01
GL_143 0 NS_143 NS_144 0 1.5156613511308689e-01
GL_144 0 NS_144 NS_143 0 -1.5156613511308689e-01
GS_143_6 0 NS_143 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 3.6604236705818273e+01
RS_146 NS_146 0 3.6604236705818266e+01
GL_145 0 NS_145 NS_146 0 1.3563092831954773e-01
GL_146 0 NS_146 NS_145 0 -1.3563092831954773e-01
GS_145_6 0 NS_145 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 2.9177663054419767e+01
RS_148 NS_148 0 2.9177663054419764e+01
GL_147 0 NS_147 NS_148 0 1.0672464725066795e-01
GL_148 0 NS_148 NS_147 0 -1.0672464725066795e-01
GS_147_6 0 NS_147 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 2.6438828877664562e+01
RS_150 NS_150 0 2.6438828877664562e+01
GL_149 0 NS_149 NS_150 0 8.4783325096234138e-02
GL_150 0 NS_150 NS_149 0 -8.4783325096234138e-02
GS_149_6 0 NS_149 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 3.2035193249046884e+01
RS_152 NS_152 0 3.2035193249046884e+01
GL_151 0 NS_151 NS_152 0 5.4984278123817384e-02
GL_152 0 NS_152 NS_151 0 -5.4984278123817384e-02
GS_151_6 0 NS_151 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 3.6868268229015122e+01
RS_154 NS_154 0 3.6868268229015115e+01
GL_153 0 NS_153 NS_154 0 3.0685149591018136e-02
GL_154 0 NS_154 NS_153 0 -3.0685149591018136e-02
GS_153_6 0 NS_153 NA_6 0 6.6612210139581451e-01
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 3.6553981154890621e+01
RS_156 NS_156 0 3.6553981154890629e+01
GL_155 0 NS_155 NS_156 0 3.8052754090332945e-03
GL_156 0 NS_156 NS_155 0 -3.8052754090332945e-03
GS_155_6 0 NS_155 NA_6 0 6.6612210139581451e-01
*
* Real pole n. 157
CS_157 NS_157 0 9.9999999999999998e-13
RS_157 NS_157 0 4.2343545449649795e+00
GS_157_7 0 NS_157 NA_7 0 6.6612210139581451e-01
*
* Real pole n. 158
CS_158 NS_158 0 9.9999999999999998e-13
RS_158 NS_158 0 3.2831077413326582e+01
GS_158_7 0 NS_158 NA_7 0 6.6612210139581451e-01
*
* Real pole n. 159
CS_159 NS_159 0 9.9999999999999998e-13
RS_159 NS_159 0 2.6080429374782270e+04
GS_159_7 0 NS_159 NA_7 0 6.6612210139581451e-01
*
* Real pole n. 160
CS_160 NS_160 0 9.9999999999999998e-13
RS_160 NS_160 0 3.7725017732018654e+02
GS_160_7 0 NS_160 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 3.3374995756891884e+01
RS_162 NS_162 0 3.3374995756891884e+01
GL_161 0 NS_161 NS_162 0 2.6701555989767023e-01
GL_162 0 NS_162 NS_161 0 -2.6701555989767023e-01
GS_161_7 0 NS_161 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 163/164
CS_163 NS_163 0 9.9999999999999998e-13
CS_164 NS_164 0 9.9999999999999998e-13
RS_163 NS_163 0 2.9295701153420790e+01
RS_164 NS_164 0 2.9295701153420794e+01
GL_163 0 NS_163 NS_164 0 2.3487955264476459e-01
GL_164 0 NS_164 NS_163 0 -2.3487955264476459e-01
GS_163_7 0 NS_163 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 2.8507729740122922e+01
RS_166 NS_166 0 2.8507729740122926e+01
GL_165 0 NS_165 NS_166 0 2.0394625738154515e-01
GL_166 0 NS_166 NS_165 0 -2.0394625738154515e-01
GS_165_7 0 NS_165 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 2.4864874006578756e+01
RS_168 NS_168 0 2.4864874006578756e+01
GL_167 0 NS_167 NS_168 0 1.7909712637378425e-01
GL_168 0 NS_168 NS_167 0 -1.7909712637378425e-01
GS_167_7 0 NS_167 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 3.3007896983248521e+01
RS_170 NS_170 0 3.3007896983248521e+01
GL_169 0 NS_169 NS_170 0 1.5156613511308689e-01
GL_170 0 NS_170 NS_169 0 -1.5156613511308689e-01
GS_169_7 0 NS_169 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 3.6604236705818273e+01
RS_172 NS_172 0 3.6604236705818266e+01
GL_171 0 NS_171 NS_172 0 1.3563092831954773e-01
GL_172 0 NS_172 NS_171 0 -1.3563092831954773e-01
GS_171_7 0 NS_171 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 2.9177663054419767e+01
RS_174 NS_174 0 2.9177663054419764e+01
GL_173 0 NS_173 NS_174 0 1.0672464725066795e-01
GL_174 0 NS_174 NS_173 0 -1.0672464725066795e-01
GS_173_7 0 NS_173 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 2.6438828877664562e+01
RS_176 NS_176 0 2.6438828877664562e+01
GL_175 0 NS_175 NS_176 0 8.4783325096234138e-02
GL_176 0 NS_176 NS_175 0 -8.4783325096234138e-02
GS_175_7 0 NS_175 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 3.2035193249046884e+01
RS_178 NS_178 0 3.2035193249046884e+01
GL_177 0 NS_177 NS_178 0 5.4984278123817384e-02
GL_178 0 NS_178 NS_177 0 -5.4984278123817384e-02
GS_177_7 0 NS_177 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 3.6868268229015122e+01
RS_180 NS_180 0 3.6868268229015115e+01
GL_179 0 NS_179 NS_180 0 3.0685149591018136e-02
GL_180 0 NS_180 NS_179 0 -3.0685149591018136e-02
GS_179_7 0 NS_179 NA_7 0 6.6612210139581451e-01
*
* Complex pair n. 181/182
CS_181 NS_181 0 9.9999999999999998e-13
CS_182 NS_182 0 9.9999999999999998e-13
RS_181 NS_181 0 3.6553981154890621e+01
RS_182 NS_182 0 3.6553981154890629e+01
GL_181 0 NS_181 NS_182 0 3.8052754090332945e-03
GL_182 0 NS_182 NS_181 0 -3.8052754090332945e-03
GS_181_7 0 NS_181 NA_7 0 6.6612210139581451e-01
*
* Real pole n. 183
CS_183 NS_183 0 9.9999999999999998e-13
RS_183 NS_183 0 4.2343545449649795e+00
GS_183_8 0 NS_183 NA_8 0 6.6612210139581451e-01
*
* Real pole n. 184
CS_184 NS_184 0 9.9999999999999998e-13
RS_184 NS_184 0 3.2831077413326582e+01
GS_184_8 0 NS_184 NA_8 0 6.6612210139581451e-01
*
* Real pole n. 185
CS_185 NS_185 0 9.9999999999999998e-13
RS_185 NS_185 0 2.6080429374782270e+04
GS_185_8 0 NS_185 NA_8 0 6.6612210139581451e-01
*
* Real pole n. 186
CS_186 NS_186 0 9.9999999999999998e-13
RS_186 NS_186 0 3.7725017732018654e+02
GS_186_8 0 NS_186 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 3.3374995756891884e+01
RS_188 NS_188 0 3.3374995756891884e+01
GL_187 0 NS_187 NS_188 0 2.6701555989767023e-01
GL_188 0 NS_188 NS_187 0 -2.6701555989767023e-01
GS_187_8 0 NS_187 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 2.9295701153420790e+01
RS_190 NS_190 0 2.9295701153420794e+01
GL_189 0 NS_189 NS_190 0 2.3487955264476459e-01
GL_190 0 NS_190 NS_189 0 -2.3487955264476459e-01
GS_189_8 0 NS_189 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 2.8507729740122922e+01
RS_192 NS_192 0 2.8507729740122926e+01
GL_191 0 NS_191 NS_192 0 2.0394625738154515e-01
GL_192 0 NS_192 NS_191 0 -2.0394625738154515e-01
GS_191_8 0 NS_191 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 2.4864874006578756e+01
RS_194 NS_194 0 2.4864874006578756e+01
GL_193 0 NS_193 NS_194 0 1.7909712637378425e-01
GL_194 0 NS_194 NS_193 0 -1.7909712637378425e-01
GS_193_8 0 NS_193 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 3.3007896983248521e+01
RS_196 NS_196 0 3.3007896983248521e+01
GL_195 0 NS_195 NS_196 0 1.5156613511308689e-01
GL_196 0 NS_196 NS_195 0 -1.5156613511308689e-01
GS_195_8 0 NS_195 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 3.6604236705818273e+01
RS_198 NS_198 0 3.6604236705818266e+01
GL_197 0 NS_197 NS_198 0 1.3563092831954773e-01
GL_198 0 NS_198 NS_197 0 -1.3563092831954773e-01
GS_197_8 0 NS_197 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 2.9177663054419767e+01
RS_200 NS_200 0 2.9177663054419764e+01
GL_199 0 NS_199 NS_200 0 1.0672464725066795e-01
GL_200 0 NS_200 NS_199 0 -1.0672464725066795e-01
GS_199_8 0 NS_199 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 201/202
CS_201 NS_201 0 9.9999999999999998e-13
CS_202 NS_202 0 9.9999999999999998e-13
RS_201 NS_201 0 2.6438828877664562e+01
RS_202 NS_202 0 2.6438828877664562e+01
GL_201 0 NS_201 NS_202 0 8.4783325096234138e-02
GL_202 0 NS_202 NS_201 0 -8.4783325096234138e-02
GS_201_8 0 NS_201 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 203/204
CS_203 NS_203 0 9.9999999999999998e-13
CS_204 NS_204 0 9.9999999999999998e-13
RS_203 NS_203 0 3.2035193249046884e+01
RS_204 NS_204 0 3.2035193249046884e+01
GL_203 0 NS_203 NS_204 0 5.4984278123817384e-02
GL_204 0 NS_204 NS_203 0 -5.4984278123817384e-02
GS_203_8 0 NS_203 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 3.6868268229015122e+01
RS_206 NS_206 0 3.6868268229015115e+01
GL_205 0 NS_205 NS_206 0 3.0685149591018136e-02
GL_206 0 NS_206 NS_205 0 -3.0685149591018136e-02
GS_205_8 0 NS_205 NA_8 0 6.6612210139581451e-01
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 3.6553981154890621e+01
RS_208 NS_208 0 3.6553981154890629e+01
GL_207 0 NS_207 NS_208 0 3.8052754090332945e-03
GL_208 0 NS_208 NS_207 0 -3.8052754090332945e-03
GS_207_8 0 NS_207 NA_8 0 6.6612210139581451e-01
*
* Real pole n. 209
CS_209 NS_209 0 9.9999999999999998e-13
RS_209 NS_209 0 4.2343545449649795e+00
GS_209_9 0 NS_209 NA_9 0 6.6612210139581451e-01
*
* Real pole n. 210
CS_210 NS_210 0 9.9999999999999998e-13
RS_210 NS_210 0 3.2831077413326582e+01
GS_210_9 0 NS_210 NA_9 0 6.6612210139581451e-01
*
* Real pole n. 211
CS_211 NS_211 0 9.9999999999999998e-13
RS_211 NS_211 0 2.6080429374782270e+04
GS_211_9 0 NS_211 NA_9 0 6.6612210139581451e-01
*
* Real pole n. 212
CS_212 NS_212 0 9.9999999999999998e-13
RS_212 NS_212 0 3.7725017732018654e+02
GS_212_9 0 NS_212 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 3.3374995756891884e+01
RS_214 NS_214 0 3.3374995756891884e+01
GL_213 0 NS_213 NS_214 0 2.6701555989767023e-01
GL_214 0 NS_214 NS_213 0 -2.6701555989767023e-01
GS_213_9 0 NS_213 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 2.9295701153420790e+01
RS_216 NS_216 0 2.9295701153420794e+01
GL_215 0 NS_215 NS_216 0 2.3487955264476459e-01
GL_216 0 NS_216 NS_215 0 -2.3487955264476459e-01
GS_215_9 0 NS_215 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 2.8507729740122922e+01
RS_218 NS_218 0 2.8507729740122926e+01
GL_217 0 NS_217 NS_218 0 2.0394625738154515e-01
GL_218 0 NS_218 NS_217 0 -2.0394625738154515e-01
GS_217_9 0 NS_217 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 2.4864874006578756e+01
RS_220 NS_220 0 2.4864874006578756e+01
GL_219 0 NS_219 NS_220 0 1.7909712637378425e-01
GL_220 0 NS_220 NS_219 0 -1.7909712637378425e-01
GS_219_9 0 NS_219 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 221/222
CS_221 NS_221 0 9.9999999999999998e-13
CS_222 NS_222 0 9.9999999999999998e-13
RS_221 NS_221 0 3.3007896983248521e+01
RS_222 NS_222 0 3.3007896983248521e+01
GL_221 0 NS_221 NS_222 0 1.5156613511308689e-01
GL_222 0 NS_222 NS_221 0 -1.5156613511308689e-01
GS_221_9 0 NS_221 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 223/224
CS_223 NS_223 0 9.9999999999999998e-13
CS_224 NS_224 0 9.9999999999999998e-13
RS_223 NS_223 0 3.6604236705818273e+01
RS_224 NS_224 0 3.6604236705818266e+01
GL_223 0 NS_223 NS_224 0 1.3563092831954773e-01
GL_224 0 NS_224 NS_223 0 -1.3563092831954773e-01
GS_223_9 0 NS_223 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 225/226
CS_225 NS_225 0 9.9999999999999998e-13
CS_226 NS_226 0 9.9999999999999998e-13
RS_225 NS_225 0 2.9177663054419767e+01
RS_226 NS_226 0 2.9177663054419764e+01
GL_225 0 NS_225 NS_226 0 1.0672464725066795e-01
GL_226 0 NS_226 NS_225 0 -1.0672464725066795e-01
GS_225_9 0 NS_225 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 2.6438828877664562e+01
RS_228 NS_228 0 2.6438828877664562e+01
GL_227 0 NS_227 NS_228 0 8.4783325096234138e-02
GL_228 0 NS_228 NS_227 0 -8.4783325096234138e-02
GS_227_9 0 NS_227 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 229/230
CS_229 NS_229 0 9.9999999999999998e-13
CS_230 NS_230 0 9.9999999999999998e-13
RS_229 NS_229 0 3.2035193249046884e+01
RS_230 NS_230 0 3.2035193249046884e+01
GL_229 0 NS_229 NS_230 0 5.4984278123817384e-02
GL_230 0 NS_230 NS_229 0 -5.4984278123817384e-02
GS_229_9 0 NS_229 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 3.6868268229015122e+01
RS_232 NS_232 0 3.6868268229015115e+01
GL_231 0 NS_231 NS_232 0 3.0685149591018136e-02
GL_232 0 NS_232 NS_231 0 -3.0685149591018136e-02
GS_231_9 0 NS_231 NA_9 0 6.6612210139581451e-01
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 3.6553981154890621e+01
RS_234 NS_234 0 3.6553981154890629e+01
GL_233 0 NS_233 NS_234 0 3.8052754090332945e-03
GL_234 0 NS_234 NS_233 0 -3.8052754090332945e-03
GS_233_9 0 NS_233 NA_9 0 6.6612210139581451e-01
*
* Real pole n. 235
CS_235 NS_235 0 9.9999999999999998e-13
RS_235 NS_235 0 4.2343545449649795e+00
GS_235_10 0 NS_235 NA_10 0 6.6612210139581451e-01
*
* Real pole n. 236
CS_236 NS_236 0 9.9999999999999998e-13
RS_236 NS_236 0 3.2831077413326582e+01
GS_236_10 0 NS_236 NA_10 0 6.6612210139581451e-01
*
* Real pole n. 237
CS_237 NS_237 0 9.9999999999999998e-13
RS_237 NS_237 0 2.6080429374782270e+04
GS_237_10 0 NS_237 NA_10 0 6.6612210139581451e-01
*
* Real pole n. 238
CS_238 NS_238 0 9.9999999999999998e-13
RS_238 NS_238 0 3.7725017732018654e+02
GS_238_10 0 NS_238 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 3.3374995756891884e+01
RS_240 NS_240 0 3.3374995756891884e+01
GL_239 0 NS_239 NS_240 0 2.6701555989767023e-01
GL_240 0 NS_240 NS_239 0 -2.6701555989767023e-01
GS_239_10 0 NS_239 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 241/242
CS_241 NS_241 0 9.9999999999999998e-13
CS_242 NS_242 0 9.9999999999999998e-13
RS_241 NS_241 0 2.9295701153420790e+01
RS_242 NS_242 0 2.9295701153420794e+01
GL_241 0 NS_241 NS_242 0 2.3487955264476459e-01
GL_242 0 NS_242 NS_241 0 -2.3487955264476459e-01
GS_241_10 0 NS_241 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 243/244
CS_243 NS_243 0 9.9999999999999998e-13
CS_244 NS_244 0 9.9999999999999998e-13
RS_243 NS_243 0 2.8507729740122922e+01
RS_244 NS_244 0 2.8507729740122926e+01
GL_243 0 NS_243 NS_244 0 2.0394625738154515e-01
GL_244 0 NS_244 NS_243 0 -2.0394625738154515e-01
GS_243_10 0 NS_243 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 245/246
CS_245 NS_245 0 9.9999999999999998e-13
CS_246 NS_246 0 9.9999999999999998e-13
RS_245 NS_245 0 2.4864874006578756e+01
RS_246 NS_246 0 2.4864874006578756e+01
GL_245 0 NS_245 NS_246 0 1.7909712637378425e-01
GL_246 0 NS_246 NS_245 0 -1.7909712637378425e-01
GS_245_10 0 NS_245 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 247/248
CS_247 NS_247 0 9.9999999999999998e-13
CS_248 NS_248 0 9.9999999999999998e-13
RS_247 NS_247 0 3.3007896983248521e+01
RS_248 NS_248 0 3.3007896983248521e+01
GL_247 0 NS_247 NS_248 0 1.5156613511308689e-01
GL_248 0 NS_248 NS_247 0 -1.5156613511308689e-01
GS_247_10 0 NS_247 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 249/250
CS_249 NS_249 0 9.9999999999999998e-13
CS_250 NS_250 0 9.9999999999999998e-13
RS_249 NS_249 0 3.6604236705818273e+01
RS_250 NS_250 0 3.6604236705818266e+01
GL_249 0 NS_249 NS_250 0 1.3563092831954773e-01
GL_250 0 NS_250 NS_249 0 -1.3563092831954773e-01
GS_249_10 0 NS_249 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 251/252
CS_251 NS_251 0 9.9999999999999998e-13
CS_252 NS_252 0 9.9999999999999998e-13
RS_251 NS_251 0 2.9177663054419767e+01
RS_252 NS_252 0 2.9177663054419764e+01
GL_251 0 NS_251 NS_252 0 1.0672464725066795e-01
GL_252 0 NS_252 NS_251 0 -1.0672464725066795e-01
GS_251_10 0 NS_251 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 253/254
CS_253 NS_253 0 9.9999999999999998e-13
CS_254 NS_254 0 9.9999999999999998e-13
RS_253 NS_253 0 2.6438828877664562e+01
RS_254 NS_254 0 2.6438828877664562e+01
GL_253 0 NS_253 NS_254 0 8.4783325096234138e-02
GL_254 0 NS_254 NS_253 0 -8.4783325096234138e-02
GS_253_10 0 NS_253 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 255/256
CS_255 NS_255 0 9.9999999999999998e-13
CS_256 NS_256 0 9.9999999999999998e-13
RS_255 NS_255 0 3.2035193249046884e+01
RS_256 NS_256 0 3.2035193249046884e+01
GL_255 0 NS_255 NS_256 0 5.4984278123817384e-02
GL_256 0 NS_256 NS_255 0 -5.4984278123817384e-02
GS_255_10 0 NS_255 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 257/258
CS_257 NS_257 0 9.9999999999999998e-13
CS_258 NS_258 0 9.9999999999999998e-13
RS_257 NS_257 0 3.6868268229015122e+01
RS_258 NS_258 0 3.6868268229015115e+01
GL_257 0 NS_257 NS_258 0 3.0685149591018136e-02
GL_258 0 NS_258 NS_257 0 -3.0685149591018136e-02
GS_257_10 0 NS_257 NA_10 0 6.6612210139581451e-01
*
* Complex pair n. 259/260
CS_259 NS_259 0 9.9999999999999998e-13
CS_260 NS_260 0 9.9999999999999998e-13
RS_259 NS_259 0 3.6553981154890621e+01
RS_260 NS_260 0 3.6553981154890629e+01
GL_259 0 NS_259 NS_260 0 3.8052754090332945e-03
GL_260 0 NS_260 NS_259 0 -3.8052754090332945e-03
GS_259_10 0 NS_259 NA_10 0 6.6612210139581451e-01
*
* Real pole n. 261
CS_261 NS_261 0 9.9999999999999998e-13
RS_261 NS_261 0 4.2343545449649795e+00
GS_261_11 0 NS_261 NA_11 0 6.6612210139581451e-01
*
* Real pole n. 262
CS_262 NS_262 0 9.9999999999999998e-13
RS_262 NS_262 0 3.2831077413326582e+01
GS_262_11 0 NS_262 NA_11 0 6.6612210139581451e-01
*
* Real pole n. 263
CS_263 NS_263 0 9.9999999999999998e-13
RS_263 NS_263 0 2.6080429374782270e+04
GS_263_11 0 NS_263 NA_11 0 6.6612210139581451e-01
*
* Real pole n. 264
CS_264 NS_264 0 9.9999999999999998e-13
RS_264 NS_264 0 3.7725017732018654e+02
GS_264_11 0 NS_264 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 265/266
CS_265 NS_265 0 9.9999999999999998e-13
CS_266 NS_266 0 9.9999999999999998e-13
RS_265 NS_265 0 3.3374995756891884e+01
RS_266 NS_266 0 3.3374995756891884e+01
GL_265 0 NS_265 NS_266 0 2.6701555989767023e-01
GL_266 0 NS_266 NS_265 0 -2.6701555989767023e-01
GS_265_11 0 NS_265 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 267/268
CS_267 NS_267 0 9.9999999999999998e-13
CS_268 NS_268 0 9.9999999999999998e-13
RS_267 NS_267 0 2.9295701153420790e+01
RS_268 NS_268 0 2.9295701153420794e+01
GL_267 0 NS_267 NS_268 0 2.3487955264476459e-01
GL_268 0 NS_268 NS_267 0 -2.3487955264476459e-01
GS_267_11 0 NS_267 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 269/270
CS_269 NS_269 0 9.9999999999999998e-13
CS_270 NS_270 0 9.9999999999999998e-13
RS_269 NS_269 0 2.8507729740122922e+01
RS_270 NS_270 0 2.8507729740122926e+01
GL_269 0 NS_269 NS_270 0 2.0394625738154515e-01
GL_270 0 NS_270 NS_269 0 -2.0394625738154515e-01
GS_269_11 0 NS_269 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 271/272
CS_271 NS_271 0 9.9999999999999998e-13
CS_272 NS_272 0 9.9999999999999998e-13
RS_271 NS_271 0 2.4864874006578756e+01
RS_272 NS_272 0 2.4864874006578756e+01
GL_271 0 NS_271 NS_272 0 1.7909712637378425e-01
GL_272 0 NS_272 NS_271 0 -1.7909712637378425e-01
GS_271_11 0 NS_271 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 273/274
CS_273 NS_273 0 9.9999999999999998e-13
CS_274 NS_274 0 9.9999999999999998e-13
RS_273 NS_273 0 3.3007896983248521e+01
RS_274 NS_274 0 3.3007896983248521e+01
GL_273 0 NS_273 NS_274 0 1.5156613511308689e-01
GL_274 0 NS_274 NS_273 0 -1.5156613511308689e-01
GS_273_11 0 NS_273 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 275/276
CS_275 NS_275 0 9.9999999999999998e-13
CS_276 NS_276 0 9.9999999999999998e-13
RS_275 NS_275 0 3.6604236705818273e+01
RS_276 NS_276 0 3.6604236705818266e+01
GL_275 0 NS_275 NS_276 0 1.3563092831954773e-01
GL_276 0 NS_276 NS_275 0 -1.3563092831954773e-01
GS_275_11 0 NS_275 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 277/278
CS_277 NS_277 0 9.9999999999999998e-13
CS_278 NS_278 0 9.9999999999999998e-13
RS_277 NS_277 0 2.9177663054419767e+01
RS_278 NS_278 0 2.9177663054419764e+01
GL_277 0 NS_277 NS_278 0 1.0672464725066795e-01
GL_278 0 NS_278 NS_277 0 -1.0672464725066795e-01
GS_277_11 0 NS_277 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 279/280
CS_279 NS_279 0 9.9999999999999998e-13
CS_280 NS_280 0 9.9999999999999998e-13
RS_279 NS_279 0 2.6438828877664562e+01
RS_280 NS_280 0 2.6438828877664562e+01
GL_279 0 NS_279 NS_280 0 8.4783325096234138e-02
GL_280 0 NS_280 NS_279 0 -8.4783325096234138e-02
GS_279_11 0 NS_279 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 281/282
CS_281 NS_281 0 9.9999999999999998e-13
CS_282 NS_282 0 9.9999999999999998e-13
RS_281 NS_281 0 3.2035193249046884e+01
RS_282 NS_282 0 3.2035193249046884e+01
GL_281 0 NS_281 NS_282 0 5.4984278123817384e-02
GL_282 0 NS_282 NS_281 0 -5.4984278123817384e-02
GS_281_11 0 NS_281 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 283/284
CS_283 NS_283 0 9.9999999999999998e-13
CS_284 NS_284 0 9.9999999999999998e-13
RS_283 NS_283 0 3.6868268229015122e+01
RS_284 NS_284 0 3.6868268229015115e+01
GL_283 0 NS_283 NS_284 0 3.0685149591018136e-02
GL_284 0 NS_284 NS_283 0 -3.0685149591018136e-02
GS_283_11 0 NS_283 NA_11 0 6.6612210139581451e-01
*
* Complex pair n. 285/286
CS_285 NS_285 0 9.9999999999999998e-13
CS_286 NS_286 0 9.9999999999999998e-13
RS_285 NS_285 0 3.6553981154890621e+01
RS_286 NS_286 0 3.6553981154890629e+01
GL_285 0 NS_285 NS_286 0 3.8052754090332945e-03
GL_286 0 NS_286 NS_285 0 -3.8052754090332945e-03
GS_285_11 0 NS_285 NA_11 0 6.6612210139581451e-01
*
* Real pole n. 287
CS_287 NS_287 0 9.9999999999999998e-13
RS_287 NS_287 0 4.2343545449649795e+00
GS_287_12 0 NS_287 NA_12 0 6.6612210139581451e-01
*
* Real pole n. 288
CS_288 NS_288 0 9.9999999999999998e-13
RS_288 NS_288 0 3.2831077413326582e+01
GS_288_12 0 NS_288 NA_12 0 6.6612210139581451e-01
*
* Real pole n. 289
CS_289 NS_289 0 9.9999999999999998e-13
RS_289 NS_289 0 2.6080429374782270e+04
GS_289_12 0 NS_289 NA_12 0 6.6612210139581451e-01
*
* Real pole n. 290
CS_290 NS_290 0 9.9999999999999998e-13
RS_290 NS_290 0 3.7725017732018654e+02
GS_290_12 0 NS_290 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 291/292
CS_291 NS_291 0 9.9999999999999998e-13
CS_292 NS_292 0 9.9999999999999998e-13
RS_291 NS_291 0 3.3374995756891884e+01
RS_292 NS_292 0 3.3374995756891884e+01
GL_291 0 NS_291 NS_292 0 2.6701555989767023e-01
GL_292 0 NS_292 NS_291 0 -2.6701555989767023e-01
GS_291_12 0 NS_291 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 293/294
CS_293 NS_293 0 9.9999999999999998e-13
CS_294 NS_294 0 9.9999999999999998e-13
RS_293 NS_293 0 2.9295701153420790e+01
RS_294 NS_294 0 2.9295701153420794e+01
GL_293 0 NS_293 NS_294 0 2.3487955264476459e-01
GL_294 0 NS_294 NS_293 0 -2.3487955264476459e-01
GS_293_12 0 NS_293 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 295/296
CS_295 NS_295 0 9.9999999999999998e-13
CS_296 NS_296 0 9.9999999999999998e-13
RS_295 NS_295 0 2.8507729740122922e+01
RS_296 NS_296 0 2.8507729740122926e+01
GL_295 0 NS_295 NS_296 0 2.0394625738154515e-01
GL_296 0 NS_296 NS_295 0 -2.0394625738154515e-01
GS_295_12 0 NS_295 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 297/298
CS_297 NS_297 0 9.9999999999999998e-13
CS_298 NS_298 0 9.9999999999999998e-13
RS_297 NS_297 0 2.4864874006578756e+01
RS_298 NS_298 0 2.4864874006578756e+01
GL_297 0 NS_297 NS_298 0 1.7909712637378425e-01
GL_298 0 NS_298 NS_297 0 -1.7909712637378425e-01
GS_297_12 0 NS_297 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 299/300
CS_299 NS_299 0 9.9999999999999998e-13
CS_300 NS_300 0 9.9999999999999998e-13
RS_299 NS_299 0 3.3007896983248521e+01
RS_300 NS_300 0 3.3007896983248521e+01
GL_299 0 NS_299 NS_300 0 1.5156613511308689e-01
GL_300 0 NS_300 NS_299 0 -1.5156613511308689e-01
GS_299_12 0 NS_299 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 301/302
CS_301 NS_301 0 9.9999999999999998e-13
CS_302 NS_302 0 9.9999999999999998e-13
RS_301 NS_301 0 3.6604236705818273e+01
RS_302 NS_302 0 3.6604236705818266e+01
GL_301 0 NS_301 NS_302 0 1.3563092831954773e-01
GL_302 0 NS_302 NS_301 0 -1.3563092831954773e-01
GS_301_12 0 NS_301 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 303/304
CS_303 NS_303 0 9.9999999999999998e-13
CS_304 NS_304 0 9.9999999999999998e-13
RS_303 NS_303 0 2.9177663054419767e+01
RS_304 NS_304 0 2.9177663054419764e+01
GL_303 0 NS_303 NS_304 0 1.0672464725066795e-01
GL_304 0 NS_304 NS_303 0 -1.0672464725066795e-01
GS_303_12 0 NS_303 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 305/306
CS_305 NS_305 0 9.9999999999999998e-13
CS_306 NS_306 0 9.9999999999999998e-13
RS_305 NS_305 0 2.6438828877664562e+01
RS_306 NS_306 0 2.6438828877664562e+01
GL_305 0 NS_305 NS_306 0 8.4783325096234138e-02
GL_306 0 NS_306 NS_305 0 -8.4783325096234138e-02
GS_305_12 0 NS_305 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 307/308
CS_307 NS_307 0 9.9999999999999998e-13
CS_308 NS_308 0 9.9999999999999998e-13
RS_307 NS_307 0 3.2035193249046884e+01
RS_308 NS_308 0 3.2035193249046884e+01
GL_307 0 NS_307 NS_308 0 5.4984278123817384e-02
GL_308 0 NS_308 NS_307 0 -5.4984278123817384e-02
GS_307_12 0 NS_307 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 309/310
CS_309 NS_309 0 9.9999999999999998e-13
CS_310 NS_310 0 9.9999999999999998e-13
RS_309 NS_309 0 3.6868268229015122e+01
RS_310 NS_310 0 3.6868268229015115e+01
GL_309 0 NS_309 NS_310 0 3.0685149591018136e-02
GL_310 0 NS_310 NS_309 0 -3.0685149591018136e-02
GS_309_12 0 NS_309 NA_12 0 6.6612210139581451e-01
*
* Complex pair n. 311/312
CS_311 NS_311 0 9.9999999999999998e-13
CS_312 NS_312 0 9.9999999999999998e-13
RS_311 NS_311 0 3.6553981154890621e+01
RS_312 NS_312 0 3.6553981154890629e+01
GL_311 0 NS_311 NS_312 0 3.8052754090332945e-03
GL_312 0 NS_312 NS_311 0 -3.8052754090332945e-03
GS_311_12 0 NS_311 NA_12 0 6.6612210139581451e-01
*
******************************


.ends
*******************
* End of subcircuit
*******************
