**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 5.0000e+10 Hz
** Order: [4 4 24] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_9_Module_wire_1mm_lowloss_85ohm
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 -4.7865465377981290e-03
GC_1_2 b_1 NI_1 NS_2 0 1.6712166530109141e-02
GC_1_3 b_1 NI_1 NS_3 0 -3.5265677044478399e-06
GC_1_4 b_1 NI_1 NS_4 0 2.9828686499955580e-08
GC_1_5 b_1 NI_1 NS_5 0 -1.0045935493791466e-09
GC_1_6 b_1 NI_1 NS_6 0 -2.0063946787977987e-06
GC_1_7 b_1 NI_1 NS_7 0 1.8824449668198545e-02
GC_1_8 b_1 NI_1 NS_8 0 5.0640142559650630e-02
GC_1_9 b_1 NI_1 NS_9 0 1.5094546986776466e-02
GC_1_10 b_1 NI_1 NS_10 0 7.1426549459003286e-02
GC_1_11 b_1 NI_1 NS_11 0 8.1524057415720219e-02
GC_1_12 b_1 NI_1 NS_12 0 4.9053274172503984e-02
GC_1_13 b_1 NI_1 NS_13 0 -2.7410735746251329e-07
GC_1_14 b_1 NI_1 NS_14 0 -6.0326930512179163e-08
GC_1_15 b_1 NI_1 NS_15 0 5.1949012719389255e-07
GC_1_16 b_1 NI_1 NS_16 0 -7.4351513903889747e-07
GC_1_17 b_1 NI_1 NS_17 0 3.9410170769459165e-07
GC_1_18 b_1 NI_1 NS_18 0 3.8363314466611478e-07
GC_1_19 b_1 NI_1 NS_19 0 1.0782291867550657e-02
GC_1_20 b_1 NI_1 NS_20 0 -2.9412988807022023e-02
GC_1_21 b_1 NI_1 NS_21 0 -1.0664358830120690e-05
GC_1_22 b_1 NI_1 NS_22 0 -6.9025041522456622e-07
GC_1_23 b_1 NI_1 NS_23 0 1.2414120994588968e-08
GC_1_24 b_1 NI_1 NS_24 0 8.5957340743521432e-06
GC_1_25 b_1 NI_1 NS_25 0 -5.1463434313970803e-02
GC_1_26 b_1 NI_1 NS_26 0 6.8753121111319593e-02
GC_1_27 b_1 NI_1 NS_27 0 -2.9076064196098976e-02
GC_1_28 b_1 NI_1 NS_28 0 -1.5435086867693890e-01
GC_1_29 b_1 NI_1 NS_29 0 -4.6621488534903310e-03
GC_1_30 b_1 NI_1 NS_30 0 -1.6535003766036616e-01
GC_1_31 b_1 NI_1 NS_31 0 4.7568108775162555e-07
GC_1_32 b_1 NI_1 NS_32 0 8.8281793835481596e-07
GC_1_33 b_1 NI_1 NS_33 0 -4.3322571947488283e-06
GC_1_34 b_1 NI_1 NS_34 0 1.0958063418161353e-07
GC_1_35 b_1 NI_1 NS_35 0 -3.3489481216933043e-06
GC_1_36 b_1 NI_1 NS_36 0 -3.5476791236984440e-06
GC_1_37 b_1 NI_1 NS_37 0 -6.0598290790652668e-04
GC_1_38 b_1 NI_1 NS_38 0 1.3722647392863136e-03
GC_1_39 b_1 NI_1 NS_39 0 -8.5960949097731986e-07
GC_1_40 b_1 NI_1 NS_40 0 -1.4388097122502816e-09
GC_1_41 b_1 NI_1 NS_41 0 -2.7334249772421357e-11
GC_1_42 b_1 NI_1 NS_42 0 -2.1412823488513985e-07
GC_1_43 b_1 NI_1 NS_43 0 -4.2068464574546898e-03
GC_1_44 b_1 NI_1 NS_44 0 1.9038017951993991e-02
GC_1_45 b_1 NI_1 NS_45 0 1.8778280881409159e-02
GC_1_46 b_1 NI_1 NS_46 0 -1.2058896275211376e-02
GC_1_47 b_1 NI_1 NS_47 0 2.1714548187059522e-03
GC_1_48 b_1 NI_1 NS_48 0 2.9269113252549217e-02
GC_1_49 b_1 NI_1 NS_49 0 -3.3659898653910109e-08
GC_1_50 b_1 NI_1 NS_50 0 -2.4511752866974977e-08
GC_1_51 b_1 NI_1 NS_51 0 8.1060534687997777e-08
GC_1_52 b_1 NI_1 NS_52 0 -4.2241276234843315e-08
GC_1_53 b_1 NI_1 NS_53 0 5.1476165046878417e-08
GC_1_54 b_1 NI_1 NS_54 0 3.1306639612583748e-08
GC_1_55 b_1 NI_1 NS_55 0 1.1707866780154507e-04
GC_1_56 b_1 NI_1 NS_56 0 -4.6241020400657564e-04
GC_1_57 b_1 NI_1 NS_57 0 3.5664998677332770e-07
GC_1_58 b_1 NI_1 NS_58 0 3.4774377331845560e-09
GC_1_59 b_1 NI_1 NS_59 0 -1.1877538574569832e-11
GC_1_60 b_1 NI_1 NS_60 0 1.2106504078955389e-07
GC_1_61 b_1 NI_1 NS_61 0 7.0283675803617461e-04
GC_1_62 b_1 NI_1 NS_62 0 -4.2878196445020490e-03
GC_1_63 b_1 NI_1 NS_63 0 -9.0099056624380110e-03
GC_1_64 b_1 NI_1 NS_64 0 -5.1462139024248902e-03
GC_1_65 b_1 NI_1 NS_65 0 1.8367936660560304e-03
GC_1_66 b_1 NI_1 NS_66 0 7.2296956128815558e-03
GC_1_67 b_1 NI_1 NS_67 0 4.0524566424039968e-09
GC_1_68 b_1 NI_1 NS_68 0 2.5486979465476586e-09
GC_1_69 b_1 NI_1 NS_69 0 1.9545768524778620e-09
GC_1_70 b_1 NI_1 NS_70 0 1.2028149427007209e-08
GC_1_71 b_1 NI_1 NS_71 0 -2.5385322697719136e-08
GC_1_72 b_1 NI_1 NS_72 0 -1.4673451662766030e-08
GC_1_73 b_1 NI_1 NS_73 0 -1.3683739784611860e-05
GC_1_74 b_1 NI_1 NS_74 0 4.5862454956669562e-05
GC_1_75 b_1 NI_1 NS_75 0 -1.4594664798258844e-08
GC_1_76 b_1 NI_1 NS_76 0 -6.5101997187818065e-10
GC_1_77 b_1 NI_1 NS_77 0 8.0662292268427709e-11
GC_1_78 b_1 NI_1 NS_78 0 -5.0747168530413411e-09
GC_1_79 b_1 NI_1 NS_79 0 1.1926470916326659e-04
GC_1_80 b_1 NI_1 NS_80 0 1.7734486113283975e-04
GC_1_81 b_1 NI_1 NS_81 0 3.0868337393563064e-04
GC_1_82 b_1 NI_1 NS_82 0 -5.1517026264686348e-04
GC_1_83 b_1 NI_1 NS_83 0 -3.8550123484002146e-04
GC_1_84 b_1 NI_1 NS_84 0 1.7218932774756520e-04
GC_1_85 b_1 NI_1 NS_85 0 -2.6650001615819164e-10
GC_1_86 b_1 NI_1 NS_86 0 -8.7560171010022071e-10
GC_1_87 b_1 NI_1 NS_87 0 -9.7850926515055483e-10
GC_1_88 b_1 NI_1 NS_88 0 3.7261673469129398e-09
GC_1_89 b_1 NI_1 NS_89 0 1.3261416225376639e-09
GC_1_90 b_1 NI_1 NS_90 0 -4.7355176712272049e-10
GC_1_91 b_1 NI_1 NS_91 0 6.5717423233210539e-06
GC_1_92 b_1 NI_1 NS_92 0 -3.4988226165527895e-06
GC_1_93 b_1 NI_1 NS_93 0 2.4262979334763084e-08
GC_1_94 b_1 NI_1 NS_94 0 6.7555753327335981e-10
GC_1_95 b_1 NI_1 NS_95 0 -8.0408494665611449e-11
GC_1_96 b_1 NI_1 NS_96 0 4.3270565343535614e-09
GC_1_97 b_1 NI_1 NS_97 0 -1.3639333441494030e-04
GC_1_98 b_1 NI_1 NS_98 0 1.8277823930736275e-04
GC_1_99 b_1 NI_1 NS_99 0 8.0660338518049994e-04
GC_1_100 b_1 NI_1 NS_100 0 2.0572608882375373e-04
GC_1_101 b_1 NI_1 NS_101 0 -5.4635656225949863e-04
GC_1_102 b_1 NI_1 NS_102 0 -9.0504419762248059e-04
GC_1_103 b_1 NI_1 NS_103 0 -1.3840410139371416e-10
GC_1_104 b_1 NI_1 NS_104 0 8.7166071980694304e-10
GC_1_105 b_1 NI_1 NS_105 0 1.8468558109725652e-09
GC_1_106 b_1 NI_1 NS_106 0 -4.9672058717753255e-09
GC_1_107 b_1 NI_1 NS_107 0 -1.0293053732673079e-09
GC_1_108 b_1 NI_1 NS_108 0 6.3126224008788411e-10
GC_1_109 b_1 NI_1 NS_109 0 1.0261216617708778e-06
GC_1_110 b_1 NI_1 NS_110 0 -6.3678978972115761e-06
GC_1_111 b_1 NI_1 NS_111 0 -3.8617175485388146e-09
GC_1_112 b_1 NI_1 NS_112 0 -2.4265030967254222e-10
GC_1_113 b_1 NI_1 NS_113 0 2.5054234697980783e-11
GC_1_114 b_1 NI_1 NS_114 0 -1.2136409174603176e-10
GC_1_115 b_1 NI_1 NS_115 0 -3.6728333809910111e-05
GC_1_116 b_1 NI_1 NS_116 0 5.6788335178666925e-05
GC_1_117 b_1 NI_1 NS_117 0 8.7836834504802823e-06
GC_1_118 b_1 NI_1 NS_118 0 1.4656168370178781e-04
GC_1_119 b_1 NI_1 NS_119 0 1.6060324238846070e-04
GC_1_120 b_1 NI_1 NS_120 0 5.6663769372135285e-05
GC_1_121 b_1 NI_1 NS_121 0 6.0601659394485999e-11
GC_1_122 b_1 NI_1 NS_122 0 -1.4093745394710007e-10
GC_1_123 b_1 NI_1 NS_123 0 -3.3707579244684988e-10
GC_1_124 b_1 NI_1 NS_124 0 1.0565795678932891e-09
GC_1_125 b_1 NI_1 NS_125 0 5.5575278555730688e-11
GC_1_126 b_1 NI_1 NS_126 0 -4.5373768002208638e-10
GC_1_127 b_1 NI_1 NS_127 0 5.0795777254334691e-06
GC_1_128 b_1 NI_1 NS_128 0 -2.0495034780533969e-05
GC_1_129 b_1 NI_1 NS_129 0 -7.3514280783932257e-10
GC_1_130 b_1 NI_1 NS_130 0 2.0742712061553730e-10
GC_1_131 b_1 NI_1 NS_131 0 -2.4670911087041540e-11
GC_1_132 b_1 NI_1 NS_132 0 6.5223519148247846e-10
GC_1_133 b_1 NI_1 NS_133 0 -1.4010400278214576e-05
GC_1_134 b_1 NI_1 NS_134 0 4.6160804333842001e-05
GC_1_135 b_1 NI_1 NS_135 0 1.4554607310930410e-04
GC_1_136 b_1 NI_1 NS_136 0 3.5634073767886241e-05
GC_1_137 b_1 NI_1 NS_137 0 -7.5467958728928197e-05
GC_1_138 b_1 NI_1 NS_138 0 -1.9906750123601782e-04
GC_1_139 b_1 NI_1 NS_139 0 1.9164604664382456e-10
GC_1_140 b_1 NI_1 NS_140 0 1.5222253685602560e-10
GC_1_141 b_1 NI_1 NS_141 0 -2.7653355800812428e-10
GC_1_142 b_1 NI_1 NS_142 0 -4.0006459054831123e-10
GC_1_143 b_1 NI_1 NS_143 0 -2.7141979702088624e-10
GC_1_144 b_1 NI_1 NS_144 0 2.8552958008527951e-10
GC_1_145 b_1 NI_1 NS_145 0 3.8927239825449180e-07
GC_1_146 b_1 NI_1 NS_146 0 -1.0156602204145936e-06
GC_1_147 b_1 NI_1 NS_147 0 -5.7479688014437815e-10
GC_1_148 b_1 NI_1 NS_148 0 -1.0307943240428172e-10
GC_1_149 b_1 NI_1 NS_149 0 8.1837463968406665e-12
GC_1_150 b_1 NI_1 NS_150 0 1.6175566693372358e-10
GC_1_151 b_1 NI_1 NS_151 0 -7.3290023295246284e-06
GC_1_152 b_1 NI_1 NS_152 0 -4.0590082157435106e-06
GC_1_153 b_1 NI_1 NS_153 0 -6.1708461647915095e-06
GC_1_154 b_1 NI_1 NS_154 0 4.5657990872758559e-06
GC_1_155 b_1 NI_1 NS_155 0 4.0300264557840970e-06
GC_1_156 b_1 NI_1 NS_156 0 2.8274381438762185e-06
GC_1_157 b_1 NI_1 NS_157 0 -1.1935950113433414e-11
GC_1_158 b_1 NI_1 NS_158 0 6.8028785277501750e-11
GC_1_159 b_1 NI_1 NS_159 0 1.8164619066710545e-10
GC_1_160 b_1 NI_1 NS_160 0 -4.3608434940568774e-10
GC_1_161 b_1 NI_1 NS_161 0 -2.6379397504985949e-11
GC_1_162 b_1 NI_1 NS_162 0 -2.3945833062785891e-10
GC_1_163 b_1 NI_1 NS_163 0 6.7099356444601829e-07
GC_1_164 b_1 NI_1 NS_164 0 -2.2973384328366014e-06
GC_1_165 b_1 NI_1 NS_165 0 -1.5909190974390131e-09
GC_1_166 b_1 NI_1 NS_166 0 5.3889759889166287e-11
GC_1_167 b_1 NI_1 NS_167 0 -7.3753147362260400e-12
GC_1_168 b_1 NI_1 NS_168 0 3.2536435323187612e-10
GC_1_169 b_1 NI_1 NS_169 0 4.0766811108705522e-06
GC_1_170 b_1 NI_1 NS_170 0 -4.1634910394737339e-06
GC_1_171 b_1 NI_1 NS_171 0 3.0280139604537012e-06
GC_1_172 b_1 NI_1 NS_172 0 -8.4376580933505429e-06
GC_1_173 b_1 NI_1 NS_173 0 -1.0871230944117084e-05
GC_1_174 b_1 NI_1 NS_174 0 -1.2340839467653628e-05
GC_1_175 b_1 NI_1 NS_175 0 6.1560076126403237e-11
GC_1_176 b_1 NI_1 NS_176 0 -1.1198994144125486e-11
GC_1_177 b_1 NI_1 NS_177 0 -5.2524152868685960e-10
GC_1_178 b_1 NI_1 NS_178 0 5.2973810639690023e-10
GC_1_179 b_1 NI_1 NS_179 0 -1.9706341172817356e-10
GC_1_180 b_1 NI_1 NS_180 0 7.7380223125124989e-12
GC_1_181 b_1 NI_1 NS_181 0 5.8596945022425887e-07
GC_1_182 b_1 NI_1 NS_182 0 -2.8556059314412193e-06
GC_1_183 b_1 NI_1 NS_183 0 1.7704154031574867e-09
GC_1_184 b_1 NI_1 NS_184 0 -6.7054019613483946e-11
GC_1_185 b_1 NI_1 NS_185 0 7.5216563176342434e-12
GC_1_186 b_1 NI_1 NS_186 0 -2.8672920896103194e-10
GC_1_187 b_1 NI_1 NS_187 0 -9.9035555185788565e-07
GC_1_188 b_1 NI_1 NS_188 0 -1.1238119875459322e-05
GC_1_189 b_1 NI_1 NS_189 0 -3.8449973488871253e-06
GC_1_190 b_1 NI_1 NS_190 0 -1.2011771404641650e-05
GC_1_191 b_1 NI_1 NS_191 0 -1.5709042024281371e-05
GC_1_192 b_1 NI_1 NS_192 0 -1.4372424485942816e-05
GC_1_193 b_1 NI_1 NS_193 0 2.7225434539004985e-12
GC_1_194 b_1 NI_1 NS_194 0 4.8461612283813171e-11
GC_1_195 b_1 NI_1 NS_195 0 -1.0541232496133611e-10
GC_1_196 b_1 NI_1 NS_196 0 9.2934561418944348e-11
GC_1_197 b_1 NI_1 NS_197 0 1.5681548503643336e-10
GC_1_198 b_1 NI_1 NS_198 0 -8.5158605070073025e-11
GC_1_199 b_1 NI_1 NS_199 0 -9.7454419163189595e-07
GC_1_200 b_1 NI_1 NS_200 0 4.1608356735359916e-06
GC_1_201 b_1 NI_1 NS_201 0 -1.1208172827678426e-09
GC_1_202 b_1 NI_1 NS_202 0 8.2924946636995707e-11
GC_1_203 b_1 NI_1 NS_203 0 -7.7974461733475224e-12
GC_1_204 b_1 NI_1 NS_204 0 1.3118859149727403e-10
GC_1_205 b_1 NI_1 NS_205 0 8.4582218013660493e-07
GC_1_206 b_1 NI_1 NS_206 0 1.3225653263079895e-05
GC_1_207 b_1 NI_1 NS_207 0 3.8098611417677385e-06
GC_1_208 b_1 NI_1 NS_208 0 1.4582517141434356e-05
GC_1_209 b_1 NI_1 NS_209 0 1.9310561717068431e-05
GC_1_210 b_1 NI_1 NS_210 0 1.9670561942202724e-05
GC_1_211 b_1 NI_1 NS_211 0 -1.5170747150491311e-11
GC_1_212 b_1 NI_1 NS_212 0 -6.4678331565679820e-11
GC_1_213 b_1 NI_1 NS_213 0 2.1121374280323579e-10
GC_1_214 b_1 NI_1 NS_214 0 -1.1076904753989782e-10
GC_1_215 b_1 NI_1 NS_215 0 -8.5473431200057612e-11
GC_1_216 b_1 NI_1 NS_216 0 1.5980371067075255e-10
GD_1_1 b_1 NI_1 NA_1 0 -9.3789092604744648e-02
GD_1_2 b_1 NI_1 NA_2 0 7.4536674973119402e-02
GD_1_3 b_1 NI_1 NA_3 0 6.2400713367368032e-03
GD_1_4 b_1 NI_1 NA_4 0 3.7902991565883109e-03
GD_1_5 b_1 NI_1 NA_5 0 6.4383450278311297e-05
GD_1_6 b_1 NI_1 NA_6 0 -3.4083347627935442e-05
GD_1_7 b_1 NI_1 NA_7 0 -5.4496394145185316e-05
GD_1_8 b_1 NI_1 NA_8 0 -1.8202757464802334e-05
GD_1_9 b_1 NI_1 NA_9 0 9.6627040244030115e-06
GD_1_10 b_1 NI_1 NA_10 0 -5.8537782160727097e-08
GD_1_11 b_1 NI_1 NA_11 0 1.3353180319101804e-05
GD_1_12 b_1 NI_1 NA_12 0 -1.5515465924102607e-05
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 1.0782410480686996e-02
GC_2_2 b_2 NI_2 NS_2 0 -2.9413305600417283e-02
GC_2_3 b_2 NI_2 NS_3 0 -1.0664792236619038e-05
GC_2_4 b_2 NI_2 NS_4 0 -6.9026185884417305e-07
GC_2_5 b_2 NI_2 NS_5 0 1.2414285312971826e-08
GC_2_6 b_2 NI_2 NS_6 0 8.5958463426413078e-06
GC_2_7 b_2 NI_2 NS_7 0 -5.1463058584844443e-02
GC_2_8 b_2 NI_2 NS_8 0 6.8753522893970534e-02
GC_2_9 b_2 NI_2 NS_9 0 -2.9075422515218115e-02
GC_2_10 b_2 NI_2 NS_10 0 -1.5435114137523198e-01
GC_2_11 b_2 NI_2 NS_11 0 -4.6623629674729444e-03
GC_2_12 b_2 NI_2 NS_12 0 -1.6535094380899537e-01
GC_2_13 b_2 NI_2 NS_13 0 4.7568788056070149e-07
GC_2_14 b_2 NI_2 NS_14 0 8.8283196705216141e-07
GC_2_15 b_2 NI_2 NS_15 0 -4.3323304344907134e-06
GC_2_16 b_2 NI_2 NS_16 0 1.0957949827620930e-07
GC_2_17 b_2 NI_2 NS_17 0 -3.3490001407832341e-06
GC_2_18 b_2 NI_2 NS_18 0 -3.5477335079791218e-06
GC_2_19 b_2 NI_2 NS_19 0 -4.7865465377251058e-03
GC_2_20 b_2 NI_2 NS_20 0 1.6712166529892217e-02
GC_2_21 b_2 NI_2 NS_21 0 -3.5265677047935449e-06
GC_2_22 b_2 NI_2 NS_22 0 2.9828686343710956e-08
GC_2_23 b_2 NI_2 NS_23 0 -1.0045935092873261e-09
GC_2_24 b_2 NI_2 NS_24 0 -2.0063946785455489e-06
GC_2_25 b_2 NI_2 NS_25 0 1.8824449668156443e-02
GC_2_26 b_2 NI_2 NS_26 0 5.0640142559262885e-02
GC_2_27 b_2 NI_2 NS_27 0 1.5094546986678739e-02
GC_2_28 b_2 NI_2 NS_28 0 7.1426549458562041e-02
GC_2_29 b_2 NI_2 NS_29 0 8.1524057415149329e-02
GC_2_30 b_2 NI_2 NS_30 0 4.9053274171792283e-02
GC_2_31 b_2 NI_2 NS_31 0 -2.7410735746156885e-07
GC_2_32 b_2 NI_2 NS_32 0 -6.0326930505102084e-08
GC_2_33 b_2 NI_2 NS_33 0 5.1949012715268090e-07
GC_2_34 b_2 NI_2 NS_34 0 -7.4351513905658013e-07
GC_2_35 b_2 NI_2 NS_35 0 3.9410170763469837e-07
GC_2_36 b_2 NI_2 NS_36 0 3.8363314435442651e-07
GC_2_37 b_2 NI_2 NS_37 0 1.1708109565208673e-04
GC_2_38 b_2 NI_2 NS_38 0 -4.6241831383685925e-04
GC_2_39 b_2 NI_2 NS_39 0 3.5664732150601587e-07
GC_2_40 b_2 NI_2 NS_40 0 3.4774181488935599e-09
GC_2_41 b_2 NI_2 NS_41 0 -1.1877247735382692e-11
GC_2_42 b_2 NI_2 NS_42 0 1.2106539863051880e-07
GC_2_43 b_2 NI_2 NS_43 0 7.0284696930866092e-04
GC_2_44 b_2 NI_2 NS_44 0 -4.2878428451726082e-03
GC_2_45 b_2 NI_2 NS_45 0 -9.0099177173569075e-03
GC_2_46 b_2 NI_2 NS_46 0 -5.1462862017371772e-03
GC_2_47 b_2 NI_2 NS_47 0 1.8367302588103561e-03
GC_2_48 b_2 NI_2 NS_48 0 7.2296615554471588e-03
GC_2_49 b_2 NI_2 NS_49 0 4.0526787785296381e-09
GC_2_50 b_2 NI_2 NS_50 0 2.5487030190121829e-09
GC_2_51 b_2 NI_2 NS_51 0 1.9540177945229166e-09
GC_2_52 b_2 NI_2 NS_52 0 1.2028729220866487e-08
GC_2_53 b_2 NI_2 NS_53 0 -2.5385461036114725e-08
GC_2_54 b_2 NI_2 NS_54 0 -1.4673550298745753e-08
GC_2_55 b_2 NI_2 NS_55 0 -6.0636875644129039e-04
GC_2_56 b_2 NI_2 NS_56 0 1.3735768115014728e-03
GC_2_57 b_2 NI_2 NS_57 0 -8.5902388733894404e-07
GC_2_58 b_2 NI_2 NS_58 0 -1.4354455574009933e-09
GC_2_59 b_2 NI_2 NS_59 0 -2.7334772697648768e-11
GC_2_60 b_2 NI_2 NS_60 0 -2.1419272170510560e-07
GC_2_61 b_2 NI_2 NS_61 0 -4.2054767110646972e-03
GC_2_62 b_2 NI_2 NS_62 0 1.9043221972858959e-02
GC_2_63 b_2 NI_2 NS_63 0 1.8780698047512562e-02
GC_2_64 b_2 NI_2 NS_64 0 -1.2054181128773839e-02
GC_2_65 b_2 NI_2 NS_65 0 2.1780333611006748e-03
GC_2_66 b_2 NI_2 NS_66 0 2.9274698322419815e-02
GC_2_67 b_2 NI_2 NS_67 0 -3.3667642354456613e-08
GC_2_68 b_2 NI_2 NS_68 0 -2.4503024043403115e-08
GC_2_69 b_2 NI_2 NS_69 0 8.1052950094942277e-08
GC_2_70 b_2 NI_2 NS_70 0 -4.2412456996812204e-08
GC_2_71 b_2 NI_2 NS_71 0 5.1503073976357350e-08
GC_2_72 b_2 NI_2 NS_72 0 3.1323534348126339e-08
GC_2_73 b_2 NI_2 NS_73 0 6.5711831312463610e-06
GC_2_74 b_2 NI_2 NS_74 0 -3.4967117490385278e-06
GC_2_75 b_2 NI_2 NS_75 0 2.4263945711147482e-08
GC_2_76 b_2 NI_2 NS_76 0 6.7556485236347844e-10
GC_2_77 b_2 NI_2 NS_77 0 -8.0408554272040409e-11
GC_2_78 b_2 NI_2 NS_78 0 4.3269205652088653e-09
GC_2_79 b_2 NI_2 NS_79 0 -1.3639461283628242e-04
GC_2_80 b_2 NI_2 NS_80 0 1.8279344955831757e-04
GC_2_81 b_2 NI_2 NS_81 0 8.0661863394303852e-04
GC_2_82 b_2 NI_2 NS_82 0 2.0572348479897722e-04
GC_2_83 b_2 NI_2 NS_83 0 -5.4635682903455987e-04
GC_2_84 b_2 NI_2 NS_84 0 -9.0504028560915283e-04
GC_2_85 b_2 NI_2 NS_85 0 -1.3851018517311760e-10
GC_2_86 b_2 NI_2 NS_86 0 8.7169044076948002e-10
GC_2_87 b_2 NI_2 NS_87 0 1.8473026916580891e-09
GC_2_88 b_2 NI_2 NS_88 0 -4.9674629176859042e-09
GC_2_89 b_2 NI_2 NS_89 0 -1.0292491196877651e-09
GC_2_90 b_2 NI_2 NS_90 0 6.3129988585486364e-10
GC_2_91 b_2 NI_2 NS_91 0 -1.3078365438743017e-05
GC_2_92 b_2 NI_2 NS_92 0 4.3753597273432148e-05
GC_2_93 b_2 NI_2 NS_93 0 -1.5372198942660393e-08
GC_2_94 b_2 NI_2 NS_94 0 -6.5434418201063975e-10
GC_2_95 b_2 NI_2 NS_95 0 8.0677079077556661e-11
GC_2_96 b_2 NI_2 NS_96 0 -4.9956381377037577e-09
GC_2_97 b_2 NI_2 NS_97 0 1.1875151156908245e-04
GC_2_98 b_2 NI_2 NS_98 0 1.7008892238497216e-04
GC_2_99 b_2 NI_2 NS_99 0 3.0495385905637894e-04
GC_2_100 b_2 NI_2 NS_100 0 -5.2260478203725274e-04
GC_2_101 b_2 NI_2 NS_101 0 -3.9414057344884664e-04
GC_2_102 b_2 NI_2 NS_102 0 1.6431869914228936e-04
GC_2_103 b_2 NI_2 NS_103 0 -2.3705730223716055e-10
GC_2_104 b_2 NI_2 NS_104 0 -8.7928231882679576e-10
GC_2_105 b_2 NI_2 NS_105 0 -1.0411019555184555e-09
GC_2_106 b_2 NI_2 NS_106 0 3.8717659985829839e-09
GC_2_107 b_2 NI_2 NS_107 0 1.2944564237383564e-09
GC_2_108 b_2 NI_2 NS_108 0 -4.9371263600189429e-10
GC_2_109 b_2 NI_2 NS_109 0 5.1102387575361105e-06
GC_2_110 b_2 NI_2 NS_110 0 -2.0595980508767141e-05
GC_2_111 b_2 NI_2 NS_111 0 -7.7535065338815083e-10
GC_2_112 b_2 NI_2 NS_112 0 2.0703880464965199e-10
GC_2_113 b_2 NI_2 NS_113 0 -2.4664140948453602e-11
GC_2_114 b_2 NI_2 NS_114 0 6.5797404362662767e-10
GC_2_115 b_2 NI_2 NS_115 0 -1.3889629173580577e-05
GC_2_116 b_2 NI_2 NS_116 0 4.5898379642033691e-05
GC_2_117 b_2 NI_2 NS_117 0 1.4542188831330818e-04
GC_2_118 b_2 NI_2 NS_118 0 3.4803298595955543e-05
GC_2_119 b_2 NI_2 NS_119 0 -7.6201453460450204e-05
GC_2_120 b_2 NI_2 NS_120 0 -1.9948388568258673e-04
GC_2_121 b_2 NI_2 NS_121 0 1.9462581418085919e-10
GC_2_122 b_2 NI_2 NS_122 0 1.5267342216832151e-10
GC_2_123 b_2 NI_2 NS_123 0 -2.8498988289114648e-10
GC_2_124 b_2 NI_2 NS_124 0 -3.9376045902798226e-10
GC_2_125 b_2 NI_2 NS_125 0 -2.7368354546716075e-10
GC_2_126 b_2 NI_2 NS_126 0 2.8376322807776944e-10
GC_2_127 b_2 NI_2 NS_127 0 1.0304670186020188e-06
GC_2_128 b_2 NI_2 NS_128 0 -6.3836436799975599e-06
GC_2_129 b_2 NI_2 NS_129 0 -3.8670306007312622e-09
GC_2_130 b_2 NI_2 NS_130 0 -2.4269284153493041e-10
GC_2_131 b_2 NI_2 NS_131 0 2.5054711783291381e-11
GC_2_132 b_2 NI_2 NS_132 0 -1.2071291267877685e-10
GC_2_133 b_2 NI_2 NS_133 0 -3.6740305593348157e-05
GC_2_134 b_2 NI_2 NS_134 0 5.6720743839828164e-05
GC_2_135 b_2 NI_2 NS_135 0 8.7520245999872645e-06
GC_2_136 b_2 NI_2 NS_136 0 1.4649196888079935e-04
GC_2_137 b_2 NI_2 NS_137 0 1.6051646263376678e-04
GC_2_138 b_2 NI_2 NS_138 0 5.6595682218046875e-05
GC_2_139 b_2 NI_2 NS_139 0 6.0843793861555569e-11
GC_2_140 b_2 NI_2 NS_140 0 -1.4081195895446384e-10
GC_2_141 b_2 NI_2 NS_141 0 -3.3787594787122105e-10
GC_2_142 b_2 NI_2 NS_142 0 1.0572116289366227e-09
GC_2_143 b_2 NI_2 NS_143 0 5.5311013342067337e-11
GC_2_144 b_2 NI_2 NS_144 0 -4.5394082896225587e-10
GC_2_145 b_2 NI_2 NS_145 0 6.7104908823048316e-07
GC_2_146 b_2 NI_2 NS_146 0 -2.2975393395064606e-06
GC_2_147 b_2 NI_2 NS_147 0 -1.5909903586403902e-09
GC_2_148 b_2 NI_2 NS_148 0 5.3888277040206272e-11
GC_2_149 b_2 NI_2 NS_149 0 -7.3752981830701296e-12
GC_2_150 b_2 NI_2 NS_150 0 3.2537974038642119e-10
GC_2_151 b_2 NI_2 NS_151 0 4.0765514432287245e-06
GC_2_152 b_2 NI_2 NS_152 0 -4.1640462436623751e-06
GC_2_153 b_2 NI_2 NS_153 0 3.0278765916453923e-06
GC_2_154 b_2 NI_2 NS_154 0 -8.4383609748999408e-06
GC_2_155 b_2 NI_2 NS_155 0 -1.0872150880383808e-05
GC_2_156 b_2 NI_2 NS_156 0 -1.2341723769055775e-05
GC_2_157 b_2 NI_2 NS_157 0 6.1561730573342052e-11
GC_2_158 b_2 NI_2 NS_158 0 -1.1197707666821573e-11
GC_2_159 b_2 NI_2 NS_159 0 -5.2525157451111569e-10
GC_2_160 b_2 NI_2 NS_160 0 5.2974150400871333e-10
GC_2_161 b_2 NI_2 NS_161 0 -1.9707045138737717e-10
GC_2_162 b_2 NI_2 NS_162 0 7.7308986573776761e-12
GC_2_163 b_2 NI_2 NS_163 0 4.0450231156575519e-07
GC_2_164 b_2 NI_2 NS_164 0 -1.0625285710591377e-06
GC_2_165 b_2 NI_2 NS_165 0 -6.0184136492519779e-10
GC_2_166 b_2 NI_2 NS_166 0 -1.0361784578982029e-10
GC_2_167 b_2 NI_2 NS_167 0 8.1965866313861958e-12
GC_2_168 b_2 NI_2 NS_168 0 1.6697163156359846e-10
GC_2_169 b_2 NI_2 NS_169 0 -7.3127907670235032e-06
GC_2_170 b_2 NI_2 NS_170 0 -4.1309640040880078e-06
GC_2_171 b_2 NI_2 NS_171 0 -6.1746465769244252e-06
GC_2_172 b_2 NI_2 NS_172 0 4.4531779061443692e-06
GC_2_173 b_2 NI_2 NS_173 0 3.8995689295721557e-06
GC_2_174 b_2 NI_2 NS_174 0 2.6656272628727077e-06
GC_2_175 b_2 NI_2 NS_175 0 -1.1522619372353912e-11
GC_2_176 b_2 NI_2 NS_176 0 6.7968294117652674e-11
GC_2_177 b_2 NI_2 NS_177 0 1.7905057087105897e-10
GC_2_178 b_2 NI_2 NS_178 0 -4.3368760539714664e-10
GC_2_179 b_2 NI_2 NS_179 0 -2.8731473623727338e-11
GC_2_180 b_2 NI_2 NS_180 0 -2.4192406761390867e-10
GC_2_181 b_2 NI_2 NS_181 0 -9.7408003267662358e-07
GC_2_182 b_2 NI_2 NS_182 0 4.1595782597732411e-06
GC_2_183 b_2 NI_2 NS_183 0 -1.1230101457792082e-09
GC_2_184 b_2 NI_2 NS_184 0 8.2869321198513029e-11
GC_2_185 b_2 NI_2 NS_185 0 -7.7963408404505366e-12
GC_2_186 b_2 NI_2 NS_186 0 1.3172460861073139e-10
GC_2_187 b_2 NI_2 NS_187 0 8.4635061412468342e-07
GC_2_188 b_2 NI_2 NS_188 0 1.3226720993935453e-05
GC_2_189 b_2 NI_2 NS_189 0 3.8130673810176548e-06
GC_2_190 b_2 NI_2 NS_190 0 1.4579715643851341e-05
GC_2_191 b_2 NI_2 NS_191 0 1.9307447860399675e-05
GC_2_192 b_2 NI_2 NS_192 0 1.9665926841288548e-05
GC_2_193 b_2 NI_2 NS_193 0 -1.5099173107863585e-11
GC_2_194 b_2 NI_2 NS_194 0 -6.4634077148166215e-11
GC_2_195 b_2 NI_2 NS_195 0 2.1080317750862075e-10
GC_2_196 b_2 NI_2 NS_196 0 -1.1068238332957600e-10
GC_2_197 b_2 NI_2 NS_197 0 -8.5719273095556411e-11
GC_2_198 b_2 NI_2 NS_198 0 1.5954466566314558e-10
GC_2_199 b_2 NI_2 NS_199 0 5.8599344741400634e-07
GC_2_200 b_2 NI_2 NS_200 0 -2.8557185776465872e-06
GC_2_201 b_2 NI_2 NS_201 0 1.7703517323275796e-09
GC_2_202 b_2 NI_2 NS_202 0 -6.7055574023739027e-11
GC_2_203 b_2 NI_2 NS_203 0 7.5216487856513055e-12
GC_2_204 b_2 NI_2 NS_204 0 -2.8671207878630399e-10
GC_2_205 b_2 NI_2 NS_205 0 -9.9060975926621147e-07
GC_2_206 b_2 NI_2 NS_206 0 -1.1239024566037076e-05
GC_2_207 b_2 NI_2 NS_207 0 -3.8455034598641233e-06
GC_2_208 b_2 NI_2 NS_208 0 -1.2012616934691704e-05
GC_2_209 b_2 NI_2 NS_209 0 -1.5710128493636216e-05
GC_2_210 b_2 NI_2 NS_210 0 -1.4373071512363962e-05
GC_2_211 b_2 NI_2 NS_211 0 2.7242231467112790e-12
GC_2_212 b_2 NI_2 NS_212 0 4.8464678376607991e-11
GC_2_213 b_2 NI_2 NS_213 0 -1.0542539833110668e-10
GC_2_214 b_2 NI_2 NS_214 0 9.2933547623341035e-11
GC_2_215 b_2 NI_2 NS_215 0 1.5680746618447291e-10
GC_2_216 b_2 NI_2 NS_216 0 -8.5166505523634738e-11
GD_2_1 b_2 NI_2 NA_1 0 7.4536168351202275e-02
GD_2_2 b_2 NI_2 NA_2 0 -9.3789092604231239e-02
GD_2_3 b_2 NI_2 NA_3 0 3.7903393781908165e-03
GD_2_4 b_2 NI_2 NA_4 0 6.2327127007393672e-03
GD_2_5 b_2 NI_2 NA_5 0 -3.4092191722670568e-05
GD_2_6 b_2 NI_2 NA_6 0 7.2422821820492618e-05
GD_2_7 b_2 NI_2 NA_7 0 -1.7748018752394321e-05
GD_2_8 b_2 NI_2 NA_8 0 -5.4411392401224562e-05
GD_2_9 b_2 NI_2 NA_9 0 -5.7714850132228616e-08
GD_2_10 b_2 NI_2 NA_10 0 9.7357563149062284e-06
GD_2_11 b_2 NI_2 NA_11 0 -1.5515985122160563e-05
GD_2_12 b_2 NI_2 NA_12 0 1.3354403657411739e-05
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 -6.0636875634466922e-04
GC_3_2 b_3 NI_3 NS_2 0 1.3735768111566543e-03
GC_3_3 b_3 NI_3 NS_3 0 -8.5902388739513535e-07
GC_3_4 b_3 NI_3 NS_4 0 -1.4354455576286112e-09
GC_3_5 b_3 NI_3 NS_5 0 -2.7334772687234125e-11
GC_3_6 b_3 NI_3 NS_6 0 -2.1419272169727367e-07
GC_3_7 b_3 NI_3 NS_7 0 -4.2054767103572536e-03
GC_3_8 b_3 NI_3 NS_8 0 1.9043221972435763e-02
GC_3_9 b_3 NI_3 NS_9 0 1.8780698047713533e-02
GC_3_10 b_3 NI_3 NS_10 0 -1.2054181129982211e-02
GC_3_11 b_3 NI_3 NS_11 0 2.1780333598461232e-03
GC_3_12 b_3 NI_3 NS_12 0 2.9274698320897328e-02
GC_3_13 b_3 NI_3 NS_13 0 -3.3667642348898674e-08
GC_3_14 b_3 NI_3 NS_14 0 -2.4503024045550231e-08
GC_3_15 b_3 NI_3 NS_15 0 8.1052950088758751e-08
GC_3_16 b_3 NI_3 NS_16 0 -4.2412456983507507e-08
GC_3_17 b_3 NI_3 NS_17 0 5.1503073973739800e-08
GC_3_18 b_3 NI_3 NS_18 0 3.1323534346362671e-08
GC_3_19 b_3 NI_3 NS_19 0 1.1707866780691721e-04
GC_3_20 b_3 NI_3 NS_20 0 -4.6241020402848195e-04
GC_3_21 b_3 NI_3 NS_21 0 3.5664998678139484e-07
GC_3_22 b_3 NI_3 NS_22 0 3.4774377332688928e-09
GC_3_23 b_3 NI_3 NS_23 0 -1.1877538575633464e-11
GC_3_24 b_3 NI_3 NS_24 0 1.2106504078807601e-07
GC_3_25 b_3 NI_3 NS_25 0 7.0283675803784590e-04
GC_3_26 b_3 NI_3 NS_26 0 -4.2878196445281028e-03
GC_3_27 b_3 NI_3 NS_27 0 -9.0099056624259079e-03
GC_3_28 b_3 NI_3 NS_28 0 -5.1462139024710174e-03
GC_3_29 b_3 NI_3 NS_29 0 1.8367936659892327e-03
GC_3_30 b_3 NI_3 NS_30 0 7.2296956127828457e-03
GC_3_31 b_3 NI_3 NS_31 0 4.0524566418956901e-09
GC_3_32 b_3 NI_3 NS_32 0 2.5486979450894868e-09
GC_3_33 b_3 NI_3 NS_33 0 1.9545768554604201e-09
GC_3_34 b_3 NI_3 NS_34 0 1.2028149426618535e-08
GC_3_35 b_3 NI_3 NS_35 0 -2.5385322697127474e-08
GC_3_36 b_3 NI_3 NS_36 0 -1.4673451662339173e-08
GC_3_37 b_3 NI_3 NS_37 0 -4.8626883259752724e-03
GC_3_38 b_3 NI_3 NS_38 0 1.6965719756401269e-02
GC_3_39 b_3 NI_3 NS_39 0 -3.4506329692844596e-06
GC_3_40 b_3 NI_3 NS_40 0 2.9325578711954448e-08
GC_3_41 b_3 NI_3 NS_41 0 -1.0119961826205942e-09
GC_3_42 b_3 NI_3 NS_42 0 -2.0011020526149260e-06
GC_3_43 b_3 NI_3 NS_43 0 1.8510240656206340e-02
GC_3_44 b_3 NI_3 NS_44 0 5.0676287657530239e-02
GC_3_45 b_3 NI_3 NS_45 0 1.4775416732760628e-02
GC_3_46 b_3 NI_3 NS_46 0 7.2026223569331180e-02
GC_3_47 b_3 NI_3 NS_47 0 8.2114599533252994e-02
GC_3_48 b_3 NI_3 NS_48 0 4.9909204215563635e-02
GC_3_49 b_3 NI_3 NS_49 0 -2.8707842539780792e-07
GC_3_50 b_3 NI_3 NS_50 0 -5.8614352254659196e-08
GC_3_51 b_3 NI_3 NS_51 0 5.7106092487621434e-07
GC_3_52 b_3 NI_3 NS_52 0 -8.2178280550852873e-07
GC_3_53 b_3 NI_3 NS_53 0 3.9091436190721690e-07
GC_3_54 b_3 NI_3 NS_54 0 3.8093864102298706e-07
GC_3_55 b_3 NI_3 NS_55 0 1.2611174725174036e-02
GC_3_56 b_3 NI_3 NS_56 0 -3.4717669517386987e-02
GC_3_57 b_3 NI_3 NS_57 0 -1.6765913514017171e-05
GC_3_58 b_3 NI_3 NS_58 0 -8.5089058310187521e-07
GC_3_59 b_3 NI_3 NS_59 0 1.4728338021106832e-08
GC_3_60 b_3 NI_3 NS_60 0 1.0166007186365942e-05
GC_3_61 b_3 NI_3 NS_61 0 -4.6985438706057495e-02
GC_3_62 b_3 NI_3 NS_62 0 6.7610304945433589e-02
GC_3_63 b_3 NI_3 NS_63 0 -2.4535617357435490e-02
GC_3_64 b_3 NI_3 NS_64 0 -1.6181720261821267e-01
GC_3_65 b_3 NI_3 NS_65 0 -1.3248647263166788e-02
GC_3_66 b_3 NI_3 NS_66 0 -1.8257613608942577e-01
GC_3_67 b_3 NI_3 NS_67 0 5.7586093799256161e-07
GC_3_68 b_3 NI_3 NS_68 0 1.0766200186064487e-06
GC_3_69 b_3 NI_3 NS_69 0 -5.4581323255530775e-06
GC_3_70 b_3 NI_3 NS_70 0 2.2863866937452269e-07
GC_3_71 b_3 NI_3 NS_71 0 -4.0768831848472039e-06
GC_3_72 b_3 NI_3 NS_72 0 -4.3109211712663880e-06
GC_3_73 b_3 NI_3 NS_73 0 -2.2359206710935147e-04
GC_3_74 b_3 NI_3 NS_74 0 6.5327047177650963e-04
GC_3_75 b_3 NI_3 NS_75 0 -1.5277950435825372e-07
GC_3_76 b_3 NI_3 NS_76 0 -6.5097059002430838e-10
GC_3_77 b_3 NI_3 NS_77 0 1.1967615935088974e-10
GC_3_78 b_3 NI_3 NS_78 0 -8.1075761199724464e-08
GC_3_79 b_3 NI_3 NS_79 0 -4.6134499543363659e-04
GC_3_80 b_3 NI_3 NS_80 0 4.9878481145899465e-03
GC_3_81 b_3 NI_3 NS_81 0 4.0331150028628370e-03
GC_3_82 b_3 NI_3 NS_82 0 -5.0048770185348547e-04
GC_3_83 b_3 NI_3 NS_83 0 2.5277456293818544e-03
GC_3_84 b_3 NI_3 NS_84 0 6.9902302348600395e-03
GC_3_85 b_3 NI_3 NS_85 0 -7.4379232386501925e-09
GC_3_86 b_3 NI_3 NS_86 0 -1.1207497198208686e-08
GC_3_87 b_3 NI_3 NS_87 0 7.8408265319679431e-09
GC_3_88 b_3 NI_3 NS_88 0 2.1821468104002567e-08
GC_3_89 b_3 NI_3 NS_89 0 2.3395567345534055e-08
GC_3_90 b_3 NI_3 NS_90 0 1.3793436735574507e-08
GC_3_91 b_3 NI_3 NS_91 0 1.3242491704093770e-04
GC_3_92 b_3 NI_3 NS_92 0 -4.8366411871300375e-04
GC_3_93 b_3 NI_3 NS_93 0 7.2243033208665290e-08
GC_3_94 b_3 NI_3 NS_94 0 5.7648710616434519e-10
GC_3_95 b_3 NI_3 NS_95 0 -1.2176376548656593e-10
GC_3_96 b_3 NI_3 NS_96 0 6.5848834543510473e-08
GC_3_97 b_3 NI_3 NS_97 0 -1.7773908794790558e-04
GC_3_98 b_3 NI_3 NS_98 0 -2.2254745015907523e-03
GC_3_99 b_3 NI_3 NS_99 0 -2.2112882456171087e-03
GC_3_100 b_3 NI_3 NS_100 0 -2.2412065124439396e-03
GC_3_101 b_3 NI_3 NS_101 0 -1.5818582732694212e-03
GC_3_102 b_3 NI_3 NS_102 0 -5.3366901910224991e-04
GC_3_103 b_3 NI_3 NS_103 0 1.3242676805379323e-09
GC_3_104 b_3 NI_3 NS_104 0 6.9372722146207733e-09
GC_3_105 b_3 NI_3 NS_105 0 9.2936715929580211e-09
GC_3_106 b_3 NI_3 NS_106 0 -2.8755168213444718e-08
GC_3_107 b_3 NI_3 NS_107 0 -1.9782456614524552e-08
GC_3_108 b_3 NI_3 NS_108 0 -1.2716700907363441e-08
GC_3_109 b_3 NI_3 NS_109 0 -1.2990464277700165e-05
GC_3_110 b_3 NI_3 NS_110 0 4.3509880019076327e-05
GC_3_111 b_3 NI_3 NS_111 0 -1.5810185763966997e-08
GC_3_112 b_3 NI_3 NS_112 0 -6.4981916496502167e-10
GC_3_113 b_3 NI_3 NS_113 0 8.0009744045139334e-11
GC_3_114 b_3 NI_3 NS_114 0 -4.9040885145742761e-09
GC_3_115 b_3 NI_3 NS_115 0 1.1939004375268689e-04
GC_3_116 b_3 NI_3 NS_116 0 1.6976512038719316e-04
GC_3_117 b_3 NI_3 NS_117 0 3.0498192253920932e-04
GC_3_118 b_3 NI_3 NS_118 0 -5.2326628672889593e-04
GC_3_119 b_3 NI_3 NS_119 0 -3.9475148092213148e-04
GC_3_120 b_3 NI_3 NS_120 0 1.6336796172319103e-04
GC_3_121 b_3 NI_3 NS_121 0 -2.3856253046178836e-10
GC_3_122 b_3 NI_3 NS_122 0 -8.7921366332752765e-10
GC_3_123 b_3 NI_3 NS_123 0 -1.0236139904153488e-09
GC_3_124 b_3 NI_3 NS_124 0 3.8234744996702970e-09
GC_3_125 b_3 NI_3 NS_125 0 1.2548481880321603e-09
GC_3_126 b_3 NI_3 NS_126 0 -5.0038262402873413e-10
GC_3_127 b_3 NI_3 NS_127 0 6.2564819578059246e-06
GC_3_128 b_3 NI_3 NS_128 0 -2.3560895237079116e-06
GC_3_129 b_3 NI_3 NS_129 0 2.4895469735885082e-08
GC_3_130 b_3 NI_3 NS_130 0 6.7282189251078040e-10
GC_3_131 b_3 NI_3 NS_131 0 -7.9766537881908715e-11
GC_3_132 b_3 NI_3 NS_132 0 4.2103474364728144e-09
GC_3_133 b_3 NI_3 NS_133 0 -1.3708369808850763e-04
GC_3_134 b_3 NI_3 NS_134 0 1.8383967135530039e-04
GC_3_135 b_3 NI_3 NS_135 0 8.0532283726682317e-04
GC_3_136 b_3 NI_3 NS_136 0 2.0770441225205586e-04
GC_3_137 b_3 NI_3 NS_137 0 -5.4316040170246393e-04
GC_3_138 b_3 NI_3 NS_138 0 -8.9973587935058088e-04
GC_3_139 b_3 NI_3 NS_139 0 -1.4772957654961670e-10
GC_3_140 b_3 NI_3 NS_140 0 8.7080771273600425e-10
GC_3_141 b_3 NI_3 NS_141 0 1.8594340082870834e-09
GC_3_142 b_3 NI_3 NS_142 0 -4.9461661422435308e-09
GC_3_143 b_3 NI_3 NS_143 0 -9.7957859381758325e-10
GC_3_144 b_3 NI_3 NS_144 0 6.4633909645210591e-10
GC_3_145 b_3 NI_3 NS_145 0 -8.0169986499449209e-07
GC_3_146 b_3 NI_3 NS_146 0 2.7307650799083838e-06
GC_3_147 b_3 NI_3 NS_147 0 -5.2077952321313074e-10
GC_3_148 b_3 NI_3 NS_148 0 -1.3300219593152615e-10
GC_3_149 b_3 NI_3 NS_149 0 1.4437311437648804e-11
GC_3_150 b_3 NI_3 NS_150 0 -3.0343762608982861e-10
GC_3_151 b_3 NI_3 NS_151 0 -1.8013126429123277e-06
GC_3_152 b_3 NI_3 NS_152 0 2.7925982229987677e-05
GC_3_153 b_3 NI_3 NS_153 0 1.0912795129530609e-05
GC_3_154 b_3 NI_3 NS_154 0 4.2540322559397984e-05
GC_3_155 b_3 NI_3 NS_155 0 4.9978014026861380e-05
GC_3_156 b_3 NI_3 NS_156 0 2.6934669267777181e-05
GC_3_157 b_3 NI_3 NS_157 0 7.0564929711755967e-11
GC_3_158 b_3 NI_3 NS_158 0 -1.8189062424113827e-10
GC_3_159 b_3 NI_3 NS_159 0 -4.0119657903600447e-10
GC_3_160 b_3 NI_3 NS_160 0 1.2111202668585052e-09
GC_3_161 b_3 NI_3 NS_161 0 1.8458101464620820e-10
GC_3_162 b_3 NI_3 NS_162 0 -1.7359411908560034e-10
GC_3_163 b_3 NI_3 NS_163 0 1.5476364182925616e-06
GC_3_164 b_3 NI_3 NS_164 0 -6.2962875331534304e-06
GC_3_165 b_3 NI_3 NS_165 0 1.2235133104465053e-10
GC_3_166 b_3 NI_3 NS_166 0 1.2886956722801027e-10
GC_3_167 b_3 NI_3 NS_167 0 -1.4440178858302458e-11
GC_3_168 b_3 NI_3 NS_168 0 3.5705197520635740e-10
GC_3_169 b_3 NI_3 NS_169 0 -6.9993933289431684e-06
GC_3_170 b_3 NI_3 NS_170 0 -7.1762888231539381e-06
GC_3_171 b_3 NI_3 NS_171 0 1.6282911358565252e-05
GC_3_172 b_3 NI_3 NS_172 0 -7.7564688156257738e-06
GC_3_173 b_3 NI_3 NS_173 0 -3.1226599586667204e-05
GC_3_174 b_3 NI_3 NS_174 0 -4.7428225172151745e-05
GC_3_175 b_3 NI_3 NS_175 0 -5.4189378623193555e-11
GC_3_176 b_3 NI_3 NS_176 0 1.7583912996407470e-10
GC_3_177 b_3 NI_3 NS_177 0 3.7769893498206312e-10
GC_3_178 b_3 NI_3 NS_178 0 -1.1564032435522056e-09
GC_3_179 b_3 NI_3 NS_179 0 -2.0765972924255901e-10
GC_3_180 b_3 NI_3 NS_180 0 1.5302906619195163e-10
GC_3_181 b_3 NI_3 NS_181 0 4.0746210733974930e-07
GC_3_182 b_3 NI_3 NS_182 0 -1.0805036659882631e-06
GC_3_183 b_3 NI_3 NS_183 0 -6.0121224378998832e-10
GC_3_184 b_3 NI_3 NS_184 0 -1.0370636439455633e-10
GC_3_185 b_3 NI_3 NS_185 0 8.2022262803007751e-12
GC_3_186 b_3 NI_3 NS_186 0 1.6745807659009921e-10
GC_3_187 b_3 NI_3 NS_187 0 -7.3117594023139070e-06
GC_3_188 b_3 NI_3 NS_188 0 -4.2280535930223904e-06
GC_3_189 b_3 NI_3 NS_189 0 -6.2102553912803706e-06
GC_3_190 b_3 NI_3 NS_190 0 4.3349178103283597e-06
GC_3_191 b_3 NI_3 NS_191 0 3.7519806082690861e-06
GC_3_192 b_3 NI_3 NS_192 0 2.5489723014392000e-06
GC_3_193 b_3 NI_3 NS_193 0 -1.1573370891636711e-11
GC_3_194 b_3 NI_3 NS_194 0 6.8390022789010385e-11
GC_3_195 b_3 NI_3 NS_195 0 1.7866341874961392e-10
GC_3_196 b_3 NI_3 NS_196 0 -4.3454381023805570e-10
GC_3_197 b_3 NI_3 NS_197 0 -2.8967394618542255e-11
GC_3_198 b_3 NI_3 NS_198 0 -2.4227178238092230e-10
GC_3_199 b_3 NI_3 NS_199 0 6.6414539997677040e-07
GC_3_200 b_3 NI_3 NS_200 0 -2.2652823003505864e-06
GC_3_201 b_3 NI_3 NS_201 0 -1.5864256251735155e-09
GC_3_202 b_3 NI_3 NS_202 0 5.4093436145299164e-11
GC_3_203 b_3 NI_3 NS_203 0 -7.3828945373005805e-12
GC_3_204 b_3 NI_3 NS_204 0 3.2373925189197344e-10
GC_3_205 b_3 NI_3 NS_205 0 4.0928296102177989e-06
GC_3_206 b_3 NI_3 NS_206 0 -3.9935320881232639e-06
GC_3_207 b_3 NI_3 NS_207 0 3.0987047498302454e-06
GC_3_208 b_3 NI_3 NS_208 0 -8.2597391007057612e-06
GC_3_209 b_3 NI_3 NS_209 0 -1.0642246301196316e-05
GC_3_210 b_3 NI_3 NS_210 0 -1.2162049103471475e-05
GC_3_211 b_3 NI_3 NS_211 0 6.1530393373177202e-11
GC_3_212 b_3 NI_3 NS_212 0 -1.1718198313874924e-11
GC_3_213 b_3 NI_3 NS_213 0 -5.2416371972375901e-10
GC_3_214 b_3 NI_3 NS_214 0 5.3037974278189149e-10
GC_3_215 b_3 NI_3 NS_215 0 -1.9630603186332797e-10
GC_3_216 b_3 NI_3 NS_216 0 8.6276851069324569e-12
GD_3_1 b_3 NI_3 NA_1 0 6.2327127007395953e-03
GD_3_2 b_3 NI_3 NA_2 0 3.7902991566286402e-03
GD_3_3 b_3 NI_3 NA_3 0 -9.3789392131004401e-02
GD_3_4 b_3 NI_3 NA_4 0 7.4456377535855225e-02
GD_3_5 b_3 NI_3 NA_5 0 -9.9162073087721262e-04
GD_3_6 b_3 NI_3 NA_6 0 2.6229987570646537e-03
GD_3_7 b_3 NI_3 NA_7 0 7.1974323158429458e-05
GD_3_8 b_3 NI_3 NA_8 0 -3.4701755055094225e-05
GD_3_9 b_3 NI_3 NA_9 0 -3.3983508248290876e-05
GD_3_10 b_3 NI_3 NA_10 0 1.8947982389611628e-05
GD_3_11 b_3 NI_3 NA_11 0 9.8463603951161484e-06
GD_3_12 b_3 NI_3 NA_12 0 -2.5590889931360315e-07
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 1.1708109564376630e-04
GC_4_2 b_4 NI_4 NS_2 0 -4.6241831380719890e-04
GC_4_3 b_4 NI_4 NS_3 0 3.5664732151082188e-07
GC_4_4 b_4 NI_4 NS_4 0 3.4774181489280930e-09
GC_4_5 b_4 NI_4 NS_5 0 -1.1877247736348004e-11
GC_4_6 b_4 NI_4 NS_6 0 1.2106539862983940e-07
GC_4_7 b_4 NI_4 NS_7 0 7.0284696924814650e-04
GC_4_8 b_4 NI_4 NS_8 0 -4.2878428451365528e-03
GC_4_9 b_4 NI_4 NS_9 0 -9.0099177173743709e-03
GC_4_10 b_4 NI_4 NS_10 0 -5.1462862016338120e-03
GC_4_11 b_4 NI_4 NS_11 0 1.8367302589177494e-03
GC_4_12 b_4 NI_4 NS_12 0 7.2296615555779032e-03
GC_4_13 b_4 NI_4 NS_13 0 4.0526787780446406e-09
GC_4_14 b_4 NI_4 NS_14 0 2.5487030191953554e-09
GC_4_15 b_4 NI_4 NS_15 0 1.9540177950582807e-09
GC_4_16 b_4 NI_4 NS_16 0 1.2028729219708990e-08
GC_4_17 b_4 NI_4 NS_17 0 -2.5385461035878589e-08
GC_4_18 b_4 NI_4 NS_18 0 -1.4673550298567307e-08
GC_4_19 b_4 NI_4 NS_19 0 -6.0598290779824383e-04
GC_4_20 b_4 NI_4 NS_20 0 1.3722647389125848e-03
GC_4_21 b_4 NI_4 NS_21 0 -8.5960949106912584e-07
GC_4_22 b_4 NI_4 NS_22 0 -1.4388097127360788e-09
GC_4_23 b_4 NI_4 NS_23 0 -2.7334249758175003e-11
GC_4_24 b_4 NI_4 NS_24 0 -2.1412823487297010e-07
GC_4_25 b_4 NI_4 NS_25 0 -4.2068464567719009e-03
GC_4_26 b_4 NI_4 NS_26 0 1.9038017951611245e-02
GC_4_27 b_4 NI_4 NS_27 0 1.8778280881652537e-02
GC_4_28 b_4 NI_4 NS_28 0 -1.2058896276377270e-02
GC_4_29 b_4 NI_4 NS_29 0 2.1714548174835454e-03
GC_4_30 b_4 NI_4 NS_30 0 2.9269113250972444e-02
GC_4_31 b_4 NI_4 NS_31 0 -3.3659898646673073e-08
GC_4_32 b_4 NI_4 NS_32 0 -2.4511752867259209e-08
GC_4_33 b_4 NI_4 NS_33 0 8.1060534674425464e-08
GC_4_34 b_4 NI_4 NS_34 0 -4.2241276218096799e-08
GC_4_35 b_4 NI_4 NS_35 0 5.1476165042444702e-08
GC_4_36 b_4 NI_4 NS_36 0 3.1306639609588944e-08
GC_4_37 b_4 NI_4 NS_37 0 1.2611136383820849e-02
GC_4_38 b_4 NI_4 NS_38 0 -3.4717584844479586e-02
GC_4_39 b_4 NI_4 NS_39 0 -1.6765740282276048e-05
GC_4_40 b_4 NI_4 NS_40 0 -8.5088586670793262e-07
GC_4_41 b_4 NI_4 NS_41 0 1.4728262665387141e-08
GC_4_42 b_4 NI_4 NS_42 0 1.0165961568991357e-05
GC_4_43 b_4 NI_4 NS_43 0 -4.6985722366427583e-02
GC_4_44 b_4 NI_4 NS_44 0 6.7609738613395462e-02
GC_4_45 b_4 NI_4 NS_45 0 -2.4536168456979913e-02
GC_4_46 b_4 NI_4 NS_46 0 -1.6181725141958922e-01
GC_4_47 b_4 NI_4 NS_47 0 -1.3248829745364022e-02
GC_4_48 b_4 NI_4 NS_48 0 -1.8257594939387672e-01
GC_4_49 b_4 NI_4 NS_49 0 5.7586032912638616e-07
GC_4_50 b_4 NI_4 NS_50 0 1.0766141356238244e-06
GC_4_51 b_4 NI_4 NS_51 0 -5.4581027524662791e-06
GC_4_52 b_4 NI_4 NS_52 0 2.2864077193343675e-07
GC_4_53 b_4 NI_4 NS_53 0 -4.0768620351751778e-06
GC_4_54 b_4 NI_4 NS_54 0 -4.3108988860352629e-06
GC_4_55 b_4 NI_4 NS_55 0 -4.8626883259710197e-03
GC_4_56 b_4 NI_4 NS_56 0 1.6965719756386666e-02
GC_4_57 b_4 NI_4 NS_57 0 -3.4506329692882238e-06
GC_4_58 b_4 NI_4 NS_58 0 2.9325578711936746e-08
GC_4_59 b_4 NI_4 NS_59 0 -1.0119961826227585e-09
GC_4_60 b_4 NI_4 NS_60 0 -2.0011020526144407e-06
GC_4_61 b_4 NI_4 NS_61 0 1.8510240656232177e-02
GC_4_62 b_4 NI_4 NS_62 0 5.0676287657515910e-02
GC_4_63 b_4 NI_4 NS_63 0 1.4775416732770332e-02
GC_4_64 b_4 NI_4 NS_64 0 7.2026223569286923e-02
GC_4_65 b_4 NI_4 NS_65 0 8.2114599533206420e-02
GC_4_66 b_4 NI_4 NS_66 0 4.9909204215502607e-02
GC_4_67 b_4 NI_4 NS_67 0 -2.8707842539751151e-07
GC_4_68 b_4 NI_4 NS_68 0 -5.8614352254655484e-08
GC_4_69 b_4 NI_4 NS_69 0 5.7106092487563857e-07
GC_4_70 b_4 NI_4 NS_70 0 -8.2178280550785089e-07
GC_4_71 b_4 NI_4 NS_71 0 3.9091436190702447e-07
GC_4_72 b_4 NI_4 NS_72 0 3.8093864102286652e-07
GC_4_73 b_4 NI_4 NS_73 0 1.3239366494649006e-04
GC_4_74 b_4 NI_4 NS_74 0 -4.8355778816134572e-04
GC_4_75 b_4 NI_4 NS_75 0 7.2278915701689853e-08
GC_4_76 b_4 NI_4 NS_76 0 5.7679787197920801e-10
GC_4_77 b_4 NI_4 NS_77 0 -1.2176774255259678e-10
GC_4_78 b_4 NI_4 NS_78 0 6.5843860469707456e-08
GC_4_79 b_4 NI_4 NS_79 0 -1.7783318424575338e-04
GC_4_80 b_4 NI_4 NS_80 0 -2.2251263872467191e-03
GC_4_81 b_4 NI_4 NS_81 0 -2.2111072263042136e-03
GC_4_82 b_4 NI_4 NS_82 0 -2.2403140914600671e-03
GC_4_83 b_4 NI_4 NS_83 0 -1.5810437559492698e-03
GC_4_84 b_4 NI_4 NS_84 0 -5.3321630765743001e-04
GC_4_85 b_4 NI_4 NS_85 0 1.3213977138885173e-09
GC_4_86 b_4 NI_4 NS_86 0 6.9371668139467860e-09
GC_4_87 b_4 NI_4 NS_87 0 9.3010342295642600e-09
GC_4_88 b_4 NI_4 NS_88 0 -2.8761363192219045e-08
GC_4_89 b_4 NI_4 NS_89 0 -1.9780396578401179e-08
GC_4_90 b_4 NI_4 NS_90 0 -1.2715079304788585e-08
GC_4_91 b_4 NI_4 NS_91 0 -2.2363248175853530e-04
GC_4_92 b_4 NI_4 NS_92 0 6.5341466351937058e-04
GC_4_93 b_4 NI_4 NS_93 0 -1.5273961825249956e-07
GC_4_94 b_4 NI_4 NS_94 0 -6.5079447719969996e-10
GC_4_95 b_4 NI_4 NS_95 0 1.1967462903414086e-10
GC_4_96 b_4 NI_4 NS_96 0 -8.1079865815348034e-08
GC_4_97 b_4 NI_4 NS_97 0 -4.6122744314804997e-04
GC_4_98 b_4 NI_4 NS_98 0 4.9884965147784710e-03
GC_4_99 b_4 NI_4 NS_99 0 4.0334339333771476e-03
GC_4_100 b_4 NI_4 NS_100 0 -4.9985991122877479e-04
GC_4_101 b_4 NI_4 NS_101 0 2.5285439398216418e-03
GC_4_102 b_4 NI_4 NS_102 0 6.9908496831149452e-03
GC_4_103 b_4 NI_4 NS_103 0 -7.4399096477826779e-09
GC_4_104 b_4 NI_4 NS_104 0 -1.1207975533300037e-08
GC_4_105 b_4 NI_4 NS_105 0 7.8472969261246859e-09
GC_4_106 b_4 NI_4 NS_106 0 2.1817007640760425e-08
GC_4_107 b_4 NI_4 NS_107 0 2.3397158971448120e-08
GC_4_108 b_4 NI_4 NS_108 0 1.3794434681988384e-08
GC_4_109 b_4 NI_4 NS_109 0 6.2533809938194054e-06
GC_4_110 b_4 NI_4 NS_110 0 -2.3445367305967620e-06
GC_4_111 b_4 NI_4 NS_111 0 2.4898512698483608e-08
GC_4_112 b_4 NI_4 NS_112 0 6.7283793529940405e-10
GC_4_113 b_4 NI_4 NS_113 0 -7.9766645295822504e-11
GC_4_114 b_4 NI_4 NS_114 0 4.2099990044708134e-09
GC_4_115 b_4 NI_4 NS_115 0 -1.3708326491444222e-04
GC_4_116 b_4 NI_4 NS_116 0 1.8387583637659538e-04
GC_4_117 b_4 NI_4 NS_117 0 8.0533408208258953e-04
GC_4_118 b_4 NI_4 NS_118 0 2.0774810288201181e-04
GC_4_119 b_4 NI_4 NS_119 0 -5.4310540531146592e-04
GC_4_120 b_4 NI_4 NS_120 0 -8.9968373095346266e-04
GC_4_121 b_4 NI_4 NS_121 0 -1.4790326283606715e-10
GC_4_122 b_4 NI_4 NS_122 0 8.7078171588710349e-10
GC_4_123 b_4 NI_4 NS_123 0 1.8598920359696891e-09
GC_4_124 b_4 NI_4 NS_124 0 -4.9466048890176315e-09
GC_4_125 b_4 NI_4 NS_125 0 -9.7944056976940514e-10
GC_4_126 b_4 NI_4 NS_126 0 6.4642666606814343e-10
GC_4_127 b_4 NI_4 NS_127 0 -1.3609002222117616e-05
GC_4_128 b_4 NI_4 NS_128 0 4.5664437320699946e-05
GC_4_129 b_4 NI_4 NS_129 0 -1.5015648345396538e-08
GC_4_130 b_4 NI_4 NS_130 0 -6.4639585047225073e-10
GC_4_131 b_4 NI_4 NS_131 0 7.9993998875343883e-11
GC_4_132 b_4 NI_4 NS_132 0 -4.9849997553681023e-09
GC_4_133 b_4 NI_4 NS_133 0 1.1994564514947637e-04
GC_4_134 b_4 NI_4 NS_134 0 1.7720715321639459e-04
GC_4_135 b_4 NI_4 NS_135 0 3.0879688681577713e-04
GC_4_136 b_4 NI_4 NS_136 0 -5.1565674750258660e-04
GC_4_137 b_4 NI_4 NS_137 0 -3.8587539985750051e-04
GC_4_138 b_4 NI_4 NS_138 0 1.7143573273994210e-04
GC_4_139 b_4 NI_4 NS_139 0 -2.6845101187407998e-10
GC_4_140 b_4 NI_4 NS_140 0 -8.7537391247304917e-10
GC_4_141 b_4 NI_4 NS_141 0 -9.6027733207034458e-10
GC_4_142 b_4 NI_4 NS_142 0 3.6739414245625351e-09
GC_4_143 b_4 NI_4 NS_143 0 1.2872832528716277e-09
GC_4_144 b_4 NI_4 NS_144 0 -4.7972492190722762e-10
GC_4_145 b_4 NI_4 NS_145 0 1.5414273439519771e-06
GC_4_146 b_4 NI_4 NS_146 0 -6.2760737915059991e-06
GC_4_147 b_4 NI_4 NS_147 0 1.3208736233924377e-10
GC_4_148 b_4 NI_4 NS_148 0 1.2903217966242287e-10
GC_4_149 b_4 NI_4 NS_149 0 -1.4443364790649296e-11
GC_4_150 b_4 NI_4 NS_150 0 3.5536535331182474e-10
GC_4_151 b_4 NI_4 NS_151 0 -7.0220257778121357e-06
GC_4_152 b_4 NI_4 NS_152 0 -7.1280529206086447e-06
GC_4_153 b_4 NI_4 NS_153 0 1.6303010788766503e-05
GC_4_154 b_4 NI_4 NS_154 0 -7.6034204704097774e-06
GC_4_155 b_4 NI_4 NS_155 0 -3.1089982587909048e-05
GC_4_156 b_4 NI_4 NS_156 0 -4.7345834308877174e-05
GC_4_157 b_4 NI_4 NS_157 0 -5.4798180522826295e-11
GC_4_158 b_4 NI_4 NS_158 0 1.7570990142140829e-10
GC_4_159 b_4 NI_4 NS_159 0 3.7966195633534773e-10
GC_4_160 b_4 NI_4 NS_160 0 -1.1576231308759438e-09
GC_4_161 b_4 NI_4 NS_161 0 -2.0690964279086397e-10
GC_4_162 b_4 NI_4 NS_162 0 1.5378523530834345e-10
GC_4_163 b_4 NI_4 NS_163 0 -8.0171136867198748e-07
GC_4_164 b_4 NI_4 NS_164 0 2.7308205519211177e-06
GC_4_165 b_4 NI_4 NS_165 0 -5.2075744271267113e-10
GC_4_166 b_4 NI_4 NS_166 0 -1.3300183420490835e-10
GC_4_167 b_4 NI_4 NS_167 0 1.4437315397803151e-11
GC_4_168 b_4 NI_4 NS_168 0 -3.0344217626950796e-10
GC_4_169 b_4 NI_4 NS_169 0 -1.8011838468522169e-06
GC_4_170 b_4 NI_4 NS_170 0 2.7926444846262050e-05
GC_4_171 b_4 NI_4 NS_171 0 1.0913058616206197e-05
GC_4_172 b_4 NI_4 NS_172 0 4.2540761936378834e-05
GC_4_173 b_4 NI_4 NS_173 0 4.9978562134236052e-05
GC_4_174 b_4 NI_4 NS_174 0 2.6934982437077549e-05
GC_4_175 b_4 NI_4 NS_175 0 7.0562614215468035e-11
GC_4_176 b_4 NI_4 NS_176 0 -1.8189059678516642e-10
GC_4_177 b_4 NI_4 NS_177 0 -4.0119182425100016e-10
GC_4_178 b_4 NI_4 NS_178 0 1.2111185518084927e-09
GC_4_179 b_4 NI_4 NS_179 0 1.8458305042405281e-10
GC_4_180 b_4 NI_4 NS_180 0 -1.7359226241488985e-10
GC_4_181 b_4 NI_4 NS_181 0 6.6412956427279364e-07
GC_4_182 b_4 NI_4 NS_182 0 -2.2652194401398076e-06
GC_4_183 b_4 NI_4 NS_183 0 -1.5864167346743775e-09
GC_4_184 b_4 NI_4 NS_184 0 5.4093612276103371e-11
GC_4_185 b_4 NI_4 NS_185 0 -7.3828932534736797e-12
GC_4_186 b_4 NI_4 NS_186 0 3.2373731834786106e-10
GC_4_187 b_4 NI_4 NS_187 0 4.0928042113082752e-06
GC_4_188 b_4 NI_4 NS_188 0 -3.9933766922049704e-06
GC_4_189 b_4 NI_4 NS_189 0 3.0987413544340247e-06
GC_4_190 b_4 NI_4 NS_190 0 -8.2595770901310379e-06
GC_4_191 b_4 NI_4 NS_191 0 -1.0642019081641338e-05
GC_4_192 b_4 NI_4 NS_192 0 -1.2161765012658572e-05
GC_4_193 b_4 NI_4 NS_193 0 6.1530274780047457e-11
GC_4_194 b_4 NI_4 NS_194 0 -1.1718474525718978e-11
GC_4_195 b_4 NI_4 NS_195 0 -5.2416217247769599e-10
GC_4_196 b_4 NI_4 NS_196 0 5.3037942008247154e-10
GC_4_197 b_4 NI_4 NS_197 0 -1.9630513334187105e-10
GC_4_198 b_4 NI_4 NS_198 0 8.6285826794268965e-12
GC_4_199 b_4 NI_4 NS_199 0 3.9250794794292441e-07
GC_4_200 b_4 NI_4 NS_200 0 -1.0348236151393933e-06
GC_4_201 b_4 NI_4 NS_201 0 -5.7480797697654443e-10
GC_4_202 b_4 NI_4 NS_202 0 -1.0318287067730907e-10
GC_4_203 b_4 NI_4 NS_203 0 8.1893937169926084e-12
GC_4_204 b_4 NI_4 NS_204 0 1.6240283667321871e-10
GC_4_205 b_4 NI_4 NS_205 0 -7.3298750323623081e-06
GC_4_206 b_4 NI_4 NS_206 0 -4.1640115958354067e-06
GC_4_207 b_4 NI_4 NS_207 0 -6.2106532648643382e-06
GC_4_208 b_4 NI_4 NS_208 0 4.4397893323355971e-06
GC_4_209 b_4 NI_4 NS_209 0 3.8725824535074292e-06
GC_4_210 b_4 NI_4 NS_210 0 2.7044156420654563e-06
GC_4_211 b_4 NI_4 NS_211 0 -1.1963601600545487e-11
GC_4_212 b_4 NI_4 NS_212 0 6.8480093006090971e-11
GC_4_213 b_4 NI_4 NS_213 0 1.8113600624298062e-10
GC_4_214 b_4 NI_4 NS_214 0 -4.3693334515538942e-10
GC_4_215 b_4 NI_4 NS_215 0 -2.6690031564613229e-11
GC_4_216 b_4 NI_4 NS_216 0 -2.3988041240838342e-10
GD_4_1 b_4 NI_4 NA_1 0 3.7903393781908165e-03
GD_4_2 b_4 NI_4 NA_2 0 6.2400713367366870e-03
GD_4_3 b_4 NI_4 NA_3 0 7.4457050476455872e-02
GD_4_4 b_4 NI_4 NA_4 0 -9.3789392131004248e-02
GD_4_5 b_4 NI_4 NA_5 0 2.6224377111535566e-03
GD_4_6 b_4 NI_4 NA_6 0 -9.9243574060401329e-04
GD_4_7 b_4 NI_4 NA_7 0 -3.4744597854691349e-05
GD_4_8 b_4 NI_4 NA_8 0 6.3682781141481622e-05
GD_4_9 b_4 NI_4 NA_9 0 1.8865361145708455e-05
GD_4_10 b_4 NI_4 NA_10 0 -3.3984119310117821e-05
GD_4_11 b_4 NI_4 NA_11 0 -2.5606532833499595e-07
GD_4_12 b_4 NI_4 NA_12 0 9.7838301411621909e-06
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 -1.3078365367187723e-05
GC_5_2 b_5 NI_5 NS_2 0 4.3753597075118879e-05
GC_5_3 b_5 NI_5 NS_3 0 -1.5372198914690025e-08
GC_5_4 b_5 NI_5 NS_4 0 -6.5434418688440374e-10
GC_5_5 b_5 NI_5 NS_5 0 8.0677078721593236e-11
GC_5_6 b_5 NI_5 NS_6 0 -4.9956381312586253e-09
GC_5_7 b_5 NI_5 NS_7 0 1.1875151188808364e-04
GC_5_8 b_5 NI_5 NS_8 0 1.7008892293002135e-04
GC_5_9 b_5 NI_5 NS_9 0 3.0495385963946026e-04
GC_5_10 b_5 NI_5 NS_10 0 -5.2260478184642134e-04
GC_5_11 b_5 NI_5 NS_11 0 -3.9414057318998806e-04
GC_5_12 b_5 NI_5 NS_12 0 1.6431869863871190e-04
GC_5_13 b_5 NI_5 NS_13 0 -2.3705728717642289e-10
GC_5_14 b_5 NI_5 NS_14 0 -8.7928232185207526e-10
GC_5_15 b_5 NI_5 NS_15 0 -1.0411019509541986e-09
GC_5_16 b_5 NI_5 NS_16 0 3.8717660430405190e-09
GC_5_17 b_5 NI_5 NS_17 0 1.2944564122635020e-09
GC_5_18 b_5 NI_5 NS_18 0 -4.9371266752411757e-10
GC_5_19 b_5 NI_5 NS_19 0 6.5717423209599140e-06
GC_5_20 b_5 NI_5 NS_20 0 -3.4988226085281561e-06
GC_5_21 b_5 NI_5 NS_21 0 2.4262979337052697e-08
GC_5_22 b_5 NI_5 NS_22 0 6.7555753328228767e-10
GC_5_23 b_5 NI_5 NS_23 0 -8.0408494665599468e-11
GC_5_24 b_5 NI_5 NS_24 0 4.3270565340613458e-09
GC_5_25 b_5 NI_5 NS_25 0 -1.3639333442874482e-04
GC_5_26 b_5 NI_5 NS_26 0 1.8277823931482946e-04
GC_5_27 b_5 NI_5 NS_27 0 8.0660338517502808e-04
GC_5_28 b_5 NI_5 NS_28 0 2.0572608884732993e-04
GC_5_29 b_5 NI_5 NS_29 0 -5.4635656223464113e-04
GC_5_30 b_5 NI_5 NS_30 0 -9.0504419758937144e-04
GC_5_31 b_5 NI_5 NS_31 0 -1.3840410156070284e-10
GC_5_32 b_5 NI_5 NS_32 0 8.7166071979194378e-10
GC_5_33 b_5 NI_5 NS_33 0 1.8468558113343487e-09
GC_5_34 b_5 NI_5 NS_34 0 -4.9672058721568998e-09
GC_5_35 b_5 NI_5 NS_35 0 -1.0293053731582052e-09
GC_5_36 b_5 NI_5 NS_36 0 6.3126224015232469e-10
GC_5_37 b_5 NI_5 NS_37 0 -2.2363248172180118e-04
GC_5_38 b_5 NI_5 NS_38 0 6.5341466339564121e-04
GC_5_39 b_5 NI_5 NS_39 0 -1.5273961829068714e-07
GC_5_40 b_5 NI_5 NS_40 0 -6.5079447739692815e-10
GC_5_41 b_5 NI_5 NS_41 0 1.1967462903762146e-10
GC_5_42 b_5 NI_5 NS_42 0 -8.1079865810432398e-08
GC_5_43 b_5 NI_5 NS_43 0 -4.6122744294295318e-04
GC_5_44 b_5 NI_5 NS_44 0 4.9884965146705434e-03
GC_5_45 b_5 NI_5 NS_45 0 4.0334339334639957e-03
GC_5_46 b_5 NI_5 NS_46 0 -4.9985991157901080e-04
GC_5_47 b_5 NI_5 NS_47 0 2.5285439394510632e-03
GC_5_48 b_5 NI_5 NS_48 0 6.9908496826111876e-03
GC_5_49 b_5 NI_5 NS_49 0 -7.4399096450958059e-09
GC_5_50 b_5 NI_5 NS_50 0 -1.1207975532879987e-08
GC_5_51 b_5 NI_5 NS_51 0 7.8472969199084666e-09
GC_5_52 b_5 NI_5 NS_52 0 2.1817007646875351e-08
GC_5_53 b_5 NI_5 NS_53 0 2.3397158969594232e-08
GC_5_54 b_5 NI_5 NS_54 0 1.3794434680795515e-08
GC_5_55 b_5 NI_5 NS_55 0 1.3242491921877406e-04
GC_5_56 b_5 NI_5 NS_56 0 -4.8366412486883448e-04
GC_5_57 b_5 NI_5 NS_57 0 7.2243028321027038e-08
GC_5_58 b_5 NI_5 NS_58 0 5.7648708570018873e-10
GC_5_59 b_5 NI_5 NS_59 0 -1.2176376529740268e-10
GC_5_60 b_5 NI_5 NS_60 0 6.5848834933224826e-08
GC_5_61 b_5 NI_5 NS_61 0 -1.7773908582146224e-04
GC_5_62 b_5 NI_5 NS_62 0 -2.2254745070497245e-03
GC_5_63 b_5 NI_5 NS_63 0 -2.2112882443942878e-03
GC_5_64 b_5 NI_5 NS_64 0 -2.2412065218593846e-03
GC_5_65 b_5 NI_5 NS_65 0 -1.5818582845621846e-03
GC_5_66 b_5 NI_5 NS_66 0 -5.3366903770264446e-04
GC_5_67 b_5 NI_5 NS_67 0 1.3242674540584287e-09
GC_5_68 b_5 NI_5 NS_68 0 6.9372728817838282e-09
GC_5_69 b_5 NI_5 NS_69 0 9.2936700044859355e-09
GC_5_70 b_5 NI_5 NS_70 0 -2.8755166423538333e-08
GC_5_71 b_5 NI_5 NS_71 0 -1.9782456762722687e-08
GC_5_72 b_5 NI_5 NS_72 0 -1.2716701007702126e-08
GC_5_73 b_5 NI_5 NS_73 0 -4.8322138401050560e-03
GC_5_74 b_5 NI_5 NS_74 0 1.6839927410549200e-02
GC_5_75 b_5 NI_5 NS_75 0 -3.4885576289392676e-06
GC_5_76 b_5 NI_5 NS_76 0 2.9143693123682918e-08
GC_5_77 b_5 NI_5 NS_77 0 -1.0018331264047442e-09
GC_5_78 b_5 NI_5 NS_78 0 -1.9968125735067089e-06
GC_5_79 b_5 NI_5 NS_79 0 1.8660666931426807e-02
GC_5_80 b_5 NI_5 NS_80 0 5.0341742983245751e-02
GC_5_81 b_5 NI_5 NS_81 0 1.4759545324540104e-02
GC_5_82 b_5 NI_5 NS_82 0 7.1489778072348298e-02
GC_5_83 b_5 NI_5 NS_83 0 8.1469900017250768e-02
GC_5_84 b_5 NI_5 NS_84 0 4.9245596332448328e-02
GC_5_85 b_5 NI_5 NS_85 0 -2.8743021846691931e-07
GC_5_86 b_5 NI_5 NS_86 0 -5.6953706962365285e-08
GC_5_87 b_5 NI_5 NS_87 0 5.7215241455416153e-07
GC_5_88 b_5 NI_5 NS_88 0 -8.2970936192604349e-07
GC_5_89 b_5 NI_5 NS_89 0 3.8940708076447761e-07
GC_5_90 b_5 NI_5 NS_90 0 3.7995942415156357e-07
GC_5_91 b_5 NI_5 NS_91 0 1.2595559251952706e-02
GC_5_92 b_5 NI_5 NS_92 0 -3.4658432696704052e-02
GC_5_93 b_5 NI_5 NS_93 0 -1.6777400680724746e-05
GC_5_94 b_5 NI_5 NS_94 0 -8.5075415211948500e-07
GC_5_95 b_5 NI_5 NS_95 0 1.4727416463639564e-08
GC_5_96 b_5 NI_5 NS_96 0 1.0163240415065454e-05
GC_5_97 b_5 NI_5 NS_97 0 -4.6901799867460722e-02
GC_5_98 b_5 NI_5 NS_98 0 6.7851984622432387e-02
GC_5_99 b_5 NI_5 NS_99 0 -2.4400432244440984e-02
GC_5_100 b_5 NI_5 NS_100 0 -1.6162327841823751e-01
GC_5_101 b_5 NI_5 NS_101 0 -1.2987354616556087e-02
GC_5_102 b_5 NI_5 NS_102 0 -1.8235267619288698e-01
GC_5_103 b_5 NI_5 NS_103 0 5.7459955593680928e-07
GC_5_104 b_5 NI_5 NS_104 0 1.0763902068039613e-06
GC_5_105 b_5 NI_5 NS_105 0 -5.4517338358574225e-06
GC_5_106 b_5 NI_5 NS_106 0 2.2107667429736568e-07
GC_5_107 b_5 NI_5 NS_107 0 -4.0754404547112319e-06
GC_5_108 b_5 NI_5 NS_108 0 -4.3104044417357537e-06
GC_5_109 b_5 NI_5 NS_109 0 -6.4982375546367849e-04
GC_5_110 b_5 NI_5 NS_110 0 1.5082834757475241e-03
GC_5_111 b_5 NI_5 NS_111 0 -7.8854179770011482e-07
GC_5_112 b_5 NI_5 NS_112 0 -1.1413279035352148e-09
GC_5_113 b_5 NI_5 NS_113 0 -3.0089389250485094e-11
GC_5_114 b_5 NI_5 NS_114 0 -2.2155990111467089e-07
GC_5_115 b_5 NI_5 NS_115 0 -4.3434184613996927e-03
GC_5_116 b_5 NI_5 NS_116 0 1.9143630618855278e-02
GC_5_117 b_5 NI_5 NS_117 0 1.8679830170594689e-02
GC_5_118 b_5 NI_5 NS_118 0 -1.1724732832404518e-02
GC_5_119 b_5 NI_5 NS_119 0 2.5507537658142065e-03
GC_5_120 b_5 NI_5 NS_120 0 2.9783263716003653e-02
GC_5_121 b_5 NI_5 NS_121 0 -3.8572889171500857e-08
GC_5_122 b_5 NI_5 NS_122 0 -2.6129286829487894e-08
GC_5_123 b_5 NI_5 NS_123 0 9.8376512132564201e-08
GC_5_124 b_5 NI_5 NS_124 0 -6.0736755715154928e-08
GC_5_125 b_5 NI_5 NS_125 0 5.4421053043725391e-08
GC_5_126 b_5 NI_5 NS_126 0 3.3115343069272144e-08
GC_5_127 b_5 NI_5 NS_127 0 1.2257943283729329e-04
GC_5_128 b_5 NI_5 NS_128 0 -4.7969203820363637e-04
GC_5_129 b_5 NI_5 NS_129 0 3.5201867675774881e-07
GC_5_130 b_5 NI_5 NS_130 0 3.6382660519985330e-09
GC_5_131 b_5 NI_5 NS_131 0 -1.2339166759156094e-11
GC_5_132 b_5 NI_5 NS_132 0 1.1983915470847397e-07
GC_5_133 b_5 NI_5 NS_133 0 7.2107242233124009e-04
GC_5_134 b_5 NI_5 NS_134 0 -4.2728279191699579e-03
GC_5_135 b_5 NI_5 NS_135 0 -8.9969966852694941e-03
GC_5_136 b_5 NI_5 NS_136 0 -5.1486263954082607e-03
GC_5_137 b_5 NI_5 NS_137 0 1.8447869489259274e-03
GC_5_138 b_5 NI_5 NS_138 0 7.1903569996370912e-03
GC_5_139 b_5 NI_5 NS_139 0 5.3585123178375480e-09
GC_5_140 b_5 NI_5 NS_140 0 1.7087696773180901e-09
GC_5_141 b_5 NI_5 NS_141 0 -2.9718376197375196e-09
GC_5_142 b_5 NI_5 NS_142 0 2.2411247258048161e-08
GC_5_143 b_5 NI_5 NS_143 0 -2.4721510618139354e-08
GC_5_144 b_5 NI_5 NS_144 0 -1.3986305852319134e-08
GC_5_145 b_5 NI_5 NS_145 0 -1.3595252233163390e-05
GC_5_146 b_5 NI_5 NS_146 0 4.5592973173014145e-05
GC_5_147 b_5 NI_5 NS_147 0 -1.5019930224481448e-08
GC_5_148 b_5 NI_5 NS_148 0 -6.4644638109903298e-10
GC_5_149 b_5 NI_5 NS_149 0 7.9994592576936558e-11
GC_5_150 b_5 NI_5 NS_150 0 -4.9840748238751341e-09
GC_5_151 b_5 NI_5 NS_151 0 1.1992735783804560e-04
GC_5_152 b_5 NI_5 NS_152 0 1.7682256064492443e-04
GC_5_153 b_5 NI_5 NS_153 0 3.0863511206745409e-04
GC_5_154 b_5 NI_5 NS_154 0 -5.1613131918464537e-04
GC_5_155 b_5 NI_5 NS_155 0 -3.8644931139917465e-04
GC_5_156 b_5 NI_5 NS_156 0 1.7101790868964331e-04
GC_5_157 b_5 NI_5 NS_157 0 -2.6793839162989381e-10
GC_5_158 b_5 NI_5 NS_158 0 -8.7398309617417848e-10
GC_5_159 b_5 NI_5 NS_159 0 -9.6236020449940535e-10
GC_5_160 b_5 NI_5 NS_160 0 3.6733300656719593e-09
GC_5_161 b_5 NI_5 NS_161 0 1.2868997046224837e-09
GC_5_162 b_5 NI_5 NS_162 0 -4.8000102618356415e-10
GC_5_163 b_5 NI_5 NS_163 0 6.2497572205673055e-06
GC_5_164 b_5 NI_5 NS_164 0 -2.3140525663473836e-06
GC_5_165 b_5 NI_5 NS_165 0 2.4895002276374942e-08
GC_5_166 b_5 NI_5 NS_166 0 6.7283313469133109e-10
GC_5_167 b_5 NI_5 NS_167 0 -7.9766204100826382e-11
GC_5_168 b_5 NI_5 NS_168 0 4.2097627111134542e-09
GC_5_169 b_5 NI_5 NS_169 0 -1.3706972091518901e-04
GC_5_170 b_5 NI_5 NS_170 0 1.8413136828360902e-04
GC_5_171 b_5 NI_5 NS_171 0 8.0544682422080231e-04
GC_5_172 b_5 NI_5 NS_172 0 2.0804712563819448e-04
GC_5_173 b_5 NI_5 NS_173 0 -5.4272486402922432e-04
GC_5_174 b_5 NI_5 NS_174 0 -8.9942561012261706e-04
GC_5_175 b_5 NI_5 NS_175 0 -1.4802286694147951e-10
GC_5_176 b_5 NI_5 NS_176 0 8.6940589169343154e-10
GC_5_177 b_5 NI_5 NS_177 0 1.8609693960234198e-09
GC_5_178 b_5 NI_5 NS_178 0 -4.9447520938130995e-09
GC_5_179 b_5 NI_5 NS_179 0 -9.7935139109024092e-10
GC_5_180 b_5 NI_5 NS_180 0 6.4646567992235579e-10
GC_5_181 b_5 NI_5 NS_181 0 1.3390392023196877e-06
GC_5_182 b_5 NI_5 NS_182 0 -7.7404820142711539e-06
GC_5_183 b_5 NI_5 NS_183 0 -3.8746466888869061e-09
GC_5_184 b_5 NI_5 NS_184 0 -2.4411479394840798e-10
GC_5_185 b_5 NI_5 NS_185 0 2.5141849853915763e-11
GC_5_186 b_5 NI_5 NS_186 0 -1.0189400453779196e-10
GC_5_187 b_5 NI_5 NS_187 0 -3.6245031099982489e-05
GC_5_188 b_5 NI_5 NS_188 0 5.2125785049946382e-05
GC_5_189 b_5 NI_5 NS_189 0 7.6021060835690356e-06
GC_5_190 b_5 NI_5 NS_190 0 1.4076152626869422e-04
GC_5_191 b_5 NI_5 NS_191 0 1.5323341884428346e-04
GC_5_192 b_5 NI_5 NS_192 0 4.9478016489837188e-05
GC_5_193 b_5 NI_5 NS_193 0 6.2298348755427034e-11
GC_5_194 b_5 NI_5 NS_194 0 -1.1932005119020389e-10
GC_5_195 b_5 NI_5 NS_195 0 -3.5791544735449363e-10
GC_5_196 b_5 NI_5 NS_196 0 1.0391252080344957e-09
GC_5_197 b_5 NI_5 NS_197 0 4.9855780172794278e-11
GC_5_198 b_5 NI_5 NS_198 0 -4.5817478979555737e-10
GC_5_199 b_5 NI_5 NS_199 0 4.4584380193701165e-06
GC_5_200 b_5 NI_5 NS_200 0 -1.7990473638426150e-05
GC_5_201 b_5 NI_5 NS_201 0 -4.6680579180436239e-10
GC_5_202 b_5 NI_5 NS_202 0 2.1056605371321810e-10
GC_5_203 b_5 NI_5 NS_203 0 -2.4757395235366436e-11
GC_5_204 b_5 NI_5 NS_204 0 6.0795985309017781e-10
GC_5_205 b_5 NI_5 NS_205 0 -1.3683880023405726e-05
GC_5_206 b_5 NI_5 NS_206 0 5.5046874711573011e-05
GC_5_207 b_5 NI_5 NS_207 0 1.4849988651770448e-04
GC_5_208 b_5 NI_5 NS_208 0 4.5509315558250131e-05
GC_5_209 b_5 NI_5 NS_209 0 -6.2796699199551406e-05
GC_5_210 b_5 NI_5 NS_210 0 -1.8722343356761671e-04
GC_5_211 b_5 NI_5 NS_211 0 1.7529360474254136e-10
GC_5_212 b_5 NI_5 NS_212 0 1.3267739172463325e-10
GC_5_213 b_5 NI_5 NS_213 0 -2.2723769274972605e-10
GC_5_214 b_5 NI_5 NS_214 0 -4.2066430109932887e-10
GC_5_215 b_5 NI_5 NS_215 0 -2.5484751318956535e-10
GC_5_216 b_5 NI_5 NS_216 0 2.9867700551396686e-10
GD_5_1 b_5 NI_5 NA_1 0 7.2422821104099283e-05
GD_5_2 b_5 NI_5 NA_2 0 -3.4083347627935442e-05
GD_5_3 b_5 NI_5 NA_3 0 -9.9243574060401828e-04
GD_5_4 b_5 NI_5 NA_4 0 2.6229987629973546e-03
GD_5_5 b_5 NI_5 NA_5 0 -9.3538553264762028e-02
GD_5_6 b_5 NI_5 NA_6 0 7.4111655686559613e-02
GD_5_7 b_5 NI_5 NA_7 0 6.1564925570875648e-03
GD_5_8 b_5 NI_5 NA_8 0 3.7689842542754214e-03
GD_5_9 b_5 NI_5 NA_9 0 6.4162387881828422e-05
GD_5_10 b_5 NI_5 NA_10 0 -3.5059837065024267e-05
GD_5_11 b_5 NI_5 NA_11 0 -4.9719336132104311e-05
GD_5_12 b_5 NI_5 NA_12 0 -2.8242996237297289e-05
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 6.5711863183111105e-06
GC_6_2 b_6 NI_6 NS_2 0 -3.4967225723075420e-06
GC_6_3 b_6 NI_6 NS_3 0 2.4263940541241598e-08
GC_6_4 b_6 NI_6 NS_4 0 6.7556484347522041e-10
GC_6_5 b_6 NI_6 NS_5 0 -8.0408554182211037e-11
GC_6_6 b_6 NI_6 NS_6 0 4.3269208271158259e-09
GC_6_7 b_6 NI_6 NS_7 0 -1.3639461183070486e-04
GC_6_8 b_6 NI_6 NS_8 0 1.8279341642053786e-04
GC_6_9 b_6 NI_6 NS_9 0 8.0661862139940399e-04
GC_6_10 b_6 NI_6 NS_10 0 2.0572344742348663e-04
GC_6_11 b_6 NI_6 NS_11 0 -5.4635687435219450e-04
GC_6_12 b_6 NI_6 NS_12 0 -9.0504032870398999e-04
GC_6_13 b_6 NI_6 NS_13 0 -1.3851006123388097e-10
GC_6_14 b_6 NI_6 NS_14 0 8.7169058698936703e-10
GC_6_15 b_6 NI_6 NS_15 0 1.8473013624120943e-09
GC_6_16 b_6 NI_6 NS_16 0 -4.9674628140791767e-09
GC_6_17 b_6 NI_6 NS_17 0 -1.0292492003308368e-09
GC_6_18 b_6 NI_6 NS_18 0 6.3129985635222012e-10
GC_6_19 b_6 NI_6 NS_19 0 -1.3683739762050597e-05
GC_6_20 b_6 NI_6 NS_20 0 4.5862454875800203e-05
GC_6_21 b_6 NI_6 NS_21 0 -1.4594664806403844e-08
GC_6_22 b_6 NI_6 NS_22 0 -6.5101996756272604e-10
GC_6_23 b_6 NI_6 NS_23 0 8.0662292415216454e-11
GC_6_24 b_6 NI_6 NS_24 0 -5.0747168616160525e-09
GC_6_25 b_6 NI_6 NS_25 0 1.1926470918773621e-04
GC_6_26 b_6 NI_6 NS_26 0 1.7734486091576193e-04
GC_6_27 b_6 NI_6 NS_27 0 3.0868337387572321e-04
GC_6_28 b_6 NI_6 NS_28 0 -5.1517026293257330e-04
GC_6_29 b_6 NI_6 NS_29 0 -3.8550123518491300e-04
GC_6_30 b_6 NI_6 NS_30 0 1.7218932740328138e-04
GC_6_31 b_6 NI_6 NS_31 0 -2.6650001444253132e-10
GC_6_32 b_6 NI_6 NS_32 0 -8.7560171014649443e-10
GC_6_33 b_6 NI_6 NS_33 0 -9.7850926728111525e-10
GC_6_34 b_6 NI_6 NS_34 0 3.7261673521121819e-09
GC_6_35 b_6 NI_6 NS_35 0 1.3261416259751091e-09
GC_6_36 b_6 NI_6 NS_36 0 -4.7355175516056252e-10
GC_6_37 b_6 NI_6 NS_37 0 1.3239366453694142e-04
GC_6_38 b_6 NI_6 NS_38 0 -4.8355778688855824e-04
GC_6_39 b_6 NI_6 NS_39 0 7.2278916321443188e-08
GC_6_40 b_6 NI_6 NS_40 0 5.7679787693009781e-10
GC_6_41 b_6 NI_6 NS_41 0 -1.2176774260190703e-10
GC_6_42 b_6 NI_6 NS_42 0 6.5843860392612528e-08
GC_6_43 b_6 NI_6 NS_43 0 -1.7783318470461558e-04
GC_6_44 b_6 NI_6 NS_44 0 -2.2251263856849423e-03
GC_6_45 b_6 NI_6 NS_45 0 -2.2111072264268286e-03
GC_6_46 b_6 NI_6 NS_46 0 -2.2403140889692111e-03
GC_6_47 b_6 NI_6 NS_47 0 -1.5810437528916044e-03
GC_6_48 b_6 NI_6 NS_48 0 -5.3321630326465133e-04
GC_6_49 b_6 NI_6 NS_49 0 1.3213976644184302e-09
GC_6_50 b_6 NI_6 NS_50 0 6.9371668040490811e-09
GC_6_51 b_6 NI_6 NS_51 0 9.3010343299289275e-09
GC_6_52 b_6 NI_6 NS_52 0 -2.8761363284020016e-08
GC_6_53 b_6 NI_6 NS_53 0 -1.9780396546415293e-08
GC_6_54 b_6 NI_6 NS_54 0 -1.2715079280015095e-08
GC_6_55 b_6 NI_6 NS_55 0 -2.2359206707011310e-04
GC_6_56 b_6 NI_6 NS_56 0 6.5327047164180987e-04
GC_6_57 b_6 NI_6 NS_57 0 -1.5277950439495732e-07
GC_6_58 b_6 NI_6 NS_58 0 -6.5097059020263156e-10
GC_6_59 b_6 NI_6 NS_59 0 1.1967615935413417e-10
GC_6_60 b_6 NI_6 NS_60 0 -8.1075761195037261e-08
GC_6_61 b_6 NI_6 NS_61 0 -4.6134499521598463e-04
GC_6_62 b_6 NI_6 NS_62 0 4.9878481144317146e-03
GC_6_63 b_6 NI_6 NS_63 0 4.0331150029301460e-03
GC_6_64 b_6 NI_6 NS_64 0 -5.0048770226916478e-04
GC_6_65 b_6 NI_6 NS_65 0 2.5277456289373879e-03
GC_6_66 b_6 NI_6 NS_66 0 6.9902302342982467e-03
GC_6_67 b_6 NI_6 NS_67 0 -7.4379232359631128e-09
GC_6_68 b_6 NI_6 NS_68 0 -1.1207497198047402e-08
GC_6_69 b_6 NI_6 NS_69 0 7.8408265262867889e-09
GC_6_70 b_6 NI_6 NS_70 0 2.1821468110209857e-08
GC_6_71 b_6 NI_6 NS_71 0 2.3395567343788661e-08
GC_6_72 b_6 NI_6 NS_72 0 1.3793436734460564e-08
GC_6_73 b_6 NI_6 NS_73 0 1.2595499050194713e-02
GC_6_74 b_6 NI_6 NS_74 0 -3.4658258700821086e-02
GC_6_75 b_6 NI_6 NS_75 0 -1.6777199855022758e-05
GC_6_76 b_6 NI_6 NS_76 0 -8.5074890194726829e-07
GC_6_77 b_6 NI_6 NS_77 0 1.4727344810596342e-08
GC_6_78 b_6 NI_6 NS_78 0 1.0163188623840127e-05
GC_6_79 b_6 NI_6 NS_79 0 -4.6901944370638424e-02
GC_6_80 b_6 NI_6 NS_80 0 6.7852014825095022e-02
GC_6_81 b_6 NI_6 NS_81 0 -2.4400579459786541e-02
GC_6_82 b_6 NI_6 NS_82 0 -1.6162304331313387e-01
GC_6_83 b_6 NI_6 NS_83 0 -1.2987090227012480e-02
GC_6_84 b_6 NI_6 NS_84 0 -1.8235212566042361e-01
GC_6_85 b_6 NI_6 NS_85 0 5.7459715165241941e-07
GC_6_86 b_6 NI_6 NS_86 0 1.0763836146787125e-06
GC_6_87 b_6 NI_6 NS_87 0 -5.4516984594420549e-06
GC_6_88 b_6 NI_6 NS_88 0 2.2107636389200749e-07
GC_6_89 b_6 NI_6 NS_89 0 -4.0754164572477468e-06
GC_6_90 b_6 NI_6 NS_90 0 -4.3103794274143807e-06
GC_6_91 b_6 NI_6 NS_91 0 -4.8322138401091126e-03
GC_6_92 b_6 NI_6 NS_92 0 1.6839927410558408e-02
GC_6_93 b_6 NI_6 NS_93 0 -3.4885576289249096e-06
GC_6_94 b_6 NI_6 NS_94 0 2.9143693123820634e-08
GC_6_95 b_6 NI_6 NS_95 0 -1.0018331264088617e-09
GC_6_96 b_6 NI_6 NS_96 0 -1.9968125735085949e-06
GC_6_97 b_6 NI_6 NS_97 0 1.8660666931443168e-02
GC_6_98 b_6 NI_6 NS_98 0 5.0341742983225572e-02
GC_6_99 b_6 NI_6 NS_99 0 1.4759545324524202e-02
GC_6_100 b_6 NI_6 NS_100 0 7.1489778072320653e-02
GC_6_101 b_6 NI_6 NS_101 0 8.1469900017227190e-02
GC_6_102 b_6 NI_6 NS_102 0 4.9245596332458480e-02
GC_6_103 b_6 NI_6 NS_103 0 -2.8743021846757047e-07
GC_6_104 b_6 NI_6 NS_104 0 -5.6953706963146018e-08
GC_6_105 b_6 NI_6 NS_105 0 5.7215241455712615e-07
GC_6_106 b_6 NI_6 NS_106 0 -8.2970936192739133e-07
GC_6_107 b_6 NI_6 NS_107 0 3.8940708076526688e-07
GC_6_108 b_6 NI_6 NS_108 0 3.7995942415219895e-07
GC_6_109 b_6 NI_6 NS_109 0 1.2258364170511770e-04
GC_6_110 b_6 NI_6 NS_110 0 -4.7970631312081648e-04
GC_6_111 b_6 NI_6 NS_111 0 3.5201421728851291e-07
GC_6_112 b_6 NI_6 NS_112 0 3.6382331994390892e-09
GC_6_113 b_6 NI_6 NS_113 0 -1.2338649439321654e-11
GC_6_114 b_6 NI_6 NS_114 0 1.1983976428987946e-07
GC_6_115 b_6 NI_6 NS_115 0 7.2108958877754230e-04
GC_6_116 b_6 NI_6 NS_116 0 -4.2728763224231091e-03
GC_6_117 b_6 NI_6 NS_117 0 -8.9970244765229836e-03
GC_6_118 b_6 NI_6 NS_118 0 -5.1487689306201848e-03
GC_6_119 b_6 NI_6 NS_119 0 1.8446620086622152e-03
GC_6_120 b_6 NI_6 NS_120 0 7.1902954169965339e-03
GC_6_121 b_6 NI_6 NS_121 0 5.3589244896294283e-09
GC_6_122 b_6 NI_6 NS_122 0 1.7087874202969563e-09
GC_6_123 b_6 NI_6 NS_123 0 -2.9727875840978656e-09
GC_6_124 b_6 NI_6 NS_124 0 2.2412183271406447e-08
GC_6_125 b_6 NI_6 NS_125 0 -2.4721744649586033e-08
GC_6_126 b_6 NI_6 NS_126 0 -1.3986471085132755e-08
GC_6_127 b_6 NI_6 NS_127 0 -6.4982386963171376e-04
GC_6_128 b_6 NI_6 NS_128 0 1.5082838515599255e-03
GC_6_129 b_6 NI_6 NS_129 0 -7.8854164035582394e-07
GC_6_130 b_6 NI_6 NS_130 0 -1.1413272092024585e-09
GC_6_131 b_6 NI_6 NS_131 0 -3.0089394923110411e-11
GC_6_132 b_6 NI_6 NS_132 0 -2.2155991723615201e-07
GC_6_133 b_6 NI_6 NS_133 0 -4.3434186031773517e-03
GC_6_134 b_6 NI_6 NS_134 0 1.9143631603052238e-02
GC_6_135 b_6 NI_6 NS_135 0 1.8679830490171564e-02
GC_6_136 b_6 NI_6 NS_136 0 -1.1724731618598499e-02
GC_6_137 b_6 NI_6 NS_137 0 2.5507552030082058e-03
GC_6_138 b_6 NI_6 NS_138 0 2.9783265166898203e-02
GC_6_139 b_6 NI_6 NS_139 0 -3.8572907509038503e-08
GC_6_140 b_6 NI_6 NS_140 0 -2.6129285726415730e-08
GC_6_141 b_6 NI_6 NS_141 0 9.8376547473574684e-08
GC_6_142 b_6 NI_6 NS_142 0 -6.0736778605672985e-08
GC_6_143 b_6 NI_6 NS_143 0 5.4421059227645422e-08
GC_6_144 b_6 NI_6 NS_144 0 3.3115346845041130e-08
GC_6_145 b_6 NI_6 NS_145 0 6.2470767217763875e-06
GC_6_146 b_6 NI_6 NS_146 0 -2.3041022057754158e-06
GC_6_147 b_6 NI_6 NS_147 0 2.4897773087797406e-08
GC_6_148 b_6 NI_6 NS_148 0 6.7284824642446328e-10
GC_6_149 b_6 NI_6 NS_149 0 -7.9766299194352200e-11
GC_6_150 b_6 NI_6 NS_150 0 4.2094381720451563e-09
GC_6_151 b_6 NI_6 NS_151 0 -1.3706989041887654e-04
GC_6_152 b_6 NI_6 NS_152 0 1.8416330744832317e-04
GC_6_153 b_6 NI_6 NS_153 0 8.0545714780458095e-04
GC_6_154 b_6 NI_6 NS_154 0 2.0808559774260639e-04
GC_6_155 b_6 NI_6 NS_155 0 -5.4267687867997987e-04
GC_6_156 b_6 NI_6 NS_156 0 -8.9938075257536831e-04
GC_6_157 b_6 NI_6 NS_157 0 -1.4819390521572134e-10
GC_6_158 b_6 NI_6 NS_158 0 8.6937252354254751e-10
GC_6_159 b_6 NI_6 NS_159 0 1.8613825513053051e-09
GC_6_160 b_6 NI_6 NS_160 0 -4.9451576607808273e-09
GC_6_161 b_6 NI_6 NS_161 0 -9.7922195171950982e-10
GC_6_162 b_6 NI_6 NS_162 0 6.4654980978562434e-10
GC_6_163 b_6 NI_6 NS_163 0 -1.2976717484184233e-05
GC_6_164 b_6 NI_6 NS_164 0 4.3440263387611889e-05
GC_6_165 b_6 NI_6 NS_165 0 -1.5814494331448843e-08
GC_6_166 b_6 NI_6 NS_166 0 -6.4986823104397051e-10
GC_6_167 b_6 NI_6 NS_167 0 8.0010305993054319e-11
GC_6_168 b_6 NI_6 NS_168 0 -4.9031448841512823e-09
GC_6_169 b_6 NI_6 NS_169 0 1.1938334132474811e-04
GC_6_170 b_6 NI_6 NS_170 0 1.6941639013043136e-04
GC_6_171 b_6 NI_6 NS_171 0 3.0484215035746497e-04
GC_6_172 b_6 NI_6 NS_172 0 -5.2370861718880691e-04
GC_6_173 b_6 NI_6 NS_173 0 -3.9528389605026672e-04
GC_6_174 b_6 NI_6 NS_174 0 1.6296889535201900e-04
GC_6_175 b_6 NI_6 NS_175 0 -2.3808620564048430e-10
GC_6_176 b_6 NI_6 NS_176 0 -8.7787697959354708e-10
GC_6_177 b_6 NI_6 NS_177 0 -1.0256008916198834e-09
GC_6_178 b_6 NI_6 NS_178 0 3.8229239096386165e-09
GC_6_179 b_6 NI_6 NS_179 0 1.2544645021937634e-09
GC_6_180 b_6 NI_6 NS_180 0 -5.0066235883652205e-10
GC_6_181 b_6 NI_6 NS_181 0 4.4889232968287804e-06
GC_6_182 b_6 NI_6 NS_182 0 -1.8090896909138476e-05
GC_6_183 b_6 NI_6 NS_183 0 -5.0679164278842060e-10
GC_6_184 b_6 NI_6 NS_184 0 2.1018088129214882e-10
GC_6_185 b_6 NI_6 NS_185 0 -2.4750708361229799e-11
GC_6_186 b_6 NI_6 NS_186 0 6.1365766451459518e-10
GC_6_187 b_6 NI_6 NS_187 0 -1.3564578292502605e-05
GC_6_188 b_6 NI_6 NS_188 0 5.4779566473945448e-05
GC_6_189 b_6 NI_6 NS_189 0 1.4837096219367659e-04
GC_6_190 b_6 NI_6 NS_190 0 4.4676736817363372e-05
GC_6_191 b_6 NI_6 NS_191 0 -6.3532199884827834e-05
GC_6_192 b_6 NI_6 NS_192 0 -1.8763781022641823e-04
GC_6_193 b_6 NI_6 NS_193 0 1.7826482449425330e-10
GC_6_194 b_6 NI_6 NS_194 0 1.3311006161359797e-10
GC_6_195 b_6 NI_6 NS_195 0 -2.3563931620349937e-10
GC_6_196 b_6 NI_6 NS_196 0 -4.1437931734307472e-10
GC_6_197 b_6 NI_6 NS_197 0 -2.5709561950322433e-10
GC_6_198 b_6 NI_6 NS_198 0 2.9692393269685765e-10
GC_6_199 b_6 NI_6 NS_199 0 1.3355195490724339e-06
GC_6_200 b_6 NI_6 NS_200 0 -7.7290133053435992e-06
GC_6_201 b_6 NI_6 NS_201 0 -3.8707216405659747e-09
GC_6_202 b_6 NI_6 NS_202 0 -2.4408415350038157e-10
GC_6_203 b_6 NI_6 NS_203 0 2.5141281247370119e-11
GC_6_204 b_6 NI_6 NS_204 0 -1.0237020675194573e-10
GC_6_205 b_6 NI_6 NS_205 0 -3.6243704103729150e-05
GC_6_206 b_6 NI_6 NS_206 0 5.2155784488651738e-05
GC_6_207 b_6 NI_6 NS_207 0 7.6127041403859016e-06
GC_6_208 b_6 NI_6 NS_208 0 1.4079630199394713e-04
GC_6_209 b_6 NI_6 NS_209 0 1.5327481378753571e-04
GC_6_210 b_6 NI_6 NS_210 0 4.9519570971493797e-05
GC_6_211 b_6 NI_6 NS_211 0 6.2161457519957826e-11
GC_6_212 b_6 NI_6 NS_212 0 -1.1934441748685021e-10
GC_6_213 b_6 NI_6 NS_213 0 -3.5746478864945607e-10
GC_6_214 b_6 NI_6 NS_214 0 1.0385955328534289e-09
GC_6_215 b_6 NI_6 NS_215 0 5.0039347016951374e-11
GC_6_216 b_6 NI_6 NS_216 0 -4.5803709786663560e-10
GD_6_1 b_6 NI_6 NA_1 0 -3.4092156140562412e-05
GD_6_2 b_6 NI_6 NA_2 0 6.4383450516593009e-05
GD_6_3 b_6 NI_6 NA_3 0 2.6224377094442356e-03
GD_6_4 b_6 NI_6 NA_4 0 -9.9162073083388595e-04
GD_6_5 b_6 NI_6 NA_5 0 7.4111664117099629e-02
GD_6_6 b_6 NI_6 NA_6 0 -9.3538553264762278e-02
GD_6_7 b_6 NI_6 NA_7 0 3.7690680881010069e-03
GD_6_8 b_6 NI_6 NA_8 0 6.1564915657368862e-03
GD_6_9 b_6 NI_6 NA_9 0 -3.5096775249106316e-05
GD_6_10 b_6 NI_6 NA_10 0 7.2404586111822453e-05
GD_6_11 b_6 NI_6 NA_11 0 -2.7783437866339298e-05
GD_6_12 b_6 NI_6 NA_12 0 -4.9753083772503213e-05
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 1.0304669723567804e-06
GC_7_2 b_7 NI_7 NS_2 0 -6.3836435845862568e-06
GC_7_3 b_7 NI_7 NS_3 0 -3.8670303712034364e-09
GC_7_4 b_7 NI_7 NS_4 0 -2.4269282911420926e-10
GC_7_5 b_7 NI_7 NS_5 0 2.5054713504031747e-11
GC_7_6 b_7 NI_7 NS_6 0 -1.2071296220481626e-10
GC_7_7 b_7 NI_7 NS_7 0 -3.6740305650376642e-05
GC_7_8 b_7 NI_7 NS_8 0 5.6720743584985061e-05
GC_7_9 b_7 NI_7 NS_9 0 8.7520244043003463e-06
GC_7_10 b_7 NI_7 NS_10 0 1.4649196866097281e-04
GC_7_11 b_7 NI_7 NS_11 0 1.6051646235341107e-04
GC_7_12 b_7 NI_7 NS_12 0 5.6595682277937065e-05
GC_7_13 b_7 NI_7 NS_13 0 6.0843776830807957e-11
GC_7_14 b_7 NI_7 NS_14 0 -1.4081195501541146e-10
GC_7_15 b_7 NI_7 NS_15 0 -3.3787590279062585e-10
GC_7_16 b_7 NI_7 NS_16 0 1.0572116408954025e-09
GC_7_17 b_7 NI_7 NS_17 0 5.5311031011767415e-11
GC_7_18 b_7 NI_7 NS_18 0 -4.5394078954224822e-10
GC_7_19 b_7 NI_7 NS_19 0 5.0795775445005959e-06
GC_7_20 b_7 NI_7 NS_20 0 -2.0495034310049820e-05
GC_7_21 b_7 NI_7 NS_21 0 -7.3514124452615235e-10
GC_7_22 b_7 NI_7 NS_22 0 2.0742717775423592e-10
GC_7_23 b_7 NI_7 NS_23 0 -2.4670911421114454e-11
GC_7_24 b_7 NI_7 NS_24 0 6.5223435357693811e-10
GC_7_25 b_7 NI_7 NS_25 0 -1.4010400342299359e-05
GC_7_26 b_7 NI_7 NS_26 0 4.6160804581011765e-05
GC_7_27 b_7 NI_7 NS_27 0 1.4554607298073702e-04
GC_7_28 b_7 NI_7 NS_28 0 3.5634074188149471e-05
GC_7_29 b_7 NI_7 NS_29 0 -7.5467958204444231e-05
GC_7_30 b_7 NI_7 NS_30 0 -1.9906750003725345e-04
GC_7_31 b_7 NI_7 NS_31 0 1.9164603618280587e-10
GC_7_32 b_7 NI_7 NS_32 0 1.5222254229657312e-10
GC_7_33 b_7 NI_7 NS_33 0 -2.7653337051258712e-10
GC_7_34 b_7 NI_7 NS_34 0 -4.0006442165505384e-10
GC_7_35 b_7 NI_7 NS_35 0 -2.7141933101619282e-10
GC_7_36 b_7 NI_7 NS_36 0 2.8552993623015319e-10
GC_7_37 b_7 NI_7 NS_37 0 -1.3609002132346642e-05
GC_7_38 b_7 NI_7 NS_38 0 4.5664436945023873e-05
GC_7_39 b_7 NI_7 NS_39 0 -1.5015648103420106e-08
GC_7_40 b_7 NI_7 NS_40 0 -6.4639584642450599e-10
GC_7_41 b_7 NI_7 NS_41 0 7.9993998293931503e-11
GC_7_42 b_7 NI_7 NS_42 0 -4.9849997937798983e-09
GC_7_43 b_7 NI_7 NS_43 0 1.1994564518704217e-04
GC_7_44 b_7 NI_7 NS_44 0 1.7720715181274318e-04
GC_7_45 b_7 NI_7 NS_45 0 3.0879688632519202e-04
GC_7_46 b_7 NI_7 NS_46 0 -5.1565674922472986e-04
GC_7_47 b_7 NI_7 NS_47 0 -3.8587540197634835e-04
GC_7_48 b_7 NI_7 NS_48 0 1.7143573088113104e-04
GC_7_49 b_7 NI_7 NS_49 0 -2.6845100659810200e-10
GC_7_50 b_7 NI_7 NS_50 0 -8.7537391230213535e-10
GC_7_51 b_7 NI_7 NS_51 0 -9.6027732947292218e-10
GC_7_52 b_7 NI_7 NS_52 0 3.6739415457743552e-09
GC_7_53 b_7 NI_7 NS_53 0 1.2872832637517833e-09
GC_7_54 b_7 NI_7 NS_54 0 -4.7972492126156001e-10
GC_7_55 b_7 NI_7 NS_55 0 6.2564823615304942e-06
GC_7_56 b_7 NI_7 NS_56 0 -2.3560903034340818e-06
GC_7_57 b_7 NI_7 NS_57 0 2.4895464732130372e-08
GC_7_58 b_7 NI_7 NS_58 0 6.7282184505874917e-10
GC_7_59 b_7 NI_7 NS_59 0 -7.9766537512302962e-11
GC_7_60 b_7 NI_7 NS_60 0 4.2103483437593610e-09
GC_7_61 b_7 NI_7 NS_61 0 -1.3708369807755347e-04
GC_7_62 b_7 NI_7 NS_62 0 1.8383967193212741e-04
GC_7_63 b_7 NI_7 NS_63 0 8.0532283779791148e-04
GC_7_64 b_7 NI_7 NS_64 0 2.0770441282950316e-04
GC_7_65 b_7 NI_7 NS_65 0 -5.4316040093594167e-04
GC_7_66 b_7 NI_7 NS_66 0 -8.9973588009620612e-04
GC_7_67 b_7 NI_7 NS_67 0 -1.4773005114757006e-10
GC_7_68 b_7 NI_7 NS_68 0 8.7080765053168708e-10
GC_7_69 b_7 NI_7 NS_69 0 1.8594330048411852e-09
GC_7_70 b_7 NI_7 NS_70 0 -4.9461662091131259e-09
GC_7_71 b_7 NI_7 NS_71 0 -9.7957896930800407e-10
GC_7_72 b_7 NI_7 NS_72 0 6.4633884882035619e-10
GC_7_73 b_7 NI_7 NS_73 0 -6.4982386964987089e-04
GC_7_74 b_7 NI_7 NS_74 0 1.5082838516261041e-03
GC_7_75 b_7 NI_7 NS_75 0 -7.8854164034857652e-07
GC_7_76 b_7 NI_7 NS_76 0 -1.1413272091866792e-09
GC_7_77 b_7 NI_7 NS_77 0 -3.0089394925295725e-11
GC_7_78 b_7 NI_7 NS_78 0 -2.2155991723723627e-07
GC_7_79 b_7 NI_7 NS_79 0 -4.3434186033222836e-03
GC_7_80 b_7 NI_7 NS_80 0 1.9143631603141486e-02
GC_7_81 b_7 NI_7 NS_81 0 1.8679830490135569e-02
GC_7_82 b_7 NI_7 NS_82 0 -1.1724731618351076e-02
GC_7_83 b_7 NI_7 NS_83 0 2.5507552032637882e-03
GC_7_84 b_7 NI_7 NS_84 0 2.9783265167198422e-02
GC_7_85 b_7 NI_7 NS_85 0 -3.8572907509973475e-08
GC_7_86 b_7 NI_7 NS_86 0 -2.6129285725782758e-08
GC_7_87 b_7 NI_7 NS_87 0 9.8376547474001523e-08
GC_7_88 b_7 NI_7 NS_88 0 -6.0736778607974718e-08
GC_7_89 b_7 NI_7 NS_89 0 5.4421059227971755e-08
GC_7_90 b_7 NI_7 NS_90 0 3.3115346845257196e-08
GC_7_91 b_7 NI_7 NS_91 0 1.2257943283893729e-04
GC_7_92 b_7 NI_7 NS_92 0 -4.7969203820931639e-04
GC_7_93 b_7 NI_7 NS_93 0 3.5201867675639456e-07
GC_7_94 b_7 NI_7 NS_94 0 3.6382660519892338e-09
GC_7_95 b_7 NI_7 NS_95 0 -1.2339166758971625e-11
GC_7_96 b_7 NI_7 NS_96 0 1.1983915470865296e-07
GC_7_97 b_7 NI_7 NS_97 0 7.2107242234162826e-04
GC_7_98 b_7 NI_7 NS_98 0 -4.2728279191757822e-03
GC_7_99 b_7 NI_7 NS_99 0 -8.9969966852657870e-03
GC_7_100 b_7 NI_7 NS_100 0 -5.1486263954260052e-03
GC_7_101 b_7 NI_7 NS_101 0 1.8447869489073196e-03
GC_7_102 b_7 NI_7 NS_102 0 7.1903569996130973e-03
GC_7_103 b_7 NI_7 NS_103 0 5.3585123179479021e-09
GC_7_104 b_7 NI_7 NS_104 0 1.7087696773120891e-09
GC_7_105 b_7 NI_7 NS_105 0 -2.9718376199364131e-09
GC_7_106 b_7 NI_7 NS_106 0 2.2411247258304971e-08
GC_7_107 b_7 NI_7 NS_107 0 -2.4721510618205382e-08
GC_7_108 b_7 NI_7 NS_108 0 -1.3986305852366707e-08
GC_7_109 b_7 NI_7 NS_109 0 -4.8318961815486195e-03
GC_7_110 b_7 NI_7 NS_110 0 1.6838946427139009e-02
GC_7_111 b_7 NI_7 NS_111 0 -3.4890861677710936e-06
GC_7_112 b_7 NI_7 NS_112 0 2.9139349562459469e-08
GC_7_113 b_7 NI_7 NS_113 0 -1.0017845007997251e-09
GC_7_114 b_7 NI_7 NS_114 0 -1.9967439769872069e-06
GC_7_115 b_7 NI_7 NS_115 0 1.8661668260788612e-02
GC_7_116 b_7 NI_7 NS_116 0 5.0341461834086866e-02
GC_7_117 b_7 NI_7 NS_117 0 1.4760431219580683e-02
GC_7_118 b_7 NI_7 NS_118 0 7.1488077085864896e-02
GC_7_119 b_7 NI_7 NS_119 0 8.1467989982105277e-02
GC_7_120 b_7 NI_7 NS_120 0 4.9242148218454601e-02
GC_7_121 b_7 NI_7 NS_121 0 -2.8739960579935276e-07
GC_7_122 b_7 NI_7 NS_122 0 -5.6935620630865208e-08
GC_7_123 b_7 NI_7 NS_123 0 5.7205423517462580e-07
GC_7_124 b_7 NI_7 NS_124 0 -8.2964255788138063e-07
GC_7_125 b_7 NI_7 NS_125 0 3.8937905046867964e-07
GC_7_126 b_7 NI_7 NS_126 0 3.7993823916868234e-07
GC_7_127 b_7 NI_7 NS_127 0 1.2588121934294004e-02
GC_7_128 b_7 NI_7 NS_128 0 -3.4636831555896024e-02
GC_7_129 b_7 NI_7 NS_129 0 -1.6752975396770956e-05
GC_7_130 b_7 NI_7 NS_130 0 -8.5012055093295780e-07
GC_7_131 b_7 NI_7 NS_131 0 1.4718624573628548e-08
GC_7_132 b_7 NI_7 NS_132 0 1.0156988988951368e-05
GC_7_133 b_7 NI_7 NS_133 0 -4.6919904890751915e-02
GC_7_134 b_7 NI_7 NS_134 0 6.7856964144494936e-02
GC_7_135 b_7 NI_7 NS_135 0 -2.4418070172235736e-02
GC_7_136 b_7 NI_7 NS_136 0 -1.6159270629212763e-01
GC_7_137 b_7 NI_7 NS_137 0 -1.2952933796106791e-02
GC_7_138 b_7 NI_7 NS_138 0 -1.8228358806847694e-01
GC_7_139 b_7 NI_7 NS_139 0 5.7422334597503098e-07
GC_7_140 b_7 NI_7 NS_140 0 1.0755743805772118e-06
GC_7_141 b_7 NI_7 NS_141 0 -5.4474327949853406e-06
GC_7_142 b_7 NI_7 NS_142 0 2.2096652345399316e-07
GC_7_143 b_7 NI_7 NS_143 0 -4.0725461826698891e-06
GC_7_144 b_7 NI_7 NS_144 0 -4.3073881444073549e-06
GC_7_145 b_7 NI_7 NS_145 0 -2.2349796860068888e-04
GC_7_146 b_7 NI_7 NS_146 0 6.5299175112532221e-04
GC_7_147 b_7 NI_7 NS_147 0 -1.5297642621090889e-07
GC_7_148 b_7 NI_7 NS_148 0 -6.5220675035394403e-10
GC_7_149 b_7 NI_7 NS_149 0 1.1968302354576163e-10
GC_7_150 b_7 NI_7 NS_150 0 -8.1050572097685793e-08
GC_7_151 b_7 NI_7 NS_151 0 -4.6083746362889614e-04
GC_7_152 b_7 NI_7 NS_152 0 4.9882322362061905e-03
GC_7_153 b_7 NI_7 NS_153 0 4.0337280091209387e-03
GC_7_154 b_7 NI_7 NS_154 0 -5.0074966247212391e-04
GC_7_155 b_7 NI_7 NS_155 0 2.5275259682582653e-03
GC_7_156 b_7 NI_7 NS_156 0 6.9892930447243836e-03
GC_7_157 b_7 NI_7 NS_157 0 -7.4263835873576243e-09
GC_7_158 b_7 NI_7 NS_158 0 -1.1198913263535639e-08
GC_7_159 b_7 NI_7 NS_159 0 7.8014494624110560e-09
GC_7_160 b_7 NI_7 NS_160 0 2.1845409484085880e-08
GC_7_161 b_7 NI_7 NS_161 0 2.3385362152775544e-08
GC_7_162 b_7 NI_7 NS_162 0 1.3786903135013470e-08
GC_7_163 b_7 NI_7 NS_163 0 1.3244052252714940e-04
GC_7_164 b_7 NI_7 NS_164 0 -4.8371347134402049e-04
GC_7_165 b_7 NI_7 NS_165 0 7.2239277594659403e-08
GC_7_166 b_7 NI_7 NS_166 0 5.7649183309694480e-10
GC_7_167 b_7 NI_7 NS_167 0 -1.2176306069741666e-10
GC_7_168 b_7 NI_7 NS_168 0 6.5848997588162048e-08
GC_7_169 b_7 NI_7 NS_169 0 -1.7772048029540162e-04
GC_7_170 b_7 NI_7 NS_170 0 -2.2254896755255055e-03
GC_7_171 b_7 NI_7 NS_171 0 -2.2112564118859802e-03
GC_7_172 b_7 NI_7 NS_172 0 -2.2412263104855685e-03
GC_7_173 b_7 NI_7 NS_173 0 -1.5818936060787219e-03
GC_7_174 b_7 NI_7 NS_174 0 -5.3381740147248613e-04
GC_7_175 b_7 NI_7 NS_175 0 1.3242086766555376e-09
GC_7_176 b_7 NI_7 NS_176 0 6.9364523309826920e-09
GC_7_177 b_7 NI_7 NS_177 0 9.2945612345419364e-09
GC_7_178 b_7 NI_7 NS_178 0 -2.8753658629631609e-08
GC_7_179 b_7 NI_7 NS_179 0 -1.9782498654623892e-08
GC_7_180 b_7 NI_7 NS_180 0 -1.2716731123341708e-08
GC_7_181 b_7 NI_7 NS_181 0 -1.2655122923688542e-05
GC_7_182 b_7 NI_7 NS_182 0 4.1969203866569938e-05
GC_7_183 b_7 NI_7 NS_183 0 -1.5475050800097794e-08
GC_7_184 b_7 NI_7 NS_184 0 -6.5458899710054915e-10
GC_7_185 b_7 NI_7 NS_185 0 8.0669248103711217e-11
GC_7_186 b_7 NI_7 NS_186 0 -4.9744620928872969e-09
GC_7_187 b_7 NI_7 NS_187 0 1.1881342708278441e-04
GC_7_188 b_7 NI_7 NS_188 0 1.6345370670485659e-04
GC_7_189 b_7 NI_7 NS_189 0 3.0273232025799433e-04
GC_7_190 b_7 NI_7 NS_190 0 -5.3028074686802863e-04
GC_7_191 b_7 NI_7 NS_191 0 -4.0384999255675636e-04
GC_7_192 b_7 NI_7 NS_192 0 1.5542131550216507e-04
GC_7_193 b_7 NI_7 NS_193 0 -2.2896668889076652e-10
GC_7_194 b_7 NI_7 NS_194 0 -8.6252774302169955e-10
GC_7_195 b_7 NI_7 NS_195 0 -1.0664715598507632e-09
GC_7_196 b_7 NI_7 NS_196 0 3.8727144738154349e-09
GC_7_197 b_7 NI_7 NS_197 0 1.2870632911978509e-09
GC_7_198 b_7 NI_7 NS_198 0 -4.9787423599968913e-10
GC_7_199 b_7 NI_7 NS_199 0 6.0001220955084397e-06
GC_7_200 b_7 NI_7 NS_200 0 -1.2007057868443140e-06
GC_7_201 b_7 NI_7 NS_201 0 2.4512811490666303e-08
GC_7_202 b_7 NI_7 NS_202 0 6.7664016595288680e-10
GC_7_203 b_7 NI_7 NS_203 0 -8.0405954235557607e-11
GC_7_204 b_7 NI_7 NS_204 0 4.2877295717343384e-09
GC_7_205 b_7 NI_7 NS_205 0 -1.3622076862102416e-04
GC_7_206 b_7 NI_7 NS_206 0 1.9072648581504271e-04
GC_7_207 b_7 NI_7 NS_207 0 8.0919478489449137e-04
GC_7_208 b_7 NI_7 NS_208 0 2.1471687001740913e-04
GC_7_209 b_7 NI_7 NS_209 0 -5.3483841130472036e-04
GC_7_210 b_7 NI_7 NS_210 0 -8.9414154534234592e-04
GC_7_211 b_7 NI_7 NS_211 0 -1.5409842707837396e-10
GC_7_212 b_7 NI_7 NS_212 0 8.5208755933434386e-10
GC_7_213 b_7 NI_7 NS_213 0 1.8956751217618269e-09
GC_7_214 b_7 NI_7 NS_214 0 -4.9875673807162502e-09
GC_7_215 b_7 NI_7 NS_215 0 -1.0147524819178614e-09
GC_7_216 b_7 NI_7 NS_216 0 6.4011215200338713e-10
GD_7_1 b_7 NI_7 NA_1 0 -5.4411392104923066e-05
GD_7_2 b_7 NI_7 NA_2 0 -1.8202757807602985e-05
GD_7_3 b_7 NI_7 NA_3 0 6.3682782755041981e-05
GD_7_4 b_7 NI_7 NA_4 0 -3.4701755552709832e-05
GD_7_5 b_7 NI_7 NA_5 0 6.1564915657370094e-03
GD_7_6 b_7 NI_7 NA_6 0 3.7689842542754214e-03
GD_7_7 b_7 NI_7 NA_7 0 -9.3538562102868372e-02
GD_7_8 b_7 NI_7 NA_8 0 7.4111657259732441e-02
GD_7_9 b_7 NI_7 NA_9 0 -9.9222315430915267e-04
GD_7_10 b_7 NI_7 NA_10 0 2.6229913124400481e-03
GD_7_11 b_7 NI_7 NA_11 0 7.9753278048827662e-05
GD_7_12 b_7 NI_7 NA_12 0 -4.3070867735153526e-05
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 5.1102384014875637e-06
GC_8_2 b_8 NI_8 NS_2 0 -2.0595979322823738e-05
GC_8_3 b_8 NI_8 NS_3 0 -7.7535052457111676e-10
GC_8_4 b_8 NI_8 NS_4 0 2.0703878608708888e-10
GC_8_5 b_8 NI_8 NS_5 0 -2.4664140735030835e-11
GC_8_6 b_8 NI_8 NS_6 0 6.5797411784114970e-10
GC_8_7 b_8 NI_8 NS_7 0 -1.3889629257204942e-05
GC_8_8 b_8 NI_8 NS_8 0 4.5898382266687387e-05
GC_8_9 b_8 NI_8 NS_9 0 1.4542188898122510e-04
GC_8_10 b_8 NI_8 NS_10 0 3.4803301862489925e-05
GC_8_11 b_8 NI_8 NS_11 0 -7.6201449394231949e-05
GC_8_12 b_8 NI_8 NS_12 0 -1.9948388116127483e-04
GC_8_13 b_8 NI_8 NS_13 0 1.9462586502391086e-10
GC_8_14 b_8 NI_8 NS_14 0 1.5267344477224127e-10
GC_8_15 b_8 NI_8 NS_15 0 -2.8498988442339304e-10
GC_8_16 b_8 NI_8 NS_16 0 -3.9376071041998142e-10
GC_8_17 b_8 NI_8 NS_17 0 -2.7368357767988939e-10
GC_8_18 b_8 NI_8 NS_18 0 2.8376315358941806e-10
GC_8_19 b_8 NI_8 NS_19 0 1.0261217058207619e-06
GC_8_20 b_8 NI_8 NS_20 0 -6.3678980462609475e-06
GC_8_21 b_8 NI_8 NS_21 0 -3.8617176025532611e-09
GC_8_22 b_8 NI_8 NS_22 0 -2.4265030883768455e-10
GC_8_23 b_8 NI_8 NS_23 0 2.5054234681972925e-11
GC_8_24 b_8 NI_8 NS_24 0 -1.2136408972714603e-10
GC_8_25 b_8 NI_8 NS_25 0 -3.6728333761013623e-05
GC_8_26 b_8 NI_8 NS_26 0 5.6788334742882460e-05
GC_8_27 b_8 NI_8 NS_27 0 8.7836833023609877e-06
GC_8_28 b_8 NI_8 NS_28 0 1.4656168315307439e-04
GC_8_29 b_8 NI_8 NS_29 0 1.6060324173963593e-04
GC_8_30 b_8 NI_8 NS_30 0 5.6663768762192843e-05
GC_8_31 b_8 NI_8 NS_31 0 6.0601689614529216e-11
GC_8_32 b_8 NI_8 NS_32 0 -1.4093745418029634e-10
GC_8_33 b_8 NI_8 NS_33 0 -3.3707578642025782e-10
GC_8_34 b_8 NI_8 NS_34 0 1.0565795747939350e-09
GC_8_35 b_8 NI_8 NS_35 0 5.5575278046807080e-11
GC_8_36 b_8 NI_8 NS_36 0 -4.5373767724120385e-10
GC_8_37 b_8 NI_8 NS_37 0 6.2533806872062627e-06
GC_8_38 b_8 NI_8 NS_38 0 -2.3445353301219446e-06
GC_8_39 b_8 NI_8 NS_39 0 2.4898512181859426e-08
GC_8_40 b_8 NI_8 NS_40 0 6.7283793532839601e-10
GC_8_41 b_8 NI_8 NS_41 0 -7.9766645288133938e-11
GC_8_42 b_8 NI_8 NS_42 0 4.2099989980728592e-09
GC_8_43 b_8 NI_8 NS_43 0 -1.3708326715750860e-04
GC_8_44 b_8 NI_8 NS_44 0 1.8387583849996072e-04
GC_8_45 b_8 NI_8 NS_45 0 8.0533408110910988e-04
GC_8_46 b_8 NI_8 NS_46 0 2.0774810816460073e-04
GC_8_47 b_8 NI_8 NS_47 0 -5.4310539915169086e-04
GC_8_48 b_8 NI_8 NS_48 0 -8.9968372355366032e-04
GC_8_49 b_8 NI_8 NS_49 0 -1.4790321422298707e-10
GC_8_50 b_8 NI_8 NS_50 0 8.7078180177712995e-10
GC_8_51 b_8 NI_8 NS_51 0 1.8598918414395046e-09
GC_8_52 b_8 NI_8 NS_52 0 -4.9466048175818895e-09
GC_8_53 b_8 NI_8 NS_53 0 -9.7944055810886917e-10
GC_8_54 b_8 NI_8 NS_54 0 6.4642667026647837e-10
GC_8_55 b_8 NI_8 NS_55 0 -1.2990464116709844e-05
GC_8_56 b_8 NI_8 NS_56 0 4.3509879534515070e-05
GC_8_57 b_8 NI_8 NS_57 0 -1.5810186317300822e-08
GC_8_58 b_8 NI_8 NS_58 0 -6.4981916984971210e-10
GC_8_59 b_8 NI_8 NS_59 0 8.0009744320667367e-11
GC_8_60 b_8 NI_8 NS_60 0 -4.9040884357677757e-09
GC_8_61 b_8 NI_8 NS_61 0 1.1939004383202923e-04
GC_8_62 b_8 NI_8 NS_62 0 1.6976511954899158e-04
GC_8_63 b_8 NI_8 NS_63 0 3.0498192237745308e-04
GC_8_64 b_8 NI_8 NS_64 0 -5.2326628782104184e-04
GC_8_65 b_8 NI_8 NS_65 0 -3.9475148225716843e-04
GC_8_66 b_8 NI_8 NS_66 0 1.6336796007807819e-04
GC_8_67 b_8 NI_8 NS_67 0 -2.3856253117889605e-10
GC_8_68 b_8 NI_8 NS_68 0 -8.7921364651012947e-10
GC_8_69 b_8 NI_8 NS_69 0 -1.0236141212608297e-09
GC_8_70 b_8 NI_8 NS_70 0 3.8234744581232532e-09
GC_8_71 b_8 NI_8 NS_71 0 1.2548481631370853e-09
GC_8_72 b_8 NI_8 NS_72 0 -5.0038263841671578e-10
GC_8_73 b_8 NI_8 NS_73 0 1.2258364182377680e-04
GC_8_74 b_8 NI_8 NS_74 0 -4.7970631352557181e-04
GC_8_75 b_8 NI_8 NS_75 0 3.5201421720605928e-07
GC_8_76 b_8 NI_8 NS_76 0 3.6382331990657226e-09
GC_8_77 b_8 NI_8 NS_77 0 -1.2338649435299493e-11
GC_8_78 b_8 NI_8 NS_78 0 1.1983976429736800e-07
GC_8_79 b_8 NI_8 NS_79 0 7.2108958910872334e-04
GC_8_80 b_8 NI_8 NS_80 0 -4.2728763228584623e-03
GC_8_81 b_8 NI_8 NS_81 0 -8.9970244763408150e-03
GC_8_82 b_8 NI_8 NS_82 0 -5.1487689315654174e-03
GC_8_83 b_8 NI_8 NS_83 0 1.8446620075343223e-03
GC_8_84 b_8 NI_8 NS_84 0 7.1902954153965160e-03
GC_8_85 b_8 NI_8 NS_85 0 5.3589244961750442e-09
GC_8_86 b_8 NI_8 NS_86 0 1.7087874159081597e-09
GC_8_87 b_8 NI_8 NS_87 0 -2.9727875906107122e-09
GC_8_88 b_8 NI_8 NS_88 0 2.2412183288370803e-08
GC_8_89 b_8 NI_8 NS_89 0 -2.4721744652408330e-08
GC_8_90 b_8 NI_8 NS_90 0 -1.3986471086995371e-08
GC_8_91 b_8 NI_8 NS_91 0 -6.4982375548483995e-04
GC_8_92 b_8 NI_8 NS_92 0 1.5082834758237283e-03
GC_8_93 b_8 NI_8 NS_93 0 -7.8854179768949895e-07
GC_8_94 b_8 NI_8 NS_94 0 -1.1413279034949805e-09
GC_8_95 b_8 NI_8 NS_95 0 -3.0089389253450013e-11
GC_8_96 b_8 NI_8 NS_96 0 -2.2155990111619444e-07
GC_8_97 b_8 NI_8 NS_97 0 -4.3434184615604937e-03
GC_8_98 b_8 NI_8 NS_98 0 1.9143630618952710e-02
GC_8_99 b_8 NI_8 NS_99 0 1.8679830170551529e-02
GC_8_100 b_8 NI_8 NS_100 0 -1.1724732832129960e-02
GC_8_101 b_8 NI_8 NS_101 0 2.5507537660986309e-03
GC_8_102 b_8 NI_8 NS_102 0 2.9783263716344030e-02
GC_8_103 b_8 NI_8 NS_103 0 -3.8572889172672026e-08
GC_8_104 b_8 NI_8 NS_104 0 -2.6129286828908054e-08
GC_8_105 b_8 NI_8 NS_105 0 9.8376512133565527e-08
GC_8_106 b_8 NI_8 NS_106 0 -6.0736755717978181e-08
GC_8_107 b_8 NI_8 NS_107 0 5.4421053044211442e-08
GC_8_108 b_8 NI_8 NS_108 0 3.3115343069603625e-08
GC_8_109 b_8 NI_8 NS_109 0 1.2588059510154282e-02
GC_8_110 b_8 NI_8 NS_110 0 -3.4636650599439898e-02
GC_8_111 b_8 NI_8 NS_111 0 -1.6752768928936892e-05
GC_8_112 b_8 NI_8 NS_112 0 -8.5011515117829390e-07
GC_8_113 b_8 NI_8 NS_113 0 1.4718550469126951e-08
GC_8_114 b_8 NI_8 NS_114 0 1.0156935749532845e-05
GC_8_115 b_8 NI_8 NS_115 0 -4.6920056639859264e-02
GC_8_116 b_8 NI_8 NS_116 0 6.7856996343655288e-02
GC_8_117 b_8 NI_8 NS_117 0 -2.4418224138739258e-02
GC_8_118 b_8 NI_8 NS_118 0 -1.6159245878739081e-01
GC_8_119 b_8 NI_8 NS_119 0 -1.2952655205655724e-02
GC_8_120 b_8 NI_8 NS_120 0 -1.8228301224487101e-01
GC_8_121 b_8 NI_8 NS_121 0 5.7422089943559151e-07
GC_8_122 b_8 NI_8 NS_122 0 1.0755676353638906e-06
GC_8_123 b_8 NI_8 NS_123 0 -5.4473964644025224e-06
GC_8_124 b_8 NI_8 NS_124 0 2.2096619761531395e-07
GC_8_125 b_8 NI_8 NS_125 0 -4.0725215149781463e-06
GC_8_126 b_8 NI_8 NS_126 0 -4.3073624244235026e-06
GC_8_127 b_8 NI_8 NS_127 0 -4.8318961817098421e-03
GC_8_128 b_8 NI_8 NS_128 0 1.6838946427584746e-02
GC_8_129 b_8 NI_8 NS_129 0 -3.4890861667113800e-06
GC_8_130 b_8 NI_8 NS_130 0 2.9139349567732286e-08
GC_8_131 b_8 NI_8 NS_131 0 -1.0017844991992228e-09
GC_8_132 b_8 NI_8 NS_132 0 -1.9967439775033981e-06
GC_8_133 b_8 NI_8 NS_133 0 1.8661668260571529e-02
GC_8_134 b_8 NI_8 NS_134 0 5.0341461834397312e-02
GC_8_135 b_8 NI_8 NS_135 0 1.4760431219427146e-02
GC_8_136 b_8 NI_8 NS_136 0 7.1488077086510018e-02
GC_8_137 b_8 NI_8 NS_137 0 8.1467989982857439e-02
GC_8_138 b_8 NI_8 NS_138 0 4.9242148219779555e-02
GC_8_139 b_8 NI_8 NS_139 0 -2.8739960579384430e-07
GC_8_140 b_8 NI_8 NS_140 0 -5.6935620651925081e-08
GC_8_141 b_8 NI_8 NS_141 0 5.7205423530211770e-07
GC_8_142 b_8 NI_8 NS_142 0 -8.2964255780129536e-07
GC_8_143 b_8 NI_8 NS_143 0 3.8937905079536712e-07
GC_8_144 b_8 NI_8 NS_144 0 3.7993823944566857e-07
GC_8_145 b_8 NI_8 NS_145 0 1.3240975272941488e-04
GC_8_146 b_8 NI_8 NS_146 0 -4.8360898983469431e-04
GC_8_147 b_8 NI_8 NS_147 0 7.2274921947849040e-08
GC_8_148 b_8 NI_8 NS_148 0 5.7680093577941563e-10
GC_8_149 b_8 NI_8 NS_149 0 -1.2176702397291079e-10
GC_8_150 b_8 NI_8 NS_150 0 6.5844045372596726e-08
GC_8_151 b_8 NI_8 NS_151 0 -1.7781545762933577e-04
GC_8_152 b_8 NI_8 NS_152 0 -2.2251465954955872e-03
GC_8_153 b_8 NI_8 NS_153 0 -2.2110764828737737e-03
GC_8_154 b_8 NI_8 NS_154 0 -2.2403402141989719e-03
GC_8_155 b_8 NI_8 NS_155 0 -1.5810875419885225e-03
GC_8_156 b_8 NI_8 NS_156 0 -5.3337321290869183e-04
GC_8_157 b_8 NI_8 NS_157 0 1.3213655315087821e-09
GC_8_158 b_8 NI_8 NS_158 0 6.9363403759806720e-09
GC_8_159 b_8 NI_8 NS_159 0 9.3019045288728721e-09
GC_8_160 b_8 NI_8 NS_160 0 -2.8759814093875733e-08
GC_8_161 b_8 NI_8 NS_161 0 -1.9780447985466340e-08
GC_8_162 b_8 NI_8 NS_162 0 -1.2715117628148823e-08
GC_8_163 b_8 NI_8 NS_163 0 -2.2345784069965644e-04
GC_8_164 b_8 NI_8 NS_164 0 6.5284991237062864e-04
GC_8_165 b_8 NI_8 NS_165 0 -1.5301568754898416e-07
GC_8_166 b_8 NI_8 NS_166 0 -6.5237658658537236e-10
GC_8_167 b_8 NI_8 NS_167 0 1.1968461273207549e-10
GC_8_168 b_8 NI_8 NS_168 0 -8.1046537779673300e-08
GC_8_169 b_8 NI_8 NS_169 0 -4.6094425156519687e-04
GC_8_170 b_8 NI_8 NS_170 0 4.9876147296234307e-03
GC_8_171 b_8 NI_8 NS_171 0 4.0334274680426914e-03
GC_8_172 b_8 NI_8 NS_172 0 -5.0135016492202603e-04
GC_8_173 b_8 NI_8 NS_173 0 2.5267637866084607e-03
GC_8_174 b_8 NI_8 NS_174 0 6.9886919109195837e-03
GC_8_175 b_8 NI_8 NS_175 0 -7.4244413319878213e-09
GC_8_176 b_8 NI_8 NS_176 0 -1.1198528770589284e-08
GC_8_177 b_8 NI_8 NS_177 0 7.7951526269503768e-09
GC_8_178 b_8 NI_8 NS_178 0 2.1849854495571797e-08
GC_8_179 b_8 NI_8 NS_179 0 2.3383806427195347e-08
GC_8_180 b_8 NI_8 NS_180 0 1.3785928646713596e-08
GC_8_181 b_8 NI_8 NS_181 0 5.9990560232303355e-06
GC_8_182 b_8 NI_8 NS_182 0 -1.1966961368629827e-06
GC_8_183 b_8 NI_8 NS_183 0 2.4514101153956619e-08
GC_8_184 b_8 NI_8 NS_184 0 6.7664907083182412e-10
GC_8_185 b_8 NI_8 NS_185 0 -8.0406027294839273e-11
GC_8_186 b_8 NI_8 NS_186 0 4.2875636336099662e-09
GC_8_187 b_8 NI_8 NS_187 0 -1.3622146005375928e-04
GC_8_188 b_8 NI_8 NS_188 0 1.9074668768451639e-04
GC_8_189 b_8 NI_8 NS_189 0 8.0921118818251959e-04
GC_8_190 b_8 NI_8 NS_190 0 2.1472039005154315e-04
GC_8_191 b_8 NI_8 NS_191 0 -5.3483054027185582e-04
GC_8_192 b_8 NI_8 NS_192 0 -8.9412916620545979e-04
GC_8_193 b_8 NI_8 NS_193 0 -1.5422750098838250e-10
GC_8_194 b_8 NI_8 NS_194 0 8.5210277780243667e-10
GC_8_195 b_8 NI_8 NS_195 0 1.8961597611353140e-09
GC_8_196 b_8 NI_8 NS_196 0 -4.9878805276413135e-09
GC_8_197 b_8 NI_8 NS_197 0 -1.0146841264980230e-09
GC_8_198 b_8 NI_8 NS_198 0 6.4015764622742048e-10
GC_8_199 b_8 NI_8 NS_199 0 -1.3260448238866919e-05
GC_8_200 b_8 NI_8 NS_200 0 4.4076051193794276e-05
GC_8_201 b_8 NI_8 NS_201 0 -1.4697575312490984e-08
GC_8_202 b_8 NI_8 NS_202 0 -6.5126883483453291e-10
GC_8_203 b_8 NI_8 NS_203 0 8.0654533072579438e-11
GC_8_204 b_8 NI_8 NS_204 0 -5.0535485724699421e-09
GC_8_205 b_8 NI_8 NS_205 0 1.1931482918384660e-04
GC_8_206 b_8 NI_8 NS_206 0 1.7067297008101047e-04
GC_8_207 b_8 NI_8 NS_207 0 3.0643937210808207e-04
GC_8_208 b_8 NI_8 NS_208 0 -5.2287913083392883e-04
GC_8_209 b_8 NI_8 NS_209 0 -3.9525301115083251e-04
GC_8_210 b_8 NI_8 NS_210 0 1.6327254253671014e-04
GC_8_211 b_8 NI_8 NS_211 0 -2.5837384380522903e-10
GC_8_212 b_8 NI_8 NS_212 0 -8.5878770704504287e-10
GC_8_213 b_8 NI_8 NS_213 0 -1.0039908515318876e-09
GC_8_214 b_8 NI_8 NS_214 0 3.7270542641301796e-09
GC_8_215 b_8 NI_8 NS_215 0 1.3187434989357310e-09
GC_8_216 b_8 NI_8 NS_216 0 -4.7771924365383472e-10
GD_8_1 b_8 NI_8 NA_1 0 -1.7748021847723683e-05
GD_8_2 b_8 NI_8 NA_2 0 -5.4496393686606360e-05
GD_8_3 b_8 NI_8 NA_3 0 -3.4744599132574246e-05
GD_8_4 b_8 NI_8 NA_4 0 7.1974324116059958e-05
GD_8_5 b_8 NI_8 NA_5 0 3.7690680884683216e-03
GD_8_6 b_8 NI_8 NA_6 0 6.1564925570876360e-03
GD_8_7 b_8 NI_8 NA_7 0 7.4111665870847013e-02
GD_8_8 b_8 NI_8 NA_8 0 -9.3538562103155254e-02
GD_8_9 b_8 NI_8 NA_9 0 2.6224374701093365e-03
GD_8_10 b_8 NI_8 NA_10 0 -9.9145202409055885e-04
GD_8_11 b_8 NI_8 NA_11 0 -4.3086487757816545e-05
GD_8_12 b_8 NI_8 NA_12 0 7.1764274680547865e-05
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 4.0450222816650316e-07
GC_9_2 b_9 NI_9 NS_2 0 -1.0625283213847504e-06
GC_9_3 b_9 NI_9 NS_3 0 -6.0184114438362729e-10
GC_9_4 b_9 NI_9 NS_4 0 -1.0361783921813655e-10
GC_9_5 b_9 NI_9 NS_5 0 8.1965865451581406e-12
GC_9_6 b_9 NI_9 NS_6 0 1.6697155184122287e-10
GC_9_7 b_9 NI_9 NS_7 0 -7.3127908439541610e-06
GC_9_8 b_9 NI_9 NS_8 0 -4.1309637563140588e-06
GC_9_9 b_9 NI_9 NS_9 0 -6.1746466264172007e-06
GC_9_10 b_9 NI_9 NS_10 0 4.4531783252914226e-06
GC_9_11 b_9 NI_9 NS_11 0 3.8995694477568330e-06
GC_9_12 b_9 NI_9 NS_12 0 2.6656280771852394e-06
GC_9_13 b_9 NI_9 NS_13 0 -1.1522618956295960e-11
GC_9_14 b_9 NI_9 NS_14 0 6.7968290519836428e-11
GC_9_15 b_9 NI_9 NS_15 0 1.7905061788373503e-10
GC_9_16 b_9 NI_9 NS_16 0 -4.3368764073670278e-10
GC_9_17 b_9 NI_9 NS_17 0 -2.8731432587041802e-11
GC_9_18 b_9 NI_9 NS_18 0 -2.4192403274099747e-10
GC_9_19 b_9 NI_9 NS_19 0 6.7099359728755802e-07
GC_9_20 b_9 NI_9 NS_20 0 -2.2973385309635845e-06
GC_9_21 b_9 NI_9 NS_21 0 -1.5909191569001149e-09
GC_9_22 b_9 NI_9 NS_22 0 5.3889760767391201e-11
GC_9_23 b_9 NI_9 NS_23 0 -7.3753147355335509e-12
GC_9_24 b_9 NI_9 NS_24 0 3.2536435900361322e-10
GC_9_25 b_9 NI_9 NS_25 0 4.0766812533278322e-06
GC_9_26 b_9 NI_9 NS_26 0 -4.1634909595177285e-06
GC_9_27 b_9 NI_9 NS_27 0 3.0280141314566035e-06
GC_9_28 b_9 NI_9 NS_28 0 -8.4376581963797428e-06
GC_9_29 b_9 NI_9 NS_29 0 -1.0871231046262227e-05
GC_9_30 b_9 NI_9 NS_30 0 -1.2340839795534475e-05
GC_9_31 b_9 NI_9 NS_31 0 6.1560074721461937e-11
GC_9_32 b_9 NI_9 NS_32 0 -1.1198981009601771e-11
GC_9_33 b_9 NI_9 NS_33 0 -5.2524154207764130e-10
GC_9_34 b_9 NI_9 NS_34 0 5.2973811855094301e-10
GC_9_35 b_9 NI_9 NS_35 0 -1.9706341588333832e-10
GC_9_36 b_9 NI_9 NS_36 0 7.7380244967553153e-12
GC_9_37 b_9 NI_9 NS_37 0 -8.0171136644906916e-07
GC_9_38 b_9 NI_9 NS_38 0 2.7308205448031111e-06
GC_9_39 b_9 NI_9 NS_39 0 -5.2075741046712989e-10
GC_9_40 b_9 NI_9 NS_40 0 -1.3300181966615424e-10
GC_9_41 b_9 NI_9 NS_41 0 1.4437314285697801e-11
GC_9_42 b_9 NI_9 NS_42 0 -3.0344221388330181e-10
GC_9_43 b_9 NI_9 NS_43 0 -1.8011838660672448e-06
GC_9_44 b_9 NI_9 NS_44 0 2.7926444815475150e-05
GC_9_45 b_9 NI_9 NS_45 0 1.0913058596048263e-05
GC_9_46 b_9 NI_9 NS_46 0 4.2540761921465972e-05
GC_9_47 b_9 NI_9 NS_47 0 4.9978562109862097e-05
GC_9_48 b_9 NI_9 NS_48 0 2.6934982417017752e-05
GC_9_49 b_9 NI_9 NS_49 0 7.0562610173281007e-11
GC_9_50 b_9 NI_9 NS_50 0 -1.8189059660204732e-10
GC_9_51 b_9 NI_9 NS_51 0 -4.0119182505195309e-10
GC_9_52 b_9 NI_9 NS_52 0 1.2111185564281583e-09
GC_9_53 b_9 NI_9 NS_53 0 1.8458306463317430e-10
GC_9_54 b_9 NI_9 NS_54 0 -1.7359222914525706e-10
GC_9_55 b_9 NI_9 NS_55 0 1.5476363541485045e-06
GC_9_56 b_9 NI_9 NS_56 0 -6.2962873467671567e-06
GC_9_57 b_9 NI_9 NS_57 0 1.2235156875331801e-10
GC_9_58 b_9 NI_9 NS_58 0 1.2886957143023071e-10
GC_9_59 b_9 NI_9 NS_59 0 -1.4440179215657743e-11
GC_9_60 b_9 NI_9 NS_60 0 3.5705193059008127e-10
GC_9_61 b_9 NI_9 NS_61 0 -6.9993933512366911e-06
GC_9_62 b_9 NI_9 NS_62 0 -7.1762885699132918e-06
GC_9_63 b_9 NI_9 NS_63 0 1.6282911379093959e-05
GC_9_64 b_9 NI_9 NS_64 0 -7.7564684847809642e-06
GC_9_65 b_9 NI_9 NS_65 0 -3.1226599171010898e-05
GC_9_66 b_9 NI_9 NS_66 0 -4.7428224579726757e-05
GC_9_67 b_9 NI_9 NS_67 0 -5.4189396076469916e-11
GC_9_68 b_9 NI_9 NS_68 0 1.7583911514789193e-10
GC_9_69 b_9 NI_9 NS_69 0 3.7769900051140900e-10
GC_9_70 b_9 NI_9 NS_70 0 -1.1564032489949419e-09
GC_9_71 b_9 NI_9 NS_71 0 -2.0765971215135720e-10
GC_9_72 b_9 NI_9 NS_72 0 1.5302908263659095e-10
GC_9_73 b_9 NI_9 NS_73 0 -1.2976717413669860e-05
GC_9_74 b_9 NI_9 NS_74 0 4.3440263131878832e-05
GC_9_75 b_9 NI_9 NS_75 0 -1.5814493950233139e-08
GC_9_76 b_9 NI_9 NS_76 0 -6.4986821482478077e-10
GC_9_77 b_9 NI_9 NS_77 0 8.0010305202962869e-11
GC_9_78 b_9 NI_9 NS_78 0 -4.9031450821602206e-09
GC_9_79 b_9 NI_9 NS_79 0 1.1938334136466629e-04
GC_9_80 b_9 NI_9 NS_80 0 1.6941638894917371e-04
GC_9_81 b_9 NI_9 NS_81 0 3.0484214976316524e-04
GC_9_82 b_9 NI_9 NS_82 0 -5.2370861836290776e-04
GC_9_83 b_9 NI_9 NS_83 0 -3.9528389742859115e-04
GC_9_84 b_9 NI_9 NS_84 0 1.6296889427873428e-04
GC_9_85 b_9 NI_9 NS_85 0 -2.3808620140304249e-10
GC_9_86 b_9 NI_9 NS_86 0 -8.7787696634648119e-10
GC_9_87 b_9 NI_9 NS_87 0 -1.0256009878306311e-09
GC_9_88 b_9 NI_9 NS_88 0 3.8229240563581506e-09
GC_9_89 b_9 NI_9 NS_89 0 1.2544645883334962e-09
GC_9_90 b_9 NI_9 NS_90 0 -5.0066228327596820e-10
GC_9_91 b_9 NI_9 NS_91 0 6.2497574398786012e-06
GC_9_92 b_9 NI_9 NS_92 0 -2.3140531313936712e-06
GC_9_93 b_9 NI_9 NS_93 0 2.4895000386000692e-08
GC_9_94 b_9 NI_9 NS_94 0 6.7283312479455150e-10
GC_9_95 b_9 NI_9 NS_95 0 -7.9766204065025035e-11
GC_9_96 b_9 NI_9 NS_96 0 4.2097631909641345e-09
GC_9_97 b_9 NI_9 NS_97 0 -1.3706972061158700e-04
GC_9_98 b_9 NI_9 NS_98 0 1.8413136807211828e-04
GC_9_99 b_9 NI_9 NS_99 0 8.0544682446989950e-04
GC_9_100 b_9 NI_9 NS_100 0 2.0804712501786314e-04
GC_9_101 b_9 NI_9 NS_101 0 -5.4272486470021363e-04
GC_9_102 b_9 NI_9 NS_102 0 -8.9942561159659122e-04
GC_9_103 b_9 NI_9 NS_103 0 -1.4802288540813254e-10
GC_9_104 b_9 NI_9 NS_104 0 8.6940592810136062e-10
GC_9_105 b_9 NI_9 NS_105 0 1.8609691736284735e-09
GC_9_106 b_9 NI_9 NS_106 0 -4.9447522741583750e-09
GC_9_107 b_9 NI_9 NS_107 0 -9.7935156409200320e-10
GC_9_108 b_9 NI_9 NS_108 0 6.4646564472003729e-10
GC_9_109 b_9 NI_9 NS_109 0 -2.2345784071681689e-04
GC_9_110 b_9 NI_9 NS_110 0 6.5284991242842236e-04
GC_9_111 b_9 NI_9 NS_111 0 -1.5301568753114477e-07
GC_9_112 b_9 NI_9 NS_112 0 -6.5237658649407830e-10
GC_9_113 b_9 NI_9 NS_113 0 1.1968461273061898e-10
GC_9_114 b_9 NI_9 NS_114 0 -8.1046537781962658e-08
GC_9_115 b_9 NI_9 NS_115 0 -4.6094425166096726e-04
GC_9_116 b_9 NI_9 NS_116 0 4.9876147296737680e-03
GC_9_117 b_9 NI_9 NS_117 0 4.0334274680020876e-03
GC_9_118 b_9 NI_9 NS_118 0 -5.0135016475853723e-04
GC_9_119 b_9 NI_9 NS_119 0 2.5267637867814473e-03
GC_9_120 b_9 NI_9 NS_120 0 6.9886919111548382e-03
GC_9_121 b_9 NI_9 NS_121 0 -7.4244413332448777e-09
GC_9_122 b_9 NI_9 NS_122 0 -1.1198528770786972e-08
GC_9_123 b_9 NI_9 NS_123 0 7.7951526298596455e-09
GC_9_124 b_9 NI_9 NS_124 0 2.1849854492710890e-08
GC_9_125 b_9 NI_9 NS_125 0 2.3383806428058533e-08
GC_9_126 b_9 NI_9 NS_126 0 1.3785928647266785e-08
GC_9_127 b_9 NI_9 NS_127 0 1.3244052261413196e-04
GC_9_128 b_9 NI_9 NS_128 0 -4.8371347151332018e-04
GC_9_129 b_9 NI_9 NS_129 0 7.2239277089269492e-08
GC_9_130 b_9 NI_9 NS_130 0 5.7649182807579015e-10
GC_9_131 b_9 NI_9 NS_131 0 -1.2176306064988837e-10
GC_9_132 b_9 NI_9 NS_132 0 6.5848997663385483e-08
GC_9_133 b_9 NI_9 NS_133 0 -1.7772048030753783e-04
GC_9_134 b_9 NI_9 NS_134 0 -2.2254896750759680e-03
GC_9_135 b_9 NI_9 NS_135 0 -2.2112564115581552e-03
GC_9_136 b_9 NI_9 NS_136 0 -2.2412263099691994e-03
GC_9_137 b_9 NI_9 NS_137 0 -1.5818936054918077e-03
GC_9_138 b_9 NI_9 NS_138 0 -5.3381740152471041e-04
GC_9_139 b_9 NI_9 NS_139 0 1.3242087257939103e-09
GC_9_140 b_9 NI_9 NS_140 0 6.9364524336066744e-09
GC_9_141 b_9 NI_9 NS_141 0 9.2945611068350155e-09
GC_9_142 b_9 NI_9 NS_142 0 -2.8753658579382617e-08
GC_9_143 b_9 NI_9 NS_143 0 -1.9782498686357935e-08
GC_9_144 b_9 NI_9 NS_144 0 -1.2716731148341543e-08
GC_9_145 b_9 NI_9 NS_145 0 -4.8625241773555183e-03
GC_9_146 b_9 NI_9 NS_146 0 1.6965213023597762e-02
GC_9_147 b_9 NI_9 NS_147 0 -3.4509061476416429e-06
GC_9_148 b_9 NI_9 NS_148 0 2.9323276789303648e-08
GC_9_149 b_9 NI_9 NS_149 0 -1.0119702753966379e-09
GC_9_150 b_9 NI_9 NS_150 0 -2.0010662620446924e-06
GC_9_151 b_9 NI_9 NS_151 0 1.8510763516702812e-02
GC_9_152 b_9 NI_9 NS_152 0 5.0676143484195357e-02
GC_9_153 b_9 NI_9 NS_153 0 1.4775875168041243e-02
GC_9_154 b_9 NI_9 NS_154 0 7.2025344573469846e-02
GC_9_155 b_9 NI_9 NS_155 0 8.2113614999496543e-02
GC_9_156 b_9 NI_9 NS_156 0 4.9907424272131976e-02
GC_9_157 b_9 NI_9 NS_157 0 -2.8706263305285930e-07
GC_9_158 b_9 NI_9 NS_158 0 -5.8605014838934107e-08
GC_9_159 b_9 NI_9 NS_159 0 5.7101018782468591e-07
GC_9_160 b_9 NI_9 NS_160 0 -8.2174834855185165e-07
GC_9_161 b_9 NI_9 NS_161 0 3.9089970822352970e-07
GC_9_162 b_9 NI_9 NS_162 0 3.8092737133258839e-07
GC_9_163 b_9 NI_9 NS_163 0 1.2607314818001382e-02
GC_9_164 b_9 NI_9 NS_164 0 -3.4706454441329998e-02
GC_9_165 b_9 NI_9 NS_165 0 -1.6753241886193218e-05
GC_9_166 b_9 NI_9 NS_166 0 -8.5056157992004944e-07
GC_9_167 b_9 NI_9 NS_167 0 1.4723737444241041e-08
GC_9_168 b_9 NI_9 NS_168 0 1.0162763294391489e-05
GC_9_169 b_9 NI_9 NS_169 0 -4.6994892158025575e-02
GC_9_170 b_9 NI_9 NS_170 0 6.7612961395024901e-02
GC_9_171 b_9 NI_9 NS_171 0 -2.4544737051546039e-02
GC_9_172 b_9 NI_9 NS_172 0 -1.6180124362427742e-01
GC_9_173 b_9 NI_9 NS_173 0 -1.3230697905623784e-02
GC_9_174 b_9 NI_9 NS_174 0 -1.8254023613301856e-01
GC_9_175 b_9 NI_9 NS_175 0 5.7566610610119728e-07
GC_9_176 b_9 NI_9 NS_176 0 1.0761968648990670e-06
GC_9_177 b_9 NI_9 NS_177 0 -5.4559011239637368e-06
GC_9_178 b_9 NI_9 NS_178 0 2.2858210761414981e-07
GC_9_179 b_9 NI_9 NS_179 0 -4.0753814072705796e-06
GC_9_180 b_9 NI_9 NS_180 0 -4.3093555882093290e-06
GC_9_181 b_9 NI_9 NS_181 0 -6.0714589214117562e-04
GC_9_182 b_9 NI_9 NS_182 0 1.3759759195824332e-03
GC_9_183 b_9 NI_9 NS_183 0 -8.5772785964701798e-07
GC_9_184 b_9 NI_9 NS_184 0 -1.4280316037494565e-09
GC_9_185 b_9 NI_9 NS_185 0 -2.7382752150965550e-11
GC_9_186 b_9 NI_9 NS_186 0 -2.1435121145938796e-07
GC_9_187 b_9 NI_9 NS_187 0 -4.2079275805202822e-03
GC_9_188 b_9 NI_9 NS_188 0 1.9043905518510422e-02
GC_9_189 b_9 NI_9 NS_189 0 1.8778530753202446e-02
GC_9_190 b_9 NI_9 NS_190 0 -1.2050033188293483e-02
GC_9_191 b_9 NI_9 NS_191 0 2.1826900266483035e-03
GC_9_192 b_9 NI_9 NS_192 0 2.9283123940223872e-02
GC_9_193 b_9 NI_9 NS_193 0 -3.3741425227195429e-08
GC_9_194 b_9 NI_9 NS_194 0 -2.4547826508540344e-08
GC_9_195 b_9 NI_9 NS_195 0 8.1296563939681722e-08
GC_9_196 b_9 NI_9 NS_196 0 -4.2574365461571661e-08
GC_9_197 b_9 NI_9 NS_197 0 5.1566298768906680e-08
GC_9_198 b_9 NI_9 NS_198 0 3.1363508263274414e-08
GC_9_199 b_9 NI_9 NS_199 0 1.1714737884190868e-04
GC_9_200 b_9 NI_9 NS_200 0 -4.6262296226664743e-04
GC_9_201 b_9 NI_9 NS_201 0 3.5654164953125905e-07
GC_9_202 b_9 NI_9 NS_202 0 3.4767317361646966e-09
GC_9_203 b_9 NI_9 NS_203 0 -1.1870736198813413e-11
GC_9_204 b_9 NI_9 NS_204 0 1.2107815938870015e-07
GC_9_205 b_9 NI_9 NS_205 0 7.0304718425388542e-04
GC_9_206 b_9 NI_9 NS_206 0 -4.2878840273526710e-03
GC_9_207 b_9 NI_9 NS_207 0 -9.0097181752555981e-03
GC_9_208 b_9 NI_9 NS_208 0 -5.1465729696761348e-03
GC_9_209 b_9 NI_9 NS_209 0 1.8363876405118908e-03
GC_9_210 b_9 NI_9 NS_210 0 7.2289510689221110e-03
GC_9_211 b_9 NI_9 NS_211 0 4.0587609512632488e-09
GC_9_212 b_9 NI_9 NS_212 0 2.5522864747852521e-09
GC_9_213 b_9 NI_9 NS_213 0 1.9345083950863041e-09
GC_9_214 b_9 NI_9 NS_214 0 1.2042396455645902e-08
GC_9_215 b_9 NI_9 NS_215 0 -2.5390538324494537e-08
GC_9_216 b_9 NI_9 NS_216 0 -1.4677008640099652e-08
GD_9_1 b_9 NI_9 NA_1 0 9.7357560231156025e-06
GD_9_2 b_9 NI_9 NA_2 0 -5.8537923115818755e-08
GD_9_3 b_9 NI_9 NA_3 0 -3.3984119262448433e-05
GD_9_4 b_9 NI_9 NA_4 0 1.8947982098009816e-05
GD_9_5 b_9 NI_9 NA_5 0 7.2404587247932187e-05
GD_9_6 b_9 NI_9 NA_6 0 -3.5059836923724487e-05
GD_9_7 b_9 NI_9 NA_7 0 -9.9145202409050659e-04
GD_9_8 b_9 NI_9 NA_8 0 2.6229913119757927e-03
GD_9_9 b_9 NI_9 NA_9 0 -9.3789405414097998e-02
GD_9_10 b_9 NI_9 NA_10 0 7.4456382656751391e-02
GD_9_11 b_9 NI_9 NA_11 0 6.2327480091610588e-03
GD_9_12 b_9 NI_9 NA_12 0 3.7902998126692548e-03
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 6.7104909040362295e-07
GC_10_2 b_10 NI_10 NS_2 0 -2.2975393229946515e-06
GC_10_3 b_10 NI_10 NS_3 0 -1.5909904472400875e-09
GC_10_4 b_10 NI_10 NS_4 0 5.3888269402360034e-11
GC_10_5 b_10 NI_10 NS_5 0 -7.3752982459193432e-12
GC_10_6 b_10 NI_10 NS_6 0 3.2537978118522007e-10
GC_10_7 b_10 NI_10 NS_7 0 4.0765517103188220e-06
GC_10_8 b_10 NI_10 NS_8 0 -4.1640455711516262e-06
GC_10_9 b_10 NI_10 NS_9 0 3.0278770838711694e-06
GC_10_10 b_10 NI_10 NS_10 0 -8.4383605848731526e-06
GC_10_11 b_10 NI_10 NS_11 0 -1.0872150345258983e-05
GC_10_12 b_10 NI_10 NS_12 0 -1.2341723616378468e-05
GC_10_13 b_10 NI_10 NS_13 0 6.1561717422595739e-11
GC_10_14 b_10 NI_10 NS_14 0 -1.1197712625369318e-11
GC_10_15 b_10 NI_10 NS_15 0 -5.2525161179638561e-10
GC_10_16 b_10 NI_10 NS_16 0 5.2974149659523726e-10
GC_10_17 b_10 NI_10 NS_17 0 -1.9707047274849773e-10
GC_10_18 b_10 NI_10 NS_18 0 7.7308633394361422e-12
GC_10_19 b_10 NI_10 NS_19 0 3.8927241323855159e-07
GC_10_20 b_10 NI_10 NS_20 0 -1.0156602593045327e-06
GC_10_21 b_10 NI_10 NS_21 0 -5.7479694200016743e-10
GC_10_22 b_10 NI_10 NS_22 0 -1.0307943300552595e-10
GC_10_23 b_10 NI_10 NS_23 0 8.1837463867978683e-12
GC_10_24 b_10 NI_10 NS_24 0 1.6175567064946581e-10
GC_10_25 b_10 NI_10 NS_25 0 -7.3290023175568516e-06
GC_10_26 b_10 NI_10 NS_26 0 -4.0590082406086083e-06
GC_10_27 b_10 NI_10 NS_27 0 -6.1708461562149952e-06
GC_10_28 b_10 NI_10 NS_28 0 4.5657990433808146e-06
GC_10_29 b_10 NI_10 NS_29 0 4.0300264050314431e-06
GC_10_30 b_10 NI_10 NS_30 0 2.8274380428784951e-06
GC_10_31 b_10 NI_10 NS_31 0 -1.1935951243841271e-11
GC_10_32 b_10 NI_10 NS_32 0 6.8028785912816850e-11
GC_10_33 b_10 NI_10 NS_33 0 1.8164615498213222e-10
GC_10_34 b_10 NI_10 NS_34 0 -4.3608435610263090e-10
GC_10_35 b_10 NI_10 NS_35 0 -2.6379398442280224e-11
GC_10_36 b_10 NI_10 NS_36 0 -2.3945833226780232e-10
GC_10_37 b_10 NI_10 NS_37 0 1.5414270286854150e-06
GC_10_38 b_10 NI_10 NS_38 0 -6.2760729160537937e-06
GC_10_39 b_10 NI_10 NS_39 0 1.3208823934427733e-10
GC_10_40 b_10 NI_10 NS_40 0 1.2903215729601963e-10
GC_10_41 b_10 NI_10 NS_41 0 -1.4443364587857641e-11
GC_10_42 b_10 NI_10 NS_42 0 3.5536541786684973e-10
GC_10_43 b_10 NI_10 NS_43 0 -7.0220260359262546e-06
GC_10_44 b_10 NI_10 NS_44 0 -7.1280520696980027e-06
GC_10_45 b_10 NI_10 NS_45 0 1.6303010717449094e-05
GC_10_46 b_10 NI_10 NS_46 0 -7.6034191659719846e-06
GC_10_47 b_10 NI_10 NS_47 0 -3.1089981034529254e-05
GC_10_48 b_10 NI_10 NS_48 0 -4.7345831765377353e-05
GC_10_49 b_10 NI_10 NS_49 0 -5.4798252063622286e-11
GC_10_50 b_10 NI_10 NS_50 0 1.7570984552652906e-10
GC_10_51 b_10 NI_10 NS_51 0 3.7966216764276289e-10
GC_10_52 b_10 NI_10 NS_52 0 -1.1576231950203590e-09
GC_10_53 b_10 NI_10 NS_53 0 -2.0690970375507239e-10
GC_10_54 b_10 NI_10 NS_54 0 1.5378512100640154e-10
GC_10_55 b_10 NI_10 NS_55 0 -8.0169988237043142e-07
GC_10_56 b_10 NI_10 NS_56 0 2.7307651291393049e-06
GC_10_57 b_10 NI_10 NS_57 0 -5.2077949140299834e-10
GC_10_58 b_10 NI_10 NS_58 0 -1.3300219605795564e-10
GC_10_59 b_10 NI_10 NS_59 0 1.4437311440500696e-11
GC_10_60 b_10 NI_10 NS_60 0 -3.0343762405432536e-10
GC_10_61 b_10 NI_10 NS_61 0 -1.8013126555606728e-06
GC_10_62 b_10 NI_10 NS_62 0 2.7925982272787971e-05
GC_10_63 b_10 NI_10 NS_63 0 1.0912795120291719e-05
GC_10_64 b_10 NI_10 NS_64 0 4.2540322631156602e-05
GC_10_65 b_10 NI_10 NS_65 0 4.9978014114617042e-05
GC_10_66 b_10 NI_10 NS_66 0 2.6934669415090535e-05
GC_10_67 b_10 NI_10 NS_67 0 7.0564923289528974e-11
GC_10_68 b_10 NI_10 NS_68 0 -1.8189062851449014e-10
GC_10_69 b_10 NI_10 NS_69 0 -4.0119657191552183e-10
GC_10_70 b_10 NI_10 NS_70 0 1.2111202563254734e-09
GC_10_71 b_10 NI_10 NS_71 0 1.8458101286471237e-10
GC_10_72 b_10 NI_10 NS_72 0 -1.7359412033107446e-10
GC_10_73 b_10 NI_10 NS_73 0 6.2470784847992300e-06
GC_10_74 b_10 NI_10 NS_74 0 -2.3041069985890719e-06
GC_10_75 b_10 NI_10 NS_75 0 2.4897760142896270e-08
GC_10_76 b_10 NI_10 NS_76 0 6.7284764328680034e-10
GC_10_77 b_10 NI_10 NS_77 0 -7.9766298446250778e-11
GC_10_78 b_10 NI_10 NS_78 0 4.2094443670091255e-09
GC_10_79 b_10 NI_10 NS_79 0 -1.3706988849886210e-04
GC_10_80 b_10 NI_10 NS_80 0 1.8416330431543919e-04
GC_10_81 b_10 NI_10 NS_81 0 8.0545714942204026e-04
GC_10_82 b_10 NI_10 NS_82 0 2.0808559140982711e-04
GC_10_83 b_10 NI_10 NS_83 0 -5.4267688617526497e-04
GC_10_84 b_10 NI_10 NS_84 0 -8.9938076638039054e-04
GC_10_85 b_10 NI_10 NS_85 0 -1.4819398513039701e-10
GC_10_86 b_10 NI_10 NS_86 0 8.6937274443357732e-10
GC_10_87 b_10 NI_10 NS_87 0 1.8613811898591580e-09
GC_10_88 b_10 NI_10 NS_88 0 -4.9451588845779512e-09
GC_10_89 b_10 NI_10 NS_89 0 -9.7922544505946375e-10
GC_10_90 b_10 NI_10 NS_90 0 6.4654579132142772e-10
GC_10_91 b_10 NI_10 NS_91 0 -1.3595252265375923e-05
GC_10_92 b_10 NI_10 NS_92 0 4.5592973334838163e-05
GC_10_93 b_10 NI_10 NS_93 0 -1.5019930431323923e-08
GC_10_94 b_10 NI_10 NS_94 0 -6.4644638273758834e-10
GC_10_95 b_10 NI_10 NS_95 0 7.9994592590083805e-11
GC_10_96 b_10 NI_10 NS_96 0 -4.9840747939464921e-09
GC_10_97 b_10 NI_10 NS_97 0 1.1992735779931157e-04
GC_10_98 b_10 NI_10 NS_98 0 1.7682256127282247e-04
GC_10_99 b_10 NI_10 NS_99 0 3.0863511228104853e-04
GC_10_100 b_10 NI_10 NS_100 0 -5.1613131842066296e-04
GC_10_101 b_10 NI_10 NS_101 0 -3.8644931045963199e-04
GC_10_102 b_10 NI_10 NS_102 0 1.7101790953782272e-04
GC_10_103 b_10 NI_10 NS_103 0 -2.6793836517100570e-10
GC_10_104 b_10 NI_10 NS_104 0 -8.7398300674065339e-10
GC_10_105 b_10 NI_10 NS_105 0 -9.6236027112918874e-10
GC_10_106 b_10 NI_10 NS_106 0 3.6733300830094019e-09
GC_10_107 b_10 NI_10 NS_107 0 1.2868996921610642e-09
GC_10_108 b_10 NI_10 NS_108 0 -4.8000103447530120e-10
GC_10_109 b_10 NI_10 NS_109 0 1.3240975244465316e-04
GC_10_110 b_10 NI_10 NS_110 0 -4.8360898895402095e-04
GC_10_111 b_10 NI_10 NS_111 0 7.2274922338357090e-08
GC_10_112 b_10 NI_10 NS_112 0 5.7680093856425637e-10
GC_10_113 b_10 NI_10 NS_113 0 -1.2176702400056837e-10
GC_10_114 b_10 NI_10 NS_114 0 6.5844045328419458e-08
GC_10_115 b_10 NI_10 NS_115 0 -1.7781545777753184e-04
GC_10_116 b_10 NI_10 NS_116 0 -2.2251465941635598e-03
GC_10_117 b_10 NI_10 NS_117 0 -2.2110764827275166e-03
GC_10_118 b_10 NI_10 NS_118 0 -2.2403402123928077e-03
GC_10_119 b_10 NI_10 NS_119 0 -1.5810875397457192e-03
GC_10_120 b_10 NI_10 NS_120 0 -5.3337320991300101e-04
GC_10_121 b_10 NI_10 NS_121 0 1.3213654894722097e-09
GC_10_122 b_10 NI_10 NS_122 0 6.9363403847693651e-09
GC_10_123 b_10 NI_10 NS_123 0 9.3019045812012425e-09
GC_10_124 b_10 NI_10 NS_124 0 -2.8759814162717403e-08
GC_10_125 b_10 NI_10 NS_125 0 -1.9780447967327702e-08
GC_10_126 b_10 NI_10 NS_126 0 -1.2715117614295912e-08
GC_10_127 b_10 NI_10 NS_127 0 -2.2349796628066024e-04
GC_10_128 b_10 NI_10 NS_128 0 6.5299174322880826e-04
GC_10_129 b_10 NI_10 NS_129 0 -1.5297642578197977e-07
GC_10_130 b_10 NI_10 NS_130 0 -6.5220673864618102e-10
GC_10_131 b_10 NI_10 NS_131 0 1.1968302352129459e-10
GC_10_132 b_10 NI_10 NS_132 0 -8.1050572289999873e-08
GC_10_133 b_10 NI_10 NS_133 0 -4.6083746142690316e-04
GC_10_134 b_10 NI_10 NS_134 0 4.9882322218590871e-03
GC_10_135 b_10 NI_10 NS_135 0 4.0337280072722656e-03
GC_10_136 b_10 NI_10 NS_136 0 -5.0074968246527883e-04
GC_10_137 b_10 NI_10 NS_137 0 2.5275259435490645e-03
GC_10_138 b_10 NI_10 NS_138 0 6.9892930145049039e-03
GC_10_139 b_10 NI_10 NS_139 0 -7.4263833898889731e-09
GC_10_140 b_10 NI_10 NS_140 0 -1.1198914380435685e-08
GC_10_141 b_10 NI_10 NS_141 0 7.8014501221587651e-09
GC_10_142 b_10 NI_10 NS_142 0 2.1845409806378677e-08
GC_10_143 b_10 NI_10 NS_143 0 2.3385362238941079e-08
GC_10_144 b_10 NI_10 NS_144 0 1.3786903194275570e-08
GC_10_145 b_10 NI_10 NS_145 0 1.2607267693462253e-02
GC_10_146 b_10 NI_10 NS_146 0 -3.4706344939961088e-02
GC_10_147 b_10 NI_10 NS_147 0 -1.6753037726520218e-05
GC_10_148 b_10 NI_10 NS_148 0 -8.5055606098946420e-07
GC_10_149 b_10 NI_10 NS_149 0 1.4723651281951992e-08
GC_10_150 b_10 NI_10 NS_150 0 1.0162709738722764e-05
GC_10_151 b_10 NI_10 NS_151 0 -4.6995196379457468e-02
GC_10_152 b_10 NI_10 NS_152 0 6.7612396120797794e-02
GC_10_153 b_10 NI_10 NS_153 0 -2.4545310444848416e-02
GC_10_154 b_10 NI_10 NS_154 0 -1.6180126302219064e-01
GC_10_155 b_10 NI_10 NS_155 0 -1.3230847882810549e-02
GC_10_156 b_10 NI_10 NS_156 0 -1.8253997408146591e-01
GC_10_157 b_10 NI_10 NS_157 0 5.7566500679306494e-07
GC_10_158 b_10 NI_10 NS_158 0 1.0761899108153395e-06
GC_10_159 b_10 NI_10 NS_159 0 -5.4558660556498877e-06
GC_10_160 b_10 NI_10 NS_160 0 2.2858409596367304e-07
GC_10_161 b_10 NI_10 NS_161 0 -4.0753565811990145e-06
GC_10_162 b_10 NI_10 NS_162 0 -4.3093294768617003e-06
GC_10_163 b_10 NI_10 NS_163 0 -4.8625241773539172e-03
GC_10_164 b_10 NI_10 NS_164 0 1.6965213023596187e-02
GC_10_165 b_10 NI_10 NS_165 0 -3.4509061476515244e-06
GC_10_166 b_10 NI_10 NS_166 0 2.9323276789306986e-08
GC_10_167 b_10 NI_10 NS_167 0 -1.0119702754068433e-09
GC_10_168 b_10 NI_10 NS_168 0 -2.0010662620436756e-06
GC_10_169 b_10 NI_10 NS_169 0 1.8510763516678318e-02
GC_10_170 b_10 NI_10 NS_170 0 5.0676143484218297e-02
GC_10_171 b_10 NI_10 NS_171 0 1.4775875168050548e-02
GC_10_172 b_10 NI_10 NS_172 0 7.2025344573511493e-02
GC_10_173 b_10 NI_10 NS_173 0 8.2113614999535706e-02
GC_10_174 b_10 NI_10 NS_174 0 4.9907424272148948e-02
GC_10_175 b_10 NI_10 NS_175 0 -2.8706263305241943e-07
GC_10_176 b_10 NI_10 NS_176 0 -5.8605014838287046e-08
GC_10_177 b_10 NI_10 NS_177 0 5.7101018782250183e-07
GC_10_178 b_10 NI_10 NS_178 0 -8.2174834855094152e-07
GC_10_179 b_10 NI_10 NS_179 0 3.9089970822309507e-07
GC_10_180 b_10 NI_10 NS_180 0 3.8092737133245112e-07
GC_10_181 b_10 NI_10 NS_181 0 1.1715003262804903e-04
GC_10_182 b_10 NI_10 NS_182 0 -4.6263179101779171e-04
GC_10_183 b_10 NI_10 NS_183 0 3.5653867165640451e-07
GC_10_184 b_10 NI_10 NS_184 0 3.4767107639531898e-09
GC_10_185 b_10 NI_10 NS_185 0 -1.1870437739671925e-11
GC_10_186 b_10 NI_10 NS_186 0 1.2107854277678194e-07
GC_10_187 b_10 NI_10 NS_187 0 7.0305739732629642e-04
GC_10_188 b_10 NI_10 NS_188 0 -4.2879088196309100e-03
GC_10_189 b_10 NI_10 NS_189 0 -9.0097307066240376e-03
GC_10_190 b_10 NI_10 NS_190 0 -5.1466471061271200e-03
GC_10_191 b_10 NI_10 NS_191 0 1.8363219535182031e-03
GC_10_192 b_10 NI_10 NS_192 0 7.2289144477589266e-03
GC_10_193 b_10 NI_10 NS_193 0 4.0590057682415761e-09
GC_10_194 b_10 NI_10 NS_194 0 2.5523055992276649e-09
GC_10_195 b_10 NI_10 NS_195 0 1.9338918151140998e-09
GC_10_196 b_10 NI_10 NS_196 0 1.2043039205112779e-08
GC_10_197 b_10 NI_10 NS_197 0 -2.5390686897210691e-08
GC_10_198 b_10 NI_10 NS_198 0 -1.4677114198394727e-08
GC_10_199 b_10 NI_10 NS_199 0 -6.0676042028037325e-04
GC_10_200 b_10 NI_10 NS_200 0 1.3746653341934624e-03
GC_10_201 b_10 NI_10 NS_201 0 -8.5831351745426601e-07
GC_10_202 b_10 NI_10 NS_202 0 -1.4313973234058509e-09
GC_10_203 b_10 NI_10 NS_203 0 -2.7382267265159473e-11
GC_10_204 b_10 NI_10 NS_204 0 -2.1428671077543280e-07
GC_10_205 b_10 NI_10 NS_205 0 -4.2092983853928758e-03
GC_10_206 b_10 NI_10 NS_206 0 1.9038706064528520e-02
GC_10_207 b_10 NI_10 NS_207 0 1.8776114831012321e-02
GC_10_208 b_10 NI_10 NS_208 0 -1.2054743222192665e-02
GC_10_209 b_10 NI_10 NS_209 0 2.1761177234677449e-03
GC_10_210 b_10 NI_10 NS_210 0 2.9277545523638697e-02
GC_10_211 b_10 NI_10 NS_211 0 -3.3733555840034811e-08
GC_10_212 b_10 NI_10 NS_212 0 -2.4556561536182975e-08
GC_10_213 b_10 NI_10 NS_213 0 8.1304153767320699e-08
GC_10_214 b_10 NI_10 NS_214 0 -4.2403234615662603e-08
GC_10_215 b_10 NI_10 NS_215 0 5.1539380829254385e-08
GC_10_216 b_10 NI_10 NS_216 0 3.1346607738466187e-08
GD_10_1 b_10 NI_10 NA_1 0 -5.7715692851269892e-08
GD_10_2 b_10 NI_10 NA_2 0 9.6627040503157213e-06
GD_10_3 b_10 NI_10 NA_3 0 1.8865360247530740e-05
GD_10_4 b_10 NI_10 NA_4 0 -3.3983508300049610e-05
GD_10_5 b_10 NI_10 NA_5 0 -3.5096772060018101e-05
GD_10_6 b_10 NI_10 NA_6 0 6.4162387199213501e-05
GD_10_7 b_10 NI_10 NA_7 0 2.6224374685507403e-03
GD_10_8 b_10 NI_10 NA_8 0 -9.9222313821831112e-04
GD_10_9 b_10 NI_10 NA_9 0 7.4457060564165178e-02
GD_10_10 b_10 NI_10 NA_10 0 -9.3789405414097818e-02
GD_10_11 b_10 NI_10 NA_11 0 3.7903418651203946e-03
GD_10_12 b_10 NI_10 NA_12 0 6.2401033715778244e-03
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 5.8599351662876957e-07
GC_11_2 b_11 NI_11 NS_2 0 -2.8557188028715044e-06
GC_11_3 b_11 NI_11 NS_3 0 1.7703516639267529e-09
GC_11_4 b_11 NI_11 NS_4 0 -6.7055574052486345e-11
GC_11_5 b_11 NI_11 NS_5 0 7.5216487137152996e-12
GC_11_6 b_11 NI_11 NS_6 0 -2.8671208732283030e-10
GC_11_7 b_11 NI_11 NS_7 0 -9.9060965130652307e-07
GC_11_8 b_11 NI_11 NS_8 0 -1.1239024882047723e-05
GC_11_9 b_11 NI_11 NS_9 0 -3.8455034358377907e-06
GC_11_10 b_11 NI_11 NS_10 0 -1.2012617478031317e-05
GC_11_11 b_11 NI_11 NS_11 0 -1.5710129155198825e-05
GC_11_12 b_11 NI_11 NS_12 0 -1.4373072368433406e-05
GC_11_13 b_11 NI_11 NS_13 0 2.7242073409567468e-12
GC_11_14 b_11 NI_11 NS_14 0 4.8464683250498086e-11
GC_11_15 b_11 NI_11 NS_15 0 -1.0542545215669699e-10
GC_11_16 b_11 NI_11 NS_16 0 9.2933564570387327e-11
GC_11_17 b_11 NI_11 NS_17 0 1.5680746627247929e-10
GC_11_18 b_11 NI_11 NS_18 0 -8.5166515356961405e-11
GC_11_19 b_11 NI_11 NS_19 0 -9.7454420465076694e-07
GC_11_20 b_11 NI_11 NS_20 0 4.1608357144702174e-06
GC_11_21 b_11 NI_11 NS_21 0 -1.1208170911508561e-09
GC_11_22 b_11 NI_11 NS_22 0 8.2924956741568467e-11
GC_11_23 b_11 NI_11 NS_23 0 -7.7974462091997435e-12
GC_11_24 b_11 NI_11 NS_24 0 1.3118852408950946e-10
GC_11_25 b_11 NI_11 NS_25 0 8.4582217121867794e-07
GC_11_26 b_11 NI_11 NS_26 0 1.3225653330554336e-05
GC_11_27 b_11 NI_11 NS_27 0 3.8098611421303986e-06
GC_11_28 b_11 NI_11 NS_28 0 1.4582517249747191e-05
GC_11_29 b_11 NI_11 NS_29 0 1.9310561854102851e-05
GC_11_30 b_11 NI_11 NS_30 0 1.9670562104515436e-05
GC_11_31 b_11 NI_11 NS_31 0 -1.5170737895296790e-11
GC_11_32 b_11 NI_11 NS_32 0 -6.4678318689623877e-11
GC_11_33 b_11 NI_11 NS_33 0 2.1121376106637269e-10
GC_11_34 b_11 NI_11 NS_34 0 -1.1076899281948695e-10
GC_11_35 b_11 NI_11 NS_35 0 -8.5473400775447523e-11
GC_11_36 b_11 NI_11 NS_36 0 1.5980375683624584e-10
GC_11_37 b_11 NI_11 NS_37 0 3.9250788939246375e-07
GC_11_38 b_11 NI_11 NS_38 0 -1.0348234494328024e-06
GC_11_39 b_11 NI_11 NS_39 0 -5.7480802916610032e-10
GC_11_40 b_11 NI_11 NS_40 0 -1.0318287873828327e-10
GC_11_41 b_11 NI_11 NS_41 0 8.1893952203640633e-12
GC_11_42 b_11 NI_11 NS_42 0 1.6240289891491812e-10
GC_11_43 b_11 NI_11 NS_43 0 -7.3298750972589444e-06
GC_11_44 b_11 NI_11 NS_44 0 -4.1640116203144945e-06
GC_11_45 b_11 NI_11 NS_45 0 -6.2106534101646233e-06
GC_11_46 b_11 NI_11 NS_46 0 4.4397894246204982e-06
GC_11_47 b_11 NI_11 NS_47 0 3.8725825732232146e-06
GC_11_48 b_11 NI_11 NS_48 0 2.7044160956719901e-06
GC_11_49 b_11 NI_11 NS_49 0 -1.1963647395351047e-11
GC_11_50 b_11 NI_11 NS_50 0 6.8480034724912576e-11
GC_11_51 b_11 NI_11 NS_51 0 1.8113597925081147e-10
GC_11_52 b_11 NI_11 NS_52 0 -4.3693339070409786e-10
GC_11_53 b_11 NI_11 NS_53 0 -2.6690058169231549e-11
GC_11_54 b_11 NI_11 NS_54 0 -2.3988044465959317e-10
GC_11_55 b_11 NI_11 NS_55 0 6.6414536849303962e-07
GC_11_56 b_11 NI_11 NS_56 0 -2.2652822376305330e-06
GC_11_57 b_11 NI_11 NS_57 0 -1.5864254264735526e-09
GC_11_58 b_11 NI_11 NS_58 0 5.4093447380226936e-11
GC_11_59 b_11 NI_11 NS_59 0 -7.3828947351132501e-12
GC_11_60 b_11 NI_11 NS_60 0 3.2373919917316196e-10
GC_11_61 b_11 NI_11 NS_61 0 4.0928293613284659e-06
GC_11_62 b_11 NI_11 NS_62 0 -3.9935326503211818e-06
GC_11_63 b_11 NI_11 NS_63 0 3.0987042875647203e-06
GC_11_64 b_11 NI_11 NS_64 0 -8.2597393682632049e-06
GC_11_65 b_11 NI_11 NS_65 0 -1.0642246681120921e-05
GC_11_66 b_11 NI_11 NS_66 0 -1.2162049038274966e-05
GC_11_67 b_11 NI_11 NS_67 0 6.1530413937145673e-11
GC_11_68 b_11 NI_11 NS_68 0 -1.1718204863877842e-11
GC_11_69 b_11 NI_11 NS_69 0 -5.2416367076875901e-10
GC_11_70 b_11 NI_11 NS_70 0 5.3037974639037820e-10
GC_11_71 b_11 NI_11 NS_71 0 -1.9630600620697532e-10
GC_11_72 b_11 NI_11 NS_72 0 8.6277375512586017e-12
GC_11_73 b_11 NI_11 NS_73 0 1.3355196328839327e-06
GC_11_74 b_11 NI_11 NS_74 0 -7.7290135864804498e-06
GC_11_75 b_11 NI_11 NS_75 0 -3.8707219108809598e-09
GC_11_76 b_11 NI_11 NS_76 0 -2.4408416564591406e-10
GC_11_77 b_11 NI_11 NS_77 0 2.5141281234588547e-11
GC_11_78 b_11 NI_11 NS_78 0 -1.0237015043767712e-10
GC_11_79 b_11 NI_11 NS_79 0 -3.6243704231856951e-05
GC_11_80 b_11 NI_11 NS_80 0 5.2155783521963840e-05
GC_11_81 b_11 NI_11 NS_81 0 7.6127037109132092e-06
GC_11_82 b_11 NI_11 NS_82 0 1.4079630107333624e-04
GC_11_83 b_11 NI_11 NS_83 0 1.5327481261126851e-04
GC_11_84 b_11 NI_11 NS_84 0 4.9519569888706793e-05
GC_11_85 b_11 NI_11 NS_85 0 6.2161467482129402e-11
GC_11_86 b_11 NI_11 NS_86 0 -1.1934444845337780e-10
GC_11_87 b_11 NI_11 NS_87 0 -3.5746489556616456e-10
GC_11_88 b_11 NI_11 NS_88 0 1.0385954787010303e-09
GC_11_89 b_11 NI_11 NS_89 0 5.0039319053567322e-11
GC_11_90 b_11 NI_11 NS_90 0 -4.5803716081382440e-10
GC_11_91 b_11 NI_11 NS_91 0 4.4584379019650565e-06
GC_11_92 b_11 NI_11 NS_92 0 -1.7990473294388364e-05
GC_11_93 b_11 NI_11 NS_93 0 -4.6680548378283724e-10
GC_11_94 b_11 NI_11 NS_94 0 2.1056605772859050e-10
GC_11_95 b_11 NI_11 NS_95 0 -2.4757395406792079e-11
GC_11_96 b_11 NI_11 NS_96 0 6.0795979404268077e-10
GC_11_97 b_11 NI_11 NS_97 0 -1.3683880474126802e-05
GC_11_98 b_11 NI_11 NS_98 0 5.5046874464740285e-05
GC_11_99 b_11 NI_11 NS_99 0 1.4849988594838596e-04
GC_11_100 b_11 NI_11 NS_100 0 4.5509315863931752e-05
GC_11_101 b_11 NI_11 NS_101 0 -6.2796698875301204e-05
GC_11_102 b_11 NI_11 NS_102 0 -1.8722343244126501e-04
GC_11_103 b_11 NI_11 NS_103 0 1.7529354234019027e-10
GC_11_104 b_11 NI_11 NS_104 0 1.3267732449348800e-10
GC_11_105 b_11 NI_11 NS_105 0 -2.2723762982055061e-10
GC_11_106 b_11 NI_11 NS_106 0 -4.2066433953060878e-10
GC_11_107 b_11 NI_11 NS_107 0 -2.5484748622363522e-10
GC_11_108 b_11 NI_11 NS_108 0 2.9867702752572345e-10
GC_11_109 b_11 NI_11 NS_109 0 -1.3260448147631601e-05
GC_11_110 b_11 NI_11 NS_110 0 4.4076050817433157e-05
GC_11_111 b_11 NI_11 NS_111 0 -1.4697575316644946e-08
GC_11_112 b_11 NI_11 NS_112 0 -6.5126882288445405e-10
GC_11_113 b_11 NI_11 NS_113 0 8.0654532504362192e-11
GC_11_114 b_11 NI_11 NS_114 0 -5.0535486116198736e-09
GC_11_115 b_11 NI_11 NS_115 0 1.1931482918595472e-04
GC_11_116 b_11 NI_11 NS_116 0 1.7067296747719839e-04
GC_11_117 b_11 NI_11 NS_117 0 3.0643937064365562e-04
GC_11_118 b_11 NI_11 NS_118 0 -5.2287913331659742e-04
GC_11_119 b_11 NI_11 NS_119 0 -3.9525301403668992e-04
GC_11_120 b_11 NI_11 NS_120 0 1.6327254070788895e-04
GC_11_121 b_11 NI_11 NS_121 0 -2.5837383887396844e-10
GC_11_122 b_11 NI_11 NS_122 0 -8.5878770716313851e-10
GC_11_123 b_11 NI_11 NS_123 0 -1.0039908558418978e-09
GC_11_124 b_11 NI_11 NS_124 0 3.7270542822885129e-09
GC_11_125 b_11 NI_11 NS_125 0 1.3187435172786510e-09
GC_11_126 b_11 NI_11 NS_126 0 -4.7771920277602417e-10
GC_11_127 b_11 NI_11 NS_127 0 6.0001220961010325e-06
GC_11_128 b_11 NI_11 NS_128 0 -1.2007057888774978e-06
GC_11_129 b_11 NI_11 NS_129 0 2.4512811490136126e-08
GC_11_130 b_11 NI_11 NS_130 0 6.7664016595104043e-10
GC_11_131 b_11 NI_11 NS_131 0 -8.0405954235565297e-11
GC_11_132 b_11 NI_11 NS_132 0 4.2877295718022152e-09
GC_11_133 b_11 NI_11 NS_133 0 -1.3622076861739398e-04
GC_11_134 b_11 NI_11 NS_134 0 1.9072648581303162e-04
GC_11_135 b_11 NI_11 NS_135 0 8.0919478489583805e-04
GC_11_136 b_11 NI_11 NS_136 0 2.1471687001120912e-04
GC_11_137 b_11 NI_11 NS_137 0 -5.3483841131123501e-04
GC_11_138 b_11 NI_11 NS_138 0 -8.9414154535085062e-04
GC_11_139 b_11 NI_11 NS_139 0 -1.5409842703791198e-10
GC_11_140 b_11 NI_11 NS_140 0 8.5208755933487378e-10
GC_11_141 b_11 NI_11 NS_141 0 1.8956751216811950e-09
GC_11_142 b_11 NI_11 NS_142 0 -4.9875673806232023e-09
GC_11_143 b_11 NI_11 NS_143 0 -1.0147524819428253e-09
GC_11_144 b_11 NI_11 NS_144 0 6.4011215198893525e-10
GC_11_145 b_11 NI_11 NS_145 0 -6.0676042028494186e-04
GC_11_146 b_11 NI_11 NS_146 0 1.3746653342055842e-03
GC_11_147 b_11 NI_11 NS_147 0 -8.5831351744235016e-07
GC_11_148 b_11 NI_11 NS_148 0 -1.4313973233811234e-09
GC_11_149 b_11 NI_11 NS_149 0 -2.7382267261591869e-11
GC_11_150 b_11 NI_11 NS_150 0 -2.1428671077666619e-07
GC_11_151 b_11 NI_11 NS_151 0 -4.2092983853895261e-03
GC_11_152 b_11 NI_11 NS_152 0 1.9038706064518289e-02
GC_11_153 b_11 NI_11 NS_153 0 1.8776114830996869e-02
GC_11_154 b_11 NI_11 NS_154 0 -1.2054743222198050e-02
GC_11_155 b_11 NI_11 NS_155 0 2.1761177234662699e-03
GC_11_156 b_11 NI_11 NS_156 0 2.9277545523667889e-02
GC_11_157 b_11 NI_11 NS_157 0 -3.3733555840636515e-08
GC_11_158 b_11 NI_11 NS_158 0 -2.4556561536787286e-08
GC_11_159 b_11 NI_11 NS_159 0 8.1304153769808831e-08
GC_11_160 b_11 NI_11 NS_160 0 -4.2403234616962878e-08
GC_11_161 b_11 NI_11 NS_161 0 5.1539380829752030e-08
GC_11_162 b_11 NI_11 NS_162 0 3.1346607738649774e-08
GC_11_163 b_11 NI_11 NS_163 0 1.1714737736095258e-04
GC_11_164 b_11 NI_11 NS_164 0 -4.6262295740927154e-04
GC_11_165 b_11 NI_11 NS_165 0 3.5654165105478963e-07
GC_11_166 b_11 NI_11 NS_166 0 3.4767317445826717e-09
GC_11_167 b_11 NI_11 NS_167 0 -1.1870736283042499e-11
GC_11_168 b_11 NI_11 NS_168 0 1.2107815922896925e-07
GC_11_169 b_11 NI_11 NS_169 0 7.0304718103259987e-04
GC_11_170 b_11 NI_11 NS_170 0 -4.2878840224376746e-03
GC_11_171 b_11 NI_11 NS_171 0 -9.0097181772219332e-03
GC_11_172 b_11 NI_11 NS_172 0 -5.1465729595455180e-03
GC_11_173 b_11 NI_11 NS_173 0 1.8363876527587087e-03
GC_11_174 b_11 NI_11 NS_174 0 7.2289510870847031e-03
GC_11_175 b_11 NI_11 NS_175 0 4.0587608400121539e-09
GC_11_176 b_11 NI_11 NS_176 0 2.5522864847883853e-09
GC_11_177 b_11 NI_11 NS_177 0 1.9345086017631886e-09
GC_11_178 b_11 NI_11 NS_178 0 1.2042396197724021e-08
GC_11_179 b_11 NI_11 NS_179 0 -2.5390538262059749e-08
GC_11_180 b_11 NI_11 NS_180 0 -1.4677008598052108e-08
GC_11_181 b_11 NI_11 NS_181 0 -4.7894741477343033e-03
GC_11_182 b_11 NI_11 NS_182 0 1.6721231895482244e-02
GC_11_183 b_11 NI_11 NS_183 0 -3.5217425139628847e-06
GC_11_184 b_11 NI_11 NS_184 0 2.9869341329959534e-08
GC_11_185 b_11 NI_11 NS_185 0 -1.0050510000652857e-09
GC_11_186 b_11 NI_11 NS_186 0 -2.0070261998670490e-06
GC_11_187 b_11 NI_11 NS_187 0 1.8815079487226709e-02
GC_11_188 b_11 NI_11 NS_188 0 5.0642922456182377e-02
GC_11_189 b_11 NI_11 NS_189 0 1.5086435845925224e-02
GC_11_190 b_11 NI_11 NS_190 0 7.1442548787440066e-02
GC_11_191 b_11 NI_11 NS_191 0 8.1541997974417441e-02
GC_11_192 b_11 NI_11 NS_192 0 4.9085291802314433e-02
GC_11_193 b_11 NI_11 NS_193 0 -2.7438712865958463e-07
GC_11_194 b_11 NI_11 NS_194 0 -6.0490113085660793e-08
GC_11_195 b_11 NI_11 NS_195 0 5.2038320036497312e-07
GC_11_196 b_11 NI_11 NS_196 0 -7.4412561535700476e-07
GC_11_197 b_11 NI_11 NS_197 0 3.9436032396737081e-07
GC_11_198 b_11 NI_11 NS_198 0 3.8383217890927020e-07
GC_11_199 b_11 NI_11 NS_199 0 1.0850981253409669e-02
GC_11_200 b_11 NI_11 NS_200 0 -2.9612919587297556e-02
GC_11_201 b_11 NI_11 NS_201 0 -1.0888096618531933e-05
GC_11_202 b_11 NI_11 NS_202 0 -6.9604747796075289e-07
GC_11_203 b_11 NI_11 NS_203 0 1.2495231273965843e-08
GC_11_204 b_11 NI_11 NS_204 0 8.6529085445556590e-06
GC_11_205 b_11 NI_11 NS_205 0 -5.1293374942927752e-02
GC_11_206 b_11 NI_11 NS_206 0 6.8705043503144020e-02
GC_11_207 b_11 NI_11 NS_207 0 -2.8913166683763536e-02
GC_11_208 b_11 NI_11 NS_208 0 -1.5463815912849158e-01
GC_11_209 b_11 NI_11 NS_209 0 -4.9850378997618235e-03
GC_11_210 b_11 NI_11 NS_210 0 -1.6599218152816389e-01
GC_11_211 b_11 NI_11 NS_211 0 4.7917150083603217e-07
GC_11_212 b_11 NI_11 NS_212 0 8.9026047260449411e-07
GC_11_213 b_11 NI_11 NS_213 0 -4.3716111455822139e-06
GC_11_214 b_11 NI_11 NS_214 0 1.1070894714174336e-07
GC_11_215 b_11 NI_11 NS_215 0 -3.3754134508189765e-06
GC_11_216 b_11 NI_11 NS_216 0 -3.5752637777674479e-06
GD_11_1 b_11 NI_11 NA_1 0 1.3354404010059112e-05
GD_11_2 b_11 NI_11 NA_2 0 -1.5515466013016709e-05
GD_11_3 b_11 NI_11 NA_3 0 9.7838301513855381e-06
GD_11_4 b_11 NI_11 NA_4 0 -2.5590821521708941e-07
GD_11_5 b_11 NI_11 NA_5 0 -4.9753082637498979e-05
GD_11_6 b_11 NI_11 NA_6 0 -2.8242995772377618e-05
GD_11_7 b_11 NI_11 NA_7 0 7.1764277194203435e-05
GD_11_8 b_11 NI_11 NA_8 0 -4.3070867735153526e-05
GD_11_9 b_11 NI_11 NA_9 0 6.2401033715774887e-03
GD_11_10 b_11 NI_11 NA_10 0 3.7902998081262174e-03
GD_11_11 b_11 NI_11 NA_11 0 -9.3789089811108631e-02
GD_11_12 b_11 NI_11 NA_12 0 7.4536667406035054e-02
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -9.7408003727919310e-07
GC_12_2 b_12 NI_12 NS_2 0 4.1595782768918854e-06
GC_12_3 b_12 NI_12 NS_3 0 -1.1230100446660965e-09
GC_12_4 b_12 NI_12 NS_4 0 8.2869325554978749e-11
GC_12_5 b_12 NI_12 NS_5 0 -7.7963410526970507e-12
GC_12_6 b_12 NI_12 NS_6 0 1.3172457631240127e-10
GC_12_7 b_12 NI_12 NS_7 0 8.4635070416212345e-07
GC_12_8 b_12 NI_12 NS_8 0 1.3226721189177532e-05
GC_12_9 b_12 NI_12 NS_9 0 3.8130675124236845e-06
GC_12_10 b_12 NI_12 NS_10 0 1.4579715766535772e-05
GC_12_11 b_12 NI_12 NS_11 0 1.9307448036928281e-05
GC_12_12 b_12 NI_12 NS_12 0 1.9665926923345126e-05
GC_12_13 b_12 NI_12 NS_13 0 -1.5099184302662235e-11
GC_12_14 b_12 NI_12 NS_14 0 -6.4634079380478948e-11
GC_12_15 b_12 NI_12 NS_15 0 2.1080319925127341e-10
GC_12_16 b_12 NI_12 NS_16 0 -1.1068236353236343e-10
GC_12_17 b_12 NI_12 NS_17 0 -8.5719261221123830e-11
GC_12_18 b_12 NI_12 NS_18 0 1.5954468157945352e-10
GC_12_19 b_12 NI_12 NS_19 0 5.8596941201015178e-07
GC_12_20 b_12 NI_12 NS_20 0 -2.8556058224307980e-06
GC_12_21 b_12 NI_12 NS_21 0 1.7704155022579094e-09
GC_12_22 b_12 NI_12 NS_22 0 -6.7054013773660450e-11
GC_12_23 b_12 NI_12 NS_23 0 7.5216562361715677e-12
GC_12_24 b_12 NI_12 NS_24 0 -2.8672924130577220e-10
GC_12_25 b_12 NI_12 NS_25 0 -9.9035559162213133e-07
GC_12_26 b_12 NI_12 NS_26 0 -1.1238119790856272e-05
GC_12_27 b_12 NI_12 NS_27 0 -3.8449973795517466e-06
GC_12_28 b_12 NI_12 NS_28 0 -1.2011771249127651e-05
GC_12_29 b_12 NI_12 NS_29 0 -1.5709041836659538e-05
GC_12_30 b_12 NI_12 NS_30 0 -1.4372424156688717e-05
GC_12_31 b_12 NI_12 NS_31 0 2.7225523038640652e-12
GC_12_32 b_12 NI_12 NS_32 0 4.8461603846966994e-11
GC_12_33 b_12 NI_12 NS_33 0 -1.0541230784015769e-10
GC_12_34 b_12 NI_12 NS_34 0 9.2934546109719611e-11
GC_12_35 b_12 NI_12 NS_35 0 1.5681550335846498e-10
GC_12_36 b_12 NI_12 NS_36 0 -8.5158576628771312e-11
GC_12_37 b_12 NI_12 NS_37 0 6.6412953826491942e-07
GC_12_38 b_12 NI_12 NS_38 0 -2.2652193686494505e-06
GC_12_39 b_12 NI_12 NS_39 0 -1.5864166454412178e-09
GC_12_40 b_12 NI_12 NS_40 0 5.4093616751522994e-11
GC_12_41 b_12 NI_12 NS_41 0 -7.3828935564380512e-12
GC_12_42 b_12 NI_12 NS_42 0 3.2373728756365922e-10
GC_12_43 b_12 NI_12 NS_43 0 4.0928043518999812e-06
GC_12_44 b_12 NI_12 NS_44 0 -3.9933763736918467e-06
GC_12_45 b_12 NI_12 NS_45 0 3.0987415603084823e-06
GC_12_46 b_12 NI_12 NS_46 0 -8.2595769316526287e-06
GC_12_47 b_12 NI_12 NS_47 0 -1.0642018845427815e-05
GC_12_48 b_12 NI_12 NS_48 0 -1.2161764829236832e-05
GC_12_49 b_12 NI_12 NS_49 0 6.1530268102773966e-11
GC_12_50 b_12 NI_12 NS_50 0 -1.1718478753821163e-11
GC_12_51 b_12 NI_12 NS_51 0 -5.2416214760218687e-10
GC_12_52 b_12 NI_12 NS_52 0 5.3037941096849133e-10
GC_12_53 b_12 NI_12 NS_53 0 -1.9630511764493030e-10
GC_12_54 b_12 NI_12 NS_54 0 8.6286024612043468e-12
GC_12_55 b_12 NI_12 NS_55 0 4.0746212568714463e-07
GC_12_56 b_12 NI_12 NS_56 0 -1.0805037158953834e-06
GC_12_57 b_12 NI_12 NS_57 0 -6.0121239297065770e-10
GC_12_58 b_12 NI_12 NS_58 0 -1.0370636878324355e-10
GC_12_59 b_12 NI_12 NS_59 0 8.2022252760456346e-12
GC_12_60 b_12 NI_12 NS_60 0 1.6745811758266334e-10
GC_12_61 b_12 NI_12 NS_61 0 -7.3117593933574441e-06
GC_12_62 b_12 NI_12 NS_62 0 -4.2280536771857507e-06
GC_12_63 b_12 NI_12 NS_63 0 -6.2102554110430477e-06
GC_12_64 b_12 NI_12 NS_64 0 4.3349177005806276e-06
GC_12_65 b_12 NI_12 NS_65 0 3.7519804780374591e-06
GC_12_66 b_12 NI_12 NS_66 0 2.5489721461894601e-06
GC_12_67 b_12 NI_12 NS_67 0 -1.1573378146508355e-11
GC_12_68 b_12 NI_12 NS_68 0 6.8390022929201226e-11
GC_12_69 b_12 NI_12 NS_69 0 1.7866336902597748e-10
GC_12_70 b_12 NI_12 NS_70 0 -4.3454381326512936e-10
GC_12_71 b_12 NI_12 NS_71 0 -2.8967414177890187e-11
GC_12_72 b_12 NI_12 NS_72 0 -2.4227180677407469e-10
GC_12_73 b_12 NI_12 NS_73 0 4.4889234398568224e-06
GC_12_74 b_12 NI_12 NS_74 0 -1.8090897376760230e-05
GC_12_75 b_12 NI_12 NS_75 0 -5.0679190160905628e-10
GC_12_76 b_12 NI_12 NS_76 0 2.1018087653962451e-10
GC_12_77 b_12 NI_12 NS_77 0 -2.4750708337632734e-11
GC_12_78 b_12 NI_12 NS_78 0 6.1365773826832188e-10
GC_12_79 b_12 NI_12 NS_79 0 -1.3564578130649979e-05
GC_12_80 b_12 NI_12 NS_80 0 5.4779565829704229e-05
GC_12_81 b_12 NI_12 NS_81 0 1.4837096224550099e-04
GC_12_82 b_12 NI_12 NS_82 0 4.4676735754534572e-05
GC_12_83 b_12 NI_12 NS_83 0 -6.3532201213046429e-05
GC_12_84 b_12 NI_12 NS_84 0 -1.8763781199191727e-04
GC_12_85 b_12 NI_12 NS_85 0 1.7826483365678780e-10
GC_12_86 b_12 NI_12 NS_86 0 1.3311006515286290e-10
GC_12_87 b_12 NI_12 NS_87 0 -2.3563934991453485e-10
GC_12_88 b_12 NI_12 NS_88 0 -4.1437930353049278e-10
GC_12_89 b_12 NI_12 NS_89 0 -2.5709565542935249e-10
GC_12_90 b_12 NI_12 NS_90 0 2.9692390596607439e-10
GC_12_91 b_12 NI_12 NS_91 0 1.3390391850501994e-06
GC_12_92 b_12 NI_12 NS_92 0 -7.7404819803201235e-06
GC_12_93 b_12 NI_12 NS_93 0 -3.8746468376827081e-09
GC_12_94 b_12 NI_12 NS_94 0 -2.4411480879633043e-10
GC_12_95 b_12 NI_12 NS_95 0 2.5141849931156409e-11
GC_12_96 b_12 NI_12 NS_96 0 -1.0189389204725251e-10
GC_12_97 b_12 NI_12 NS_97 0 -3.6245031269110127e-05
GC_12_98 b_12 NI_12 NS_98 0 5.2125784371440330e-05
GC_12_99 b_12 NI_12 NS_99 0 7.6021055494084750e-06
GC_12_100 b_12 NI_12 NS_100 0 1.4076152582916527e-04
GC_12_101 b_12 NI_12 NS_101 0 1.5323341831752934e-04
GC_12_102 b_12 NI_12 NS_102 0 4.9478016486416937e-05
GC_12_103 b_12 NI_12 NS_103 0 6.2298357841092054e-11
GC_12_104 b_12 NI_12 NS_104 0 -1.1932006108488397e-10
GC_12_105 b_12 NI_12 NS_105 0 -3.5791540070686572e-10
GC_12_106 b_12 NI_12 NS_106 0 1.0391251590689022e-09
GC_12_107 b_12 NI_12 NS_107 0 4.9855717621526005e-11
GC_12_108 b_12 NI_12 NS_108 0 -4.5817487404215792e-10
GC_12_109 b_12 NI_12 NS_109 0 5.9990566143326606e-06
GC_12_110 b_12 NI_12 NS_110 0 -1.1966985884043141e-06
GC_12_111 b_12 NI_12 NS_111 0 2.4514104334414259e-08
GC_12_112 b_12 NI_12 NS_112 0 6.7664913384540011e-10
GC_12_113 b_12 NI_12 NS_113 0 -8.0406027761895871e-11
GC_12_114 b_12 NI_12 NS_114 0 4.2875625146223765e-09
GC_12_115 b_12 NI_12 NS_115 0 -1.3622145998226382e-04
GC_12_116 b_12 NI_12 NS_116 0 1.9074668011898285e-04
GC_12_117 b_12 NI_12 NS_117 0 8.0921118582710989e-04
GC_12_118 b_12 NI_12 NS_118 0 2.1472038095280612e-04
GC_12_119 b_12 NI_12 NS_119 0 -5.3483055169574131e-04
GC_12_120 b_12 NI_12 NS_120 0 -8.9412917747181298e-04
GC_12_121 b_12 NI_12 NS_121 0 -1.5422765424595003e-10
GC_12_122 b_12 NI_12 NS_122 0 8.5210227168310199e-10
GC_12_123 b_12 NI_12 NS_123 0 1.8961601134564764e-09
GC_12_124 b_12 NI_12 NS_124 0 -4.9878803313819615e-09
GC_12_125 b_12 NI_12 NS_125 0 -1.0146836318618536e-09
GC_12_126 b_12 NI_12 NS_126 0 6.4015799221464667e-10
GC_12_127 b_12 NI_12 NS_127 0 -1.2655122938975591e-05
GC_12_128 b_12 NI_12 NS_128 0 4.1969203911094902e-05
GC_12_129 b_12 NI_12 NS_129 0 -1.5475050713847621e-08
GC_12_130 b_12 NI_12 NS_130 0 -6.5458898469368048e-10
GC_12_131 b_12 NI_12 NS_131 0 8.0669247534678500e-11
GC_12_132 b_12 NI_12 NS_132 0 -4.9744621424605511e-09
GC_12_133 b_12 NI_12 NS_133 0 1.1881342706323334e-04
GC_12_134 b_12 NI_12 NS_134 0 1.6345370675851010e-04
GC_12_135 b_12 NI_12 NS_135 0 3.0273232025576776e-04
GC_12_136 b_12 NI_12 NS_136 0 -5.3028074678107269e-04
GC_12_137 b_12 NI_12 NS_137 0 -4.0384999245408318e-04
GC_12_138 b_12 NI_12 NS_138 0 1.5542131564728288e-04
GC_12_139 b_12 NI_12 NS_139 0 -2.2896668868368914e-10
GC_12_140 b_12 NI_12 NS_140 0 -8.6252774463404982e-10
GC_12_141 b_12 NI_12 NS_141 0 -1.0664715499387909e-09
GC_12_142 b_12 NI_12 NS_142 0 3.8727144796673969e-09
GC_12_143 b_12 NI_12 NS_143 0 1.2870633136821934e-09
GC_12_144 b_12 NI_12 NS_144 0 -4.9787419256907865e-10
GC_12_145 b_12 NI_12 NS_145 0 1.1715003186506469e-04
GC_12_146 b_12 NI_12 NS_146 0 -4.6263178872032388e-04
GC_12_147 b_12 NI_12 NS_147 0 3.5653867287386937e-07
GC_12_148 b_12 NI_12 NS_148 0 3.4767107719523936e-09
GC_12_149 b_12 NI_12 NS_149 0 -1.1870437822590819e-11
GC_12_150 b_12 NI_12 NS_150 0 1.2107854262941925e-07
GC_12_151 b_12 NI_12 NS_151 0 7.0305739463262778e-04
GC_12_152 b_12 NI_12 NS_152 0 -4.2879088211702646e-03
GC_12_153 b_12 NI_12 NS_153 0 -9.0097307104426184e-03
GC_12_154 b_12 NI_12 NS_154 0 -5.1466471039655886e-03
GC_12_155 b_12 NI_12 NS_155 0 1.8363219559824795e-03
GC_12_156 b_12 NI_12 NS_156 0 7.2289144554878388e-03
GC_12_157 b_12 NI_12 NS_157 0 4.0590056914778968e-09
GC_12_158 b_12 NI_12 NS_158 0 2.5523055621577758e-09
GC_12_159 b_12 NI_12 NS_159 0 1.9338920384270956e-09
GC_12_160 b_12 NI_12 NS_160 0 1.2043039037528786e-08
GC_12_161 b_12 NI_12 NS_161 0 -2.5390686838875886e-08
GC_12_162 b_12 NI_12 NS_162 0 -1.4677114158259819e-08
GC_12_163 b_12 NI_12 NS_163 0 -6.0714589214531543e-04
GC_12_164 b_12 NI_12 NS_164 0 1.3759759195925850e-03
GC_12_165 b_12 NI_12 NS_165 0 -8.5772785963412286e-07
GC_12_166 b_12 NI_12 NS_166 0 -1.4280316037120561e-09
GC_12_167 b_12 NI_12 NS_167 0 -2.7382752147589900e-11
GC_12_168 b_12 NI_12 NS_168 0 -2.1435121146076394e-07
GC_12_169 b_12 NI_12 NS_169 0 -4.2079275805101419e-03
GC_12_170 b_12 NI_12 NS_170 0 1.9043905518495784e-02
GC_12_171 b_12 NI_12 NS_171 0 1.8778530753187726e-02
GC_12_172 b_12 NI_12 NS_172 0 -1.2050033188310090e-02
GC_12_173 b_12 NI_12 NS_173 0 2.1826900266355320e-03
GC_12_174 b_12 NI_12 NS_174 0 2.9283123940241910e-02
GC_12_175 b_12 NI_12 NS_175 0 -3.3741425227792627e-08
GC_12_176 b_12 NI_12 NS_176 0 -2.4547826509216362e-08
GC_12_177 b_12 NI_12 NS_177 0 8.1296563942339738e-08
GC_12_178 b_12 NI_12 NS_178 0 -4.2574365462842614e-08
GC_12_179 b_12 NI_12 NS_179 0 5.1566298769467681e-08
GC_12_180 b_12 NI_12 NS_180 0 3.1363508263516884e-08
GC_12_181 b_12 NI_12 NS_181 0 1.0851108981875789e-02
GC_12_182 b_12 NI_12 NS_182 0 -2.9613262495104469e-02
GC_12_183 b_12 NI_12 NS_183 0 -1.0888561530805789e-05
GC_12_184 b_12 NI_12 NS_184 0 -6.9605973491380587e-07
GC_12_185 b_12 NI_12 NS_185 0 1.2495406330252362e-08
GC_12_186 b_12 NI_12 NS_186 0 8.6530288767533445e-06
GC_12_187 b_12 NI_12 NS_187 0 -5.1292982245432536e-02
GC_12_188 b_12 NI_12 NS_188 0 6.8705434572019441e-02
GC_12_189 b_12 NI_12 NS_189 0 -2.8912508781474930e-02
GC_12_190 b_12 NI_12 NS_190 0 -1.5463846793044189e-01
GC_12_191 b_12 NI_12 NS_191 0 -4.9852937500885824e-03
GC_12_192 b_12 NI_12 NS_192 0 -1.6599316864634245e-01
GC_12_193 b_12 NI_12 NS_193 0 4.7917880819059967e-07
GC_12_194 b_12 NI_12 NS_194 0 8.9027560937444183e-07
GC_12_195 b_12 NI_12 NS_195 0 -4.3716899890095664e-06
GC_12_196 b_12 NI_12 NS_196 0 1.1070795194436870e-07
GC_12_197 b_12 NI_12 NS_197 0 -3.3754692040236320e-06
GC_12_198 b_12 NI_12 NS_198 0 -3.5753220432498962e-06
GC_12_199 b_12 NI_12 NS_199 0 -4.7894741477349399e-03
GC_12_200 b_12 NI_12 NS_200 0 1.6721231895481539e-02
GC_12_201 b_12 NI_12 NS_201 0 -3.5217425139558022e-06
GC_12_202 b_12 NI_12 NS_202 0 2.9869341330020878e-08
GC_12_203 b_12 NI_12 NS_203 0 -1.0050510000658381e-09
GC_12_204 b_12 NI_12 NS_204 0 -2.0070261998679719e-06
GC_12_205 b_12 NI_12 NS_205 0 1.8815079487248188e-02
GC_12_206 b_12 NI_12 NS_206 0 5.0642922456163572e-02
GC_12_207 b_12 NI_12 NS_207 0 1.5086435845919644e-02
GC_12_208 b_12 NI_12 NS_208 0 7.1442548787403443e-02
GC_12_209 b_12 NI_12 NS_209 0 8.1541997974382316e-02
GC_12_210 b_12 NI_12 NS_210 0 4.9085291802293936e-02
GC_12_211 b_12 NI_12 NS_211 0 -2.7438712865987003e-07
GC_12_212 b_12 NI_12 NS_212 0 -6.0490113086140492e-08
GC_12_213 b_12 NI_12 NS_213 0 5.2038320036656279e-07
GC_12_214 b_12 NI_12 NS_214 0 -7.4412561535754728e-07
GC_12_215 b_12 NI_12 NS_215 0 3.9436032396776982e-07
GC_12_216 b_12 NI_12 NS_216 0 3.8383217890957768e-07
GD_12_1 b_12 NI_12 NA_1 0 -1.5515985395771453e-05
GD_12_2 b_12 NI_12 NA_2 0 1.3353180228019851e-05
GD_12_3 b_12 NI_12 NA_3 0 -2.5606573167412140e-07
GD_12_4 b_12 NI_12 NA_4 0 9.8463604899017610e-06
GD_12_5 b_12 NI_12 NA_5 0 -2.7783437097327603e-05
GD_12_6 b_12 NI_12 NA_6 0 -4.9719335398735772e-05
GD_12_7 b_12 NI_12 NA_7 0 -4.3086478925310096e-05
GD_12_8 b_12 NI_12 NA_8 0 7.9753277994871176e-05
GD_12_9 b_12 NI_12 NA_9 0 3.7903418676586594e-03
GD_12_10 b_12 NI_12 NA_10 0 6.2327480091603320e-03
GD_12_11 b_12 NI_12 NA_11 0 7.4536168576468234e-02
GD_12_12 b_12 NI_12 NA_12 0 -9.3789089811108700e-02
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 8.5062695981493661e+00
GS_1_1 0 NS_1 NA_1 0 9.8455044987356888e-01
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 6.6124413087934162e+00
GS_2_1 0 NS_2 NA_1 0 9.8455044987356888e-01
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-13
RS_3 NS_3 0 5.0191788921294943e+01
GS_3_1 0 NS_3 NA_1 0 9.8455044987356888e-01
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-13
RS_4 NS_4 0 1.2665334842050991e+03
GS_4_1 0 NS_4 NA_1 0 9.8455044987356888e-01
*
* Real pole n. 5
CS_5 NS_5 0 9.9999999999999998e-13
RS_5 NS_5 0 1.4009873029214565e+04
GS_5_1 0 NS_5 NA_1 0 9.8455044987356888e-01
*
* Real pole n. 6
CS_6 NS_6 0 9.9999999999999998e-13
RS_6 NS_6 0 2.6077399387449515e+02
GS_6_1 0 NS_6 NA_1 0 9.8455044987356888e-01
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 5.1178878130294372e+00
RS_8 NS_8 0 5.1178878130294372e+00
GL_7 0 NS_7 NS_8 0 6.0508395241620216e-01
GL_8 0 NS_8 NS_7 0 -6.0508395241620216e-01
GS_7_1 0 NS_7 NA_1 0 9.8455044987356888e-01
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 3.7089246454198972e+00
RS_10 NS_10 0 3.7089246454198967e+00
GL_9 0 NS_9 NS_10 0 3.0956092481489988e-01
GL_10 0 NS_10 NS_9 0 -3.0956092481489988e-01
GS_9_1 0 NS_9 NA_1 0 9.8455044987356888e-01
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 3.7950611064409761e+00
RS_12 NS_12 0 3.7950611064409765e+00
GL_11 0 NS_11 NS_12 0 1.0768516390617248e-01
GL_12 0 NS_12 NS_11 0 -1.0768516390617248e-01
GS_11_1 0 NS_11 NA_1 0 9.8455044987356888e-01
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 2.7209036367703328e+02
RS_14 NS_14 0 2.7209036367703322e+02
GL_13 0 NS_13 NS_14 0 6.1072499247316107e-02
GL_14 0 NS_14 NS_13 0 -6.1072499247316107e-02
GS_13_1 0 NS_13 NA_1 0 9.8455044987356888e-01
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 1.1531527114161022e+02
RS_16 NS_16 0 1.1531527114161022e+02
GL_15 0 NS_15 NS_16 0 2.9421516884318294e-02
GL_16 0 NS_16 NS_15 0 -2.9421516884318294e-02
GS_15_1 0 NS_15 NA_1 0 9.8455044987356888e-01
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 6.1076117465889047e+02
RS_18 NS_18 0 6.1076117465889035e+02
GL_17 0 NS_17 NS_18 0 9.2445115841435419e-04
GL_18 0 NS_18 NS_17 0 -9.2445115841435419e-04
GS_17_1 0 NS_17 NA_1 0 9.8455044987356888e-01
*
* Real pole n. 19
CS_19 NS_19 0 9.9999999999999998e-13
RS_19 NS_19 0 8.5062695981493661e+00
GS_19_2 0 NS_19 NA_2 0 9.8455044987356888e-01
*
* Real pole n. 20
CS_20 NS_20 0 9.9999999999999998e-13
RS_20 NS_20 0 6.6124413087934162e+00
GS_20_2 0 NS_20 NA_2 0 9.8455044987356888e-01
*
* Real pole n. 21
CS_21 NS_21 0 9.9999999999999998e-13
RS_21 NS_21 0 5.0191788921294943e+01
GS_21_2 0 NS_21 NA_2 0 9.8455044987356888e-01
*
* Real pole n. 22
CS_22 NS_22 0 9.9999999999999998e-13
RS_22 NS_22 0 1.2665334842050991e+03
GS_22_2 0 NS_22 NA_2 0 9.8455044987356888e-01
*
* Real pole n. 23
CS_23 NS_23 0 9.9999999999999998e-13
RS_23 NS_23 0 1.4009873029214565e+04
GS_23_2 0 NS_23 NA_2 0 9.8455044987356888e-01
*
* Real pole n. 24
CS_24 NS_24 0 9.9999999999999998e-13
RS_24 NS_24 0 2.6077399387449515e+02
GS_24_2 0 NS_24 NA_2 0 9.8455044987356888e-01
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 5.1178878130294372e+00
RS_26 NS_26 0 5.1178878130294372e+00
GL_25 0 NS_25 NS_26 0 6.0508395241620216e-01
GL_26 0 NS_26 NS_25 0 -6.0508395241620216e-01
GS_25_2 0 NS_25 NA_2 0 9.8455044987356888e-01
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 3.7089246454198972e+00
RS_28 NS_28 0 3.7089246454198967e+00
GL_27 0 NS_27 NS_28 0 3.0956092481489988e-01
GL_28 0 NS_28 NS_27 0 -3.0956092481489988e-01
GS_27_2 0 NS_27 NA_2 0 9.8455044987356888e-01
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 3.7950611064409761e+00
RS_30 NS_30 0 3.7950611064409765e+00
GL_29 0 NS_29 NS_30 0 1.0768516390617248e-01
GL_30 0 NS_30 NS_29 0 -1.0768516390617248e-01
GS_29_2 0 NS_29 NA_2 0 9.8455044987356888e-01
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 2.7209036367703328e+02
RS_32 NS_32 0 2.7209036367703322e+02
GL_31 0 NS_31 NS_32 0 6.1072499247316107e-02
GL_32 0 NS_32 NS_31 0 -6.1072499247316107e-02
GS_31_2 0 NS_31 NA_2 0 9.8455044987356888e-01
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 1.1531527114161022e+02
RS_34 NS_34 0 1.1531527114161022e+02
GL_33 0 NS_33 NS_34 0 2.9421516884318294e-02
GL_34 0 NS_34 NS_33 0 -2.9421516884318294e-02
GS_33_2 0 NS_33 NA_2 0 9.8455044987356888e-01
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 6.1076117465889047e+02
RS_36 NS_36 0 6.1076117465889035e+02
GL_35 0 NS_35 NS_36 0 9.2445115841435419e-04
GL_36 0 NS_36 NS_35 0 -9.2445115841435419e-04
GS_35_2 0 NS_35 NA_2 0 9.8455044987356888e-01
*
* Real pole n. 37
CS_37 NS_37 0 9.9999999999999998e-13
RS_37 NS_37 0 8.5062695981493661e+00
GS_37_3 0 NS_37 NA_3 0 9.8455044987356888e-01
*
* Real pole n. 38
CS_38 NS_38 0 9.9999999999999998e-13
RS_38 NS_38 0 6.6124413087934162e+00
GS_38_3 0 NS_38 NA_3 0 9.8455044987356888e-01
*
* Real pole n. 39
CS_39 NS_39 0 9.9999999999999998e-13
RS_39 NS_39 0 5.0191788921294943e+01
GS_39_3 0 NS_39 NA_3 0 9.8455044987356888e-01
*
* Real pole n. 40
CS_40 NS_40 0 9.9999999999999998e-13
RS_40 NS_40 0 1.2665334842050991e+03
GS_40_3 0 NS_40 NA_3 0 9.8455044987356888e-01
*
* Real pole n. 41
CS_41 NS_41 0 9.9999999999999998e-13
RS_41 NS_41 0 1.4009873029214565e+04
GS_41_3 0 NS_41 NA_3 0 9.8455044987356888e-01
*
* Real pole n. 42
CS_42 NS_42 0 9.9999999999999998e-13
RS_42 NS_42 0 2.6077399387449515e+02
GS_42_3 0 NS_42 NA_3 0 9.8455044987356888e-01
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 5.1178878130294372e+00
RS_44 NS_44 0 5.1178878130294372e+00
GL_43 0 NS_43 NS_44 0 6.0508395241620216e-01
GL_44 0 NS_44 NS_43 0 -6.0508395241620216e-01
GS_43_3 0 NS_43 NA_3 0 9.8455044987356888e-01
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 3.7089246454198972e+00
RS_46 NS_46 0 3.7089246454198967e+00
GL_45 0 NS_45 NS_46 0 3.0956092481489988e-01
GL_46 0 NS_46 NS_45 0 -3.0956092481489988e-01
GS_45_3 0 NS_45 NA_3 0 9.8455044987356888e-01
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 3.7950611064409761e+00
RS_48 NS_48 0 3.7950611064409765e+00
GL_47 0 NS_47 NS_48 0 1.0768516390617248e-01
GL_48 0 NS_48 NS_47 0 -1.0768516390617248e-01
GS_47_3 0 NS_47 NA_3 0 9.8455044987356888e-01
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 2.7209036367703328e+02
RS_50 NS_50 0 2.7209036367703322e+02
GL_49 0 NS_49 NS_50 0 6.1072499247316107e-02
GL_50 0 NS_50 NS_49 0 -6.1072499247316107e-02
GS_49_3 0 NS_49 NA_3 0 9.8455044987356888e-01
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 1.1531527114161022e+02
RS_52 NS_52 0 1.1531527114161022e+02
GL_51 0 NS_51 NS_52 0 2.9421516884318294e-02
GL_52 0 NS_52 NS_51 0 -2.9421516884318294e-02
GS_51_3 0 NS_51 NA_3 0 9.8455044987356888e-01
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 6.1076117465889047e+02
RS_54 NS_54 0 6.1076117465889035e+02
GL_53 0 NS_53 NS_54 0 9.2445115841435419e-04
GL_54 0 NS_54 NS_53 0 -9.2445115841435419e-04
GS_53_3 0 NS_53 NA_3 0 9.8455044987356888e-01
*
* Real pole n. 55
CS_55 NS_55 0 9.9999999999999998e-13
RS_55 NS_55 0 8.5062695981493661e+00
GS_55_4 0 NS_55 NA_4 0 9.8455044987356888e-01
*
* Real pole n. 56
CS_56 NS_56 0 9.9999999999999998e-13
RS_56 NS_56 0 6.6124413087934162e+00
GS_56_4 0 NS_56 NA_4 0 9.8455044987356888e-01
*
* Real pole n. 57
CS_57 NS_57 0 9.9999999999999998e-13
RS_57 NS_57 0 5.0191788921294943e+01
GS_57_4 0 NS_57 NA_4 0 9.8455044987356888e-01
*
* Real pole n. 58
CS_58 NS_58 0 9.9999999999999998e-13
RS_58 NS_58 0 1.2665334842050991e+03
GS_58_4 0 NS_58 NA_4 0 9.8455044987356888e-01
*
* Real pole n. 59
CS_59 NS_59 0 9.9999999999999998e-13
RS_59 NS_59 0 1.4009873029214565e+04
GS_59_4 0 NS_59 NA_4 0 9.8455044987356888e-01
*
* Real pole n. 60
CS_60 NS_60 0 9.9999999999999998e-13
RS_60 NS_60 0 2.6077399387449515e+02
GS_60_4 0 NS_60 NA_4 0 9.8455044987356888e-01
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 5.1178878130294372e+00
RS_62 NS_62 0 5.1178878130294372e+00
GL_61 0 NS_61 NS_62 0 6.0508395241620216e-01
GL_62 0 NS_62 NS_61 0 -6.0508395241620216e-01
GS_61_4 0 NS_61 NA_4 0 9.8455044987356888e-01
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 3.7089246454198972e+00
RS_64 NS_64 0 3.7089246454198967e+00
GL_63 0 NS_63 NS_64 0 3.0956092481489988e-01
GL_64 0 NS_64 NS_63 0 -3.0956092481489988e-01
GS_63_4 0 NS_63 NA_4 0 9.8455044987356888e-01
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 3.7950611064409761e+00
RS_66 NS_66 0 3.7950611064409765e+00
GL_65 0 NS_65 NS_66 0 1.0768516390617248e-01
GL_66 0 NS_66 NS_65 0 -1.0768516390617248e-01
GS_65_4 0 NS_65 NA_4 0 9.8455044987356888e-01
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 2.7209036367703328e+02
RS_68 NS_68 0 2.7209036367703322e+02
GL_67 0 NS_67 NS_68 0 6.1072499247316107e-02
GL_68 0 NS_68 NS_67 0 -6.1072499247316107e-02
GS_67_4 0 NS_67 NA_4 0 9.8455044987356888e-01
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 1.1531527114161022e+02
RS_70 NS_70 0 1.1531527114161022e+02
GL_69 0 NS_69 NS_70 0 2.9421516884318294e-02
GL_70 0 NS_70 NS_69 0 -2.9421516884318294e-02
GS_69_4 0 NS_69 NA_4 0 9.8455044987356888e-01
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 6.1076117465889047e+02
RS_72 NS_72 0 6.1076117465889035e+02
GL_71 0 NS_71 NS_72 0 9.2445115841435419e-04
GL_72 0 NS_72 NS_71 0 -9.2445115841435419e-04
GS_71_4 0 NS_71 NA_4 0 9.8455044987356888e-01
*
* Real pole n. 73
CS_73 NS_73 0 9.9999999999999998e-13
RS_73 NS_73 0 8.5062695981493661e+00
GS_73_5 0 NS_73 NA_5 0 9.8455044987356888e-01
*
* Real pole n. 74
CS_74 NS_74 0 9.9999999999999998e-13
RS_74 NS_74 0 6.6124413087934162e+00
GS_74_5 0 NS_74 NA_5 0 9.8455044987356888e-01
*
* Real pole n. 75
CS_75 NS_75 0 9.9999999999999998e-13
RS_75 NS_75 0 5.0191788921294943e+01
GS_75_5 0 NS_75 NA_5 0 9.8455044987356888e-01
*
* Real pole n. 76
CS_76 NS_76 0 9.9999999999999998e-13
RS_76 NS_76 0 1.2665334842050991e+03
GS_76_5 0 NS_76 NA_5 0 9.8455044987356888e-01
*
* Real pole n. 77
CS_77 NS_77 0 9.9999999999999998e-13
RS_77 NS_77 0 1.4009873029214565e+04
GS_77_5 0 NS_77 NA_5 0 9.8455044987356888e-01
*
* Real pole n. 78
CS_78 NS_78 0 9.9999999999999998e-13
RS_78 NS_78 0 2.6077399387449515e+02
GS_78_5 0 NS_78 NA_5 0 9.8455044987356888e-01
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 5.1178878130294372e+00
RS_80 NS_80 0 5.1178878130294372e+00
GL_79 0 NS_79 NS_80 0 6.0508395241620216e-01
GL_80 0 NS_80 NS_79 0 -6.0508395241620216e-01
GS_79_5 0 NS_79 NA_5 0 9.8455044987356888e-01
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 3.7089246454198972e+00
RS_82 NS_82 0 3.7089246454198967e+00
GL_81 0 NS_81 NS_82 0 3.0956092481489988e-01
GL_82 0 NS_82 NS_81 0 -3.0956092481489988e-01
GS_81_5 0 NS_81 NA_5 0 9.8455044987356888e-01
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 3.7950611064409761e+00
RS_84 NS_84 0 3.7950611064409765e+00
GL_83 0 NS_83 NS_84 0 1.0768516390617248e-01
GL_84 0 NS_84 NS_83 0 -1.0768516390617248e-01
GS_83_5 0 NS_83 NA_5 0 9.8455044987356888e-01
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 2.7209036367703328e+02
RS_86 NS_86 0 2.7209036367703322e+02
GL_85 0 NS_85 NS_86 0 6.1072499247316107e-02
GL_86 0 NS_86 NS_85 0 -6.1072499247316107e-02
GS_85_5 0 NS_85 NA_5 0 9.8455044987356888e-01
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 1.1531527114161022e+02
RS_88 NS_88 0 1.1531527114161022e+02
GL_87 0 NS_87 NS_88 0 2.9421516884318294e-02
GL_88 0 NS_88 NS_87 0 -2.9421516884318294e-02
GS_87_5 0 NS_87 NA_5 0 9.8455044987356888e-01
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 6.1076117465889047e+02
RS_90 NS_90 0 6.1076117465889035e+02
GL_89 0 NS_89 NS_90 0 9.2445115841435419e-04
GL_90 0 NS_90 NS_89 0 -9.2445115841435419e-04
GS_89_5 0 NS_89 NA_5 0 9.8455044987356888e-01
*
* Real pole n. 91
CS_91 NS_91 0 9.9999999999999998e-13
RS_91 NS_91 0 8.5062695981493661e+00
GS_91_6 0 NS_91 NA_6 0 9.8455044987356888e-01
*
* Real pole n. 92
CS_92 NS_92 0 9.9999999999999998e-13
RS_92 NS_92 0 6.6124413087934162e+00
GS_92_6 0 NS_92 NA_6 0 9.8455044987356888e-01
*
* Real pole n. 93
CS_93 NS_93 0 9.9999999999999998e-13
RS_93 NS_93 0 5.0191788921294943e+01
GS_93_6 0 NS_93 NA_6 0 9.8455044987356888e-01
*
* Real pole n. 94
CS_94 NS_94 0 9.9999999999999998e-13
RS_94 NS_94 0 1.2665334842050991e+03
GS_94_6 0 NS_94 NA_6 0 9.8455044987356888e-01
*
* Real pole n. 95
CS_95 NS_95 0 9.9999999999999998e-13
RS_95 NS_95 0 1.4009873029214565e+04
GS_95_6 0 NS_95 NA_6 0 9.8455044987356888e-01
*
* Real pole n. 96
CS_96 NS_96 0 9.9999999999999998e-13
RS_96 NS_96 0 2.6077399387449515e+02
GS_96_6 0 NS_96 NA_6 0 9.8455044987356888e-01
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 5.1178878130294372e+00
RS_98 NS_98 0 5.1178878130294372e+00
GL_97 0 NS_97 NS_98 0 6.0508395241620216e-01
GL_98 0 NS_98 NS_97 0 -6.0508395241620216e-01
GS_97_6 0 NS_97 NA_6 0 9.8455044987356888e-01
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 3.7089246454198972e+00
RS_100 NS_100 0 3.7089246454198967e+00
GL_99 0 NS_99 NS_100 0 3.0956092481489988e-01
GL_100 0 NS_100 NS_99 0 -3.0956092481489988e-01
GS_99_6 0 NS_99 NA_6 0 9.8455044987356888e-01
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 3.7950611064409761e+00
RS_102 NS_102 0 3.7950611064409765e+00
GL_101 0 NS_101 NS_102 0 1.0768516390617248e-01
GL_102 0 NS_102 NS_101 0 -1.0768516390617248e-01
GS_101_6 0 NS_101 NA_6 0 9.8455044987356888e-01
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 2.7209036367703328e+02
RS_104 NS_104 0 2.7209036367703322e+02
GL_103 0 NS_103 NS_104 0 6.1072499247316107e-02
GL_104 0 NS_104 NS_103 0 -6.1072499247316107e-02
GS_103_6 0 NS_103 NA_6 0 9.8455044987356888e-01
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 1.1531527114161022e+02
RS_106 NS_106 0 1.1531527114161022e+02
GL_105 0 NS_105 NS_106 0 2.9421516884318294e-02
GL_106 0 NS_106 NS_105 0 -2.9421516884318294e-02
GS_105_6 0 NS_105 NA_6 0 9.8455044987356888e-01
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 6.1076117465889047e+02
RS_108 NS_108 0 6.1076117465889035e+02
GL_107 0 NS_107 NS_108 0 9.2445115841435419e-04
GL_108 0 NS_108 NS_107 0 -9.2445115841435419e-04
GS_107_6 0 NS_107 NA_6 0 9.8455044987356888e-01
*
* Real pole n. 109
CS_109 NS_109 0 9.9999999999999998e-13
RS_109 NS_109 0 8.5062695981493661e+00
GS_109_7 0 NS_109 NA_7 0 9.8455044987356888e-01
*
* Real pole n. 110
CS_110 NS_110 0 9.9999999999999998e-13
RS_110 NS_110 0 6.6124413087934162e+00
GS_110_7 0 NS_110 NA_7 0 9.8455044987356888e-01
*
* Real pole n. 111
CS_111 NS_111 0 9.9999999999999998e-13
RS_111 NS_111 0 5.0191788921294943e+01
GS_111_7 0 NS_111 NA_7 0 9.8455044987356888e-01
*
* Real pole n. 112
CS_112 NS_112 0 9.9999999999999998e-13
RS_112 NS_112 0 1.2665334842050991e+03
GS_112_7 0 NS_112 NA_7 0 9.8455044987356888e-01
*
* Real pole n. 113
CS_113 NS_113 0 9.9999999999999998e-13
RS_113 NS_113 0 1.4009873029214565e+04
GS_113_7 0 NS_113 NA_7 0 9.8455044987356888e-01
*
* Real pole n. 114
CS_114 NS_114 0 9.9999999999999998e-13
RS_114 NS_114 0 2.6077399387449515e+02
GS_114_7 0 NS_114 NA_7 0 9.8455044987356888e-01
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 5.1178878130294372e+00
RS_116 NS_116 0 5.1178878130294372e+00
GL_115 0 NS_115 NS_116 0 6.0508395241620216e-01
GL_116 0 NS_116 NS_115 0 -6.0508395241620216e-01
GS_115_7 0 NS_115 NA_7 0 9.8455044987356888e-01
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 3.7089246454198972e+00
RS_118 NS_118 0 3.7089246454198967e+00
GL_117 0 NS_117 NS_118 0 3.0956092481489988e-01
GL_118 0 NS_118 NS_117 0 -3.0956092481489988e-01
GS_117_7 0 NS_117 NA_7 0 9.8455044987356888e-01
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 3.7950611064409761e+00
RS_120 NS_120 0 3.7950611064409765e+00
GL_119 0 NS_119 NS_120 0 1.0768516390617248e-01
GL_120 0 NS_120 NS_119 0 -1.0768516390617248e-01
GS_119_7 0 NS_119 NA_7 0 9.8455044987356888e-01
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 2.7209036367703328e+02
RS_122 NS_122 0 2.7209036367703322e+02
GL_121 0 NS_121 NS_122 0 6.1072499247316107e-02
GL_122 0 NS_122 NS_121 0 -6.1072499247316107e-02
GS_121_7 0 NS_121 NA_7 0 9.8455044987356888e-01
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 1.1531527114161022e+02
RS_124 NS_124 0 1.1531527114161022e+02
GL_123 0 NS_123 NS_124 0 2.9421516884318294e-02
GL_124 0 NS_124 NS_123 0 -2.9421516884318294e-02
GS_123_7 0 NS_123 NA_7 0 9.8455044987356888e-01
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 6.1076117465889047e+02
RS_126 NS_126 0 6.1076117465889035e+02
GL_125 0 NS_125 NS_126 0 9.2445115841435419e-04
GL_126 0 NS_126 NS_125 0 -9.2445115841435419e-04
GS_125_7 0 NS_125 NA_7 0 9.8455044987356888e-01
*
* Real pole n. 127
CS_127 NS_127 0 9.9999999999999998e-13
RS_127 NS_127 0 8.5062695981493661e+00
GS_127_8 0 NS_127 NA_8 0 9.8455044987356888e-01
*
* Real pole n. 128
CS_128 NS_128 0 9.9999999999999998e-13
RS_128 NS_128 0 6.6124413087934162e+00
GS_128_8 0 NS_128 NA_8 0 9.8455044987356888e-01
*
* Real pole n. 129
CS_129 NS_129 0 9.9999999999999998e-13
RS_129 NS_129 0 5.0191788921294943e+01
GS_129_8 0 NS_129 NA_8 0 9.8455044987356888e-01
*
* Real pole n. 130
CS_130 NS_130 0 9.9999999999999998e-13
RS_130 NS_130 0 1.2665334842050991e+03
GS_130_8 0 NS_130 NA_8 0 9.8455044987356888e-01
*
* Real pole n. 131
CS_131 NS_131 0 9.9999999999999998e-13
RS_131 NS_131 0 1.4009873029214565e+04
GS_131_8 0 NS_131 NA_8 0 9.8455044987356888e-01
*
* Real pole n. 132
CS_132 NS_132 0 9.9999999999999998e-13
RS_132 NS_132 0 2.6077399387449515e+02
GS_132_8 0 NS_132 NA_8 0 9.8455044987356888e-01
*
* Complex pair n. 133/134
CS_133 NS_133 0 9.9999999999999998e-13
CS_134 NS_134 0 9.9999999999999998e-13
RS_133 NS_133 0 5.1178878130294372e+00
RS_134 NS_134 0 5.1178878130294372e+00
GL_133 0 NS_133 NS_134 0 6.0508395241620216e-01
GL_134 0 NS_134 NS_133 0 -6.0508395241620216e-01
GS_133_8 0 NS_133 NA_8 0 9.8455044987356888e-01
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 3.7089246454198972e+00
RS_136 NS_136 0 3.7089246454198967e+00
GL_135 0 NS_135 NS_136 0 3.0956092481489988e-01
GL_136 0 NS_136 NS_135 0 -3.0956092481489988e-01
GS_135_8 0 NS_135 NA_8 0 9.8455044987356888e-01
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 3.7950611064409761e+00
RS_138 NS_138 0 3.7950611064409765e+00
GL_137 0 NS_137 NS_138 0 1.0768516390617248e-01
GL_138 0 NS_138 NS_137 0 -1.0768516390617248e-01
GS_137_8 0 NS_137 NA_8 0 9.8455044987356888e-01
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 2.7209036367703328e+02
RS_140 NS_140 0 2.7209036367703322e+02
GL_139 0 NS_139 NS_140 0 6.1072499247316107e-02
GL_140 0 NS_140 NS_139 0 -6.1072499247316107e-02
GS_139_8 0 NS_139 NA_8 0 9.8455044987356888e-01
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 1.1531527114161022e+02
RS_142 NS_142 0 1.1531527114161022e+02
GL_141 0 NS_141 NS_142 0 2.9421516884318294e-02
GL_142 0 NS_142 NS_141 0 -2.9421516884318294e-02
GS_141_8 0 NS_141 NA_8 0 9.8455044987356888e-01
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 6.1076117465889047e+02
RS_144 NS_144 0 6.1076117465889035e+02
GL_143 0 NS_143 NS_144 0 9.2445115841435419e-04
GL_144 0 NS_144 NS_143 0 -9.2445115841435419e-04
GS_143_8 0 NS_143 NA_8 0 9.8455044987356888e-01
*
* Real pole n. 145
CS_145 NS_145 0 9.9999999999999998e-13
RS_145 NS_145 0 8.5062695981493661e+00
GS_145_9 0 NS_145 NA_9 0 9.8455044987356888e-01
*
* Real pole n. 146
CS_146 NS_146 0 9.9999999999999998e-13
RS_146 NS_146 0 6.6124413087934162e+00
GS_146_9 0 NS_146 NA_9 0 9.8455044987356888e-01
*
* Real pole n. 147
CS_147 NS_147 0 9.9999999999999998e-13
RS_147 NS_147 0 5.0191788921294943e+01
GS_147_9 0 NS_147 NA_9 0 9.8455044987356888e-01
*
* Real pole n. 148
CS_148 NS_148 0 9.9999999999999998e-13
RS_148 NS_148 0 1.2665334842050991e+03
GS_148_9 0 NS_148 NA_9 0 9.8455044987356888e-01
*
* Real pole n. 149
CS_149 NS_149 0 9.9999999999999998e-13
RS_149 NS_149 0 1.4009873029214565e+04
GS_149_9 0 NS_149 NA_9 0 9.8455044987356888e-01
*
* Real pole n. 150
CS_150 NS_150 0 9.9999999999999998e-13
RS_150 NS_150 0 2.6077399387449515e+02
GS_150_9 0 NS_150 NA_9 0 9.8455044987356888e-01
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 5.1178878130294372e+00
RS_152 NS_152 0 5.1178878130294372e+00
GL_151 0 NS_151 NS_152 0 6.0508395241620216e-01
GL_152 0 NS_152 NS_151 0 -6.0508395241620216e-01
GS_151_9 0 NS_151 NA_9 0 9.8455044987356888e-01
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 3.7089246454198972e+00
RS_154 NS_154 0 3.7089246454198967e+00
GL_153 0 NS_153 NS_154 0 3.0956092481489988e-01
GL_154 0 NS_154 NS_153 0 -3.0956092481489988e-01
GS_153_9 0 NS_153 NA_9 0 9.8455044987356888e-01
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 3.7950611064409761e+00
RS_156 NS_156 0 3.7950611064409765e+00
GL_155 0 NS_155 NS_156 0 1.0768516390617248e-01
GL_156 0 NS_156 NS_155 0 -1.0768516390617248e-01
GS_155_9 0 NS_155 NA_9 0 9.8455044987356888e-01
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 2.7209036367703328e+02
RS_158 NS_158 0 2.7209036367703322e+02
GL_157 0 NS_157 NS_158 0 6.1072499247316107e-02
GL_158 0 NS_158 NS_157 0 -6.1072499247316107e-02
GS_157_9 0 NS_157 NA_9 0 9.8455044987356888e-01
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 1.1531527114161022e+02
RS_160 NS_160 0 1.1531527114161022e+02
GL_159 0 NS_159 NS_160 0 2.9421516884318294e-02
GL_160 0 NS_160 NS_159 0 -2.9421516884318294e-02
GS_159_9 0 NS_159 NA_9 0 9.8455044987356888e-01
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 6.1076117465889047e+02
RS_162 NS_162 0 6.1076117465889035e+02
GL_161 0 NS_161 NS_162 0 9.2445115841435419e-04
GL_162 0 NS_162 NS_161 0 -9.2445115841435419e-04
GS_161_9 0 NS_161 NA_9 0 9.8455044987356888e-01
*
* Real pole n. 163
CS_163 NS_163 0 9.9999999999999998e-13
RS_163 NS_163 0 8.5062695981493661e+00
GS_163_10 0 NS_163 NA_10 0 9.8455044987356888e-01
*
* Real pole n. 164
CS_164 NS_164 0 9.9999999999999998e-13
RS_164 NS_164 0 6.6124413087934162e+00
GS_164_10 0 NS_164 NA_10 0 9.8455044987356888e-01
*
* Real pole n. 165
CS_165 NS_165 0 9.9999999999999998e-13
RS_165 NS_165 0 5.0191788921294943e+01
GS_165_10 0 NS_165 NA_10 0 9.8455044987356888e-01
*
* Real pole n. 166
CS_166 NS_166 0 9.9999999999999998e-13
RS_166 NS_166 0 1.2665334842050991e+03
GS_166_10 0 NS_166 NA_10 0 9.8455044987356888e-01
*
* Real pole n. 167
CS_167 NS_167 0 9.9999999999999998e-13
RS_167 NS_167 0 1.4009873029214565e+04
GS_167_10 0 NS_167 NA_10 0 9.8455044987356888e-01
*
* Real pole n. 168
CS_168 NS_168 0 9.9999999999999998e-13
RS_168 NS_168 0 2.6077399387449515e+02
GS_168_10 0 NS_168 NA_10 0 9.8455044987356888e-01
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 5.1178878130294372e+00
RS_170 NS_170 0 5.1178878130294372e+00
GL_169 0 NS_169 NS_170 0 6.0508395241620216e-01
GL_170 0 NS_170 NS_169 0 -6.0508395241620216e-01
GS_169_10 0 NS_169 NA_10 0 9.8455044987356888e-01
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 3.7089246454198972e+00
RS_172 NS_172 0 3.7089246454198967e+00
GL_171 0 NS_171 NS_172 0 3.0956092481489988e-01
GL_172 0 NS_172 NS_171 0 -3.0956092481489988e-01
GS_171_10 0 NS_171 NA_10 0 9.8455044987356888e-01
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 3.7950611064409761e+00
RS_174 NS_174 0 3.7950611064409765e+00
GL_173 0 NS_173 NS_174 0 1.0768516390617248e-01
GL_174 0 NS_174 NS_173 0 -1.0768516390617248e-01
GS_173_10 0 NS_173 NA_10 0 9.8455044987356888e-01
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 2.7209036367703328e+02
RS_176 NS_176 0 2.7209036367703322e+02
GL_175 0 NS_175 NS_176 0 6.1072499247316107e-02
GL_176 0 NS_176 NS_175 0 -6.1072499247316107e-02
GS_175_10 0 NS_175 NA_10 0 9.8455044987356888e-01
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 1.1531527114161022e+02
RS_178 NS_178 0 1.1531527114161022e+02
GL_177 0 NS_177 NS_178 0 2.9421516884318294e-02
GL_178 0 NS_178 NS_177 0 -2.9421516884318294e-02
GS_177_10 0 NS_177 NA_10 0 9.8455044987356888e-01
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 6.1076117465889047e+02
RS_180 NS_180 0 6.1076117465889035e+02
GL_179 0 NS_179 NS_180 0 9.2445115841435419e-04
GL_180 0 NS_180 NS_179 0 -9.2445115841435419e-04
GS_179_10 0 NS_179 NA_10 0 9.8455044987356888e-01
*
* Real pole n. 181
CS_181 NS_181 0 9.9999999999999998e-13
RS_181 NS_181 0 8.5062695981493661e+00
GS_181_11 0 NS_181 NA_11 0 9.8455044987356888e-01
*
* Real pole n. 182
CS_182 NS_182 0 9.9999999999999998e-13
RS_182 NS_182 0 6.6124413087934162e+00
GS_182_11 0 NS_182 NA_11 0 9.8455044987356888e-01
*
* Real pole n. 183
CS_183 NS_183 0 9.9999999999999998e-13
RS_183 NS_183 0 5.0191788921294943e+01
GS_183_11 0 NS_183 NA_11 0 9.8455044987356888e-01
*
* Real pole n. 184
CS_184 NS_184 0 9.9999999999999998e-13
RS_184 NS_184 0 1.2665334842050991e+03
GS_184_11 0 NS_184 NA_11 0 9.8455044987356888e-01
*
* Real pole n. 185
CS_185 NS_185 0 9.9999999999999998e-13
RS_185 NS_185 0 1.4009873029214565e+04
GS_185_11 0 NS_185 NA_11 0 9.8455044987356888e-01
*
* Real pole n. 186
CS_186 NS_186 0 9.9999999999999998e-13
RS_186 NS_186 0 2.6077399387449515e+02
GS_186_11 0 NS_186 NA_11 0 9.8455044987356888e-01
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 5.1178878130294372e+00
RS_188 NS_188 0 5.1178878130294372e+00
GL_187 0 NS_187 NS_188 0 6.0508395241620216e-01
GL_188 0 NS_188 NS_187 0 -6.0508395241620216e-01
GS_187_11 0 NS_187 NA_11 0 9.8455044987356888e-01
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 3.7089246454198972e+00
RS_190 NS_190 0 3.7089246454198967e+00
GL_189 0 NS_189 NS_190 0 3.0956092481489988e-01
GL_190 0 NS_190 NS_189 0 -3.0956092481489988e-01
GS_189_11 0 NS_189 NA_11 0 9.8455044987356888e-01
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 3.7950611064409761e+00
RS_192 NS_192 0 3.7950611064409765e+00
GL_191 0 NS_191 NS_192 0 1.0768516390617248e-01
GL_192 0 NS_192 NS_191 0 -1.0768516390617248e-01
GS_191_11 0 NS_191 NA_11 0 9.8455044987356888e-01
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 2.7209036367703328e+02
RS_194 NS_194 0 2.7209036367703322e+02
GL_193 0 NS_193 NS_194 0 6.1072499247316107e-02
GL_194 0 NS_194 NS_193 0 -6.1072499247316107e-02
GS_193_11 0 NS_193 NA_11 0 9.8455044987356888e-01
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 1.1531527114161022e+02
RS_196 NS_196 0 1.1531527114161022e+02
GL_195 0 NS_195 NS_196 0 2.9421516884318294e-02
GL_196 0 NS_196 NS_195 0 -2.9421516884318294e-02
GS_195_11 0 NS_195 NA_11 0 9.8455044987356888e-01
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 6.1076117465889047e+02
RS_198 NS_198 0 6.1076117465889035e+02
GL_197 0 NS_197 NS_198 0 9.2445115841435419e-04
GL_198 0 NS_198 NS_197 0 -9.2445115841435419e-04
GS_197_11 0 NS_197 NA_11 0 9.8455044987356888e-01
*
* Real pole n. 199
CS_199 NS_199 0 9.9999999999999998e-13
RS_199 NS_199 0 8.5062695981493661e+00
GS_199_12 0 NS_199 NA_12 0 9.8455044987356888e-01
*
* Real pole n. 200
CS_200 NS_200 0 9.9999999999999998e-13
RS_200 NS_200 0 6.6124413087934162e+00
GS_200_12 0 NS_200 NA_12 0 9.8455044987356888e-01
*
* Real pole n. 201
CS_201 NS_201 0 9.9999999999999998e-13
RS_201 NS_201 0 5.0191788921294943e+01
GS_201_12 0 NS_201 NA_12 0 9.8455044987356888e-01
*
* Real pole n. 202
CS_202 NS_202 0 9.9999999999999998e-13
RS_202 NS_202 0 1.2665334842050991e+03
GS_202_12 0 NS_202 NA_12 0 9.8455044987356888e-01
*
* Real pole n. 203
CS_203 NS_203 0 9.9999999999999998e-13
RS_203 NS_203 0 1.4009873029214565e+04
GS_203_12 0 NS_203 NA_12 0 9.8455044987356888e-01
*
* Real pole n. 204
CS_204 NS_204 0 9.9999999999999998e-13
RS_204 NS_204 0 2.6077399387449515e+02
GS_204_12 0 NS_204 NA_12 0 9.8455044987356888e-01
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 5.1178878130294372e+00
RS_206 NS_206 0 5.1178878130294372e+00
GL_205 0 NS_205 NS_206 0 6.0508395241620216e-01
GL_206 0 NS_206 NS_205 0 -6.0508395241620216e-01
GS_205_12 0 NS_205 NA_12 0 9.8455044987356888e-01
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 3.7089246454198972e+00
RS_208 NS_208 0 3.7089246454198967e+00
GL_207 0 NS_207 NS_208 0 3.0956092481489988e-01
GL_208 0 NS_208 NS_207 0 -3.0956092481489988e-01
GS_207_12 0 NS_207 NA_12 0 9.8455044987356888e-01
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 3.7950611064409761e+00
RS_210 NS_210 0 3.7950611064409765e+00
GL_209 0 NS_209 NS_210 0 1.0768516390617248e-01
GL_210 0 NS_210 NS_209 0 -1.0768516390617248e-01
GS_209_12 0 NS_209 NA_12 0 9.8455044987356888e-01
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 2.7209036367703328e+02
RS_212 NS_212 0 2.7209036367703322e+02
GL_211 0 NS_211 NS_212 0 6.1072499247316107e-02
GL_212 0 NS_212 NS_211 0 -6.1072499247316107e-02
GS_211_12 0 NS_211 NA_12 0 9.8455044987356888e-01
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 1.1531527114161022e+02
RS_214 NS_214 0 1.1531527114161022e+02
GL_213 0 NS_213 NS_214 0 2.9421516884318294e-02
GL_214 0 NS_214 NS_213 0 -2.9421516884318294e-02
GS_213_12 0 NS_213 NA_12 0 9.8455044987356888e-01
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 6.1076117465889047e+02
RS_216 NS_216 0 6.1076117465889035e+02
GL_215 0 NS_215 NS_216 0 9.2445115841435419e-04
GL_216 0 NS_216 NS_215 0 -9.2445115841435419e-04
GS_215_12 0 NS_215 NA_12 0 9.8455044987356888e-01
*
******************************


.ends
*******************
* End of subcircuit
*******************
