**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [6 4 36] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_6_LGA
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 6.3409394050007090e-02
GC_1_2 b_1 NI_1 NS_2 0 -1.2379524327476145e-03
GC_1_3 b_1 NI_1 NS_3 0 4.6073378398346465e-02
GC_1_4 b_1 NI_1 NS_4 0 -5.0065076530390717e-02
GC_1_5 b_1 NI_1 NS_5 0 -2.9926551457762534e-03
GC_1_6 b_1 NI_1 NS_6 0 -1.8501879444927753e-03
GC_1_7 b_1 NI_1 NS_7 0 -4.0119655192179986e-04
GC_1_8 b_1 NI_1 NS_8 0 -1.2256490973020472e-05
GC_1_9 b_1 NI_1 NS_9 0 -1.2531312099263711e-02
GC_1_10 b_1 NI_1 NS_10 0 1.6865019365300767e-02
GC_1_11 b_1 NI_1 NS_11 0 -7.4538663120960293e-05
GC_1_12 b_1 NI_1 NS_12 0 -9.6345032008630799e-05
GC_1_13 b_1 NI_1 NS_13 0 -3.9674262974394012e-02
GC_1_14 b_1 NI_1 NS_14 0 -7.0594357554221762e-04
GC_1_15 b_1 NI_1 NS_15 0 -4.5249135453259130e-05
GC_1_16 b_1 NI_1 NS_16 0 -3.6856301740939378e-05
GC_1_17 b_1 NI_1 NS_17 0 -5.7965869313555383e-05
GC_1_18 b_1 NI_1 NS_18 0 -2.4216504921878857e-05
GC_1_19 b_1 NI_1 NS_19 0 -5.8473332391373344e-05
GC_1_20 b_1 NI_1 NS_20 0 4.1298008549675723e-06
GC_1_21 b_1 NI_1 NS_21 0 -4.1026641164075056e-05
GC_1_22 b_1 NI_1 NS_22 0 -2.9404242648457732e-05
GC_1_23 b_1 NI_1 NS_23 0 -7.3052264697329727e-03
GC_1_24 b_1 NI_1 NS_24 0 1.0271366626290341e-02
GC_1_25 b_1 NI_1 NS_25 0 -3.6739400340659445e-04
GC_1_26 b_1 NI_1 NS_26 0 -1.1862329580617369e-03
GC_1_27 b_1 NI_1 NS_27 0 1.6159917242791061e-04
GC_1_28 b_1 NI_1 NS_28 0 -1.1332102644453174e-03
GC_1_29 b_1 NI_1 NS_29 0 9.0710692897574309e-05
GC_1_30 b_1 NI_1 NS_30 0 3.0720445250427176e-05
GC_1_31 b_1 NI_1 NS_31 0 1.6338475847260477e-04
GC_1_32 b_1 NI_1 NS_32 0 -8.6688481201208445e-05
GC_1_33 b_1 NI_1 NS_33 0 4.4769602124791053e-06
GC_1_34 b_1 NI_1 NS_34 0 -1.0966912483294991e-04
GC_1_35 b_1 NI_1 NS_35 0 5.9570127056589263e-05
GC_1_36 b_1 NI_1 NS_36 0 1.2301645595262591e-05
GC_1_37 b_1 NI_1 NS_37 0 -1.6823342962559893e-05
GC_1_38 b_1 NI_1 NS_38 0 1.1009882901711967e-05
GC_1_39 b_1 NI_1 NS_39 0 1.0650907369936303e-02
GC_1_40 b_1 NI_1 NS_40 0 1.8827176324940039e-03
GC_1_41 b_1 NI_1 NS_41 0 2.3026429658907610e-02
GC_1_42 b_1 NI_1 NS_42 0 -4.8878704631495889e-03
GC_1_43 b_1 NI_1 NS_43 0 1.5236725319327622e-03
GC_1_44 b_1 NI_1 NS_44 0 -3.7328947839356246e-04
GC_1_45 b_1 NI_1 NS_45 0 1.5101632490463804e-04
GC_1_46 b_1 NI_1 NS_46 0 -8.9723266115792266e-05
GC_1_47 b_1 NI_1 NS_47 0 2.8807388984512936e-02
GC_1_48 b_1 NI_1 NS_48 0 6.2177155832794434e-03
GC_1_49 b_1 NI_1 NS_49 0 8.4526510529554514e-05
GC_1_50 b_1 NI_1 NS_50 0 9.8787536491944268e-05
GC_1_51 b_1 NI_1 NS_51 0 -3.7001712283476651e-02
GC_1_52 b_1 NI_1 NS_52 0 2.4514955521278782e-02
GC_1_53 b_1 NI_1 NS_53 0 2.0118713930660446e-05
GC_1_54 b_1 NI_1 NS_54 0 -1.9169926178054439e-05
GC_1_55 b_1 NI_1 NS_55 0 -2.1327609641753493e-05
GC_1_56 b_1 NI_1 NS_56 0 2.3716206545073458e-05
GC_1_57 b_1 NI_1 NS_57 0 3.4203801545744422e-06
GC_1_58 b_1 NI_1 NS_58 0 -4.2893814670879836e-06
GC_1_59 b_1 NI_1 NS_59 0 -8.0155204785734154e-05
GC_1_60 b_1 NI_1 NS_60 0 -3.1763228423879869e-05
GC_1_61 b_1 NI_1 NS_61 0 -4.8797181912797853e-03
GC_1_62 b_1 NI_1 NS_62 0 5.0548261556877276e-03
GC_1_63 b_1 NI_1 NS_63 0 -1.3089892711484965e-05
GC_1_64 b_1 NI_1 NS_64 0 -1.0262745314332819e-03
GC_1_65 b_1 NI_1 NS_65 0 8.3613929690514230e-05
GC_1_66 b_1 NI_1 NS_66 0 -7.1118247421535772e-04
GC_1_67 b_1 NI_1 NS_67 0 8.3565504555772302e-05
GC_1_68 b_1 NI_1 NS_68 0 9.2884968394408188e-05
GC_1_69 b_1 NI_1 NS_69 0 1.7747120583700733e-04
GC_1_70 b_1 NI_1 NS_70 0 5.4669582647738854e-05
GC_1_71 b_1 NI_1 NS_71 0 8.8939812219624901e-05
GC_1_72 b_1 NI_1 NS_72 0 -1.7282694505556612e-05
GC_1_73 b_1 NI_1 NS_73 0 1.6069616271231483e-05
GC_1_74 b_1 NI_1 NS_74 0 1.0946235620283329e-04
GC_1_75 b_1 NI_1 NS_75 0 3.2579973535145607e-05
GC_1_76 b_1 NI_1 NS_76 0 3.8085187297403361e-07
GC_1_77 b_1 NI_1 NS_77 0 -1.0704833817444821e-02
GC_1_78 b_1 NI_1 NS_78 0 -1.2959578050847700e-03
GC_1_79 b_1 NI_1 NS_79 0 7.4730685754213037e-03
GC_1_80 b_1 NI_1 NS_80 0 2.6999598521385577e-02
GC_1_81 b_1 NI_1 NS_81 0 -6.6139802310007166e-04
GC_1_82 b_1 NI_1 NS_82 0 8.1781311449083307e-04
GC_1_83 b_1 NI_1 NS_83 0 -1.4920222909183846e-04
GC_1_84 b_1 NI_1 NS_84 0 2.1318936273700449e-04
GC_1_85 b_1 NI_1 NS_85 0 1.1678198801964796e-02
GC_1_86 b_1 NI_1 NS_86 0 2.6150106747549279e-02
GC_1_87 b_1 NI_1 NS_87 0 -8.0788403086348411e-05
GC_1_88 b_1 NI_1 NS_88 0 -9.4560221926931736e-05
GC_1_89 b_1 NI_1 NS_89 0 2.5073251329049893e-02
GC_1_90 b_1 NI_1 NS_90 0 -1.8648166809013798e-02
GC_1_91 b_1 NI_1 NS_91 0 -2.0425432789350248e-05
GC_1_92 b_1 NI_1 NS_92 0 4.3970970783254755e-05
GC_1_93 b_1 NI_1 NS_93 0 -4.9911093016427707e-05
GC_1_94 b_1 NI_1 NS_94 0 3.8562923245575451e-05
GC_1_95 b_1 NI_1 NS_95 0 -7.9760337451183677e-05
GC_1_96 b_1 NI_1 NS_96 0 2.6368965399389159e-05
GC_1_97 b_1 NI_1 NS_97 0 -4.7376855356545164e-05
GC_1_98 b_1 NI_1 NS_98 0 -2.0609916030783225e-05
GC_1_99 b_1 NI_1 NS_99 0 -6.8818992432827337e-03
GC_1_100 b_1 NI_1 NS_100 0 9.5613655517597339e-03
GC_1_101 b_1 NI_1 NS_101 0 -4.4134715143751761e-04
GC_1_102 b_1 NI_1 NS_102 0 -8.7287213952908979e-04
GC_1_103 b_1 NI_1 NS_103 0 9.9826580140823242e-05
GC_1_104 b_1 NI_1 NS_104 0 -8.0633012442567578e-04
GC_1_105 b_1 NI_1 NS_105 0 -5.8180413954773205e-05
GC_1_106 b_1 NI_1 NS_106 0 1.1744433098889590e-04
GC_1_107 b_1 NI_1 NS_107 0 3.3429252365941907e-05
GC_1_108 b_1 NI_1 NS_108 0 -2.5162636003712549e-05
GC_1_109 b_1 NI_1 NS_109 0 1.0933256797598855e-05
GC_1_110 b_1 NI_1 NS_110 0 -4.1734037718263358e-05
GC_1_111 b_1 NI_1 NS_111 0 3.3589445116990426e-05
GC_1_112 b_1 NI_1 NS_112 0 4.6712129804751619e-05
GC_1_113 b_1 NI_1 NS_113 0 -3.0245274965552642e-06
GC_1_114 b_1 NI_1 NS_114 0 -2.1823156734097347e-05
GC_1_115 b_1 NI_1 NS_115 0 4.6918996303763789e-02
GC_1_116 b_1 NI_1 NS_116 0 9.5175003908571254e-04
GC_1_117 b_1 NI_1 NS_117 0 -2.3991815423288865e-02
GC_1_118 b_1 NI_1 NS_118 0 -8.5613364136407754e-03
GC_1_119 b_1 NI_1 NS_119 0 3.3749504296659973e-04
GC_1_120 b_1 NI_1 NS_120 0 2.3567729855460939e-04
GC_1_121 b_1 NI_1 NS_121 0 6.0091159007593968e-05
GC_1_122 b_1 NI_1 NS_122 0 -3.0968443300845738e-05
GC_1_123 b_1 NI_1 NS_123 0 -2.2167859133124423e-02
GC_1_124 b_1 NI_1 NS_124 0 -3.9930126250198192e-02
GC_1_125 b_1 NI_1 NS_125 0 5.7345741813366296e-05
GC_1_126 b_1 NI_1 NS_126 0 8.9687003769448319e-05
GC_1_127 b_1 NI_1 NS_127 0 1.4218144553906589e-02
GC_1_128 b_1 NI_1 NS_128 0 -6.1773959939576371e-03
GC_1_129 b_1 NI_1 NS_129 0 -1.5276087199723002e-05
GC_1_130 b_1 NI_1 NS_130 0 2.5154329590049305e-06
GC_1_131 b_1 NI_1 NS_131 0 -4.3516903537862830e-05
GC_1_132 b_1 NI_1 NS_132 0 2.9770762275706330e-05
GC_1_133 b_1 NI_1 NS_133 0 -4.5496413678883696e-05
GC_1_134 b_1 NI_1 NS_134 0 -6.6928898341052905e-06
GC_1_135 b_1 NI_1 NS_135 0 -8.4995362453942343e-05
GC_1_136 b_1 NI_1 NS_136 0 -2.9800897348258094e-05
GC_1_137 b_1 NI_1 NS_137 0 -7.3286419760752930e-03
GC_1_138 b_1 NI_1 NS_138 0 7.5406808639995188e-03
GC_1_139 b_1 NI_1 NS_139 0 1.2005299355973576e-05
GC_1_140 b_1 NI_1 NS_140 0 -1.1072893023910293e-03
GC_1_141 b_1 NI_1 NS_141 0 3.2176174986001566e-04
GC_1_142 b_1 NI_1 NS_142 0 -7.7197315295882900e-04
GC_1_143 b_1 NI_1 NS_143 0 -1.0165011229349856e-04
GC_1_144 b_1 NI_1 NS_144 0 1.0155342936533567e-04
GC_1_145 b_1 NI_1 NS_145 0 4.1726959517787869e-05
GC_1_146 b_1 NI_1 NS_146 0 2.0460240106657596e-05
GC_1_147 b_1 NI_1 NS_147 0 3.8728392779762029e-05
GC_1_148 b_1 NI_1 NS_148 0 -3.3021358330545765e-05
GC_1_149 b_1 NI_1 NS_149 0 2.7863663045171219e-06
GC_1_150 b_1 NI_1 NS_150 0 5.7341013921523302e-05
GC_1_151 b_1 NI_1 NS_151 0 2.3794412432357431e-06
GC_1_152 b_1 NI_1 NS_152 0 -1.1728646503574080e-05
GC_1_153 b_1 NI_1 NS_153 0 -3.2188801210878498e-02
GC_1_154 b_1 NI_1 NS_154 0 -1.1241405309017781e-03
GC_1_155 b_1 NI_1 NS_155 0 1.4244167656580932e-02
GC_1_156 b_1 NI_1 NS_156 0 1.8916724866412500e-02
GC_1_157 b_1 NI_1 NS_157 0 1.9076681024447683e-04
GC_1_158 b_1 NI_1 NS_158 0 3.5721267304668213e-06
GC_1_159 b_1 NI_1 NS_159 0 -9.0201098687638803e-05
GC_1_160 b_1 NI_1 NS_160 0 1.0889445360337820e-04
GC_1_161 b_1 NI_1 NS_161 0 9.8052455155111795e-03
GC_1_162 b_1 NI_1 NS_162 0 1.0291667833388661e-02
GC_1_163 b_1 NI_1 NS_163 0 -2.7827928302149400e-05
GC_1_164 b_1 NI_1 NS_164 0 1.8957874277442287e-06
GC_1_165 b_1 NI_1 NS_165 0 1.4131971102857729e-02
GC_1_166 b_1 NI_1 NS_166 0 -1.5304046184102820e-02
GC_1_167 b_1 NI_1 NS_167 0 -1.0284047090093823e-05
GC_1_168 b_1 NI_1 NS_168 0 2.2017342491942941e-05
GC_1_169 b_1 NI_1 NS_169 0 -3.1579080361274381e-05
GC_1_170 b_1 NI_1 NS_170 0 4.0468757340660636e-05
GC_1_171 b_1 NI_1 NS_171 0 1.7174472671103824e-05
GC_1_172 b_1 NI_1 NS_172 0 1.6685482562742546e-05
GC_1_173 b_1 NI_1 NS_173 0 1.0878146744810198e-05
GC_1_174 b_1 NI_1 NS_174 0 1.4951767979893850e-06
GC_1_175 b_1 NI_1 NS_175 0 -2.8644479843243750e-03
GC_1_176 b_1 NI_1 NS_176 0 4.9853452530148074e-03
GC_1_177 b_1 NI_1 NS_177 0 -5.2683169013240225e-04
GC_1_178 b_1 NI_1 NS_178 0 -8.2190136274773418e-04
GC_1_179 b_1 NI_1 NS_179 0 -1.3725038526491877e-04
GC_1_180 b_1 NI_1 NS_180 0 -7.8407212946381686e-04
GC_1_181 b_1 NI_1 NS_181 0 -9.6729348161980018e-06
GC_1_182 b_1 NI_1 NS_182 0 2.8515155242716709e-04
GC_1_183 b_1 NI_1 NS_183 0 -4.5413575980261187e-05
GC_1_184 b_1 NI_1 NS_184 0 1.0551725753051919e-04
GC_1_185 b_1 NI_1 NS_185 0 2.6488977630058210e-06
GC_1_186 b_1 NI_1 NS_186 0 7.9233770939662348e-05
GC_1_187 b_1 NI_1 NS_187 0 8.1010313841314534e-05
GC_1_188 b_1 NI_1 NS_188 0 9.7842348544995982e-05
GC_1_189 b_1 NI_1 NS_189 0 -2.6828637035585078e-05
GC_1_190 b_1 NI_1 NS_190 0 -4.0184060664876233e-05
GC_1_191 b_1 NI_1 NS_191 0 2.4178326584252253e-03
GC_1_192 b_1 NI_1 NS_192 0 1.2757471181307502e-03
GC_1_193 b_1 NI_1 NS_193 0 -4.4337191139083637e-03
GC_1_194 b_1 NI_1 NS_194 0 6.6354183585103435e-03
GC_1_195 b_1 NI_1 NS_195 0 -6.2658384800678066e-05
GC_1_196 b_1 NI_1 NS_196 0 -1.6625398041982380e-04
GC_1_197 b_1 NI_1 NS_197 0 -2.6207852308386311e-05
GC_1_198 b_1 NI_1 NS_198 0 -5.0791884244800923e-06
GC_1_199 b_1 NI_1 NS_199 0 -4.1617461402393384e-03
GC_1_200 b_1 NI_1 NS_200 0 -2.2673697139994884e-03
GC_1_201 b_1 NI_1 NS_201 0 3.9083015204156583e-05
GC_1_202 b_1 NI_1 NS_202 0 3.7325123546996073e-06
GC_1_203 b_1 NI_1 NS_203 0 9.5292113965731538e-03
GC_1_204 b_1 NI_1 NS_204 0 -5.1998320189605412e-03
GC_1_205 b_1 NI_1 NS_205 0 -7.5097917316433048e-06
GC_1_206 b_1 NI_1 NS_206 0 -4.8420226051586350e-07
GC_1_207 b_1 NI_1 NS_207 0 -1.9775251951928636e-05
GC_1_208 b_1 NI_1 NS_208 0 1.5570491630930006e-05
GC_1_209 b_1 NI_1 NS_209 0 1.8954086279978643e-05
GC_1_210 b_1 NI_1 NS_210 0 -1.2690666474478618e-05
GC_1_211 b_1 NI_1 NS_211 0 -7.5635491711978307e-06
GC_1_212 b_1 NI_1 NS_212 0 2.9259148356205519e-06
GC_1_213 b_1 NI_1 NS_213 0 -1.3630737497482672e-03
GC_1_214 b_1 NI_1 NS_214 0 2.6990652204350219e-03
GC_1_215 b_1 NI_1 NS_215 0 -3.1433243388243797e-04
GC_1_216 b_1 NI_1 NS_216 0 -5.7769938275662716e-04
GC_1_217 b_1 NI_1 NS_217 0 -7.8696851711446968e-05
GC_1_218 b_1 NI_1 NS_218 0 -5.9334478062514123e-04
GC_1_219 b_1 NI_1 NS_219 0 -5.5416326010870961e-05
GC_1_220 b_1 NI_1 NS_220 0 1.9006851331876691e-04
GC_1_221 b_1 NI_1 NS_221 0 -9.2353665730955797e-05
GC_1_222 b_1 NI_1 NS_222 0 -8.7763326963737179e-05
GC_1_223 b_1 NI_1 NS_223 0 -7.7298046790358146e-05
GC_1_224 b_1 NI_1 NS_224 0 1.6349453087673841e-05
GC_1_225 b_1 NI_1 NS_225 0 6.5680326140255964e-05
GC_1_226 b_1 NI_1 NS_226 0 9.3310826033092458e-05
GC_1_227 b_1 NI_1 NS_227 0 -3.2476573043885679e-06
GC_1_228 b_1 NI_1 NS_228 0 -4.9509390879380475e-05
GC_1_229 b_1 NI_1 NS_229 0 -1.4590837568084696e-02
GC_1_230 b_1 NI_1 NS_230 0 -9.7658014189895494e-04
GC_1_231 b_1 NI_1 NS_231 0 2.8849302026386536e-03
GC_1_232 b_1 NI_1 NS_232 0 1.0660660547352525e-02
GC_1_233 b_1 NI_1 NS_233 0 2.8907803126399650e-04
GC_1_234 b_1 NI_1 NS_234 0 -3.1791246069200554e-04
GC_1_235 b_1 NI_1 NS_235 0 5.7955616305363761e-05
GC_1_236 b_1 NI_1 NS_236 0 -8.9854426092035584e-06
GC_1_237 b_1 NI_1 NS_237 0 4.5969205200758912e-03
GC_1_238 b_1 NI_1 NS_238 0 -1.0911706460923903e-03
GC_1_239 b_1 NI_1 NS_239 0 -1.6371468497657230e-05
GC_1_240 b_1 NI_1 NS_240 0 3.5436566821676679e-06
GC_1_241 b_1 NI_1 NS_241 0 8.0996293001833249e-03
GC_1_242 b_1 NI_1 NS_242 0 -7.9714428752573341e-03
GC_1_243 b_1 NI_1 NS_243 0 -1.0753767815149645e-05
GC_1_244 b_1 NI_1 NS_244 0 2.8766925558150364e-06
GC_1_245 b_1 NI_1 NS_245 0 -1.7133419281552935e-05
GC_1_246 b_1 NI_1 NS_246 0 2.9860485477361859e-05
GC_1_247 b_1 NI_1 NS_247 0 3.7297981409058403e-05
GC_1_248 b_1 NI_1 NS_248 0 1.4573857699229308e-05
GC_1_249 b_1 NI_1 NS_249 0 2.3374805911718736e-06
GC_1_250 b_1 NI_1 NS_250 0 1.1095401964979381e-05
GC_1_251 b_1 NI_1 NS_251 0 2.6655517752210414e-04
GC_1_252 b_1 NI_1 NS_252 0 2.8026211158875465e-03
GC_1_253 b_1 NI_1 NS_253 0 -4.8457496582264602e-04
GC_1_254 b_1 NI_1 NS_254 0 -4.4664101027849529e-04
GC_1_255 b_1 NI_1 NS_255 0 -2.4747836630911941e-04
GC_1_256 b_1 NI_1 NS_256 0 -3.9012679990455728e-04
GC_1_257 b_1 NI_1 NS_257 0 -8.7730796227172034e-05
GC_1_258 b_1 NI_1 NS_258 0 3.5207486229409742e-04
GC_1_259 b_1 NI_1 NS_259 0 -2.8764843259068368e-05
GC_1_260 b_1 NI_1 NS_260 0 4.6273964386944755e-05
GC_1_261 b_1 NI_1 NS_261 0 1.2080181515046684e-05
GC_1_262 b_1 NI_1 NS_262 0 4.9148839024000083e-06
GC_1_263 b_1 NI_1 NS_263 0 -1.5959633396132440e-05
GC_1_264 b_1 NI_1 NS_264 0 8.6850608606439561e-05
GC_1_265 b_1 NI_1 NS_265 0 7.4548889640918308e-06
GC_1_266 b_1 NI_1 NS_266 0 -1.1847656711697213e-05
GC_1_267 b_1 NI_1 NS_267 0 7.8599479261189167e-03
GC_1_268 b_1 NI_1 NS_268 0 1.1231864585735762e-03
GC_1_269 b_1 NI_1 NS_269 0 -8.2824915266546655e-03
GC_1_270 b_1 NI_1 NS_270 0 7.9313933431573516e-03
GC_1_271 b_1 NI_1 NS_271 0 -3.4439967074084312e-05
GC_1_272 b_1 NI_1 NS_272 0 -2.6131151974763449e-04
GC_1_273 b_1 NI_1 NS_273 0 3.8416003344253910e-05
GC_1_274 b_1 NI_1 NS_274 0 -1.9606227953378973e-05
GC_1_275 b_1 NI_1 NS_275 0 -1.1516219355582908e-03
GC_1_276 b_1 NI_1 NS_276 0 6.1451470750385449e-03
GC_1_277 b_1 NI_1 NS_277 0 2.7448858624557906e-05
GC_1_278 b_1 NI_1 NS_278 0 -1.0352181883514750e-06
GC_1_279 b_1 NI_1 NS_279 0 7.4351566029204758e-03
GC_1_280 b_1 NI_1 NS_280 0 -2.8371018056722007e-03
GC_1_281 b_1 NI_1 NS_281 0 7.3953960816620329e-07
GC_1_282 b_1 NI_1 NS_282 0 -7.0799338589079926e-06
GC_1_283 b_1 NI_1 NS_283 0 -1.1393145065014159e-05
GC_1_284 b_1 NI_1 NS_284 0 1.0296265425555772e-05
GC_1_285 b_1 NI_1 NS_285 0 2.1143878849388985e-05
GC_1_286 b_1 NI_1 NS_286 0 6.8779692203848365e-06
GC_1_287 b_1 NI_1 NS_287 0 -1.7141447257151437e-05
GC_1_288 b_1 NI_1 NS_288 0 9.5060533966882349e-06
GC_1_289 b_1 NI_1 NS_289 0 -5.1234239053487109e-04
GC_1_290 b_1 NI_1 NS_290 0 2.3448483710771296e-03
GC_1_291 b_1 NI_1 NS_291 0 -2.2839666310580484e-04
GC_1_292 b_1 NI_1 NS_292 0 -4.3182061719659469e-04
GC_1_293 b_1 NI_1 NS_293 0 -4.1587821827057640e-05
GC_1_294 b_1 NI_1 NS_294 0 -3.8978878656681273e-04
GC_1_295 b_1 NI_1 NS_295 0 -1.7937842475420284e-04
GC_1_296 b_1 NI_1 NS_296 0 2.4930704561710931e-04
GC_1_297 b_1 NI_1 NS_297 0 -6.5062380817462628e-05
GC_1_298 b_1 NI_1 NS_298 0 -1.7574977819482310e-05
GC_1_299 b_1 NI_1 NS_299 0 1.4897702923055356e-05
GC_1_300 b_1 NI_1 NS_300 0 1.0950305803272533e-05
GC_1_301 b_1 NI_1 NS_301 0 -3.9188049967716994e-05
GC_1_302 b_1 NI_1 NS_302 0 6.8775857610461940e-05
GC_1_303 b_1 NI_1 NS_303 0 1.3676319918399610e-05
GC_1_304 b_1 NI_1 NS_304 0 -1.2746500661368081e-05
GC_1_305 b_1 NI_1 NS_305 0 1.1317842816901506e-02
GC_1_306 b_1 NI_1 NS_306 0 -7.4996207040337482e-04
GC_1_307 b_1 NI_1 NS_307 0 -1.1349910223059577e-02
GC_1_308 b_1 NI_1 NS_308 0 6.3516962073581094e-03
GC_1_309 b_1 NI_1 NS_309 0 4.2981257075341118e-04
GC_1_310 b_1 NI_1 NS_310 0 -6.0569244353291484e-04
GC_1_311 b_1 NI_1 NS_311 0 1.5495003777453659e-04
GC_1_312 b_1 NI_1 NS_312 0 -1.5851039650095333e-04
GC_1_313 b_1 NI_1 NS_313 0 7.1864019018527431e-04
GC_1_314 b_1 NI_1 NS_314 0 -4.9678850074451695e-03
GC_1_315 b_1 NI_1 NS_315 0 -1.9006975163588711e-05
GC_1_316 b_1 NI_1 NS_316 0 3.9729466145524387e-05
GC_1_317 b_1 NI_1 NS_317 0 7.1329690637405609e-03
GC_1_318 b_1 NI_1 NS_318 0 1.0861131294561425e-03
GC_1_319 b_1 NI_1 NS_319 0 -2.6156636600684902e-05
GC_1_320 b_1 NI_1 NS_320 0 1.0729429812939124e-05
GC_1_321 b_1 NI_1 NS_321 0 -2.8017547864817243e-05
GC_1_322 b_1 NI_1 NS_322 0 3.9785812126366603e-05
GC_1_323 b_1 NI_1 NS_323 0 1.3432538663544377e-04
GC_1_324 b_1 NI_1 NS_324 0 -1.0815750296379228e-06
GC_1_325 b_1 NI_1 NS_325 0 4.4661568918835692e-05
GC_1_326 b_1 NI_1 NS_326 0 3.4175001552559253e-05
GC_1_327 b_1 NI_1 NS_327 0 -1.1001497359123921e-03
GC_1_328 b_1 NI_1 NS_328 0 1.2466325849872632e-03
GC_1_329 b_1 NI_1 NS_329 0 -1.4387294016977414e-04
GC_1_330 b_1 NI_1 NS_330 0 -5.6899665343646520e-04
GC_1_331 b_1 NI_1 NS_331 0 9.2176360397452624e-05
GC_1_332 b_1 NI_1 NS_332 0 -3.2726721037370512e-04
GC_1_333 b_1 NI_1 NS_333 0 -1.3793729808534387e-04
GC_1_334 b_1 NI_1 NS_334 0 2.1575652889225126e-04
GC_1_335 b_1 NI_1 NS_335 0 -2.8127143661438519e-05
GC_1_336 b_1 NI_1 NS_336 0 -6.3699364273830624e-05
GC_1_337 b_1 NI_1 NS_337 0 -2.8324407138860249e-05
GC_1_338 b_1 NI_1 NS_338 0 3.5070484897085010e-05
GC_1_339 b_1 NI_1 NS_339 0 -3.5357334491426649e-06
GC_1_340 b_1 NI_1 NS_340 0 7.1642898604165080e-05
GC_1_341 b_1 NI_1 NS_341 0 1.7217128791756168e-05
GC_1_342 b_1 NI_1 NS_342 0 -2.3061900704197748e-05
GC_1_343 b_1 NI_1 NS_343 0 9.4377489885013790e-03
GC_1_344 b_1 NI_1 NS_344 0 7.6168678886991636e-04
GC_1_345 b_1 NI_1 NS_345 0 -7.2020937236107162e-03
GC_1_346 b_1 NI_1 NS_346 0 9.2330377661732947e-04
GC_1_347 b_1 NI_1 NS_347 0 8.7783499637153383e-05
GC_1_348 b_1 NI_1 NS_348 0 -1.4228469608315301e-04
GC_1_349 b_1 NI_1 NS_349 0 6.1952679154929580e-05
GC_1_350 b_1 NI_1 NS_350 0 -4.5139144264482775e-05
GC_1_351 b_1 NI_1 NS_351 0 -1.0154978327770192e-03
GC_1_352 b_1 NI_1 NS_352 0 5.0973672206220417e-03
GC_1_353 b_1 NI_1 NS_353 0 2.2250669753009084e-05
GC_1_354 b_1 NI_1 NS_354 0 -3.3073376518780374e-05
GC_1_355 b_1 NI_1 NS_355 0 2.4283165962179650e-03
GC_1_356 b_1 NI_1 NS_356 0 2.4954725882599146e-03
GC_1_357 b_1 NI_1 NS_357 0 -1.1169593771853770e-05
GC_1_358 b_1 NI_1 NS_358 0 2.0638576206109754e-05
GC_1_359 b_1 NI_1 NS_359 0 -2.9919691003254073e-05
GC_1_360 b_1 NI_1 NS_360 0 3.3750716271744255e-05
GC_1_361 b_1 NI_1 NS_361 0 6.9109447238761723e-05
GC_1_362 b_1 NI_1 NS_362 0 -8.2386287700561847e-06
GC_1_363 b_1 NI_1 NS_363 0 3.7904461026536230e-05
GC_1_364 b_1 NI_1 NS_364 0 3.0649327973390549e-05
GC_1_365 b_1 NI_1 NS_365 0 -5.5283374971222456e-04
GC_1_366 b_1 NI_1 NS_366 0 6.0956695598034629e-04
GC_1_367 b_1 NI_1 NS_367 0 7.5289815548352609e-05
GC_1_368 b_1 NI_1 NS_368 0 -5.9359535494219015e-04
GC_1_369 b_1 NI_1 NS_369 0 -1.1399785794970051e-05
GC_1_370 b_1 NI_1 NS_370 0 -3.1204729850078147e-04
GC_1_371 b_1 NI_1 NS_371 0 -1.4002721937395512e-04
GC_1_372 b_1 NI_1 NS_372 0 1.5161204844804386e-04
GC_1_373 b_1 NI_1 NS_373 0 -1.5366906868318875e-05
GC_1_374 b_1 NI_1 NS_374 0 3.9513429811979284e-06
GC_1_375 b_1 NI_1 NS_375 0 -1.2900963988652920e-05
GC_1_376 b_1 NI_1 NS_376 0 5.9710543632293013e-05
GC_1_377 b_1 NI_1 NS_377 0 1.0584966502936365e-05
GC_1_378 b_1 NI_1 NS_378 0 -1.4312604221007201e-05
GC_1_379 b_1 NI_1 NS_379 0 -1.3643748884979131e-05
GC_1_380 b_1 NI_1 NS_380 0 9.2972711127377677e-07
GC_1_381 b_1 NI_1 NS_381 0 8.5419941104449941e-03
GC_1_382 b_1 NI_1 NS_382 0 -4.9689569339204421e-04
GC_1_383 b_1 NI_1 NS_383 0 -6.6708855844563623e-03
GC_1_384 b_1 NI_1 NS_384 0 3.0245285987089568e-03
GC_1_385 b_1 NI_1 NS_385 0 4.1886245843274590e-05
GC_1_386 b_1 NI_1 NS_386 0 -2.6208377348180464e-05
GC_1_387 b_1 NI_1 NS_387 0 1.7916193879894353e-04
GC_1_388 b_1 NI_1 NS_388 0 -1.6276076715084978e-04
GC_1_389 b_1 NI_1 NS_389 0 -1.1767213761023893e-04
GC_1_390 b_1 NI_1 NS_390 0 -4.2758636550417140e-03
GC_1_391 b_1 NI_1 NS_391 0 -1.6650486615285754e-05
GC_1_392 b_1 NI_1 NS_392 0 3.6525990696184113e-05
GC_1_393 b_1 NI_1 NS_393 0 2.4608527846076687e-03
GC_1_394 b_1 NI_1 NS_394 0 7.9712738294196082e-04
GC_1_395 b_1 NI_1 NS_395 0 -4.0241120619459865e-06
GC_1_396 b_1 NI_1 NS_396 0 1.0939495429389081e-05
GC_1_397 b_1 NI_1 NS_397 0 1.0195199248034885e-05
GC_1_398 b_1 NI_1 NS_398 0 2.1819517184922678e-05
GC_1_399 b_1 NI_1 NS_399 0 1.3691765670682061e-04
GC_1_400 b_1 NI_1 NS_400 0 -1.9802455018768589e-05
GC_1_401 b_1 NI_1 NS_401 0 3.3573864028800613e-05
GC_1_402 b_1 NI_1 NS_402 0 2.3801831435226048e-05
GC_1_403 b_1 NI_1 NS_403 0 2.5634821791055255e-04
GC_1_404 b_1 NI_1 NS_404 0 1.1310494063061702e-04
GC_1_405 b_1 NI_1 NS_405 0 -2.0051874928366851e-04
GC_1_406 b_1 NI_1 NS_406 0 -2.4647001502487370e-04
GC_1_407 b_1 NI_1 NS_407 0 2.8763905312154228e-05
GC_1_408 b_1 NI_1 NS_408 0 6.7724777813653306e-05
GC_1_409 b_1 NI_1 NS_409 0 -9.6072245079193076e-05
GC_1_410 b_1 NI_1 NS_410 0 2.0919693422001724e-04
GC_1_411 b_1 NI_1 NS_411 0 8.5561778943220123e-06
GC_1_412 b_1 NI_1 NS_412 0 -7.2599888897102057e-05
GC_1_413 b_1 NI_1 NS_413 0 1.7602840319329817e-06
GC_1_414 b_1 NI_1 NS_414 0 7.5003810095596724e-05
GC_1_415 b_1 NI_1 NS_415 0 -2.2611990802127010e-05
GC_1_416 b_1 NI_1 NS_416 0 -1.9114435409901747e-05
GC_1_417 b_1 NI_1 NS_417 0 1.0465183154318432e-05
GC_1_418 b_1 NI_1 NS_418 0 6.6404457612953573e-06
GC_1_419 b_1 NI_1 NS_419 0 -1.2388777377791134e-03
GC_1_420 b_1 NI_1 NS_420 0 5.1570779410900860e-04
GC_1_421 b_1 NI_1 NS_421 0 -6.5345123656219343e-04
GC_1_422 b_1 NI_1 NS_422 0 -9.2586254206822836e-04
GC_1_423 b_1 NI_1 NS_423 0 -9.1862157244503330e-05
GC_1_424 b_1 NI_1 NS_424 0 2.2352116033090086e-04
GC_1_425 b_1 NI_1 NS_425 0 7.3111175376819822e-05
GC_1_426 b_1 NI_1 NS_426 0 -1.0500395908718404e-05
GC_1_427 b_1 NI_1 NS_427 0 2.7462077488182804e-05
GC_1_428 b_1 NI_1 NS_428 0 4.5900424685715330e-03
GC_1_429 b_1 NI_1 NS_429 0 1.9614335606212422e-05
GC_1_430 b_1 NI_1 NS_430 0 -3.2331328643351105e-05
GC_1_431 b_1 NI_1 NS_431 0 4.1682482618242872e-04
GC_1_432 b_1 NI_1 NS_432 0 2.0360928778539403e-04
GC_1_433 b_1 NI_1 NS_433 0 5.9368288029028471e-06
GC_1_434 b_1 NI_1 NS_434 0 3.3468415382194080e-05
GC_1_435 b_1 NI_1 NS_435 0 -5.4464038262793241e-07
GC_1_436 b_1 NI_1 NS_436 0 3.3307342287631789e-05
GC_1_437 b_1 NI_1 NS_437 0 8.3237861023324378e-05
GC_1_438 b_1 NI_1 NS_438 0 1.5055238942432173e-07
GC_1_439 b_1 NI_1 NS_439 0 2.7190034221547944e-05
GC_1_440 b_1 NI_1 NS_440 0 2.6244531516631304e-05
GC_1_441 b_1 NI_1 NS_441 0 -2.5006515524590909e-05
GC_1_442 b_1 NI_1 NS_442 0 4.9807465442752404e-04
GC_1_443 b_1 NI_1 NS_443 0 9.8187510865033233e-05
GC_1_444 b_1 NI_1 NS_444 0 -4.7653960398673785e-04
GC_1_445 b_1 NI_1 NS_445 0 -1.0709213354238736e-05
GC_1_446 b_1 NI_1 NS_446 0 -1.2070415055190458e-04
GC_1_447 b_1 NI_1 NS_447 0 -1.9293921916005067e-04
GC_1_448 b_1 NI_1 NS_448 0 1.7760718034843127e-04
GC_1_449 b_1 NI_1 NS_449 0 3.9441088389546425e-05
GC_1_450 b_1 NI_1 NS_450 0 -4.2471877949187512e-05
GC_1_451 b_1 NI_1 NS_451 0 -4.4345429089529055e-05
GC_1_452 b_1 NI_1 NS_452 0 6.7680638143282563e-05
GC_1_453 b_1 NI_1 NS_453 0 7.0036416828120619e-06
GC_1_454 b_1 NI_1 NS_454 0 -4.1817353351585225e-05
GC_1_455 b_1 NI_1 NS_455 0 -1.3573710407840314e-06
GC_1_456 b_1 NI_1 NS_456 0 1.1220227395361187e-05
GD_1_1 b_1 NI_1 NA_1 0 -7.9874683997289128e-02
GD_1_2 b_1 NI_1 NA_2 0 -3.3257000726479913e-02
GD_1_3 b_1 NI_1 NA_3 0 -2.6417015392010114e-02
GD_1_4 b_1 NI_1 NA_4 0 -5.6184608176892319e-03
GD_1_5 b_1 NI_1 NA_5 0 -6.7857744185622270e-03
GD_1_6 b_1 NI_1 NA_6 0 -2.7828060221248680e-03
GD_1_7 b_1 NI_1 NA_7 0 -2.5259571609359084e-03
GD_1_8 b_1 NI_1 NA_8 0 -5.6753042802240219e-03
GD_1_9 b_1 NI_1 NA_9 0 -6.0496873434184298e-03
GD_1_10 b_1 NI_1 NA_10 0 -3.2463454549814131e-03
GD_1_11 b_1 NI_1 NA_11 0 -3.5471208340938300e-03
GD_1_12 b_1 NI_1 NA_12 0 1.1841434918443481e-03
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 1.0651026835158717e-02
GC_2_2 b_2 NI_2 NS_2 0 1.8827170391979937e-03
GC_2_3 b_2 NI_2 NS_3 0 2.3026350423349454e-02
GC_2_4 b_2 NI_2 NS_4 0 -4.8878978634441577e-03
GC_2_5 b_2 NI_2 NS_5 0 1.5236754000792926e-03
GC_2_6 b_2 NI_2 NS_6 0 -3.7328940244383445e-04
GC_2_7 b_2 NI_2 NS_7 0 1.5101682698137964e-04
GC_2_8 b_2 NI_2 NS_8 0 -8.9723492575311819e-05
GC_2_9 b_2 NI_2 NS_9 0 2.8807374754398336e-02
GC_2_10 b_2 NI_2 NS_10 0 6.2176936377808540e-03
GC_2_11 b_2 NI_2 NS_11 0 8.4526490686065439e-05
GC_2_12 b_2 NI_2 NS_12 0 9.8787522729438837e-05
GC_2_13 b_2 NI_2 NS_13 0 -3.7001701453448547e-02
GC_2_14 b_2 NI_2 NS_14 0 2.4515003681792394e-02
GC_2_15 b_2 NI_2 NS_15 0 2.0118864998413178e-05
GC_2_16 b_2 NI_2 NS_16 0 -1.9169979416647599e-05
GC_2_17 b_2 NI_2 NS_17 0 -2.1327513113687770e-05
GC_2_18 b_2 NI_2 NS_18 0 2.3716191240720035e-05
GC_2_19 b_2 NI_2 NS_19 0 3.4204263628804247e-06
GC_2_20 b_2 NI_2 NS_20 0 -4.2893575245951021e-06
GC_2_21 b_2 NI_2 NS_21 0 -8.0155204973828825e-05
GC_2_22 b_2 NI_2 NS_22 0 -3.1763208047225851e-05
GC_2_23 b_2 NI_2 NS_23 0 -4.8797289508780723e-03
GC_2_24 b_2 NI_2 NS_24 0 5.0548175694464870e-03
GC_2_25 b_2 NI_2 NS_25 0 -1.3088355165743692e-05
GC_2_26 b_2 NI_2 NS_26 0 -1.0262738814007728e-03
GC_2_27 b_2 NI_2 NS_27 0 8.3615905412129092e-05
GC_2_28 b_2 NI_2 NS_28 0 -7.1118197270883586e-04
GC_2_29 b_2 NI_2 NS_29 0 8.3565615787569282e-05
GC_2_30 b_2 NI_2 NS_30 0 9.2884544729550950e-05
GC_2_31 b_2 NI_2 NS_31 0 1.7747114393865698e-04
GC_2_32 b_2 NI_2 NS_32 0 5.4669583069097508e-05
GC_2_33 b_2 NI_2 NS_33 0 8.8939885053881363e-05
GC_2_34 b_2 NI_2 NS_34 0 -1.7282773760459312e-05
GC_2_35 b_2 NI_2 NS_35 0 1.6069802497437007e-05
GC_2_36 b_2 NI_2 NS_36 0 1.0946227546055804e-04
GC_2_37 b_2 NI_2 NS_37 0 3.2579922699029806e-05
GC_2_38 b_2 NI_2 NS_38 0 3.8080050508583096e-07
GC_2_39 b_2 NI_2 NS_39 0 1.0269859825691248e-01
GC_2_40 b_2 NI_2 NS_40 0 -1.3843636239412353e-03
GC_2_41 b_2 NI_2 NS_41 0 1.4724669215979468e-02
GC_2_42 b_2 NI_2 NS_42 0 -3.8986387026068013e-02
GC_2_43 b_2 NI_2 NS_43 0 2.4406911341859922e-04
GC_2_44 b_2 NI_2 NS_44 0 -5.7344901555439779e-04
GC_2_45 b_2 NI_2 NS_45 0 2.1849303016131576e-06
GC_2_46 b_2 NI_2 NS_46 0 -3.7498357030497566e-05
GC_2_47 b_2 NI_2 NS_47 0 -1.2396669483318419e-02
GC_2_48 b_2 NI_2 NS_48 0 1.3466713538117887e-02
GC_2_49 b_2 NI_2 NS_49 0 -6.2083838767553373e-05
GC_2_50 b_2 NI_2 NS_50 0 -8.5183635054604742e-05
GC_2_51 b_2 NI_2 NS_51 0 -1.8686313439370831e-02
GC_2_52 b_2 NI_2 NS_52 0 8.7865116922901682e-03
GC_2_53 b_2 NI_2 NS_53 0 -4.9905605293764151e-05
GC_2_54 b_2 NI_2 NS_54 0 1.6002353110674100e-07
GC_2_55 b_2 NI_2 NS_55 0 -2.7249946770514102e-05
GC_2_56 b_2 NI_2 NS_56 0 3.4010383258287460e-05
GC_2_57 b_2 NI_2 NS_57 0 1.3984969137274758e-05
GC_2_58 b_2 NI_2 NS_58 0 -2.0166333257834389e-06
GC_2_59 b_2 NI_2 NS_59 0 -1.3322024959410271e-04
GC_2_60 b_2 NI_2 NS_60 0 -4.5558303683665563e-05
GC_2_61 b_2 NI_2 NS_61 0 -6.2845415145934159e-03
GC_2_62 b_2 NI_2 NS_62 0 6.6893970822377094e-03
GC_2_63 b_2 NI_2 NS_63 0 3.2684831302101723e-04
GC_2_64 b_2 NI_2 NS_64 0 -1.2753569874515052e-03
GC_2_65 b_2 NI_2 NS_65 0 2.4279717222351927e-04
GC_2_66 b_2 NI_2 NS_66 0 -8.7905290495073160e-04
GC_2_67 b_2 NI_2 NS_67 0 -6.1476723768741424e-06
GC_2_68 b_2 NI_2 NS_68 0 3.1828548347910570e-05
GC_2_69 b_2 NI_2 NS_69 0 5.2678862353003275e-05
GC_2_70 b_2 NI_2 NS_70 0 1.5743795175319599e-04
GC_2_71 b_2 NI_2 NS_71 0 8.5557767581250264e-05
GC_2_72 b_2 NI_2 NS_72 0 5.3330247578275053e-05
GC_2_73 b_2 NI_2 NS_73 0 -1.1728960696203093e-05
GC_2_74 b_2 NI_2 NS_74 0 7.0741612908760141e-05
GC_2_75 b_2 NI_2 NS_75 0 1.8032532010913246e-07
GC_2_76 b_2 NI_2 NS_76 0 9.4614517145977879e-07
GC_2_77 b_2 NI_2 NS_77 0 4.4906646503149003e-02
GC_2_78 b_2 NI_2 NS_78 0 1.0098540319137892e-03
GC_2_79 b_2 NI_2 NS_79 0 -3.3448160768010562e-02
GC_2_80 b_2 NI_2 NS_80 0 -9.6425326836972157e-03
GC_2_81 b_2 NI_2 NS_81 0 -7.3728499014054632e-04
GC_2_82 b_2 NI_2 NS_82 0 -5.8861728127255915e-05
GC_2_83 b_2 NI_2 NS_83 0 -5.4327280889544964e-05
GC_2_84 b_2 NI_2 NS_84 0 9.3904588989898905e-07
GC_2_85 b_2 NI_2 NS_85 0 -2.2113167281513916e-02
GC_2_86 b_2 NI_2 NS_86 0 -4.0057244045921134e-02
GC_2_87 b_2 NI_2 NS_87 0 5.8191133235432072e-05
GC_2_88 b_2 NI_2 NS_88 0 8.6733333291950595e-05
GC_2_89 b_2 NI_2 NS_89 0 1.9374089560457695e-02
GC_2_90 b_2 NI_2 NS_90 0 -4.8949123496303650e-03
GC_2_91 b_2 NI_2 NS_91 0 -1.1448432147835330e-05
GC_2_92 b_2 NI_2 NS_92 0 -6.8727804184841458e-06
GC_2_93 b_2 NI_2 NS_93 0 -4.8172302928197696e-05
GC_2_94 b_2 NI_2 NS_94 0 4.1741281785086407e-05
GC_2_95 b_2 NI_2 NS_95 0 -1.0562297738045195e-05
GC_2_96 b_2 NI_2 NS_96 0 -1.3324055153591920e-05
GC_2_97 b_2 NI_2 NS_97 0 -7.3175484945249230e-05
GC_2_98 b_2 NI_2 NS_98 0 -2.4624261359288859e-05
GC_2_99 b_2 NI_2 NS_99 0 -6.6072909017288531e-03
GC_2_100 b_2 NI_2 NS_100 0 7.3716077301789109e-03
GC_2_101 b_2 NI_2 NS_101 0 -9.3846437015536561e-05
GC_2_102 b_2 NI_2 NS_102 0 -9.5569058241785519e-04
GC_2_103 b_2 NI_2 NS_103 0 2.3931078919401522e-04
GC_2_104 b_2 NI_2 NS_104 0 -7.1252240520128544e-04
GC_2_105 b_2 NI_2 NS_105 0 -7.2488112916791817e-05
GC_2_106 b_2 NI_2 NS_106 0 7.5916825465962250e-05
GC_2_107 b_2 NI_2 NS_107 0 3.6331488394681978e-05
GC_2_108 b_2 NI_2 NS_108 0 1.1184717393855726e-05
GC_2_109 b_2 NI_2 NS_109 0 4.2164067419478642e-05
GC_2_110 b_2 NI_2 NS_110 0 -1.8490159448206894e-05
GC_2_111 b_2 NI_2 NS_111 0 6.3580639750910700e-06
GC_2_112 b_2 NI_2 NS_112 0 6.6122090833454299e-05
GC_2_113 b_2 NI_2 NS_113 0 1.5455521458592374e-06
GC_2_114 b_2 NI_2 NS_114 0 -2.6659176082446626e-06
GC_2_115 b_2 NI_2 NS_115 0 2.7843718933642184e-02
GC_2_116 b_2 NI_2 NS_116 0 -1.3958882137996955e-03
GC_2_117 b_2 NI_2 NS_117 0 -1.8781833740685743e-02
GC_2_118 b_2 NI_2 NS_118 0 1.5374934639103325e-03
GC_2_119 b_2 NI_2 NS_119 0 -1.1052374501098765e-04
GC_2_120 b_2 NI_2 NS_120 0 8.6907220341963598e-06
GC_2_121 b_2 NI_2 NS_121 0 -6.8244063814531573e-05
GC_2_122 b_2 NI_2 NS_122 0 8.9280080623942200e-05
GC_2_123 b_2 NI_2 NS_123 0 5.5126314557419577e-03
GC_2_124 b_2 NI_2 NS_124 0 2.1162901512775043e-02
GC_2_125 b_2 NI_2 NS_125 0 -6.4492432675637416e-05
GC_2_126 b_2 NI_2 NS_126 0 -8.5830346877220859e-05
GC_2_127 b_2 NI_2 NS_127 0 1.2318223227272794e-02
GC_2_128 b_2 NI_2 NS_128 0 2.0662887039058085e-03
GC_2_129 b_2 NI_2 NS_129 0 -4.1391239936346504e-05
GC_2_130 b_2 NI_2 NS_130 0 5.8552806532566784e-05
GC_2_131 b_2 NI_2 NS_131 0 -4.3606452443289284e-05
GC_2_132 b_2 NI_2 NS_132 0 5.0319220168712435e-05
GC_2_133 b_2 NI_2 NS_133 0 1.2460970498963716e-06
GC_2_134 b_2 NI_2 NS_134 0 -6.0395013970604174e-06
GC_2_135 b_2 NI_2 NS_135 0 -1.3967199906119788e-04
GC_2_136 b_2 NI_2 NS_136 0 -3.6578396108286973e-05
GC_2_137 b_2 NI_2 NS_137 0 -7.6749529260695696e-03
GC_2_138 b_2 NI_2 NS_138 0 5.7994706364983360e-03
GC_2_139 b_2 NI_2 NS_139 0 4.3794498101753300e-04
GC_2_140 b_2 NI_2 NS_140 0 -1.0747401656436518e-03
GC_2_141 b_2 NI_2 NS_141 0 4.3551852783254820e-04
GC_2_142 b_2 NI_2 NS_142 0 -7.2205130692936498e-04
GC_2_143 b_2 NI_2 NS_143 0 -1.0782302552584957e-04
GC_2_144 b_2 NI_2 NS_144 0 5.0009078055113034e-05
GC_2_145 b_2 NI_2 NS_145 0 6.2085875786300695e-06
GC_2_146 b_2 NI_2 NS_146 0 4.6956380856858470e-05
GC_2_147 b_2 NI_2 NS_147 0 4.8375767663846462e-05
GC_2_148 b_2 NI_2 NS_148 0 3.9594008367703881e-06
GC_2_149 b_2 NI_2 NS_149 0 -8.2439516759388127e-06
GC_2_150 b_2 NI_2 NS_150 0 5.8701658958189134e-05
GC_2_151 b_2 NI_2 NS_151 0 -4.5287747262386293e-06
GC_2_152 b_2 NI_2 NS_152 0 -1.2267366418168520e-05
GC_2_153 b_2 NI_2 NS_153 0 2.4454542388991023e-02
GC_2_154 b_2 NI_2 NS_154 0 1.2486812281270114e-03
GC_2_155 b_2 NI_2 NS_155 0 -1.3688565839528283e-02
GC_2_156 b_2 NI_2 NS_156 0 7.3662054352561391e-03
GC_2_157 b_2 NI_2 NS_157 0 -1.1679029918811092e-04
GC_2_158 b_2 NI_2 NS_158 0 2.5932176926355500e-04
GC_2_159 b_2 NI_2 NS_159 0 1.5402650893642064e-05
GC_2_160 b_2 NI_2 NS_160 0 -6.3259751201254547e-05
GC_2_161 b_2 NI_2 NS_161 0 -7.5914573390637877e-03
GC_2_162 b_2 NI_2 NS_162 0 -6.6537181025567056e-03
GC_2_163 b_2 NI_2 NS_163 0 3.1118477861073515e-05
GC_2_164 b_2 NI_2 NS_164 0 3.6341371599101956e-06
GC_2_165 b_2 NI_2 NS_165 0 1.2578555437239430e-02
GC_2_166 b_2 NI_2 NS_166 0 -4.1410771229659820e-03
GC_2_167 b_2 NI_2 NS_167 0 2.4606981013310094e-05
GC_2_168 b_2 NI_2 NS_168 0 -2.1105028301260717e-05
GC_2_169 b_2 NI_2 NS_169 0 -2.2598965846465716e-05
GC_2_170 b_2 NI_2 NS_170 0 5.8673631689935920e-05
GC_2_171 b_2 NI_2 NS_171 0 8.5325412911728244e-06
GC_2_172 b_2 NI_2 NS_172 0 1.9647298769095240e-06
GC_2_173 b_2 NI_2 NS_173 0 1.9206357364165006e-05
GC_2_174 b_2 NI_2 NS_174 0 3.2121239509603164e-06
GC_2_175 b_2 NI_2 NS_175 0 -3.8538054948637915e-03
GC_2_176 b_2 NI_2 NS_176 0 4.4434809101242265e-03
GC_2_177 b_2 NI_2 NS_177 0 -1.9679972603884986e-04
GC_2_178 b_2 NI_2 NS_178 0 -1.0660725520377935e-03
GC_2_179 b_2 NI_2 NS_179 0 -3.1095791846252190e-05
GC_2_180 b_2 NI_2 NS_180 0 -7.9284534773663585e-04
GC_2_181 b_2 NI_2 NS_181 0 -6.7900369287862846e-05
GC_2_182 b_2 NI_2 NS_182 0 2.3103621851552962e-04
GC_2_183 b_2 NI_2 NS_183 0 -1.0971167505116470e-04
GC_2_184 b_2 NI_2 NS_184 0 1.3590007494779571e-05
GC_2_185 b_2 NI_2 NS_185 0 -2.9430444933014041e-05
GC_2_186 b_2 NI_2 NS_186 0 5.8691885455844515e-05
GC_2_187 b_2 NI_2 NS_187 0 1.7815950424658677e-05
GC_2_188 b_2 NI_2 NS_188 0 1.5427058602861282e-04
GC_2_189 b_2 NI_2 NS_189 0 2.2686109950368386e-05
GC_2_190 b_2 NI_2 NS_190 0 2.1521631059979744e-05
GC_2_191 b_2 NI_2 NS_191 0 -1.6742568955586727e-02
GC_2_192 b_2 NI_2 NS_192 0 -1.1938106668352906e-03
GC_2_193 b_2 NI_2 NS_193 0 6.4186937867928096e-04
GC_2_194 b_2 NI_2 NS_194 0 1.0394551550417779e-02
GC_2_195 b_2 NI_2 NS_195 0 -1.8237192011791927e-04
GC_2_196 b_2 NI_2 NS_196 0 2.2337638669260171e-05
GC_2_197 b_2 NI_2 NS_197 0 -4.1233071539963545e-05
GC_2_198 b_2 NI_2 NS_198 0 -1.4491997418321080e-05
GC_2_199 b_2 NI_2 NS_199 0 7.5915543081407633e-03
GC_2_200 b_2 NI_2 NS_200 0 7.4925433398412237e-03
GC_2_201 b_2 NI_2 NS_201 0 -2.9456128702818613e-05
GC_2_202 b_2 NI_2 NS_202 0 -2.2041775846189952e-06
GC_2_203 b_2 NI_2 NS_203 0 1.2167654123172222e-02
GC_2_204 b_2 NI_2 NS_204 0 -6.7260140255376551e-03
GC_2_205 b_2 NI_2 NS_205 0 -1.4499698140497847e-05
GC_2_206 b_2 NI_2 NS_206 0 1.2139487942276129e-05
GC_2_207 b_2 NI_2 NS_207 0 -2.2658310814780305e-05
GC_2_208 b_2 NI_2 NS_208 0 2.7670794889029227e-05
GC_2_209 b_2 NI_2 NS_209 0 5.6745626273946885e-06
GC_2_210 b_2 NI_2 NS_210 0 -2.9482193272391084e-06
GC_2_211 b_2 NI_2 NS_211 0 -1.2771765753973611e-05
GC_2_212 b_2 NI_2 NS_212 0 5.7272882978034620e-06
GC_2_213 b_2 NI_2 NS_213 0 -2.6452180020804738e-03
GC_2_214 b_2 NI_2 NS_214 0 3.9280347521953567e-03
GC_2_215 b_2 NI_2 NS_215 0 -1.1065005979964606e-04
GC_2_216 b_2 NI_2 NS_216 0 -8.0410134233353488e-04
GC_2_217 b_2 NI_2 NS_217 0 5.5549458767874146e-05
GC_2_218 b_2 NI_2 NS_218 0 -6.7263713999161673e-04
GC_2_219 b_2 NI_2 NS_219 0 -9.8895828297210017e-05
GC_2_220 b_2 NI_2 NS_220 0 1.2941608284195967e-04
GC_2_221 b_2 NI_2 NS_221 0 1.1506404187529180e-07
GC_2_222 b_2 NI_2 NS_222 0 -1.2995263167945992e-04
GC_2_223 b_2 NI_2 NS_223 0 -2.6014687576196976e-05
GC_2_224 b_2 NI_2 NS_224 0 -4.9425742033245981e-05
GC_2_225 b_2 NI_2 NS_225 0 1.2024231891020202e-05
GC_2_226 b_2 NI_2 NS_226 0 1.1972742707531927e-04
GC_2_227 b_2 NI_2 NS_227 0 4.5968119243747581e-06
GC_2_228 b_2 NI_2 NS_228 0 1.2806494658002612e-05
GC_2_229 b_2 NI_2 NS_229 0 9.5796389711342682e-03
GC_2_230 b_2 NI_2 NS_230 0 1.1362924778278486e-03
GC_2_231 b_2 NI_2 NS_231 0 -9.1221717804130485e-03
GC_2_232 b_2 NI_2 NS_232 0 5.8762828187022102e-03
GC_2_233 b_2 NI_2 NS_233 0 5.8317042738960229e-05
GC_2_234 b_2 NI_2 NS_234 0 6.7266207274294722e-05
GC_2_235 b_2 NI_2 NS_235 0 4.8865310625932813e-06
GC_2_236 b_2 NI_2 NS_236 0 -6.6602248437735862e-05
GC_2_237 b_2 NI_2 NS_237 0 -1.1382651407322937e-03
GC_2_238 b_2 NI_2 NS_238 0 6.6170851859905519e-03
GC_2_239 b_2 NI_2 NS_239 0 2.1092243425458295e-05
GC_2_240 b_2 NI_2 NS_240 0 7.7624736406749301e-07
GC_2_241 b_2 NI_2 NS_241 0 7.6360801543900875e-03
GC_2_242 b_2 NI_2 NS_242 0 -9.9564076348239439e-04
GC_2_243 b_2 NI_2 NS_243 0 1.3548793480422770e-05
GC_2_244 b_2 NI_2 NS_244 0 -1.8040049903969937e-05
GC_2_245 b_2 NI_2 NS_245 0 -6.0788991279168812e-06
GC_2_246 b_2 NI_2 NS_246 0 4.8589452208827620e-05
GC_2_247 b_2 NI_2 NS_247 0 1.0144236048381345e-05
GC_2_248 b_2 NI_2 NS_248 0 5.0180362389180876e-06
GC_2_249 b_2 NI_2 NS_249 0 6.2466725930924349e-06
GC_2_250 b_2 NI_2 NS_250 0 1.8153583468823333e-05
GC_2_251 b_2 NI_2 NS_251 0 -1.3092308746739103e-03
GC_2_252 b_2 NI_2 NS_252 0 2.3539156458999670e-03
GC_2_253 b_2 NI_2 NS_253 0 -1.6271075622619673e-04
GC_2_254 b_2 NI_2 NS_254 0 -6.2410897866869844e-04
GC_2_255 b_2 NI_2 NS_255 0 -4.0202186006690152e-05
GC_2_256 b_2 NI_2 NS_256 0 -4.2849986525718084e-04
GC_2_257 b_2 NI_2 NS_257 0 -8.5911754021258827e-05
GC_2_258 b_2 NI_2 NS_258 0 2.5324857045888166e-04
GC_2_259 b_2 NI_2 NS_259 0 -5.2747907154711885e-05
GC_2_260 b_2 NI_2 NS_260 0 2.7784937560626351e-06
GC_2_261 b_2 NI_2 NS_261 0 1.1869385762332296e-05
GC_2_262 b_2 NI_2 NS_262 0 8.1580037638937585e-06
GC_2_263 b_2 NI_2 NS_263 0 1.7327773768508060e-05
GC_2_264 b_2 NI_2 NS_264 0 6.5323310906497268e-05
GC_2_265 b_2 NI_2 NS_265 0 -1.3441274571298048e-05
GC_2_266 b_2 NI_2 NS_266 0 -2.4890686839644642e-05
GC_2_267 b_2 NI_2 NS_267 0 -1.9134560293949446e-02
GC_2_268 b_2 NI_2 NS_268 0 -1.0287198775640112e-03
GC_2_269 b_2 NI_2 NS_269 0 3.5560768603972595e-03
GC_2_270 b_2 NI_2 NS_270 0 8.3936877055946491e-03
GC_2_271 b_2 NI_2 NS_271 0 2.4696697697747810e-05
GC_2_272 b_2 NI_2 NS_272 0 -9.1459255127580310e-05
GC_2_273 b_2 NI_2 NS_273 0 -4.5822662576773147e-05
GC_2_274 b_2 NI_2 NS_274 0 1.8035066379807503e-05
GC_2_275 b_2 NI_2 NS_275 0 4.9834326711422896e-03
GC_2_276 b_2 NI_2 NS_276 0 -1.0725222150016968e-03
GC_2_277 b_2 NI_2 NS_277 0 -2.0578140971306858e-05
GC_2_278 b_2 NI_2 NS_278 0 2.5749804406711746e-06
GC_2_279 b_2 NI_2 NS_279 0 9.3384561337339321e-03
GC_2_280 b_2 NI_2 NS_280 0 -7.4119342946753208e-03
GC_2_281 b_2 NI_2 NS_281 0 9.0336914351127627e-07
GC_2_282 b_2 NI_2 NS_282 0 2.6095597491587582e-05
GC_2_283 b_2 NI_2 NS_283 0 -1.5577205468935963e-05
GC_2_284 b_2 NI_2 NS_284 0 2.6682605100473874e-05
GC_2_285 b_2 NI_2 NS_285 0 4.6317129973240880e-06
GC_2_286 b_2 NI_2 NS_286 0 1.1814747731537416e-07
GC_2_287 b_2 NI_2 NS_287 0 -2.7670353228714959e-05
GC_2_288 b_2 NI_2 NS_288 0 1.5730623088292574e-05
GC_2_289 b_2 NI_2 NS_289 0 -1.7663235038365521e-03
GC_2_290 b_2 NI_2 NS_290 0 3.2729911000229078e-03
GC_2_291 b_2 NI_2 NS_291 0 -1.9692568078135887e-05
GC_2_292 b_2 NI_2 NS_292 0 -5.6526298717673909e-04
GC_2_293 b_2 NI_2 NS_293 0 1.3175389445692890e-04
GC_2_294 b_2 NI_2 NS_294 0 -4.6464838391093767e-04
GC_2_295 b_2 NI_2 NS_295 0 -1.6935564120636214e-04
GC_2_296 b_2 NI_2 NS_296 0 1.6192707574590965e-04
GC_2_297 b_2 NI_2 NS_297 0 -3.0382540455613861e-05
GC_2_298 b_2 NI_2 NS_298 0 -5.4079138851963173e-05
GC_2_299 b_2 NI_2 NS_299 0 7.2707235170291237e-06
GC_2_300 b_2 NI_2 NS_300 0 4.8476181956317214e-06
GC_2_301 b_2 NI_2 NS_301 0 -9.8043959587319445e-06
GC_2_302 b_2 NI_2 NS_302 0 5.4741398347935594e-05
GC_2_303 b_2 NI_2 NS_303 0 -1.3757194825962334e-06
GC_2_304 b_2 NI_2 NS_304 0 -2.8254052199654990e-05
GC_2_305 b_2 NI_2 NS_305 0 -6.7357232759896156e-03
GC_2_306 b_2 NI_2 NS_306 0 8.2734121436904128e-04
GC_2_307 b_2 NI_2 NS_307 0 1.0004315217329105e-03
GC_2_308 b_2 NI_2 NS_308 0 -9.2292144513046043e-03
GC_2_309 b_2 NI_2 NS_309 0 -3.7287836685008902e-06
GC_2_310 b_2 NI_2 NS_310 0 8.0043120315762028e-04
GC_2_311 b_2 NI_2 NS_311 0 3.8383367919482954e-05
GC_2_312 b_2 NI_2 NS_312 0 1.3981017585489706e-04
GC_2_313 b_2 NI_2 NS_313 0 2.1086382287467965e-05
GC_2_314 b_2 NI_2 NS_314 0 7.0555614226072792e-03
GC_2_315 b_2 NI_2 NS_315 0 2.2150447888279270e-05
GC_2_316 b_2 NI_2 NS_316 0 -3.1865270908716176e-05
GC_2_317 b_2 NI_2 NS_317 0 2.8333542137604296e-04
GC_2_318 b_2 NI_2 NS_318 0 3.7445470254451429e-03
GC_2_319 b_2 NI_2 NS_319 0 4.8671961674401152e-05
GC_2_320 b_2 NI_2 NS_320 0 6.0519232473996767e-05
GC_2_321 b_2 NI_2 NS_321 0 -1.5301173500985719e-05
GC_2_322 b_2 NI_2 NS_322 0 8.8606389873236056e-05
GC_2_323 b_2 NI_2 NS_323 0 1.8994469683077860e-05
GC_2_324 b_2 NI_2 NS_324 0 2.0650507818271372e-05
GC_2_325 b_2 NI_2 NS_325 0 7.3548906828309446e-05
GC_2_326 b_2 NI_2 NS_326 0 5.0569622273354552e-05
GC_2_327 b_2 NI_2 NS_327 0 -1.5520411258263291e-03
GC_2_328 b_2 NI_2 NS_328 0 9.3337436845366458e-05
GC_2_329 b_2 NI_2 NS_329 0 2.2341481457431928e-04
GC_2_330 b_2 NI_2 NS_330 0 -5.9917206203754180e-04
GC_2_331 b_2 NI_2 NS_331 0 1.8599270753850099e-04
GC_2_332 b_2 NI_2 NS_332 0 -2.9580291672337994e-04
GC_2_333 b_2 NI_2 NS_333 0 -1.2185274120640143e-04
GC_2_334 b_2 NI_2 NS_334 0 1.6010820550193576e-04
GC_2_335 b_2 NI_2 NS_335 0 2.5411978782271468e-05
GC_2_336 b_2 NI_2 NS_336 0 -6.7810943980528080e-05
GC_2_337 b_2 NI_2 NS_337 0 -2.6913840633104730e-05
GC_2_338 b_2 NI_2 NS_338 0 6.8258138824941862e-06
GC_2_339 b_2 NI_2 NS_339 0 -3.1762236799811244e-05
GC_2_340 b_2 NI_2 NS_340 0 6.7559223982036729e-05
GC_2_341 b_2 NI_2 NS_341 0 5.8011170330429400e-06
GC_2_342 b_2 NI_2 NS_342 0 6.4624222089377477e-07
GC_2_343 b_2 NI_2 NS_343 0 7.7922810071475350e-03
GC_2_344 b_2 NI_2 NS_344 0 -8.1321772808482537e-04
GC_2_345 b_2 NI_2 NS_345 0 -7.5105718574250508e-03
GC_2_346 b_2 NI_2 NS_346 0 -4.0557208720238070e-03
GC_2_347 b_2 NI_2 NS_347 0 1.0926908815040627e-04
GC_2_348 b_2 NI_2 NS_348 0 2.0190860866914820e-04
GC_2_349 b_2 NI_2 NS_349 0 3.4349253885962620e-05
GC_2_350 b_2 NI_2 NS_350 0 9.5203017138084629e-05
GC_2_351 b_2 NI_2 NS_351 0 -2.0548214717297356e-04
GC_2_352 b_2 NI_2 NS_352 0 -6.8745975272847043e-03
GC_2_353 b_2 NI_2 NS_353 0 -2.3831861460607272e-05
GC_2_354 b_2 NI_2 NS_354 0 2.8334784450190213e-05
GC_2_355 b_2 NI_2 NS_355 0 3.9174412781514158e-03
GC_2_356 b_2 NI_2 NS_356 0 5.0602839171838389e-03
GC_2_357 b_2 NI_2 NS_357 0 5.7307274923675275e-05
GC_2_358 b_2 NI_2 NS_358 0 5.4375089253430649e-05
GC_2_359 b_2 NI_2 NS_359 0 -1.4927697411173972e-05
GC_2_360 b_2 NI_2 NS_360 0 6.5501188112214873e-05
GC_2_361 b_2 NI_2 NS_361 0 1.3431919042343565e-05
GC_2_362 b_2 NI_2 NS_362 0 1.5206285027272250e-05
GC_2_363 b_2 NI_2 NS_363 0 6.0601833385788017e-05
GC_2_364 b_2 NI_2 NS_364 0 4.6012916425120759e-05
GC_2_365 b_2 NI_2 NS_365 0 -2.2718081459470159e-03
GC_2_366 b_2 NI_2 NS_366 0 3.9767442761518045e-04
GC_2_367 b_2 NI_2 NS_367 0 3.8241881849600295e-04
GC_2_368 b_2 NI_2 NS_368 0 -6.7399738082608157e-04
GC_2_369 b_2 NI_2 NS_369 0 1.6608857738253005e-04
GC_2_370 b_2 NI_2 NS_370 0 -3.6132906695310086e-04
GC_2_371 b_2 NI_2 NS_371 0 -1.2799432439965694e-04
GC_2_372 b_2 NI_2 NS_372 0 9.4648912295661655e-05
GC_2_373 b_2 NI_2 NS_373 0 -2.1317665689589989e-05
GC_2_374 b_2 NI_2 NS_374 0 -7.8120499537232875e-06
GC_2_375 b_2 NI_2 NS_375 0 -4.4546725441746127e-05
GC_2_376 b_2 NI_2 NS_376 0 1.0523822276958472e-05
GC_2_377 b_2 NI_2 NS_377 0 3.0892428542550562e-05
GC_2_378 b_2 NI_2 NS_378 0 -2.8813279633652060e-06
GC_2_379 b_2 NI_2 NS_379 0 7.5762539436130283e-06
GC_2_380 b_2 NI_2 NS_380 0 1.6180155687220631e-06
GC_2_381 b_2 NI_2 NS_381 0 -6.0891644580837187e-03
GC_2_382 b_2 NI_2 NS_382 0 5.1284647626996212e-04
GC_2_383 b_2 NI_2 NS_383 0 2.0297249605622596e-03
GC_2_384 b_2 NI_2 NS_384 0 -7.2133164204792703e-03
GC_2_385 b_2 NI_2 NS_385 0 1.6452870892688431e-05
GC_2_386 b_2 NI_2 NS_386 0 3.8607085645534444e-04
GC_2_387 b_2 NI_2 NS_387 0 6.7672575239282911e-06
GC_2_388 b_2 NI_2 NS_388 0 1.6247950466898373e-04
GC_2_389 b_2 NI_2 NS_389 0 -6.3362370656991083e-05
GC_2_390 b_2 NI_2 NS_390 0 4.4581827383140408e-03
GC_2_391 b_2 NI_2 NS_391 0 1.8118271791205940e-05
GC_2_392 b_2 NI_2 NS_392 0 -3.1341299908877874e-05
GC_2_393 b_2 NI_2 NS_393 0 -1.8163961246184209e-03
GC_2_394 b_2 NI_2 NS_394 0 2.2732331889647878e-03
GC_2_395 b_2 NI_2 NS_395 0 1.5960019179492392e-05
GC_2_396 b_2 NI_2 NS_396 0 6.2604102593316992e-05
GC_2_397 b_2 NI_2 NS_397 0 2.2757009225522485e-05
GC_2_398 b_2 NI_2 NS_398 0 3.8454740021755051e-05
GC_2_399 b_2 NI_2 NS_399 0 1.5255512051063282e-05
GC_2_400 b_2 NI_2 NS_400 0 1.1679489898863155e-05
GC_2_401 b_2 NI_2 NS_401 0 5.7222165608991990e-05
GC_2_402 b_2 NI_2 NS_402 0 3.4478833742332644e-05
GC_2_403 b_2 NI_2 NS_403 0 -2.1949629061749276e-04
GC_2_404 b_2 NI_2 NS_404 0 -4.2444969104626131e-04
GC_2_405 b_2 NI_2 NS_405 0 7.1381891954491129e-05
GC_2_406 b_2 NI_2 NS_406 0 -3.0009897917500193e-04
GC_2_407 b_2 NI_2 NS_407 0 1.0856582869410921e-04
GC_2_408 b_2 NI_2 NS_408 0 -1.0593351885154416e-05
GC_2_409 b_2 NI_2 NS_409 0 -7.5738490590704548e-05
GC_2_410 b_2 NI_2 NS_410 0 1.5424521762712900e-04
GC_2_411 b_2 NI_2 NS_411 0 5.0741669282899014e-05
GC_2_412 b_2 NI_2 NS_412 0 -3.6179183789107997e-05
GC_2_413 b_2 NI_2 NS_413 0 -5.7671963375390980e-05
GC_2_414 b_2 NI_2 NS_414 0 4.0656272831485748e-05
GC_2_415 b_2 NI_2 NS_415 0 -2.2724833986002238e-05
GC_2_416 b_2 NI_2 NS_416 0 -4.9982670859545206e-05
GC_2_417 b_2 NI_2 NS_417 0 3.6063592699771421e-06
GC_2_418 b_2 NI_2 NS_418 0 3.9597869406959149e-06
GC_2_419 b_2 NI_2 NS_419 0 6.3440071676991033e-03
GC_2_420 b_2 NI_2 NS_420 0 -5.5836183856769147e-04
GC_2_421 b_2 NI_2 NS_421 0 -5.2521164479901157e-03
GC_2_422 b_2 NI_2 NS_422 0 -4.4858401717756740e-03
GC_2_423 b_2 NI_2 NS_423 0 8.0082659816472072e-05
GC_2_424 b_2 NI_2 NS_424 0 8.9791422255136423e-05
GC_2_425 b_2 NI_2 NS_425 0 -5.5764321987182278e-06
GC_2_426 b_2 NI_2 NS_426 0 1.2806677172180346e-04
GC_2_427 b_2 NI_2 NS_427 0 -7.8554240246968927e-04
GC_2_428 b_2 NI_2 NS_428 0 -5.9315531719057847e-03
GC_2_429 b_2 NI_2 NS_429 0 -2.0761637562601214e-05
GC_2_430 b_2 NI_2 NS_430 0 2.6683474468596911e-05
GC_2_431 b_2 NI_2 NS_431 0 1.9552758909398968e-03
GC_2_432 b_2 NI_2 NS_432 0 4.1917737609174733e-03
GC_2_433 b_2 NI_2 NS_433 0 3.8972294983543728e-05
GC_2_434 b_2 NI_2 NS_434 0 5.5701416210861472e-05
GC_2_435 b_2 NI_2 NS_435 0 1.2633121127726174e-05
GC_2_436 b_2 NI_2 NS_436 0 4.0861767815829384e-05
GC_2_437 b_2 NI_2 NS_437 0 1.1063491219519908e-05
GC_2_438 b_2 NI_2 NS_438 0 8.6024052662507949e-06
GC_2_439 b_2 NI_2 NS_439 0 4.6828918939163682e-05
GC_2_440 b_2 NI_2 NS_440 0 3.9094885225908928e-05
GC_2_441 b_2 NI_2 NS_441 0 -1.8761000853194201e-03
GC_2_442 b_2 NI_2 NS_442 0 1.1362116912694472e-04
GC_2_443 b_2 NI_2 NS_443 0 4.4578106744120515e-04
GC_2_444 b_2 NI_2 NS_444 0 -5.3002153439179144e-04
GC_2_445 b_2 NI_2 NS_445 0 2.3017488978325885e-04
GC_2_446 b_2 NI_2 NS_446 0 -2.2603774462416135e-04
GC_2_447 b_2 NI_2 NS_447 0 -1.6770892489566933e-04
GC_2_448 b_2 NI_2 NS_448 0 9.9080396311860709e-05
GC_2_449 b_2 NI_2 NS_449 0 4.4992876413129622e-05
GC_2_450 b_2 NI_2 NS_450 0 3.5275462039524061e-06
GC_2_451 b_2 NI_2 NS_451 0 -7.5820246047620960e-05
GC_2_452 b_2 NI_2 NS_452 0 -7.5056908702646344e-06
GC_2_453 b_2 NI_2 NS_453 0 2.5240953737656808e-05
GC_2_454 b_2 NI_2 NS_454 0 -7.2476864272677340e-05
GC_2_455 b_2 NI_2 NS_455 0 -2.9013162033531307e-06
GC_2_456 b_2 NI_2 NS_456 0 9.9041084060414563e-06
GD_2_1 b_2 NI_2 NA_1 0 -3.3257023698683996e-02
GD_2_2 b_2 NI_2 NA_2 0 -1.4455964424875617e-01
GD_2_3 b_2 NI_2 NA_3 0 5.6270751421489225e-03
GD_2_4 b_2 NI_2 NA_4 0 -1.2289446340743537e-02
GD_2_5 b_2 NI_2 NA_5 0 -1.2140451874073427e-02
GD_2_6 b_2 NI_2 NA_6 0 2.3087122746019009e-04
GD_2_7 b_2 NI_2 NA_7 0 -6.3704395317998319e-03
GD_2_8 b_2 NI_2 NA_8 0 3.0898996475311933e-03
GD_2_9 b_2 NI_2 NA_9 0 5.6987502162232570e-03
GD_2_10 b_2 NI_2 NA_10 0 -8.2353152620211504e-04
GD_2_11 b_2 NI_2 NA_11 0 5.6421802316679896e-03
GD_2_12 b_2 NI_2 NA_12 0 2.7983352121760125e-04
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 -1.0704681850964588e-02
GC_3_2 b_3 NI_3 NS_2 0 -1.2959594644571470e-03
GC_3_3 b_3 NI_3 NS_3 0 7.4730742017340510e-03
GC_3_4 b_3 NI_3 NS_4 0 2.6999431900822386e-02
GC_3_5 b_3 NI_3 NS_5 0 -6.6140035530856808e-04
GC_3_6 b_3 NI_3 NS_6 0 8.1782028166218644e-04
GC_3_7 b_3 NI_3 NS_7 0 -1.4920215600097052e-04
GC_3_8 b_3 NI_3 NS_8 0 2.1319085796439209e-04
GC_3_9 b_3 NI_3 NS_9 0 1.1678156967848278e-02
GC_3_10 b_3 NI_3 NS_10 0 2.6150037192165878e-02
GC_3_11 b_3 NI_3 NS_11 0 -8.0788508449279451e-05
GC_3_12 b_3 NI_3 NS_12 0 -9.4560313484867990e-05
GC_3_13 b_3 NI_3 NS_13 0 2.5073142883660200e-02
GC_3_14 b_3 NI_3 NS_14 0 -1.8648045323804863e-02
GC_3_15 b_3 NI_3 NS_15 0 -2.0425501146832069e-05
GC_3_16 b_3 NI_3 NS_16 0 4.3971487278065076e-05
GC_3_17 b_3 NI_3 NS_17 0 -4.9911196231412579e-05
GC_3_18 b_3 NI_3 NS_18 0 3.8563287793189700e-05
GC_3_19 b_3 NI_3 NS_19 0 -7.9760517317430858e-05
GC_3_20 b_3 NI_3 NS_20 0 2.6369130322289026e-05
GC_3_21 b_3 NI_3 NS_21 0 -4.7376974584809137e-05
GC_3_22 b_3 NI_3 NS_22 0 -2.0609936695758527e-05
GC_3_23 b_3 NI_3 NS_23 0 -6.8818927436894101e-03
GC_3_24 b_3 NI_3 NS_24 0 9.5613042878111548e-03
GC_3_25 b_3 NI_3 NS_25 0 -4.4134657446301645e-04
GC_3_26 b_3 NI_3 NS_26 0 -8.7286341438918744e-04
GC_3_27 b_3 NI_3 NS_27 0 9.9830121451865205e-05
GC_3_28 b_3 NI_3 NS_28 0 -8.0632018496186268e-04
GC_3_29 b_3 NI_3 NS_29 0 -5.8178333247594773e-05
GC_3_30 b_3 NI_3 NS_30 0 1.1744348332144341e-04
GC_3_31 b_3 NI_3 NS_31 0 3.3429064622996049e-05
GC_3_32 b_3 NI_3 NS_32 0 -2.5162915829746015e-05
GC_3_33 b_3 NI_3 NS_33 0 1.0933833225394028e-05
GC_3_34 b_3 NI_3 NS_34 0 -4.1733939952106521e-05
GC_3_35 b_3 NI_3 NS_35 0 3.3590246626076253e-05
GC_3_36 b_3 NI_3 NS_36 0 4.6712634622684172e-05
GC_3_37 b_3 NI_3 NS_37 0 -3.0244461079648822e-06
GC_3_38 b_3 NI_3 NS_38 0 -2.1823476107113957e-05
GC_3_39 b_3 NI_3 NS_39 0 4.4906524709699830e-02
GC_3_40 b_3 NI_3 NS_40 0 1.0098525506197231e-03
GC_3_41 b_3 NI_3 NS_41 0 -3.3448062304904443e-02
GC_3_42 b_3 NI_3 NS_42 0 -9.6429770387188272e-03
GC_3_43 b_3 NI_3 NS_43 0 -7.3728142209322214e-04
GC_3_44 b_3 NI_3 NS_44 0 -5.8838409351743835e-05
GC_3_45 b_3 NI_3 NS_45 0 -5.4324950167565800e-05
GC_3_46 b_3 NI_3 NS_46 0 9.4252371060680118e-07
GC_3_47 b_3 NI_3 NS_47 0 -2.2113205446758433e-02
GC_3_48 b_3 NI_3 NS_48 0 -4.0057309013534603e-02
GC_3_49 b_3 NI_3 NS_49 0 5.8191013215202335e-05
GC_3_50 b_3 NI_3 NS_50 0 8.6733251543189650e-05
GC_3_51 b_3 NI_3 NS_51 0 1.9373910007621949e-02
GC_3_52 b_3 NI_3 NS_52 0 -4.8947103127041716e-03
GC_3_53 b_3 NI_3 NS_53 0 -1.1447868069283763e-05
GC_3_54 b_3 NI_3 NS_54 0 -6.8716234407741745e-06
GC_3_55 b_3 NI_3 NS_55 0 -4.8172060157989754e-05
GC_3_56 b_3 NI_3 NS_56 0 4.1742097087426085e-05
GC_3_57 b_3 NI_3 NS_57 0 -1.0562437020223788e-05
GC_3_58 b_3 NI_3 NS_58 0 -1.3323581308037021e-05
GC_3_59 b_3 NI_3 NS_59 0 -7.3175692870212651e-05
GC_3_60 b_3 NI_3 NS_60 0 -2.4624194764561782e-05
GC_3_61 b_3 NI_3 NS_61 0 -6.6073021380898180e-03
GC_3_62 b_3 NI_3 NS_62 0 7.3715092934020041e-03
GC_3_63 b_3 NI_3 NS_63 0 -9.3841681206298223e-05
GC_3_64 b_3 NI_3 NS_64 0 -9.5567640518198348e-04
GC_3_65 b_3 NI_3 NS_65 0 2.3932178861085904e-04
GC_3_66 b_3 NI_3 NS_66 0 -7.1250796299871183e-04
GC_3_67 b_3 NI_3 NS_67 0 -7.2485163648864392e-05
GC_3_68 b_3 NI_3 NS_68 0 7.5914125620751870e-05
GC_3_69 b_3 NI_3 NS_69 0 3.6331100555874799e-05
GC_3_70 b_3 NI_3 NS_70 0 1.1184527308445452e-05
GC_3_71 b_3 NI_3 NS_71 0 4.2164787321537011e-05
GC_3_72 b_3 NI_3 NS_72 0 -1.8490448746398975e-05
GC_3_73 b_3 NI_3 NS_73 0 6.3597562817980098e-06
GC_3_74 b_3 NI_3 NS_74 0 6.6122113904655471e-05
GC_3_75 b_3 NI_3 NS_75 0 1.5453082186584917e-06
GC_3_76 b_3 NI_3 NS_76 0 -2.6664366792046222e-06
GC_3_77 b_3 NI_3 NS_77 0 6.6606101853789276e-02
GC_3_78 b_3 NI_3 NS_78 0 -1.8596527420712806e-03
GC_3_79 b_3 NI_3 NS_79 0 4.2158912071745692e-02
GC_3_80 b_3 NI_3 NS_80 0 -5.7701895728679280e-02
GC_3_81 b_3 NI_3 NS_81 0 -2.5022598192966984e-03
GC_3_82 b_3 NI_3 NS_82 0 -1.2989178264627684e-03
GC_3_83 b_3 NI_3 NS_83 0 -2.6498991653036119e-04
GC_3_84 b_3 NI_3 NS_84 0 5.5845218106659522e-05
GC_3_85 b_3 NI_3 NS_85 0 -1.1424835958712435e-02
GC_3_86 b_3 NI_3 NS_86 0 1.4108438539785304e-02
GC_3_87 b_3 NI_3 NS_87 0 -8.3316832387310121e-05
GC_3_88 b_3 NI_3 NS_88 0 -8.6827701420409724e-05
GC_3_89 b_3 NI_3 NS_89 0 -4.2211884260027761e-02
GC_3_90 b_3 NI_3 NS_90 0 1.0192815168473436e-02
GC_3_91 b_3 NI_3 NS_91 0 -4.6770668127562852e-05
GC_3_92 b_3 NI_3 NS_92 0 2.8512334422299287e-06
GC_3_93 b_3 NI_3 NS_93 0 -4.9985447068182472e-05
GC_3_94 b_3 NI_3 NS_94 0 3.2499089495302356e-06
GC_3_95 b_3 NI_3 NS_95 0 -7.6695781434477954e-05
GC_3_96 b_3 NI_3 NS_96 0 8.7612531029906057e-06
GC_3_97 b_3 NI_3 NS_97 0 -3.7898790028009018e-05
GC_3_98 b_3 NI_3 NS_98 0 -1.2363490220127685e-05
GC_3_99 b_3 NI_3 NS_99 0 -6.0322621419373543e-03
GC_3_100 b_3 NI_3 NS_100 0 4.1405922839926265e-03
GC_3_101 b_3 NI_3 NS_101 0 -2.7932461976897682e-04
GC_3_102 b_3 NI_3 NS_102 0 -6.6715835036612852e-04
GC_3_103 b_3 NI_3 NS_103 0 1.6676411602262531e-04
GC_3_104 b_3 NI_3 NS_104 0 -3.7344415342631604e-04
GC_3_105 b_3 NI_3 NS_105 0 -2.6712314293978512e-05
GC_3_106 b_3 NI_3 NS_106 0 8.0305445263952998e-05
GC_3_107 b_3 NI_3 NS_107 0 1.3314594566707635e-05
GC_3_108 b_3 NI_3 NS_108 0 -6.6794329646864792e-06
GC_3_109 b_3 NI_3 NS_109 0 5.0978830146351878e-06
GC_3_110 b_3 NI_3 NS_110 0 -6.1094837012586557e-06
GC_3_111 b_3 NI_3 NS_111 0 2.9195806747337765e-05
GC_3_112 b_3 NI_3 NS_112 0 7.1804835072878691e-05
GC_3_113 b_3 NI_3 NS_113 0 1.4898004285097515e-05
GC_3_114 b_3 NI_3 NS_114 0 -4.3393384713785649e-06
GC_3_115 b_3 NI_3 NS_115 0 1.5561470136141379e-02
GC_3_116 b_3 NI_3 NS_116 0 2.3525604000369476e-03
GC_3_117 b_3 NI_3 NS_117 0 2.2368783366066954e-02
GC_3_118 b_3 NI_3 NS_118 0 -1.2322490941452886e-02
GC_3_119 b_3 NI_3 NS_119 0 1.6215800158972330e-03
GC_3_120 b_3 NI_3 NS_120 0 -2.7837981311646870e-06
GC_3_121 b_3 NI_3 NS_121 0 1.3580151628676663e-04
GC_3_122 b_3 NI_3 NS_122 0 -7.5900375214469956e-05
GC_3_123 b_3 NI_3 NS_123 0 2.6760681353034124e-02
GC_3_124 b_3 NI_3 NS_124 0 6.1411247052310693e-03
GC_3_125 b_3 NI_3 NS_125 0 8.6757877783889245e-05
GC_3_126 b_3 NI_3 NS_126 0 8.8881632568016880e-05
GC_3_127 b_3 NI_3 NS_127 0 -3.9846377957156551e-02
GC_3_128 b_3 NI_3 NS_128 0 3.2317948155332628e-02
GC_3_129 b_3 NI_3 NS_129 0 2.2692107417156738e-05
GC_3_130 b_3 NI_3 NS_130 0 -1.3835185064836411e-05
GC_3_131 b_3 NI_3 NS_131 0 -1.4139493326641673e-05
GC_3_132 b_3 NI_3 NS_132 0 4.7844126970344467e-05
GC_3_133 b_3 NI_3 NS_133 0 -3.9590749021016725e-05
GC_3_134 b_3 NI_3 NS_134 0 -1.4241313405124700e-06
GC_3_135 b_3 NI_3 NS_135 0 -7.7823806696017620e-05
GC_3_136 b_3 NI_3 NS_136 0 -1.2126489985072138e-05
GC_3_137 b_3 NI_3 NS_137 0 -4.4817924492654600e-03
GC_3_138 b_3 NI_3 NS_138 0 6.3341778695482330e-04
GC_3_139 b_3 NI_3 NS_139 0 6.5595598708235859e-05
GC_3_140 b_3 NI_3 NS_140 0 -6.1039593076298525e-04
GC_3_141 b_3 NI_3 NS_141 0 2.0984700851322646e-04
GC_3_142 b_3 NI_3 NS_142 0 -2.0542529227859599e-04
GC_3_143 b_3 NI_3 NS_143 0 -4.4171046195198384e-05
GC_3_144 b_3 NI_3 NS_144 0 9.9930131290435094e-05
GC_3_145 b_3 NI_3 NS_145 0 2.7338245132940085e-05
GC_3_146 b_3 NI_3 NS_146 0 -7.2405168557233018e-08
GC_3_147 b_3 NI_3 NS_147 0 8.5936546713256282e-06
GC_3_148 b_3 NI_3 NS_148 0 1.9876329190240162e-05
GC_3_149 b_3 NI_3 NS_149 0 -1.3005387985890481e-05
GC_3_150 b_3 NI_3 NS_150 0 8.9884533517700567e-05
GC_3_151 b_3 NI_3 NS_151 0 1.9836994168841216e-05
GC_3_152 b_3 NI_3 NS_152 0 6.9973566617936380e-06
GC_3_153 b_3 NI_3 NS_153 0 4.5060895564114512e-03
GC_3_154 b_3 NI_3 NS_154 0 -1.5161834916055620e-03
GC_3_155 b_3 NI_3 NS_155 0 -3.1876384006868856e-03
GC_3_156 b_3 NI_3 NS_156 0 1.2275667149333827e-02
GC_3_157 b_3 NI_3 NS_157 0 -1.8297922411956104e-03
GC_3_158 b_3 NI_3 NS_158 0 2.5881345541045424e-05
GC_3_159 b_3 NI_3 NS_159 0 -1.6147441999403713e-04
GC_3_160 b_3 NI_3 NS_160 0 1.1411986136583047e-04
GC_3_161 b_3 NI_3 NS_161 0 5.7952619563784724e-03
GC_3_162 b_3 NI_3 NS_162 0 1.2293736651129131e-02
GC_3_163 b_3 NI_3 NS_163 0 -2.8792122053087890e-05
GC_3_164 b_3 NI_3 NS_164 0 1.1372782261889673e-07
GC_3_165 b_3 NI_3 NS_165 0 8.9702102942032531e-03
GC_3_166 b_3 NI_3 NS_166 0 -5.7599962658150556e-03
GC_3_167 b_3 NI_3 NS_167 0 -3.7184124550029336e-05
GC_3_168 b_3 NI_3 NS_168 0 3.3446472557227593e-05
GC_3_169 b_3 NI_3 NS_169 0 -3.8535095149713117e-05
GC_3_170 b_3 NI_3 NS_170 0 2.2278526263268568e-05
GC_3_171 b_3 NI_3 NS_171 0 1.9407199382852936e-05
GC_3_172 b_3 NI_3 NS_172 0 1.0714834519466659e-05
GC_3_173 b_3 NI_3 NS_173 0 1.1993563997259345e-05
GC_3_174 b_3 NI_3 NS_174 0 -3.5757068152724232e-08
GC_3_175 b_3 NI_3 NS_175 0 -5.7537980374954799e-03
GC_3_176 b_3 NI_3 NS_176 0 2.1098232424589460e-03
GC_3_177 b_3 NI_3 NS_177 0 -3.1259017676491641e-04
GC_3_178 b_3 NI_3 NS_178 0 -6.8342915179026779e-04
GC_3_179 b_3 NI_3 NS_179 0 2.2150067316064725e-04
GC_3_180 b_3 NI_3 NS_180 0 -4.2000032046220892e-04
GC_3_181 b_3 NI_3 NS_181 0 -6.5848411145599454e-06
GC_3_182 b_3 NI_3 NS_182 0 1.2313043764053928e-04
GC_3_183 b_3 NI_3 NS_183 0 -2.5752875144234834e-06
GC_3_184 b_3 NI_3 NS_184 0 2.0294137681833097e-05
GC_3_185 b_3 NI_3 NS_185 0 1.3236524368379479e-05
GC_3_186 b_3 NI_3 NS_186 0 3.4588771292081454e-05
GC_3_187 b_3 NI_3 NS_187 0 1.0389569179946272e-04
GC_3_188 b_3 NI_3 NS_188 0 1.1134558779096595e-04
GC_3_189 b_3 NI_3 NS_189 0 3.9781291236035462e-05
GC_3_190 b_3 NI_3 NS_190 0 -2.8747291313757968e-05
GC_3_191 b_3 NI_3 NS_191 0 -2.8440426196980489e-02
GC_3_192 b_3 NI_3 NS_192 0 1.4955254069561829e-03
GC_3_193 b_3 NI_3 NS_193 0 1.8245902112039723e-02
GC_3_194 b_3 NI_3 NS_194 0 5.3009871234334224e-03
GC_3_195 b_3 NI_3 NS_195 0 -4.5207070062066448e-05
GC_3_196 b_3 NI_3 NS_196 0 -2.7706599786253490e-04
GC_3_197 b_3 NI_3 NS_197 0 -3.9818197437925530e-05
GC_3_198 b_3 NI_3 NS_198 0 -2.6414770037396725e-06
GC_3_199 b_3 NI_3 NS_199 0 -7.1108117226173278e-03
GC_3_200 b_3 NI_3 NS_200 0 -1.1194010191108980e-02
GC_3_201 b_3 NI_3 NS_201 0 3.5138933100393476e-05
GC_3_202 b_3 NI_3 NS_202 0 1.6781560606055262e-06
GC_3_203 b_3 NI_3 NS_203 0 7.2416927278247173e-03
GC_3_204 b_3 NI_3 NS_204 0 -1.6740673387206178e-02
GC_3_205 b_3 NI_3 NS_205 0 -1.3406920523299379e-05
GC_3_206 b_3 NI_3 NS_206 0 2.0210504239078913e-06
GC_3_207 b_3 NI_3 NS_207 0 -1.5958746898574912e-05
GC_3_208 b_3 NI_3 NS_208 0 2.4838767145589127e-05
GC_3_209 b_3 NI_3 NS_209 0 1.9781110397687088e-05
GC_3_210 b_3 NI_3 NS_210 0 -1.0052051305303814e-05
GC_3_211 b_3 NI_3 NS_211 0 -7.0407200288778764e-06
GC_3_212 b_3 NI_3 NS_212 0 3.3239720747350653e-06
GC_3_213 b_3 NI_3 NS_213 0 -2.9707678301838913e-03
GC_3_214 b_3 NI_3 NS_214 0 1.8890857251166596e-03
GC_3_215 b_3 NI_3 NS_215 0 -2.5723518054770062e-04
GC_3_216 b_3 NI_3 NS_216 0 -4.5693203037823016e-04
GC_3_217 b_3 NI_3 NS_217 0 1.0925348306816711e-04
GC_3_218 b_3 NI_3 NS_218 0 -3.1933876293255135e-04
GC_3_219 b_3 NI_3 NS_219 0 -1.7160005617579076e-05
GC_3_220 b_3 NI_3 NS_220 0 1.0940520918402217e-04
GC_3_221 b_3 NI_3 NS_221 0 -1.6800228241282233e-05
GC_3_222 b_3 NI_3 NS_222 0 -1.6651600071906611e-05
GC_3_223 b_3 NI_3 NS_223 0 -2.6023894632015375e-05
GC_3_224 b_3 NI_3 NS_224 0 1.0672966907649938e-05
GC_3_225 b_3 NI_3 NS_225 0 6.7047450895425798e-05
GC_3_226 b_3 NI_3 NS_226 0 1.1878474537778141e-04
GC_3_227 b_3 NI_3 NS_227 0 3.5665740396047320e-05
GC_3_228 b_3 NI_3 NS_228 0 -7.8251457793689218e-06
GC_3_229 b_3 NI_3 NS_229 0 -1.4948017766284372e-02
GC_3_230 b_3 NI_3 NS_230 0 -1.3192713761394793e-03
GC_3_231 b_3 NI_3 NS_231 0 7.3862161179905012e-03
GC_3_232 b_3 NI_3 NS_232 0 1.1632343778996985e-02
GC_3_233 b_3 NI_3 NS_233 0 2.7340006042463852e-04
GC_3_234 b_3 NI_3 NS_234 0 4.0314908824793310e-04
GC_3_235 b_3 NI_3 NS_235 0 1.1059666623179773e-04
GC_3_236 b_3 NI_3 NS_236 0 4.2664863610202207e-05
GC_3_237 b_3 NI_3 NS_237 0 6.4062900599206945e-03
GC_3_238 b_3 NI_3 NS_238 0 3.6842934933914353e-03
GC_3_239 b_3 NI_3 NS_239 0 -1.5916876310250524e-05
GC_3_240 b_3 NI_3 NS_240 0 4.5527931143405005e-06
GC_3_241 b_3 NI_3 NS_241 0 9.7027177669886406e-03
GC_3_242 b_3 NI_3 NS_242 0 -8.5819153170080143e-03
GC_3_243 b_3 NI_3 NS_243 0 4.8955247916163264e-06
GC_3_244 b_3 NI_3 NS_244 0 3.5544419888274422e-05
GC_3_245 b_3 NI_3 NS_245 0 -1.5892054008526519e-05
GC_3_246 b_3 NI_3 NS_246 0 3.3464478089959288e-05
GC_3_247 b_3 NI_3 NS_247 0 3.6536330073564866e-05
GC_3_248 b_3 NI_3 NS_248 0 1.9463727086717439e-05
GC_3_249 b_3 NI_3 NS_249 0 2.2067150694022008e-06
GC_3_250 b_3 NI_3 NS_250 0 8.5370296821321266e-06
GC_3_251 b_3 NI_3 NS_251 0 -2.3718837144697060e-03
GC_3_252 b_3 NI_3 NS_252 0 2.7402844495118118e-03
GC_3_253 b_3 NI_3 NS_253 0 -4.5188458691674009e-04
GC_3_254 b_3 NI_3 NS_254 0 -4.1350548986594815e-04
GC_3_255 b_3 NI_3 NS_255 0 1.8328015060189662e-04
GC_3_256 b_3 NI_3 NS_256 0 -1.5940858077979626e-04
GC_3_257 b_3 NI_3 NS_257 0 2.1629688028155075e-05
GC_3_258 b_3 NI_3 NS_258 0 5.3189190037861575e-05
GC_3_259 b_3 NI_3 NS_259 0 9.8538940677037747e-06
GC_3_260 b_3 NI_3 NS_260 0 1.0981182936876578e-05
GC_3_261 b_3 NI_3 NS_261 0 2.1316943952602712e-06
GC_3_262 b_3 NI_3 NS_262 0 8.8400938155602974e-06
GC_3_263 b_3 NI_3 NS_263 0 4.7644421354593692e-05
GC_3_264 b_3 NI_3 NS_264 0 1.4609958694066851e-05
GC_3_265 b_3 NI_3 NS_265 0 7.0911202418817103e-06
GC_3_266 b_3 NI_3 NS_266 0 1.0019305693948721e-05
GC_3_267 b_3 NI_3 NS_267 0 7.3104217103036918e-03
GC_3_268 b_3 NI_3 NS_268 0 1.3556885265617162e-03
GC_3_269 b_3 NI_3 NS_269 0 -6.4265947678699359e-03
GC_3_270 b_3 NI_3 NS_270 0 2.9715965024843011e-03
GC_3_271 b_3 NI_3 NS_271 0 1.1175177558875330e-04
GC_3_272 b_3 NI_3 NS_272 0 5.3070637155521688e-05
GC_3_273 b_3 NI_3 NS_273 0 4.3956277825056672e-05
GC_3_274 b_3 NI_3 NS_274 0 1.5663055606532026e-05
GC_3_275 b_3 NI_3 NS_275 0 -5.9821366734605858e-03
GC_3_276 b_3 NI_3 NS_276 0 -3.4130491553683593e-03
GC_3_277 b_3 NI_3 NS_277 0 2.3284912115420031e-05
GC_3_278 b_3 NI_3 NS_278 0 -2.9307845829947819e-06
GC_3_279 b_3 NI_3 NS_279 0 9.0967949640132061e-03
GC_3_280 b_3 NI_3 NS_280 0 -4.9039973251783090e-03
GC_3_281 b_3 NI_3 NS_281 0 -4.2591984207099640e-06
GC_3_282 b_3 NI_3 NS_282 0 -6.9905740101868910e-06
GC_3_283 b_3 NI_3 NS_283 0 -1.2409485950598228e-05
GC_3_284 b_3 NI_3 NS_284 0 2.4964446591694486e-05
GC_3_285 b_3 NI_3 NS_285 0 1.6655983009916094e-05
GC_3_286 b_3 NI_3 NS_286 0 1.0331552051605511e-05
GC_3_287 b_3 NI_3 NS_287 0 -1.4970442595091787e-05
GC_3_288 b_3 NI_3 NS_288 0 8.5888361977921238e-06
GC_3_289 b_3 NI_3 NS_289 0 -2.9815518731719343e-03
GC_3_290 b_3 NI_3 NS_290 0 2.3381436983940223e-03
GC_3_291 b_3 NI_3 NS_291 0 -2.4069950423775578e-04
GC_3_292 b_3 NI_3 NS_292 0 -4.0204184320256616e-04
GC_3_293 b_3 NI_3 NS_293 0 2.3789943584122717e-04
GC_3_294 b_3 NI_3 NS_294 0 -8.6088512456372835e-05
GC_3_295 b_3 NI_3 NS_295 0 8.8884883363267850e-06
GC_3_296 b_3 NI_3 NS_296 0 5.1375945636707423e-05
GC_3_297 b_3 NI_3 NS_297 0 -6.7249131821953211e-06
GC_3_298 b_3 NI_3 NS_298 0 6.5463160187938975e-06
GC_3_299 b_3 NI_3 NS_299 0 2.0543311480822612e-06
GC_3_300 b_3 NI_3 NS_300 0 1.1084769599205269e-05
GC_3_301 b_3 NI_3 NS_301 0 4.1187077294028590e-05
GC_3_302 b_3 NI_3 NS_302 0 4.8813604262794629e-05
GC_3_303 b_3 NI_3 NS_303 0 2.7085557451036663e-06
GC_3_304 b_3 NI_3 NS_304 0 8.0924743441852937e-06
GC_3_305 b_3 NI_3 NS_305 0 4.2068036937810182e-03
GC_3_306 b_3 NI_3 NS_306 0 -1.1129306956504492e-03
GC_3_307 b_3 NI_3 NS_307 0 -8.5750552783475896e-03
GC_3_308 b_3 NI_3 NS_308 0 5.7767737563639635e-03
GC_3_309 b_3 NI_3 NS_309 0 6.9631319080159105e-04
GC_3_310 b_3 NI_3 NS_310 0 -2.2696042693939235e-04
GC_3_311 b_3 NI_3 NS_311 0 1.9031237966730098e-04
GC_3_312 b_3 NI_3 NS_312 0 -1.4908496501221010e-04
GC_3_313 b_3 NI_3 NS_313 0 2.5814892054433765e-03
GC_3_314 b_3 NI_3 NS_314 0 -4.7567022160007197e-03
GC_3_315 b_3 NI_3 NS_315 0 -2.0078537943419071e-05
GC_3_316 b_3 NI_3 NS_316 0 3.9966635342827634e-05
GC_3_317 b_3 NI_3 NS_317 0 8.5037799733264658e-03
GC_3_318 b_3 NI_3 NS_318 0 2.2810147627120828e-03
GC_3_319 b_3 NI_3 NS_319 0 -4.9935696308283221e-06
GC_3_320 b_3 NI_3 NS_320 0 -6.8608044681368265e-06
GC_3_321 b_3 NI_3 NS_321 0 -2.8732365987755220e-05
GC_3_322 b_3 NI_3 NS_322 0 4.8234639121804423e-05
GC_3_323 b_3 NI_3 NS_323 0 1.4192797579230530e-04
GC_3_324 b_3 NI_3 NS_324 0 1.0455909756373402e-05
GC_3_325 b_3 NI_3 NS_325 0 4.1046196925288603e-05
GC_3_326 b_3 NI_3 NS_326 0 2.4656114265454384e-05
GC_3_327 b_3 NI_3 NS_327 0 -2.1812877531420085e-03
GC_3_328 b_3 NI_3 NS_328 0 -3.9476920145216008e-04
GC_3_329 b_3 NI_3 NS_329 0 -1.6432094993911963e-04
GC_3_330 b_3 NI_3 NS_330 0 -4.2855393041127182e-04
GC_3_331 b_3 NI_3 NS_331 0 2.7431666799524113e-04
GC_3_332 b_3 NI_3 NS_332 0 1.6459640897784651e-05
GC_3_333 b_3 NI_3 NS_333 0 3.1323472931801677e-06
GC_3_334 b_3 NI_3 NS_334 0 4.9385217175849348e-05
GC_3_335 b_3 NI_3 NS_335 0 -9.3997374082604348e-06
GC_3_336 b_3 NI_3 NS_336 0 -1.9125057791591320e-05
GC_3_337 b_3 NI_3 NS_337 0 -1.6170017475823874e-05
GC_3_338 b_3 NI_3 NS_338 0 2.0283489069341708e-05
GC_3_339 b_3 NI_3 NS_339 0 -4.4479676696203584e-06
GC_3_340 b_3 NI_3 NS_340 0 6.6246351851705624e-05
GC_3_341 b_3 NI_3 NS_341 0 1.9521404550133195e-05
GC_3_342 b_3 NI_3 NS_342 0 8.2199732886348492e-06
GC_3_343 b_3 NI_3 NS_343 0 1.3481328046554159e-02
GC_3_344 b_3 NI_3 NS_344 0 1.1270842129977668e-03
GC_3_345 b_3 NI_3 NS_345 0 -9.5721589624651240e-03
GC_3_346 b_3 NI_3 NS_346 0 1.2007819604415056e-03
GC_3_347 b_3 NI_3 NS_347 0 2.3592480766022224e-04
GC_3_348 b_3 NI_3 NS_348 0 -2.1851919121074870e-04
GC_3_349 b_3 NI_3 NS_349 0 6.7386663253362058e-05
GC_3_350 b_3 NI_3 NS_350 0 -6.1487116857180402e-05
GC_3_351 b_3 NI_3 NS_351 0 -2.0750350794418605e-03
GC_3_352 b_3 NI_3 NS_352 0 5.6028640793807476e-03
GC_3_353 b_3 NI_3 NS_353 0 2.3440942412942161e-05
GC_3_354 b_3 NI_3 NS_354 0 -3.3427809773325065e-05
GC_3_355 b_3 NI_3 NS_355 0 3.6182047877074191e-03
GC_3_356 b_3 NI_3 NS_356 0 4.4649912564169187e-03
GC_3_357 b_3 NI_3 NS_357 0 -1.7556360514813792e-05
GC_3_358 b_3 NI_3 NS_358 0 -9.8179956495864785e-06
GC_3_359 b_3 NI_3 NS_359 0 -2.2334661783348113e-05
GC_3_360 b_3 NI_3 NS_360 0 4.2470990826086385e-05
GC_3_361 b_3 NI_3 NS_361 0 7.6370079295239851e-05
GC_3_362 b_3 NI_3 NS_362 0 -2.4913237405453439e-06
GC_3_363 b_3 NI_3 NS_363 0 3.5651920604191791e-05
GC_3_364 b_3 NI_3 NS_364 0 2.3031375813404204e-05
GC_3_365 b_3 NI_3 NS_365 0 -1.3672004813282065e-03
GC_3_366 b_3 NI_3 NS_366 0 -7.7233658135993088e-04
GC_3_367 b_3 NI_3 NS_367 0 4.7760374525386131e-05
GC_3_368 b_3 NI_3 NS_368 0 -4.3130410095207258e-04
GC_3_369 b_3 NI_3 NS_369 0 1.3790554808191946e-04
GC_3_370 b_3 NI_3 NS_370 0 2.0906214225556120e-05
GC_3_371 b_3 NI_3 NS_371 0 2.5085064784756686e-05
GC_3_372 b_3 NI_3 NS_372 0 4.9385198824265207e-05
GC_3_373 b_3 NI_3 NS_373 0 -6.1958532220649337e-06
GC_3_374 b_3 NI_3 NS_374 0 -3.0095791723437575e-06
GC_3_375 b_3 NI_3 NS_375 0 -1.0205870719126389e-05
GC_3_376 b_3 NI_3 NS_376 0 2.1584018502838159e-05
GC_3_377 b_3 NI_3 NS_377 0 2.8935657045633514e-05
GC_3_378 b_3 NI_3 NS_378 0 3.0485874864880066e-06
GC_3_379 b_3 NI_3 NS_379 0 4.7198241320282562e-06
GC_3_380 b_3 NI_3 NS_380 0 -9.0579207748312065e-06
GC_3_381 b_3 NI_3 NS_381 0 1.7525377343270115e-02
GC_3_382 b_3 NI_3 NS_382 0 -8.1893414815559630e-04
GC_3_383 b_3 NI_3 NS_383 0 -1.4206778699395071e-02
GC_3_384 b_3 NI_3 NS_384 0 2.3392006311431838e-03
GC_3_385 b_3 NI_3 NS_385 0 7.4477722613787087e-04
GC_3_386 b_3 NI_3 NS_386 0 -3.6149687201366288e-04
GC_3_387 b_3 NI_3 NS_387 0 1.8738085918008229e-04
GC_3_388 b_3 NI_3 NS_388 0 -2.1661032666624354e-04
GC_3_389 b_3 NI_3 NS_389 0 -6.6974295438135701e-04
GC_3_390 b_3 NI_3 NS_390 0 -7.4150387757149182e-03
GC_3_391 b_3 NI_3 NS_391 0 -1.8566596287886362e-05
GC_3_392 b_3 NI_3 NS_392 0 3.7166816428163102e-05
GC_3_393 b_3 NI_3 NS_393 0 4.6433006821784070e-03
GC_3_394 b_3 NI_3 NS_394 0 4.4301281856072286e-03
GC_3_395 b_3 NI_3 NS_395 0 2.2013953639515894e-05
GC_3_396 b_3 NI_3 NS_396 0 -4.2412697254144368e-05
GC_3_397 b_3 NI_3 NS_397 0 9.7578150376899501e-06
GC_3_398 b_3 NI_3 NS_398 0 3.8359175161763285e-05
GC_3_399 b_3 NI_3 NS_399 0 1.4627979004854465e-04
GC_3_400 b_3 NI_3 NS_400 0 -6.4987412868448097e-06
GC_3_401 b_3 NI_3 NS_401 0 3.0306555441855254e-05
GC_3_402 b_3 NI_3 NS_402 0 1.7091778218305186e-05
GC_3_403 b_3 NI_3 NS_403 0 -8.3197585136561049e-04
GC_3_404 b_3 NI_3 NS_404 0 -6.9563961115966060e-04
GC_3_405 b_3 NI_3 NS_405 0 -2.3649277676255080e-04
GC_3_406 b_3 NI_3 NS_406 0 -1.4542364418863242e-04
GC_3_407 b_3 NI_3 NS_407 0 2.9862105075121692e-04
GC_3_408 b_3 NI_3 NS_408 0 3.2664844928297543e-04
GC_3_409 b_3 NI_3 NS_409 0 7.2063527462695162e-05
GC_3_410 b_3 NI_3 NS_410 0 -3.4202645749685490e-05
GC_3_411 b_3 NI_3 NS_411 0 -2.0604166123517850e-05
GC_3_412 b_3 NI_3 NS_412 0 -2.6419109265893614e-05
GC_3_413 b_3 NI_3 NS_413 0 -8.1636158091461836e-06
GC_3_414 b_3 NI_3 NS_414 0 3.0365278384817353e-05
GC_3_415 b_3 NI_3 NS_415 0 -4.2276686866260388e-05
GC_3_416 b_3 NI_3 NS_416 0 -1.6526209492136316e-05
GC_3_417 b_3 NI_3 NS_417 0 1.1539291060814884e-06
GC_3_418 b_3 NI_3 NS_418 0 2.4982398010172180e-06
GC_3_419 b_3 NI_3 NS_419 0 7.3339002936033690e-03
GC_3_420 b_3 NI_3 NS_420 0 8.2243802221426340e-04
GC_3_421 b_3 NI_3 NS_421 0 -7.3854133629246170e-03
GC_3_422 b_3 NI_3 NS_422 0 1.6955082414941403e-03
GC_3_423 b_3 NI_3 NS_423 0 1.4765721368394010e-04
GC_3_424 b_3 NI_3 NS_424 0 -9.3134188719072358e-05
GC_3_425 b_3 NI_3 NS_425 0 6.8656667420131343e-05
GC_3_426 b_3 NI_3 NS_426 0 -6.8102334879647321e-05
GC_3_427 b_3 NI_3 NS_427 0 -3.6468522902273395e-04
GC_3_428 b_3 NI_3 NS_428 0 6.6707450435927185e-03
GC_3_429 b_3 NI_3 NS_429 0 2.0794163365064540e-05
GC_3_430 b_3 NI_3 NS_430 0 -3.2738974849129796e-05
GC_3_431 b_3 NI_3 NS_431 0 3.6219183327026398e-03
GC_3_432 b_3 NI_3 NS_432 0 2.6309979245972052e-03
GC_3_433 b_3 NI_3 NS_433 0 4.4586111898706023e-06
GC_3_434 b_3 NI_3 NS_434 0 -2.3074139388097791e-05
GC_3_435 b_3 NI_3 NS_435 0 -2.4885326796411735e-06
GC_3_436 b_3 NI_3 NS_436 0 4.5350783949399271e-05
GC_3_437 b_3 NI_3 NS_437 0 8.7426863685381256e-05
GC_3_438 b_3 NI_3 NS_438 0 6.9923407306235968e-06
GC_3_439 b_3 NI_3 NS_439 0 2.5887689063646546e-05
GC_3_440 b_3 NI_3 NS_440 0 1.9262438384381482e-05
GC_3_441 b_3 NI_3 NS_441 0 -1.2001191538979384e-03
GC_3_442 b_3 NI_3 NS_442 0 -2.2059217680719405e-04
GC_3_443 b_3 NI_3 NS_443 0 1.5451408941152281e-05
GC_3_444 b_3 NI_3 NS_444 0 -3.6371147009630462e-04
GC_3_445 b_3 NI_3 NS_445 0 1.9751354701732102e-04
GC_3_446 b_3 NI_3 NS_446 0 2.3879414573204830e-04
GC_3_447 b_3 NI_3 NS_447 0 6.3161919347452496e-05
GC_3_448 b_3 NI_3 NS_448 0 7.5036489340181022e-06
GC_3_449 b_3 NI_3 NS_449 0 -5.0935499325381707e-06
GC_3_450 b_3 NI_3 NS_450 0 -2.8261365960472175e-05
GC_3_451 b_3 NI_3 NS_451 0 -2.3421894916712890e-05
GC_3_452 b_3 NI_3 NS_452 0 1.8312310269507989e-05
GC_3_453 b_3 NI_3 NS_453 0 -1.4242404113050274e-05
GC_3_454 b_3 NI_3 NS_454 0 -4.4665022531166332e-05
GC_3_455 b_3 NI_3 NS_455 0 -2.1349478536523089e-06
GC_3_456 b_3 NI_3 NS_456 0 -1.4680732568770215e-06
GD_3_1 b_3 NI_3 NA_1 0 -2.6417047654601858e-02
GD_3_2 b_3 NI_3 NA_2 0 5.6273026377701308e-03
GD_3_3 b_3 NI_3 NA_3 0 -7.8088306178392297e-02
GD_3_4 b_3 NI_3 NA_4 0 -3.3552893402017982e-02
GD_3_5 b_3 NI_3 NA_5 0 7.1967619955791277e-05
GD_3_6 b_3 NI_3 NA_6 0 9.4839467656445721e-03
GD_3_7 b_3 NI_3 NA_7 0 -9.2751569968421346e-03
GD_3_8 b_3 NI_3 NA_8 0 -2.1883799587090950e-03
GD_3_9 b_3 NI_3 NA_9 0 -5.1206640902632140e-03
GD_3_10 b_3 NI_3 NA_10 0 -5.0829306474011841e-03
GD_3_11 b_3 NI_3 NA_11 0 -5.8234465193401572e-03
GD_3_12 b_3 NI_3 NA_12 0 -2.6553122869846682e-03
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 4.6919127373847312e-02
GC_4_2 b_4 NI_4 NS_2 0 9.5176128559025899e-04
GC_4_3 b_4 NI_4 NS_3 0 -2.3992666956204868e-02
GC_4_4 b_4 NI_4 NS_4 0 -8.5599133551307743e-03
GC_4_5 b_4 NI_4 NS_5 0 3.3753035542260660e-04
GC_4_6 b_4 NI_4 NS_6 0 2.3559976929710775e-04
GC_4_7 b_4 NI_4 NS_7 0 6.0091679574396042e-05
GC_4_8 b_4 NI_4 NS_8 0 -3.0984343937678305e-05
GC_4_9 b_4 NI_4 NS_9 0 -2.2167639469028982e-02
GC_4_10 b_4 NI_4 NS_10 0 -3.9929711504899879e-02
GC_4_11 b_4 NI_4 NS_11 0 5.7346320174944333e-05
GC_4_12 b_4 NI_4 NS_12 0 8.9687751204336634e-05
GC_4_13 b_4 NI_4 NS_13 0 1.4219187577189801e-02
GC_4_14 b_4 NI_4 NS_14 0 -6.1780281854255043e-03
GC_4_15 b_4 NI_4 NS_15 0 -1.5275074692200343e-05
GC_4_16 b_4 NI_4 NS_16 0 2.5103270749082782e-06
GC_4_17 b_4 NI_4 NS_17 0 -4.3515637965323777e-05
GC_4_18 b_4 NI_4 NS_18 0 2.9767339110445096e-05
GC_4_19 b_4 NI_4 NS_19 0 -4.5494630241995746e-05
GC_4_20 b_4 NI_4 NS_20 0 -6.6942863219384272e-06
GC_4_21 b_4 NI_4 NS_21 0 -8.4994318081807522e-05
GC_4_22 b_4 NI_4 NS_22 0 -2.9800616736493228e-05
GC_4_23 b_4 NI_4 NS_23 0 -7.3287528063583629e-03
GC_4_24 b_4 NI_4 NS_24 0 7.5411413511547835e-03
GC_4_25 b_4 NI_4 NS_25 0 1.2010039973311187e-05
GC_4_26 b_4 NI_4 NS_26 0 -1.1073634674601668e-03
GC_4_27 b_4 NI_4 NS_27 0 3.2173367976664986e-04
GC_4_28 b_4 NI_4 NS_28 0 -7.7206066505325582e-04
GC_4_29 b_4 NI_4 NS_29 0 -1.0166881702227544e-04
GC_4_30 b_4 NI_4 NS_30 0 1.0156219640060589e-04
GC_4_31 b_4 NI_4 NS_31 0 4.1728445253213813e-05
GC_4_32 b_4 NI_4 NS_32 0 2.0461670769346953e-05
GC_4_33 b_4 NI_4 NS_33 0 3.8724779207608156e-05
GC_4_34 b_4 NI_4 NS_34 0 -3.3021069759367554e-05
GC_4_35 b_4 NI_4 NS_35 0 2.7785496594916103e-06
GC_4_36 b_4 NI_4 NS_36 0 5.7339003651090390e-05
GC_4_37 b_4 NI_4 NS_37 0 2.3799277754344639e-06
GC_4_38 b_4 NI_4 NS_38 0 -1.1726083761419066e-05
GC_4_39 b_4 NI_4 NS_39 0 2.7839475463308443e-02
GC_4_40 b_4 NI_4 NS_40 0 -1.3958640395799323e-03
GC_4_41 b_4 NI_4 NS_41 0 -1.8779537642344721e-02
GC_4_42 b_4 NI_4 NS_42 0 1.5397658801355218e-03
GC_4_43 b_4 NI_4 NS_43 0 -1.1059695070343961e-04
GC_4_44 b_4 NI_4 NS_44 0 8.6291017897882681e-06
GC_4_45 b_4 NI_4 NS_45 0 -6.8260359162762682e-05
GC_4_46 b_4 NI_4 NS_46 0 8.9272551414701438e-05
GC_4_47 b_4 NI_4 NS_47 0 5.5133180419014082e-03
GC_4_48 b_4 NI_4 NS_48 0 2.1163950755365288e-02
GC_4_49 b_4 NI_4 NS_49 0 -6.4490927816608076e-05
GC_4_50 b_4 NI_4 NS_50 0 -8.5829429650404929e-05
GC_4_51 b_4 NI_4 NS_51 0 1.2318662983425504e-02
GC_4_52 b_4 NI_4 NS_52 0 2.0639247945742926e-03
GC_4_53 b_4 NI_4 NS_53 0 -4.1395918242371461e-05
GC_4_54 b_4 NI_4 NS_54 0 5.8549107171423182e-05
GC_4_55 b_4 NI_4 NS_55 0 -4.3609242235206579e-05
GC_4_56 b_4 NI_4 NS_56 0 5.0315936712891865e-05
GC_4_57 b_4 NI_4 NS_57 0 1.2457632930921660e-06
GC_4_58 b_4 NI_4 NS_58 0 -6.0421725522354234e-06
GC_4_59 b_4 NI_4 NS_59 0 -1.3967100896159759e-04
GC_4_60 b_4 NI_4 NS_60 0 -3.6579218568410465e-05
GC_4_61 b_4 NI_4 NS_61 0 -7.6746471231996984e-03
GC_4_62 b_4 NI_4 NS_62 0 5.8001420728070359e-03
GC_4_63 b_4 NI_4 NS_63 0 4.3788338047868287e-04
GC_4_64 b_4 NI_4 NS_64 0 -1.0748139498922310e-03
GC_4_65 b_4 NI_4 NS_65 0 4.3543311621031502e-04
GC_4_66 b_4 NI_4 NS_66 0 -7.2211581308820392e-04
GC_4_67 b_4 NI_4 NS_67 0 -1.0783462589033617e-04
GC_4_68 b_4 NI_4 NS_68 0 5.0025721202538719e-05
GC_4_69 b_4 NI_4 NS_69 0 6.2107792484727410e-06
GC_4_70 b_4 NI_4 NS_70 0 4.6958543158612597e-05
GC_4_71 b_4 NI_4 NS_71 0 4.8370292792911104e-05
GC_4_72 b_4 NI_4 NS_72 0 3.9597819339822975e-06
GC_4_73 b_4 NI_4 NS_73 0 -8.2515854531982019e-06
GC_4_74 b_4 NI_4 NS_74 0 5.8699291828585211e-05
GC_4_75 b_4 NI_4 NS_75 0 -4.5289690832266719e-06
GC_4_76 b_4 NI_4 NS_76 0 -1.2264286024171700e-05
GC_4_77 b_4 NI_4 NS_77 0 1.5561535113461153e-02
GC_4_78 b_4 NI_4 NS_78 0 2.3525586844203232e-03
GC_4_79 b_4 NI_4 NS_79 0 2.2368779242911044e-02
GC_4_80 b_4 NI_4 NS_80 0 -1.2322543112868404e-02
GC_4_81 b_4 NI_4 NS_81 0 1.6215823412790175e-03
GC_4_82 b_4 NI_4 NS_82 0 -2.7839373382255668e-06
GC_4_83 b_4 NI_4 NS_83 0 1.3580162328290509e-04
GC_4_84 b_4 NI_4 NS_84 0 -7.5901001688784045e-05
GC_4_85 b_4 NI_4 NS_85 0 2.6760656876423306e-02
GC_4_86 b_4 NI_4 NS_86 0 6.1410744770937341e-03
GC_4_87 b_4 NI_4 NS_87 0 8.6757846627514971e-05
GC_4_88 b_4 NI_4 NS_88 0 8.8881550163818303e-05
GC_4_89 b_4 NI_4 NS_89 0 -3.9846440159693200e-02
GC_4_90 b_4 NI_4 NS_90 0 3.2317970201151014e-02
GC_4_91 b_4 NI_4 NS_91 0 2.2692020679981069e-05
GC_4_92 b_4 NI_4 NS_92 0 -1.3835406684620439e-05
GC_4_93 b_4 NI_4 NS_93 0 -1.4139593307438484e-05
GC_4_94 b_4 NI_4 NS_94 0 4.7843999159320008e-05
GC_4_95 b_4 NI_4 NS_95 0 -3.9590794883970337e-05
GC_4_96 b_4 NI_4 NS_96 0 -1.4242202553660717e-06
GC_4_97 b_4 NI_4 NS_97 0 -7.7823797377817762e-05
GC_4_98 b_4 NI_4 NS_98 0 -1.2126538347049535e-05
GC_4_99 b_4 NI_4 NS_99 0 -4.4817679341380189e-03
GC_4_100 b_4 NI_4 NS_100 0 6.3339902679701110e-04
GC_4_101 b_4 NI_4 NS_101 0 6.5591687505585261e-05
GC_4_102 b_4 NI_4 NS_102 0 -6.1039377259711636e-04
GC_4_103 b_4 NI_4 NS_103 0 2.0984265486842117e-04
GC_4_104 b_4 NI_4 NS_104 0 -2.0542007757407230e-04
GC_4_105 b_4 NI_4 NS_105 0 -4.4169702476647744e-05
GC_4_106 b_4 NI_4 NS_106 0 9.9931131039498984e-05
GC_4_107 b_4 NI_4 NS_107 0 2.7338247364133861e-05
GC_4_108 b_4 NI_4 NS_108 0 -7.2668200941554158e-08
GC_4_109 b_4 NI_4 NS_109 0 8.5939849745777291e-06
GC_4_110 b_4 NI_4 NS_110 0 1.9876655237163336e-05
GC_4_111 b_4 NI_4 NS_111 0 -1.3005229628870387e-05
GC_4_112 b_4 NI_4 NS_112 0 8.9885364093955856e-05
GC_4_113 b_4 NI_4 NS_113 0 1.9837254252271187e-05
GC_4_114 b_4 NI_4 NS_114 0 6.9971855102738481e-06
GC_4_115 b_4 NI_4 NS_115 0 9.8043580091702220e-02
GC_4_116 b_4 NI_4 NS_116 0 -1.8367183290063664e-03
GC_4_117 b_4 NI_4 NS_117 0 1.7955814645363864e-02
GC_4_118 b_4 NI_4 NS_118 0 -5.0948487344290791e-02
GC_4_119 b_4 NI_4 NS_119 0 -3.5626000233128638e-04
GC_4_120 b_4 NI_4 NS_120 0 -3.8658160975358491e-04
GC_4_121 b_4 NI_4 NS_121 0 -1.2125382946232493e-04
GC_4_122 b_4 NI_4 NS_122 0 1.0423694285421428e-04
GC_4_123 b_4 NI_4 NS_123 0 -1.1845690340497204e-02
GC_4_124 b_4 NI_4 NS_124 0 1.1394038466349536e-02
GC_4_125 b_4 NI_4 NS_125 0 -6.6531804575227084e-05
GC_4_126 b_4 NI_4 NS_126 0 -8.1262271817991044e-05
GC_4_127 b_4 NI_4 NS_127 0 -2.1831485901718739e-02
GC_4_128 b_4 NI_4 NS_128 0 1.8158037338174369e-02
GC_4_129 b_4 NI_4 NS_129 0 -1.4925618919911080e-05
GC_4_130 b_4 NI_4 NS_130 0 6.4038151234227574e-05
GC_4_131 b_4 NI_4 NS_131 0 -4.8318541948246338e-05
GC_4_132 b_4 NI_4 NS_132 0 5.1152942071440491e-05
GC_4_133 b_4 NI_4 NS_133 0 -2.1538275200022546e-05
GC_4_134 b_4 NI_4 NS_134 0 -2.0205282511321205e-05
GC_4_135 b_4 NI_4 NS_135 0 -1.4276655566447988e-04
GC_4_136 b_4 NI_4 NS_136 0 -2.5701107182892560e-05
GC_4_137 b_4 NI_4 NS_137 0 -7.2370446538658527e-03
GC_4_138 b_4 NI_4 NS_138 0 2.5292978300149871e-03
GC_4_139 b_4 NI_4 NS_139 0 5.2572408516181714e-04
GC_4_140 b_4 NI_4 NS_140 0 -8.3116327662294341e-04
GC_4_141 b_4 NI_4 NS_141 0 5.3798034793098499e-04
GC_4_142 b_4 NI_4 NS_142 0 -3.8037564501477099e-04
GC_4_143 b_4 NI_4 NS_143 0 -1.0008261595386718e-04
GC_4_144 b_4 NI_4 NS_144 0 6.7176725037724745e-06
GC_4_145 b_4 NI_4 NS_145 0 2.4910935670555588e-06
GC_4_146 b_4 NI_4 NS_146 0 2.4027297197282188e-05
GC_4_147 b_4 NI_4 NS_147 0 1.4812397001371312e-05
GC_4_148 b_4 NI_4 NS_148 0 -3.1049215823952830e-06
GC_4_149 b_4 NI_4 NS_149 0 3.3478373711044112e-07
GC_4_150 b_4 NI_4 NS_150 0 3.9957266258935144e-05
GC_4_151 b_4 NI_4 NS_151 0 2.2818741462120951e-06
GC_4_152 b_4 NI_4 NS_152 0 8.9896796379643049e-07
GC_4_153 b_4 NI_4 NS_153 0 -2.0035670469729271e-02
GC_4_154 b_4 NI_4 NS_154 0 1.4593307372057357e-03
GC_4_155 b_4 NI_4 NS_155 0 1.0614493483473332e-02
GC_4_156 b_4 NI_4 NS_156 0 5.6714270219198996e-03
GC_4_157 b_4 NI_4 NS_157 0 1.2764118262547649e-04
GC_4_158 b_4 NI_4 NS_158 0 -2.6431000337993595e-04
GC_4_159 b_4 NI_4 NS_159 0 1.2508782086370244e-05
GC_4_160 b_4 NI_4 NS_160 0 -5.4172026598897153e-05
GC_4_161 b_4 NI_4 NS_161 0 -7.2699213836575766e-03
GC_4_162 b_4 NI_4 NS_162 0 -1.1536139719330056e-02
GC_4_163 b_4 NI_4 NS_163 0 3.0182592421165198e-05
GC_4_164 b_4 NI_4 NS_164 0 2.1998449675091230e-06
GC_4_165 b_4 NI_4 NS_165 0 1.2426228602227633e-02
GC_4_166 b_4 NI_4 NS_166 0 -1.3289797349668519e-02
GC_4_167 b_4 NI_4 NS_167 0 2.0653160871448705e-06
GC_4_168 b_4 NI_4 NS_168 0 -3.3527094974695920e-05
GC_4_169 b_4 NI_4 NS_169 0 -1.6132441297694090e-05
GC_4_170 b_4 NI_4 NS_170 0 5.6883239251661415e-05
GC_4_171 b_4 NI_4 NS_171 0 1.1337735981200587e-05
GC_4_172 b_4 NI_4 NS_172 0 1.4504949532664673e-05
GC_4_173 b_4 NI_4 NS_173 0 1.7896341490689035e-05
GC_4_174 b_4 NI_4 NS_174 0 1.5775395738684515e-06
GC_4_175 b_4 NI_4 NS_175 0 -5.6019377053605620e-03
GC_4_176 b_4 NI_4 NS_176 0 2.4609818413827422e-03
GC_4_177 b_4 NI_4 NS_177 0 -1.3607005632946824e-05
GC_4_178 b_4 NI_4 NS_178 0 -9.6373545753760596e-04
GC_4_179 b_4 NI_4 NS_179 0 3.4062317337936850e-04
GC_4_180 b_4 NI_4 NS_180 0 -5.2564405498662314e-04
GC_4_181 b_4 NI_4 NS_181 0 -9.1034649259009602e-05
GC_4_182 b_4 NI_4 NS_182 0 1.0867439092676586e-04
GC_4_183 b_4 NI_4 NS_183 0 -2.0153398784339018e-05
GC_4_184 b_4 NI_4 NS_184 0 3.2347234607583745e-06
GC_4_185 b_4 NI_4 NS_185 0 -7.8511747159023816e-06
GC_4_186 b_4 NI_4 NS_186 0 3.7488165521422805e-05
GC_4_187 b_4 NI_4 NS_187 0 3.6430057801658379e-05
GC_4_188 b_4 NI_4 NS_188 0 9.8694386645948915e-05
GC_4_189 b_4 NI_4 NS_189 0 2.4461548192623889e-05
GC_4_190 b_4 NI_4 NS_190 0 1.0555730541233868e-05
GC_4_191 b_4 NI_4 NS_191 0 -1.2534824971609012e-02
GC_4_192 b_4 NI_4 NS_192 0 -1.4706205380383196e-03
GC_4_193 b_4 NI_4 NS_193 0 7.0059989811682944e-03
GC_4_194 b_4 NI_4 NS_194 0 2.7492836220017899e-02
GC_4_195 b_4 NI_4 NS_195 0 -1.6242137895639691e-04
GC_4_196 b_4 NI_4 NS_196 0 1.8915911459731530e-04
GC_4_197 b_4 NI_4 NS_197 0 -4.6484458819859653e-05
GC_4_198 b_4 NI_4 NS_198 0 8.3393055467316869e-06
GC_4_199 b_4 NI_4 NS_199 0 7.3644626241614192e-03
GC_4_200 b_4 NI_4 NS_200 0 1.0677150415539795e-02
GC_4_201 b_4 NI_4 NS_201 0 -3.0034943539550572e-05
GC_4_202 b_4 NI_4 NS_202 0 -2.0695110074233992e-06
GC_4_203 b_4 NI_4 NS_203 0 1.6169394045068879e-02
GC_4_204 b_4 NI_4 NS_204 0 -1.6385215542641943e-02
GC_4_205 b_4 NI_4 NS_205 0 -4.0272626007263166e-06
GC_4_206 b_4 NI_4 NS_206 0 1.3209470123038189e-05
GC_4_207 b_4 NI_4 NS_207 0 -2.0938316090952148e-05
GC_4_208 b_4 NI_4 NS_208 0 3.0007504226957177e-05
GC_4_209 b_4 NI_4 NS_209 0 1.5415374377871610e-05
GC_4_210 b_4 NI_4 NS_210 0 -3.3136325377485663e-06
GC_4_211 b_4 NI_4 NS_211 0 -1.2480182453756805e-05
GC_4_212 b_4 NI_4 NS_212 0 7.0579895032194905e-06
GC_4_213 b_4 NI_4 NS_213 0 -4.4794724676983930e-03
GC_4_214 b_4 NI_4 NS_214 0 2.4824772529016669e-03
GC_4_215 b_4 NI_4 NS_215 0 2.3593440684799642e-05
GC_4_216 b_4 NI_4 NS_216 0 -7.3604910781945119e-04
GC_4_217 b_4 NI_4 NS_217 0 3.2318711253247748e-04
GC_4_218 b_4 NI_4 NS_218 0 -4.2596650881757142e-04
GC_4_219 b_4 NI_4 NS_219 0 -7.6483039520775100e-05
GC_4_220 b_4 NI_4 NS_220 0 6.3434746411563758e-05
GC_4_221 b_4 NI_4 NS_221 0 6.4447379048771329e-06
GC_4_222 b_4 NI_4 NS_222 0 -3.1301308876755557e-05
GC_4_223 b_4 NI_4 NS_223 0 -1.9256528925134617e-05
GC_4_224 b_4 NI_4 NS_224 0 -9.9542971839817198e-06
GC_4_225 b_4 NI_4 NS_225 0 3.1384183995652512e-05
GC_4_226 b_4 NI_4 NS_226 0 9.2400992443839033e-05
GC_4_227 b_4 NI_4 NS_227 0 6.8903114826811804e-06
GC_4_228 b_4 NI_4 NS_228 0 1.2902967411347314e-05
GC_4_229 b_4 NI_4 NS_229 0 1.9130359166861562e-02
GC_4_230 b_4 NI_4 NS_230 0 1.3328305569640852e-03
GC_4_231 b_4 NI_4 NS_231 0 -1.3763866685470675e-02
GC_4_232 b_4 NI_4 NS_232 0 6.4266279069840407e-03
GC_4_233 b_4 NI_4 NS_233 0 -3.0887858368990517e-04
GC_4_234 b_4 NI_4 NS_234 0 -7.8654110272255624e-05
GC_4_235 b_4 NI_4 NS_235 0 -1.5354420210778312e-05
GC_4_236 b_4 NI_4 NS_236 0 4.3643102468817935e-06
GC_4_237 b_4 NI_4 NS_237 0 -4.6960859607423329e-03
GC_4_238 b_4 NI_4 NS_238 0 -9.2005629073209187e-04
GC_4_239 b_4 NI_4 NS_239 0 1.8350415813166972e-05
GC_4_240 b_4 NI_4 NS_240 0 -1.1971018778149051e-06
GC_4_241 b_4 NI_4 NS_241 0 1.1931221008111483e-02
GC_4_242 b_4 NI_4 NS_242 0 9.1680587288840937e-04
GC_4_243 b_4 NI_4 NS_243 0 -5.8841228751965271e-06
GC_4_244 b_4 NI_4 NS_244 0 -1.2517919957750394e-05
GC_4_245 b_4 NI_4 NS_245 0 -5.3815079433978825e-06
GC_4_246 b_4 NI_4 NS_246 0 4.8503016863926067e-05
GC_4_247 b_4 NI_4 NS_247 0 1.9597962587899650e-05
GC_4_248 b_4 NI_4 NS_248 0 1.8926779670178877e-05
GC_4_249 b_4 NI_4 NS_249 0 6.6641883469380487e-06
GC_4_250 b_4 NI_4 NS_250 0 1.6179055606982627e-05
GC_4_251 b_4 NI_4 NS_251 0 -3.7345114169495706e-03
GC_4_252 b_4 NI_4 NS_252 0 1.7252111619755013e-03
GC_4_253 b_4 NI_4 NS_253 0 -1.0800770270966602e-04
GC_4_254 b_4 NI_4 NS_254 0 -6.4700242367403307e-04
GC_4_255 b_4 NI_4 NS_255 0 3.6371088684654515e-04
GC_4_256 b_4 NI_4 NS_256 0 -1.9916813687558265e-04
GC_4_257 b_4 NI_4 NS_257 0 -1.4364771327033621e-05
GC_4_258 b_4 NI_4 NS_258 0 3.8404787527145181e-05
GC_4_259 b_4 NI_4 NS_259 0 4.2524663475881360e-06
GC_4_260 b_4 NI_4 NS_260 0 3.7457259807944993e-06
GC_4_261 b_4 NI_4 NS_261 0 1.6994719530176405e-06
GC_4_262 b_4 NI_4 NS_262 0 1.2189476331216937e-05
GC_4_263 b_4 NI_4 NS_263 0 5.0773367030474986e-05
GC_4_264 b_4 NI_4 NS_264 0 1.6475193085531410e-05
GC_4_265 b_4 NI_4 NS_265 0 1.9251367005941875e-05
GC_4_266 b_4 NI_4 NS_266 0 -5.1456149593696851e-06
GC_4_267 b_4 NI_4 NS_267 0 -5.0911851467856401e-04
GC_4_268 b_4 NI_4 NS_268 0 -1.3150661066003268e-03
GC_4_269 b_4 NI_4 NS_269 0 -7.4775209488115646e-03
GC_4_270 b_4 NI_4 NS_270 0 8.3599321011363949e-03
GC_4_271 b_4 NI_4 NS_271 0 -3.8139728648420845e-05
GC_4_272 b_4 NI_4 NS_272 0 -1.0974052103016518e-04
GC_4_273 b_4 NI_4 NS_273 0 -7.0940489324140880e-05
GC_4_274 b_4 NI_4 NS_274 0 2.3385953009516426e-05
GC_4_275 b_4 NI_4 NS_275 0 5.1211658790088288e-03
GC_4_276 b_4 NI_4 NS_276 0 2.8106007916322007e-03
GC_4_277 b_4 NI_4 NS_277 0 -2.0552463019362003e-05
GC_4_278 b_4 NI_4 NS_278 0 3.4759025367565706e-06
GC_4_279 b_4 NI_4 NS_279 0 1.3221020690775772e-02
GC_4_280 b_4 NI_4 NS_280 0 -1.5087973317154991e-03
GC_4_281 b_4 NI_4 NS_281 0 7.1085394267377465e-06
GC_4_282 b_4 NI_4 NS_282 0 2.1873811424425415e-05
GC_4_283 b_4 NI_4 NS_283 0 -1.8966277065103165e-05
GC_4_284 b_4 NI_4 NS_284 0 2.6956884359927100e-05
GC_4_285 b_4 NI_4 NS_285 0 7.8609016108513716e-06
GC_4_286 b_4 NI_4 NS_286 0 6.4804586560800370e-06
GC_4_287 b_4 NI_4 NS_287 0 -2.6456423642127941e-05
GC_4_288 b_4 NI_4 NS_288 0 1.7036421850240315e-05
GC_4_289 b_4 NI_4 NS_289 0 -4.3092817223783549e-03
GC_4_290 b_4 NI_4 NS_290 0 1.8529488361891445e-03
GC_4_291 b_4 NI_4 NS_291 0 5.7629121689363948e-05
GC_4_292 b_4 NI_4 NS_292 0 -5.4673622385314612e-04
GC_4_293 b_4 NI_4 NS_293 0 4.2508607862702083e-04
GC_4_294 b_4 NI_4 NS_294 0 -1.1110195524313521e-04
GC_4_295 b_4 NI_4 NS_295 0 -2.5197959201782553e-05
GC_4_296 b_4 NI_4 NS_296 0 1.6542407805451387e-05
GC_4_297 b_4 NI_4 NS_297 0 -2.0510479226684266e-06
GC_4_298 b_4 NI_4 NS_298 0 3.3908260639912644e-06
GC_4_299 b_4 NI_4 NS_299 0 -5.3559763722397920e-06
GC_4_300 b_4 NI_4 NS_300 0 3.9830858152951054e-06
GC_4_301 b_4 NI_4 NS_301 0 4.4739359821733816e-05
GC_4_302 b_4 NI_4 NS_302 0 4.1455587144330194e-05
GC_4_303 b_4 NI_4 NS_303 0 1.4547330729881639e-05
GC_4_304 b_4 NI_4 NS_304 0 3.0054277005848408e-06
GC_4_305 b_4 NI_4 NS_305 0 7.1472150851992836e-03
GC_4_306 b_4 NI_4 NS_306 0 1.1225186662247957e-03
GC_4_307 b_4 NI_4 NS_307 0 -5.9685683038411498e-03
GC_4_308 b_4 NI_4 NS_308 0 -5.5599321762797686e-03
GC_4_309 b_4 NI_4 NS_309 0 3.1555631237049168e-05
GC_4_310 b_4 NI_4 NS_310 0 5.9865779209178783e-04
GC_4_311 b_4 NI_4 NS_311 0 9.9759941213428530e-05
GC_4_312 b_4 NI_4 NS_312 0 1.6334924121177700e-04
GC_4_313 b_4 NI_4 NS_313 0 -1.7806242108917274e-03
GC_4_314 b_4 NI_4 NS_314 0 5.9238112962446089e-03
GC_4_315 b_4 NI_4 NS_315 0 2.3591994345211412e-05
GC_4_316 b_4 NI_4 NS_316 0 -3.1794463558692192e-05
GC_4_317 b_4 NI_4 NS_317 0 3.0199869153953733e-03
GC_4_318 b_4 NI_4 NS_318 0 6.4399065245807343e-03
GC_4_319 b_4 NI_4 NS_319 0 5.2755118938959639e-05
GC_4_320 b_4 NI_4 NS_320 0 3.7785189041957657e-05
GC_4_321 b_4 NI_4 NS_321 0 -9.9972050366250254e-06
GC_4_322 b_4 NI_4 NS_322 0 8.0791512556076202e-05
GC_4_323 b_4 NI_4 NS_323 0 7.8379289960351888e-05
GC_4_324 b_4 NI_4 NS_324 0 4.6936558466998651e-05
GC_4_325 b_4 NI_4 NS_325 0 7.5986280731443070e-05
GC_4_326 b_4 NI_4 NS_326 0 4.3037383680433549e-05
GC_4_327 b_4 NI_4 NS_327 0 -2.5617263524957260e-03
GC_4_328 b_4 NI_4 NS_328 0 -1.1726539335751138e-03
GC_4_329 b_4 NI_4 NS_329 0 2.3700157428163378e-04
GC_4_330 b_4 NI_4 NS_330 0 -5.3062440631404409e-04
GC_4_331 b_4 NI_4 NS_331 0 4.1876568704281254e-04
GC_4_332 b_4 NI_4 NS_332 0 1.5535740294293775e-05
GC_4_333 b_4 NI_4 NS_333 0 -2.5761398422320329e-05
GC_4_334 b_4 NI_4 NS_334 0 2.0424411724927748e-05
GC_4_335 b_4 NI_4 NS_335 0 4.6496891432508097e-06
GC_4_336 b_4 NI_4 NS_336 0 -2.3589851182262126e-05
GC_4_337 b_4 NI_4 NS_337 0 -2.3101857116910918e-05
GC_4_338 b_4 NI_4 NS_338 0 7.3311628752537926e-06
GC_4_339 b_4 NI_4 NS_339 0 -1.2044539605439503e-05
GC_4_340 b_4 NI_4 NS_340 0 4.6556743356284547e-05
GC_4_341 b_4 NI_4 NS_341 0 7.2528852563680345e-06
GC_4_342 b_4 NI_4 NS_342 0 7.5927200224405962e-06
GC_4_343 b_4 NI_4 NS_343 0 9.8336321653813320e-03
GC_4_344 b_4 NI_4 NS_344 0 -1.1184869009313318e-03
GC_4_345 b_4 NI_4 NS_345 0 -8.9642364590077090e-03
GC_4_346 b_4 NI_4 NS_346 0 -2.7023361803908169e-03
GC_4_347 b_4 NI_4 NS_347 0 1.4215319858091851e-04
GC_4_348 b_4 NI_4 NS_348 0 1.7288217914313480e-04
GC_4_349 b_4 NI_4 NS_349 0 4.9934645038850926e-05
GC_4_350 b_4 NI_4 NS_350 0 9.8026996190157437e-05
GC_4_351 b_4 NI_4 NS_351 0 8.0738604502419531e-04
GC_4_352 b_4 NI_4 NS_352 0 -6.7270844052737663e-03
GC_4_353 b_4 NI_4 NS_353 0 -2.5664904564046002e-05
GC_4_354 b_4 NI_4 NS_354 0 2.8406610907864808e-05
GC_4_355 b_4 NI_4 NS_355 0 4.4520290119373874e-03
GC_4_356 b_4 NI_4 NS_356 0 6.7709037688819581e-03
GC_4_357 b_4 NI_4 NS_357 0 5.8580230428704517e-05
GC_4_358 b_4 NI_4 NS_358 0 2.6942073968152455e-05
GC_4_359 b_4 NI_4 NS_359 0 -1.7983154095332710e-05
GC_4_360 b_4 NI_4 NS_360 0 5.9731569334913837e-05
GC_4_361 b_4 NI_4 NS_361 0 4.6612506329265923e-05
GC_4_362 b_4 NI_4 NS_362 0 2.1553341635066680e-05
GC_4_363 b_4 NI_4 NS_363 0 6.5181178097810816e-05
GC_4_364 b_4 NI_4 NS_364 0 4.0000024227891676e-05
GC_4_365 b_4 NI_4 NS_365 0 -2.5410391417517299e-03
GC_4_366 b_4 NI_4 NS_366 0 -8.8531441627227837e-04
GC_4_367 b_4 NI_4 NS_367 0 3.9371123602443457e-04
GC_4_368 b_4 NI_4 NS_368 0 -5.3416580537802107e-04
GC_4_369 b_4 NI_4 NS_369 0 3.0599247685533652e-04
GC_4_370 b_4 NI_4 NS_370 0 -6.9971817136506068e-05
GC_4_371 b_4 NI_4 NS_371 0 -1.5587966367397177e-05
GC_4_372 b_4 NI_4 NS_372 0 1.8615201994975526e-05
GC_4_373 b_4 NI_4 NS_373 0 -1.0442488319560312e-05
GC_4_374 b_4 NI_4 NS_374 0 -8.9638509501228088e-06
GC_4_375 b_4 NI_4 NS_375 0 -2.0186857436072775e-05
GC_4_376 b_4 NI_4 NS_376 0 5.7590465644353844e-06
GC_4_377 b_4 NI_4 NS_377 0 2.4797825657315856e-05
GC_4_378 b_4 NI_4 NS_378 0 -3.3068032826975199e-06
GC_4_379 b_4 NI_4 NS_379 0 4.5253060894046565e-06
GC_4_380 b_4 NI_4 NS_380 0 6.8548358867702993e-06
GC_4_381 b_4 NI_4 NS_381 0 3.3126580564993712e-03
GC_4_382 b_4 NI_4 NS_382 0 7.6895886508722292e-04
GC_4_383 b_4 NI_4 NS_383 0 -4.0804260401456332e-03
GC_4_384 b_4 NI_4 NS_384 0 -4.7421793880034974e-03
GC_4_385 b_4 NI_4 NS_385 0 1.2052536297039802e-04
GC_4_386 b_4 NI_4 NS_386 0 4.2767871864461617e-04
GC_4_387 b_4 NI_4 NS_387 0 7.2140366031770375e-05
GC_4_388 b_4 NI_4 NS_388 0 1.5686264324504281e-04
GC_4_389 b_4 NI_4 NS_389 0 -7.2547612127391297e-04
GC_4_390 b_4 NI_4 NS_390 0 5.5616551947612431e-03
GC_4_391 b_4 NI_4 NS_391 0 1.9791493396002807e-05
GC_4_392 b_4 NI_4 NS_392 0 -3.1303820293091504e-05
GC_4_393 b_4 NI_4 NS_393 0 1.0265404969344262e-03
GC_4_394 b_4 NI_4 NS_394 0 4.0272092022370486e-03
GC_4_395 b_4 NI_4 NS_395 0 4.0325300129274763e-05
GC_4_396 b_4 NI_4 NS_396 0 6.4029914807755555e-05
GC_4_397 b_4 NI_4 NS_397 0 2.0007417484900495e-05
GC_4_398 b_4 NI_4 NS_398 0 3.5171255456699630e-05
GC_4_399 b_4 NI_4 NS_399 0 8.1185152423089588e-05
GC_4_400 b_4 NI_4 NS_400 0 3.3200216653401512e-05
GC_4_401 b_4 NI_4 NS_401 0 5.8665202487005904e-05
GC_4_402 b_4 NI_4 NS_402 0 2.8730280484681946e-05
GC_4_403 b_4 NI_4 NS_403 0 -1.1141916443758568e-03
GC_4_404 b_4 NI_4 NS_404 0 -6.3143374115006258e-04
GC_4_405 b_4 NI_4 NS_405 0 7.1121207277703167e-06
GC_4_406 b_4 NI_4 NS_406 0 -2.8415384159584194e-04
GC_4_407 b_4 NI_4 NS_407 0 3.5994503781373036e-04
GC_4_408 b_4 NI_4 NS_408 0 2.2121722074209938e-04
GC_4_409 b_4 NI_4 NS_409 0 4.4364865662524394e-05
GC_4_410 b_4 NI_4 NS_410 0 -3.9892007488008156e-05
GC_4_411 b_4 NI_4 NS_411 0 -1.1723747284862296e-05
GC_4_412 b_4 NI_4 NS_412 0 -2.6256864935517516e-05
GC_4_413 b_4 NI_4 NS_413 0 -3.0778159430076734e-05
GC_4_414 b_4 NI_4 NS_414 0 1.5045833997344051e-05
GC_4_415 b_4 NI_4 NS_415 0 -3.4281907276244604e-05
GC_4_416 b_4 NI_4 NS_416 0 -3.5248830760730619e-05
GC_4_417 b_4 NI_4 NS_417 0 -1.7825890530566488e-06
GC_4_418 b_4 NI_4 NS_418 0 2.4531373826550789e-06
GC_4_419 b_4 NI_4 NS_419 0 1.7604561611477318e-02
GC_4_420 b_4 NI_4 NS_420 0 -8.5633053374368020e-04
GC_4_421 b_4 NI_4 NS_421 0 -1.2299225185066182e-02
GC_4_422 b_4 NI_4 NS_422 0 -4.1211586009423859e-03
GC_4_423 b_4 NI_4 NS_423 0 2.8176433330138204e-04
GC_4_424 b_4 NI_4 NS_424 0 3.6195172054022825e-06
GC_4_425 b_4 NI_4 NS_425 0 4.2441195419836321e-05
GC_4_426 b_4 NI_4 NS_426 0 8.1711280744908309e-05
GC_4_427 b_4 NI_4 NS_427 0 -1.4405655414025491e-03
GC_4_428 b_4 NI_4 NS_428 0 -8.7482324247992720e-03
GC_4_429 b_4 NI_4 NS_429 0 -2.3899059120750954e-05
GC_4_430 b_4 NI_4 NS_430 0 2.6164874676344089e-05
GC_4_431 b_4 NI_4 NS_431 0 3.3222408043386618e-03
GC_4_432 b_4 NI_4 NS_432 0 7.6831006887890648e-03
GC_4_433 b_4 NI_4 NS_433 0 5.0517566270597170e-05
GC_4_434 b_4 NI_4 NS_434 0 3.7503027517118321e-05
GC_4_435 b_4 NI_4 NS_435 0 5.7796799496596912e-06
GC_4_436 b_4 NI_4 NS_436 0 3.3711667839095640e-05
GC_4_437 b_4 NI_4 NS_437 0 4.9011863328642214e-05
GC_4_438 b_4 NI_4 NS_438 0 2.3614345214009293e-05
GC_4_439 b_4 NI_4 NS_439 0 5.0474990901939018e-05
GC_4_440 b_4 NI_4 NS_440 0 3.4328939939131784e-05
GC_4_441 b_4 NI_4 NS_441 0 -2.4659189725312215e-03
GC_4_442 b_4 NI_4 NS_442 0 -9.0314464321207977e-04
GC_4_443 b_4 NI_4 NS_443 0 3.9476995679493072e-04
GC_4_444 b_4 NI_4 NS_444 0 -4.2264569727751066e-04
GC_4_445 b_4 NI_4 NS_445 0 3.9089256950085863e-04
GC_4_446 b_4 NI_4 NS_446 0 1.3971471141324966e-04
GC_4_447 b_4 NI_4 NS_447 0 2.7987697142160299e-05
GC_4_448 b_4 NI_4 NS_448 0 -2.7292501782942819e-05
GC_4_449 b_4 NI_4 NS_449 0 -1.9097389732225489e-06
GC_4_450 b_4 NI_4 NS_450 0 -2.3373059358173929e-05
GC_4_451 b_4 NI_4 NS_451 0 -3.4922858381742214e-05
GC_4_452 b_4 NI_4 NS_452 0 -1.2539818387071247e-05
GC_4_453 b_4 NI_4 NS_453 0 1.0813713335780564e-06
GC_4_454 b_4 NI_4 NS_454 0 -6.3106678387416515e-05
GC_4_455 b_4 NI_4 NS_455 0 -1.0039102459864398e-05
GC_4_456 b_4 NI_4 NS_456 0 1.9683235781641156e-06
GD_4_1 b_4 NI_4 NA_1 0 -5.6186933756573109e-03
GD_4_2 b_4 NI_4 NA_2 0 -1.2288969999712913e-02
GD_4_3 b_4 NI_4 NA_3 0 -3.3552874461844677e-02
GD_4_4 b_4 NI_4 NA_4 0 -1.3769270927850905e-01
GD_4_5 b_4 NI_4 NA_5 0 6.4943145781561030e-03
GD_4_6 b_4 NI_4 NA_6 0 -9.2660573097538626e-03
GD_4_7 b_4 NI_4 NA_7 0 -8.9590849593405852e-03
GD_4_8 b_4 NI_4 NA_8 0 -4.7772772154668214e-03
GD_4_9 b_4 NI_4 NA_9 0 -1.8005646268776751e-03
GD_4_10 b_4 NI_4 NA_10 0 -2.8725201887023926e-03
GD_4_11 b_4 NI_4 NA_11 0 3.3123630071309413e-04
GD_4_12 b_4 NI_4 NA_12 0 -3.7050046791482446e-03
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 -3.2188609940924165e-02
GC_5_2 b_5 NI_5 NS_2 0 -1.1241411422738617e-03
GC_5_3 b_5 NI_5 NS_3 0 1.4244074681588533e-02
GC_5_4 b_5 NI_5 NS_4 0 1.8916722587216793e-02
GC_5_5 b_5 NI_5 NS_5 0 1.9076761456581848e-04
GC_5_6 b_5 NI_5 NS_6 0 3.5707262347837249e-06
GC_5_7 b_5 NI_5 NS_7 0 -9.0201031552596364e-05
GC_5_8 b_5 NI_5 NS_8 0 1.0889426335286105e-04
GC_5_9 b_5 NI_5 NS_9 0 9.8052259639964268e-03
GC_5_10 b_5 NI_5 NS_10 0 1.0291639721377657e-02
GC_5_11 b_5 NI_5 NS_11 0 -2.7827964707820751e-05
GC_5_12 b_5 NI_5 NS_12 0 1.8957671828089657e-06
GC_5_13 b_5 NI_5 NS_13 0 1.4131979803259044e-02
GC_5_14 b_5 NI_5 NS_14 0 -1.5303989922202853e-02
GC_5_15 b_5 NI_5 NS_15 0 -1.0284019776289655e-05
GC_5_16 b_5 NI_5 NS_16 0 2.2017310516186893e-05
GC_5_17 b_5 NI_5 NS_17 0 -3.1579056750460644e-05
GC_5_18 b_5 NI_5 NS_18 0 4.0468751764191472e-05
GC_5_19 b_5 NI_5 NS_19 0 1.7174483114844532e-05
GC_5_20 b_5 NI_5 NS_20 0 1.6685494845769982e-05
GC_5_21 b_5 NI_5 NS_21 0 1.0878141402056503e-05
GC_5_22 b_5 NI_5 NS_22 0 1.4951846063462488e-06
GC_5_23 b_5 NI_5 NS_23 0 -2.8644565407466025e-03
GC_5_24 b_5 NI_5 NS_24 0 4.9853307115217743e-03
GC_5_25 b_5 NI_5 NS_25 0 -5.2683096210683240e-04
GC_5_26 b_5 NI_5 NS_26 0 -8.2189971428641177e-04
GC_5_27 b_5 NI_5 NS_27 0 -1.3724840103427013e-04
GC_5_28 b_5 NI_5 NS_28 0 -7.8406967165332029e-04
GC_5_29 b_5 NI_5 NS_29 0 -9.6723649118608906e-06
GC_5_30 b_5 NI_5 NS_30 0 2.8515103100041413e-04
GC_5_31 b_5 NI_5 NS_31 0 -4.5413688115043922e-05
GC_5_32 b_5 NI_5 NS_32 0 1.0551722622461470e-04
GC_5_33 b_5 NI_5 NS_33 0 2.6490771633808862e-06
GC_5_34 b_5 NI_5 NS_34 0 7.9233666957986376e-05
GC_5_35 b_5 NI_5 NS_35 0 8.1010689014677533e-05
GC_5_36 b_5 NI_5 NS_36 0 9.7842365271812312e-05
GC_5_37 b_5 NI_5 NS_37 0 -2.6828682464833609e-05
GC_5_38 b_5 NI_5 NS_38 0 -4.0184188143575101e-05
GC_5_39 b_5 NI_5 NS_39 0 2.4454348158521298e-02
GC_5_40 b_5 NI_5 NS_40 0 1.2486815810610354e-03
GC_5_41 b_5 NI_5 NS_41 0 -1.3688454755995500e-02
GC_5_42 b_5 NI_5 NS_42 0 7.3661800987242319e-03
GC_5_43 b_5 NI_5 NS_43 0 -1.1679165318766710e-04
GC_5_44 b_5 NI_5 NS_44 0 2.5932399137972440e-04
GC_5_45 b_5 NI_5 NS_45 0 1.5402499417100325e-05
GC_5_46 b_5 NI_5 NS_46 0 -6.3259379556975637e-05
GC_5_47 b_5 NI_5 NS_47 0 -7.5914435504750351e-03
GC_5_48 b_5 NI_5 NS_48 0 -6.6537006025656695e-03
GC_5_49 b_5 NI_5 NS_49 0 3.1118498134875778e-05
GC_5_50 b_5 NI_5 NS_50 0 3.6341372720391568e-06
GC_5_51 b_5 NI_5 NS_51 0 1.2578518379711816e-02
GC_5_52 b_5 NI_5 NS_52 0 -4.1411239937955953e-03
GC_5_53 b_5 NI_5 NS_53 0 2.4606908253049502e-05
GC_5_54 b_5 NI_5 NS_54 0 -2.1104939970747678e-05
GC_5_55 b_5 NI_5 NS_55 0 -2.2599031608687512e-05
GC_5_56 b_5 NI_5 NS_56 0 5.8673672355875923e-05
GC_5_57 b_5 NI_5 NS_57 0 8.5324930982652706e-06
GC_5_58 b_5 NI_5 NS_58 0 1.9647239601634948e-06
GC_5_59 b_5 NI_5 NS_59 0 1.9206348877525660e-05
GC_5_60 b_5 NI_5 NS_60 0 3.2121051339309392e-06
GC_5_61 b_5 NI_5 NS_61 0 -3.8537879320889325e-03
GC_5_62 b_5 NI_5 NS_62 0 4.4434855000057265e-03
GC_5_63 b_5 NI_5 NS_63 0 -1.9680181710594617e-04
GC_5_64 b_5 NI_5 NS_64 0 -1.0660731315447129e-03
GC_5_65 b_5 NI_5 NS_65 0 -3.1099379868919342e-05
GC_5_66 b_5 NI_5 NS_66 0 -7.9284528820855124e-04
GC_5_67 b_5 NI_5 NS_67 0 -6.7900293262539480e-05
GC_5_68 b_5 NI_5 NS_68 0 2.3103711627005653e-04
GC_5_69 b_5 NI_5 NS_69 0 -1.0971160918811682e-04
GC_5_70 b_5 NI_5 NS_70 0 1.3589898841079413e-05
GC_5_71 b_5 NI_5 NS_71 0 -2.9430401830494346e-05
GC_5_72 b_5 NI_5 NS_72 0 5.8692114281503816e-05
GC_5_73 b_5 NI_5 NS_73 0 1.7815692125030416e-05
GC_5_74 b_5 NI_5 NS_74 0 1.5427097662887586e-04
GC_5_75 b_5 NI_5 NS_75 0 2.2686283159317014e-05
GC_5_76 b_5 NI_5 NS_76 0 2.1521656213092206e-05
GC_5_77 b_5 NI_5 NS_77 0 4.5064432844739433e-03
GC_5_78 b_5 NI_5 NS_78 0 -1.5161842820128264e-03
GC_5_79 b_5 NI_5 NS_79 0 -3.1878412900292652e-03
GC_5_80 b_5 NI_5 NS_80 0 1.2275614044657384e-02
GC_5_81 b_5 NI_5 NS_81 0 -1.8297885256241665e-03
GC_5_82 b_5 NI_5 NS_82 0 2.5881265512628487e-05
GC_5_83 b_5 NI_5 NS_83 0 -1.6147372056975353e-04
GC_5_84 b_5 NI_5 NS_84 0 1.1411979583934238e-04
GC_5_85 b_5 NI_5 NS_85 0 5.7952270889066806e-03
GC_5_86 b_5 NI_5 NS_86 0 1.2293691673864975e-02
GC_5_87 b_5 NI_5 NS_87 0 -2.8792193821524475e-05
GC_5_88 b_5 NI_5 NS_88 0 1.1372384341312716e-07
GC_5_89 b_5 NI_5 NS_89 0 8.9702420325768438e-03
GC_5_90 b_5 NI_5 NS_90 0 -5.7598530741420663e-03
GC_5_91 b_5 NI_5 NS_91 0 -3.7183897247743984e-05
GC_5_92 b_5 NI_5 NS_92 0 3.3446557141808482e-05
GC_5_93 b_5 NI_5 NS_93 0 -3.8534926743974517e-05
GC_5_94 b_5 NI_5 NS_94 0 2.2278618707086340e-05
GC_5_95 b_5 NI_5 NS_95 0 1.9407250563538656e-05
GC_5_96 b_5 NI_5 NS_96 0 1.0714939197344284e-05
GC_5_97 b_5 NI_5 NS_97 0 1.1993530649067441e-05
GC_5_98 b_5 NI_5 NS_98 0 -3.5715233255700609e-08
GC_5_99 b_5 NI_5 NS_99 0 -5.7538337419544899e-03
GC_5_100 b_5 NI_5 NS_100 0 2.1097898965913415e-03
GC_5_101 b_5 NI_5 NS_101 0 -3.1258481279634680e-04
GC_5_102 b_5 NI_5 NS_102 0 -6.8342497832974834e-04
GC_5_103 b_5 NI_5 NS_103 0 2.2150903299974510e-04
GC_5_104 b_5 NI_5 NS_104 0 -4.1999781065975951e-04
GC_5_105 b_5 NI_5 NS_105 0 -6.5845652761748762e-06
GC_5_106 b_5 NI_5 NS_106 0 1.2312863182342996e-04
GC_5_107 b_5 NI_5 NS_107 0 -2.5755654752893903e-06
GC_5_108 b_5 NI_5 NS_108 0 2.0294108925430954e-05
GC_5_109 b_5 NI_5 NS_109 0 1.3236893545785511e-05
GC_5_110 b_5 NI_5 NS_110 0 3.4588457200605095e-05
GC_5_111 b_5 NI_5 NS_111 0 1.0389627029598681e-04
GC_5_112 b_5 NI_5 NS_112 0 1.1134551856410321e-04
GC_5_113 b_5 NI_5 NS_113 0 3.9781210455771548e-05
GC_5_114 b_5 NI_5 NS_114 0 -2.8747568179879574e-05
GC_5_115 b_5 NI_5 NS_115 0 -2.0035663582701861e-02
GC_5_116 b_5 NI_5 NS_116 0 1.4593311508336298e-03
GC_5_117 b_5 NI_5 NS_117 0 1.0614461340308863e-02
GC_5_118 b_5 NI_5 NS_118 0 5.6714359347324892e-03
GC_5_119 b_5 NI_5 NS_119 0 1.2764290092259875e-04
GC_5_120 b_5 NI_5 NS_120 0 -2.6431052939663099e-04
GC_5_121 b_5 NI_5 NS_121 0 1.2509029245858092e-05
GC_5_122 b_5 NI_5 NS_122 0 -5.4172245288426027e-05
GC_5_123 b_5 NI_5 NS_123 0 -7.2699166510390252e-03
GC_5_124 b_5 NI_5 NS_124 0 -1.1536128320930488e-02
GC_5_125 b_5 NI_5 NS_125 0 3.0182600896341904e-05
GC_5_126 b_5 NI_5 NS_126 0 2.1998720226874446e-06
GC_5_127 b_5 NI_5 NS_127 0 1.2426257173336275e-02
GC_5_128 b_5 NI_5 NS_128 0 -1.3289792670160862e-02
GC_5_129 b_5 NI_5 NS_129 0 2.0654070795333374e-06
GC_5_130 b_5 NI_5 NS_130 0 -3.3527152609981780e-05
GC_5_131 b_5 NI_5 NS_131 0 -1.6132375550712491e-05
GC_5_132 b_5 NI_5 NS_132 0 5.6883207325629840e-05
GC_5_133 b_5 NI_5 NS_133 0 1.1337775794674097e-05
GC_5_134 b_5 NI_5 NS_134 0 1.4504956278311124e-05
GC_5_135 b_5 NI_5 NS_135 0 1.7896347193775126e-05
GC_5_136 b_5 NI_5 NS_136 0 1.5775577172305905e-06
GC_5_137 b_5 NI_5 NS_137 0 -5.6019487919096705e-03
GC_5_138 b_5 NI_5 NS_138 0 2.4609883936632820e-03
GC_5_139 b_5 NI_5 NS_139 0 -1.3605136234008256e-05
GC_5_140 b_5 NI_5 NS_140 0 -9.6373654975666389e-04
GC_5_141 b_5 NI_5 NS_141 0 3.4062455650546301e-04
GC_5_142 b_5 NI_5 NS_142 0 -5.2564669896894604e-04
GC_5_143 b_5 NI_5 NS_143 0 -9.1035344214105175e-05
GC_5_144 b_5 NI_5 NS_144 0 1.0867423692988449e-04
GC_5_145 b_5 NI_5 NS_145 0 -2.0153426630066478e-05
GC_5_146 b_5 NI_5 NS_146 0 3.2347638426712531e-06
GC_5_147 b_5 NI_5 NS_147 0 -7.8511936989643895e-06
GC_5_148 b_5 NI_5 NS_148 0 3.7488089962831026e-05
GC_5_149 b_5 NI_5 NS_149 0 3.6429825957811233e-05
GC_5_150 b_5 NI_5 NS_150 0 9.8694348427627178e-05
GC_5_151 b_5 NI_5 NS_151 0 2.4461626030860162e-05
GC_5_152 b_5 NI_5 NS_152 0 1.0555740420350450e-05
GC_5_153 b_5 NI_5 NS_153 0 1.0483741453438788e-01
GC_5_154 b_5 NI_5 NS_154 0 -1.7510761253956514e-03
GC_5_155 b_5 NI_5 NS_155 0 2.2541871142914126e-02
GC_5_156 b_5 NI_5 NS_156 0 -5.9733810413013261e-02
GC_5_157 b_5 NI_5 NS_157 0 -2.6797480673720177e-03
GC_5_158 b_5 NI_5 NS_158 0 -1.7340556930886362e-03
GC_5_159 b_5 NI_5 NS_159 0 -1.7225682177880210e-04
GC_5_160 b_5 NI_5 NS_160 0 -4.5890097297390762e-05
GC_5_161 b_5 NI_5 NS_161 0 -1.9514783906589603e-02
GC_5_162 b_5 NI_5 NS_162 0 -3.8543947173349810e-03
GC_5_163 b_5 NI_5 NS_163 0 -1.1151134492359333e-05
GC_5_164 b_5 NI_5 NS_164 0 5.8769291484556053e-06
GC_5_165 b_5 NI_5 NS_165 0 -4.0581134971731193e-02
GC_5_166 b_5 NI_5 NS_166 0 1.5921822284479231e-02
GC_5_167 b_5 NI_5 NS_167 0 -4.4242723560094328e-05
GC_5_168 b_5 NI_5 NS_168 0 6.3912118527452604e-06
GC_5_169 b_5 NI_5 NS_169 0 -3.8200376817975742e-05
GC_5_170 b_5 NI_5 NS_170 0 -3.2601645574327765e-06
GC_5_171 b_5 NI_5 NS_171 0 1.5273406979473963e-05
GC_5_172 b_5 NI_5 NS_172 0 -2.8651142167052884e-05
GC_5_173 b_5 NI_5 NS_173 0 5.6701141093741137e-06
GC_5_174 b_5 NI_5 NS_174 0 -8.5678685907581652e-07
GC_5_175 b_5 NI_5 NS_175 0 -5.4319995733546405e-03
GC_5_176 b_5 NI_5 NS_176 0 6.6587378656452808e-03
GC_5_177 b_5 NI_5 NS_177 0 -5.7831641411607080e-04
GC_5_178 b_5 NI_5 NS_178 0 -8.8591560683603827e-04
GC_5_179 b_5 NI_5 NS_179 0 2.0854794333113912e-04
GC_5_180 b_5 NI_5 NS_180 0 -8.0977722036954783e-04
GC_5_181 b_5 NI_5 NS_181 0 -4.7303477398816352e-05
GC_5_182 b_5 NI_5 NS_182 0 1.6431673173012364e-04
GC_5_183 b_5 NI_5 NS_183 0 3.9251141569449339e-06
GC_5_184 b_5 NI_5 NS_184 0 -8.5165130119916580e-05
GC_5_185 b_5 NI_5 NS_185 0 -2.0202272364499099e-05
GC_5_186 b_5 NI_5 NS_186 0 -3.2028374035704413e-05
GC_5_187 b_5 NI_5 NS_187 0 2.6873351988991742e-04
GC_5_188 b_5 NI_5 NS_188 0 8.6840364952453717e-05
GC_5_189 b_5 NI_5 NS_189 0 5.7214859690624296e-05
GC_5_190 b_5 NI_5 NS_190 0 -1.4240547152782413e-04
GC_5_191 b_5 NI_5 NS_191 0 -2.1746091852982256e-02
GC_5_192 b_5 NI_5 NS_192 0 2.3989607795563885e-03
GC_5_193 b_5 NI_5 NS_193 0 3.8826022878741422e-02
GC_5_194 b_5 NI_5 NS_194 0 -5.8367941703060672e-03
GC_5_195 b_5 NI_5 NS_195 0 9.1004746075298187e-04
GC_5_196 b_5 NI_5 NS_196 0 5.6568921314958994e-05
GC_5_197 b_5 NI_5 NS_197 0 4.1683557152023526e-05
GC_5_198 b_5 NI_5 NS_198 0 -7.4943000074461154e-06
GC_5_199 b_5 NI_5 NS_199 0 3.6784461623194382e-02
GC_5_200 b_5 NI_5 NS_200 0 2.6844189169821366e-02
GC_5_201 b_5 NI_5 NS_201 0 2.9071482500662762e-05
GC_5_202 b_5 NI_5 NS_202 0 2.8922352306317376e-06
GC_5_203 b_5 NI_5 NS_203 0 -4.2909210338046726e-02
GC_5_204 b_5 NI_5 NS_204 0 2.1736260016364684e-02
GC_5_205 b_5 NI_5 NS_205 0 2.5193832521323326e-06
GC_5_206 b_5 NI_5 NS_206 0 1.0165715639576446e-05
GC_5_207 b_5 NI_5 NS_207 0 -9.0834705199573567e-07
GC_5_208 b_5 NI_5 NS_208 0 4.2851571564127299e-05
GC_5_209 b_5 NI_5 NS_209 0 1.4262710929610972e-07
GC_5_210 b_5 NI_5 NS_210 0 2.4290384054909198e-06
GC_5_211 b_5 NI_5 NS_211 0 7.4505434836659962e-09
GC_5_212 b_5 NI_5 NS_212 0 1.3773392229147214e-06
GC_5_213 b_5 NI_5 NS_213 0 -1.4314936939014964e-03
GC_5_214 b_5 NI_5 NS_214 0 4.2304686037950897e-03
GC_5_215 b_5 NI_5 NS_215 0 -4.5169652475186487e-04
GC_5_216 b_5 NI_5 NS_216 0 -4.4265618181612020e-04
GC_5_217 b_5 NI_5 NS_217 0 2.0189360588628803e-05
GC_5_218 b_5 NI_5 NS_218 0 -4.7709425684660048e-04
GC_5_219 b_5 NI_5 NS_219 0 -1.5235434419512792e-05
GC_5_220 b_5 NI_5 NS_220 0 1.7022656918999767e-04
GC_5_221 b_5 NI_5 NS_221 0 1.0710117278457285e-04
GC_5_222 b_5 NI_5 NS_222 0 1.2874331430818116e-05
GC_5_223 b_5 NI_5 NS_223 0 2.8948695804092154e-05
GC_5_224 b_5 NI_5 NS_224 0 -1.3241370916578563e-06
GC_5_225 b_5 NI_5 NS_225 0 2.0427669689658258e-04
GC_5_226 b_5 NI_5 NS_226 0 1.6541931560344397e-04
GC_5_227 b_5 NI_5 NS_227 0 1.0472499216285785e-04
GC_5_228 b_5 NI_5 NS_228 0 -7.7255481270301651e-05
GC_5_229 b_5 NI_5 NS_229 0 2.6549362019154799e-02
GC_5_230 b_5 NI_5 NS_230 0 -1.4757316747489766e-03
GC_5_231 b_5 NI_5 NS_231 0 -6.1702228278182995e-03
GC_5_232 b_5 NI_5 NS_232 0 1.9721088126745955e-02
GC_5_233 b_5 NI_5 NS_233 0 -1.4237726332678449e-04
GC_5_234 b_5 NI_5 NS_234 0 1.0296482848257775e-03
GC_5_235 b_5 NI_5 NS_235 0 1.2376695541811662e-04
GC_5_236 b_5 NI_5 NS_236 0 6.8549750727094541e-05
GC_5_237 b_5 NI_5 NS_237 0 2.4207816608074386e-03
GC_5_238 b_5 NI_5 NS_238 0 6.0131159060295104e-03
GC_5_239 b_5 NI_5 NS_239 0 -9.5944277535622988e-06
GC_5_240 b_5 NI_5 NS_240 0 1.4384920318016200e-06
GC_5_241 b_5 NI_5 NS_241 0 1.6850247302030014e-02
GC_5_242 b_5 NI_5 NS_242 0 -1.2034517353050393e-02
GC_5_243 b_5 NI_5 NS_243 0 5.6718140009897957e-06
GC_5_244 b_5 NI_5 NS_244 0 5.8071306111465379e-05
GC_5_245 b_5 NI_5 NS_245 0 -2.5091115538714552e-05
GC_5_246 b_5 NI_5 NS_246 0 4.1322833174306703e-05
GC_5_247 b_5 NI_5 NS_247 0 -2.2209790748164933e-06
GC_5_248 b_5 NI_5 NS_248 0 -1.1921723681695547e-05
GC_5_249 b_5 NI_5 NS_249 0 -2.8885979573306900e-06
GC_5_250 b_5 NI_5 NS_250 0 -3.8370744317080833e-06
GC_5_251 b_5 NI_5 NS_251 0 -3.6728429658018590e-03
GC_5_252 b_5 NI_5 NS_252 0 8.2084668503622938e-03
GC_5_253 b_5 NI_5 NS_253 0 -7.3829747115306075e-04
GC_5_254 b_5 NI_5 NS_254 0 -5.4548774159952310e-04
GC_5_255 b_5 NI_5 NS_255 0 2.4647908320391969e-04
GC_5_256 b_5 NI_5 NS_256 0 -5.9445175398261350e-04
GC_5_257 b_5 NI_5 NS_257 0 -6.5440352510381600e-05
GC_5_258 b_5 NI_5 NS_258 0 1.1352041079629130e-05
GC_5_259 b_5 NI_5 NS_259 0 7.0688898452147361e-06
GC_5_260 b_5 NI_5 NS_260 0 -6.3151254820958109e-05
GC_5_261 b_5 NI_5 NS_261 0 2.8909377182584398e-05
GC_5_262 b_5 NI_5 NS_262 0 1.0865101692403229e-05
GC_5_263 b_5 NI_5 NS_263 0 3.0539045481804466e-05
GC_5_264 b_5 NI_5 NS_264 0 -4.8049224593056311e-05
GC_5_265 b_5 NI_5 NS_265 0 2.5508888091815403e-05
GC_5_266 b_5 NI_5 NS_266 0 3.9156863379882083e-05
GC_5_267 b_5 NI_5 NS_267 0 -2.4971594576457343e-03
GC_5_268 b_5 NI_5 NS_268 0 1.1659585035991103e-03
GC_5_269 b_5 NI_5 NS_269 0 1.4959099837819664e-03
GC_5_270 b_5 NI_5 NS_270 0 -6.3560605622840528e-03
GC_5_271 b_5 NI_5 NS_271 0 -5.5644224687339383e-05
GC_5_272 b_5 NI_5 NS_272 0 7.7035156092209334e-04
GC_5_273 b_5 NI_5 NS_273 0 3.6592463717765451e-05
GC_5_274 b_5 NI_5 NS_274 0 9.7290367293024634e-05
GC_5_275 b_5 NI_5 NS_275 0 -1.2769222814613505e-02
GC_5_276 b_5 NI_5 NS_276 0 -1.9886361806241395e-02
GC_5_277 b_5 NI_5 NS_277 0 -7.7311559703026935e-07
GC_5_278 b_5 NI_5 NS_278 0 -4.9343589355615095e-06
GC_5_279 b_5 NI_5 NS_279 0 7.6752981653354811e-03
GC_5_280 b_5 NI_5 NS_280 0 -1.7877396024429611e-02
GC_5_281 b_5 NI_5 NS_281 0 -1.7263460496868343e-05
GC_5_282 b_5 NI_5 NS_282 0 8.4620317381809730e-06
GC_5_283 b_5 NI_5 NS_283 0 -2.0330356811530423e-05
GC_5_284 b_5 NI_5 NS_284 0 4.7619475121230945e-05
GC_5_285 b_5 NI_5 NS_285 0 -6.0876428658247271e-06
GC_5_286 b_5 NI_5 NS_286 0 -3.4050066576581987e-06
GC_5_287 b_5 NI_5 NS_287 0 3.9523536010655239e-07
GC_5_288 b_5 NI_5 NS_288 0 -5.6837396071609503e-06
GC_5_289 b_5 NI_5 NS_289 0 -3.8285643593890650e-03
GC_5_290 b_5 NI_5 NS_290 0 8.7866670661717189e-03
GC_5_291 b_5 NI_5 NS_291 0 -5.2098947272650705e-04
GC_5_292 b_5 NI_5 NS_292 0 -5.8846887537936294e-04
GC_5_293 b_5 NI_5 NS_293 0 3.7055993748796900e-04
GC_5_294 b_5 NI_5 NS_294 0 -5.3886174612955903e-04
GC_5_295 b_5 NI_5 NS_295 0 -7.1652385380499957e-05
GC_5_296 b_5 NI_5 NS_296 0 -1.4463440516835607e-05
GC_5_297 b_5 NI_5 NS_297 0 6.0196290187172629e-05
GC_5_298 b_5 NI_5 NS_298 0 -2.0499867398563269e-05
GC_5_299 b_5 NI_5 NS_299 0 1.4083624100949393e-05
GC_5_300 b_5 NI_5 NS_300 0 2.2907342498772090e-05
GC_5_301 b_5 NI_5 NS_301 0 5.9660379448098215e-05
GC_5_302 b_5 NI_5 NS_302 0 -2.4588159612687504e-05
GC_5_303 b_5 NI_5 NS_303 0 -1.2181378269507771e-06
GC_5_304 b_5 NI_5 NS_304 0 4.4775901322060367e-05
GC_5_305 b_5 NI_5 NS_305 0 -1.8458925845428638e-02
GC_5_306 b_5 NI_5 NS_306 0 -1.2992290564723162e-03
GC_5_307 b_5 NI_5 NS_307 0 6.6809226242653570e-03
GC_5_308 b_5 NI_5 NS_308 0 1.1259900496311382e-02
GC_5_309 b_5 NI_5 NS_309 0 6.4840651454294853e-04
GC_5_310 b_5 NI_5 NS_310 0 7.7943220436935893e-04
GC_5_311 b_5 NI_5 NS_311 0 2.0724746381684190e-04
GC_5_312 b_5 NI_5 NS_312 0 -8.8605741386969025e-05
GC_5_313 b_5 NI_5 NS_313 0 6.8036075074580388e-03
GC_5_314 b_5 NI_5 NS_314 0 4.2615357388301103e-03
GC_5_315 b_5 NI_5 NS_315 0 -1.0369083900238884e-05
GC_5_316 b_5 NI_5 NS_316 0 5.9758407061885098e-07
GC_5_317 b_5 NI_5 NS_317 0 1.2412878327471455e-02
GC_5_318 b_5 NI_5 NS_318 0 -9.3232862864907860e-03
GC_5_319 b_5 NI_5 NS_319 0 5.0525964234738531e-06
GC_5_320 b_5 NI_5 NS_320 0 -1.1262583771150057e-05
GC_5_321 b_5 NI_5 NS_321 0 -3.8782804968951341e-05
GC_5_322 b_5 NI_5 NS_322 0 6.8361224231757529e-05
GC_5_323 b_5 NI_5 NS_323 0 -5.0518954995744676e-06
GC_5_324 b_5 NI_5 NS_324 0 -3.5392454933187993e-05
GC_5_325 b_5 NI_5 NS_325 0 -1.0250098299392103e-05
GC_5_326 b_5 NI_5 NS_326 0 -7.7962653455294070e-07
GC_5_327 b_5 NI_5 NS_327 0 -3.9060016505965355e-03
GC_5_328 b_5 NI_5 NS_328 0 3.3805662267721039e-03
GC_5_329 b_5 NI_5 NS_329 0 -3.3049643347509713e-04
GC_5_330 b_5 NI_5 NS_330 0 -5.6535717591216803e-04
GC_5_331 b_5 NI_5 NS_331 0 4.1296284708627385e-04
GC_5_332 b_5 NI_5 NS_332 0 -2.7805008541931193e-04
GC_5_333 b_5 NI_5 NS_333 0 -4.7328204886957191e-05
GC_5_334 b_5 NI_5 NS_334 0 1.8363638381430021e-05
GC_5_335 b_5 NI_5 NS_335 0 3.0442594215134486e-05
GC_5_336 b_5 NI_5 NS_336 0 2.3585013782290456e-05
GC_5_337 b_5 NI_5 NS_337 0 9.3128699326932609e-06
GC_5_338 b_5 NI_5 NS_338 0 -8.5490219973064937e-06
GC_5_339 b_5 NI_5 NS_339 0 2.5838969170324509e-05
GC_5_340 b_5 NI_5 NS_340 0 1.0007706260401648e-04
GC_5_341 b_5 NI_5 NS_341 0 6.1105743962887475e-05
GC_5_342 b_5 NI_5 NS_342 0 3.5030306594745207e-06
GC_5_343 b_5 NI_5 NS_343 0 1.0944576073872817e-02
GC_5_344 b_5 NI_5 NS_344 0 1.3496442904264068e-03
GC_5_345 b_5 NI_5 NS_345 0 -1.2355860376009584e-02
GC_5_346 b_5 NI_5 NS_346 0 2.0266715960675602e-03
GC_5_347 b_5 NI_5 NS_347 0 3.0286230347337982e-04
GC_5_348 b_5 NI_5 NS_348 0 -5.5943784402189350e-05
GC_5_349 b_5 NI_5 NS_349 0 7.4864717977725159e-05
GC_5_350 b_5 NI_5 NS_350 0 -6.3940601230532158e-05
GC_5_351 b_5 NI_5 NS_351 0 -4.2789902167527892e-03
GC_5_352 b_5 NI_5 NS_352 0 -5.6125858829747066e-04
GC_5_353 b_5 NI_5 NS_353 0 1.3780800100462177e-05
GC_5_354 b_5 NI_5 NS_354 0 2.2699521906947812e-06
GC_5_355 b_5 NI_5 NS_355 0 1.1409484792164587e-02
GC_5_356 b_5 NI_5 NS_356 0 1.6020733974489859e-03
GC_5_357 b_5 NI_5 NS_357 0 -2.1548214845832227e-05
GC_5_358 b_5 NI_5 NS_358 0 -3.1646757726260136e-05
GC_5_359 b_5 NI_5 NS_359 0 -1.7189091486872813e-05
GC_5_360 b_5 NI_5 NS_360 0 5.5921613234506654e-05
GC_5_361 b_5 NI_5 NS_361 0 1.1204464866154965e-06
GC_5_362 b_5 NI_5 NS_362 0 -1.8508488977215644e-05
GC_5_363 b_5 NI_5 NS_363 0 -7.9308748792240137e-06
GC_5_364 b_5 NI_5 NS_364 0 -5.7422302193997429e-07
GC_5_365 b_5 NI_5 NS_365 0 -3.7107829393811490e-03
GC_5_366 b_5 NI_5 NS_366 0 1.3307656008600670e-03
GC_5_367 b_5 NI_5 NS_367 0 5.5059173873492814e-06
GC_5_368 b_5 NI_5 NS_368 0 -6.2286923541341366e-04
GC_5_369 b_5 NI_5 NS_369 0 3.2649451316424513e-04
GC_5_370 b_5 NI_5 NS_370 0 -1.7113251511873836e-04
GC_5_371 b_5 NI_5 NS_371 0 1.8901940948911067e-05
GC_5_372 b_5 NI_5 NS_372 0 -8.2996580858078914e-06
GC_5_373 b_5 NI_5 NS_373 0 8.1960824268637938e-06
GC_5_374 b_5 NI_5 NS_374 0 -1.1917994092277191e-05
GC_5_375 b_5 NI_5 NS_375 0 -2.2656754353297768e-05
GC_5_376 b_5 NI_5 NS_376 0 -1.3419957833285681e-05
GC_5_377 b_5 NI_5 NS_377 0 6.4455687308701074e-05
GC_5_378 b_5 NI_5 NS_378 0 -5.1900271486757277e-05
GC_5_379 b_5 NI_5 NS_379 0 -1.9762695379737338e-05
GC_5_380 b_5 NI_5 NS_380 0 -4.2242085176098725e-05
GC_5_381 b_5 NI_5 NS_381 0 -1.2243440229192524e-02
GC_5_382 b_5 NI_5 NS_382 0 -1.0230968241244801e-03
GC_5_383 b_5 NI_5 NS_383 0 -5.2687458351901705e-04
GC_5_384 b_5 NI_5 NS_384 0 7.4680608131642351e-03
GC_5_385 b_5 NI_5 NS_385 0 1.0116743672013504e-03
GC_5_386 b_5 NI_5 NS_386 0 -7.4477842525016983e-05
GC_5_387 b_5 NI_5 NS_387 0 1.4568483107349207e-04
GC_5_388 b_5 NI_5 NS_388 0 -1.9821030766074621e-04
GC_5_389 b_5 NI_5 NS_389 0 3.9935588764083716e-03
GC_5_390 b_5 NI_5 NS_390 0 -2.3501735701699786e-03
GC_5_391 b_5 NI_5 NS_391 0 -1.1344459234568547e-05
GC_5_392 b_5 NI_5 NS_392 0 -2.1422768023557226e-06
GC_5_393 b_5 NI_5 NS_393 0 8.1839985058773379e-03
GC_5_394 b_5 NI_5 NS_394 0 -5.2425631452285579e-03
GC_5_395 b_5 NI_5 NS_395 0 2.9233137916905286e-05
GC_5_396 b_5 NI_5 NS_396 0 -7.8957672134465635e-05
GC_5_397 b_5 NI_5 NS_397 0 3.9330158180892534e-06
GC_5_398 b_5 NI_5 NS_398 0 5.2531850614590770e-05
GC_5_399 b_5 NI_5 NS_399 0 -1.3963028610001260e-05
GC_5_400 b_5 NI_5 NS_400 0 -3.7407663895300018e-05
GC_5_401 b_5 NI_5 NS_401 0 -8.1075976549025850e-06
GC_5_402 b_5 NI_5 NS_402 0 -3.9234609059649420e-07
GC_5_403 b_5 NI_5 NS_403 0 -1.0696833689533500e-03
GC_5_404 b_5 NI_5 NS_404 0 1.6545890592747675e-03
GC_5_405 b_5 NI_5 NS_405 0 -3.1129580040031564e-04
GC_5_406 b_5 NI_5 NS_406 0 -1.3497337035769325e-04
GC_5_407 b_5 NI_5 NS_407 0 4.6296705848246063e-04
GC_5_408 b_5 NI_5 NS_408 0 8.7032318273398918e-05
GC_5_409 b_5 NI_5 NS_409 0 8.1032182733006911e-06
GC_5_410 b_5 NI_5 NS_410 0 -1.2224610060496431e-04
GC_5_411 b_5 NI_5 NS_411 0 -1.0120764239074905e-05
GC_5_412 b_5 NI_5 NS_412 0 5.3253368083855083e-05
GC_5_413 b_5 NI_5 NS_413 0 -2.8254812270746803e-05
GC_5_414 b_5 NI_5 NS_414 0 -1.6647623889960553e-05
GC_5_415 b_5 NI_5 NS_415 0 -1.0520165056382719e-04
GC_5_416 b_5 NI_5 NS_416 0 -2.4069789331625161e-06
GC_5_417 b_5 NI_5 NS_417 0 -2.8863529551486811e-06
GC_5_418 b_5 NI_5 NS_418 0 1.4300261671492734e-05
GC_5_419 b_5 NI_5 NS_419 0 2.4018928091190203e-02
GC_5_420 b_5 NI_5 NS_420 0 1.1010201037260727e-03
GC_5_421 b_5 NI_5 NS_421 0 -1.9026933839991909e-02
GC_5_422 b_5 NI_5 NS_422 0 7.3243369711151049e-03
GC_5_423 b_5 NI_5 NS_423 0 3.8568776199776080e-04
GC_5_424 b_5 NI_5 NS_424 0 -5.4604611787761523e-04
GC_5_425 b_5 NI_5 NS_425 0 5.4855736756652366e-05
GC_5_426 b_5 NI_5 NS_426 0 -1.2298791074429714e-04
GC_5_427 b_5 NI_5 NS_427 0 -2.3024289516938045e-03
GC_5_428 b_5 NI_5 NS_428 0 4.9587873680959436e-03
GC_5_429 b_5 NI_5 NS_429 0 1.3957690699997629e-05
GC_5_430 b_5 NI_5 NS_430 0 3.3805925059044064e-06
GC_5_431 b_5 NI_5 NS_431 0 1.0233658323616524e-02
GC_5_432 b_5 NI_5 NS_432 0 3.6585487134749230e-03
GC_5_433 b_5 NI_5 NS_433 0 5.4703207254008622e-06
GC_5_434 b_5 NI_5 NS_434 0 -7.3520293694205688e-05
GC_5_435 b_5 NI_5 NS_435 0 2.3385122554214987e-06
GC_5_436 b_5 NI_5 NS_436 0 5.4777984409509516e-05
GC_5_437 b_5 NI_5 NS_437 0 -1.5234496894889409e-06
GC_5_438 b_5 NI_5 NS_438 0 -2.2211163334934944e-05
GC_5_439 b_5 NI_5 NS_439 0 -7.1498529527242076e-06
GC_5_440 b_5 NI_5 NS_440 0 -1.1896445747343180e-07
GC_5_441 b_5 NI_5 NS_441 0 -2.9511948100472201e-03
GC_5_442 b_5 NI_5 NS_442 0 9.2746862587667729e-04
GC_5_443 b_5 NI_5 NS_443 0 4.8661853580650417e-05
GC_5_444 b_5 NI_5 NS_444 0 -4.2792047793059553e-04
GC_5_445 b_5 NI_5 NS_445 0 4.7332672641533298e-04
GC_5_446 b_5 NI_5 NS_446 0 1.3517647890072166e-04
GC_5_447 b_5 NI_5 NS_447 0 7.2380783382189435e-05
GC_5_448 b_5 NI_5 NS_448 0 -9.4996062333991413e-05
GC_5_449 b_5 NI_5 NS_449 0 -3.6983211374651785e-05
GC_5_450 b_5 NI_5 NS_450 0 2.9796025086453457e-05
GC_5_451 b_5 NI_5 NS_451 0 -1.3266229775825231e-05
GC_5_452 b_5 NI_5 NS_452 0 -3.7228691682927443e-05
GC_5_453 b_5 NI_5 NS_453 0 -4.8364343126400997e-05
GC_5_454 b_5 NI_5 NS_454 0 -6.2144443960398033e-05
GC_5_455 b_5 NI_5 NS_455 0 -1.4212768011268579e-05
GC_5_456 b_5 NI_5 NS_456 0 -1.2310036531374020e-05
GD_5_1 b_5 NI_5 NA_1 0 -6.7858544798315963e-03
GD_5_2 b_5 NI_5 NA_2 0 -1.2140357211764532e-02
GD_5_3 b_5 NI_5 NA_3 0 7.1846922445859270e-05
GD_5_4 b_5 NI_5 NA_4 0 6.4943179521555656e-03
GD_5_5 b_5 NI_5 NA_5 0 -8.9663376891664079e-02
GD_5_6 b_5 NI_5 NA_6 0 -2.3084949215942872e-02
GD_5_7 b_5 NI_5 NA_7 0 -3.4465407382335209e-02
GD_5_8 b_5 NI_5 NA_8 0 1.0065939315554979e-02
GD_5_9 b_5 NI_5 NA_9 0 -7.3343710144443000e-03
GD_5_10 b_5 NI_5 NA_10 0 -3.1501632733959973e-03
GD_5_11 b_5 NI_5 NA_11 0 -4.7349435278623076e-04
GD_5_12 b_5 NI_5 NA_12 0 -1.0633091615751069e-02
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 2.4178360865711175e-03
GC_6_2 b_6 NI_6 NS_2 0 1.2757473058295056e-03
GC_6_3 b_6 NI_6 NS_3 0 -4.4337225936820117e-03
GC_6_4 b_6 NI_6 NS_4 0 6.6354211154788416e-03
GC_6_5 b_6 NI_6 NS_5 0 -6.2658676922004882e-05
GC_6_6 b_6 NI_6 NS_6 0 -1.6625360027838266e-04
GC_6_7 b_6 NI_6 NS_7 0 -2.6207789803272999e-05
GC_6_8 b_6 NI_6 NS_8 0 -5.0790761141216481e-06
GC_6_9 b_6 NI_6 NS_9 0 -4.1617445949706450e-03
GC_6_10 b_6 NI_6 NS_10 0 -2.2673655156195014e-03
GC_6_11 b_6 NI_6 NS_11 0 3.9083015268570613e-05
GC_6_12 b_6 NI_6 NS_12 0 3.7325207341679119e-06
GC_6_13 b_6 NI_6 NS_13 0 9.5292179931826641e-03
GC_6_14 b_6 NI_6 NS_14 0 -5.1998294790768654e-03
GC_6_15 b_6 NI_6 NS_15 0 -7.5097632703969989e-06
GC_6_16 b_6 NI_6 NS_16 0 -4.8417069305130071e-07
GC_6_17 b_6 NI_6 NS_17 0 -1.9775231522449371e-05
GC_6_18 b_6 NI_6 NS_18 0 1.5570511141690434e-05
GC_6_19 b_6 NI_6 NS_19 0 1.8954093548947453e-05
GC_6_20 b_6 NI_6 NS_20 0 -1.2690652052064905e-05
GC_6_21 b_6 NI_6 NS_21 0 -7.5635512779553380e-06
GC_6_22 b_6 NI_6 NS_22 0 2.9259218824340466e-06
GC_6_23 b_6 NI_6 NS_23 0 -1.3630774666985822e-03
GC_6_24 b_6 NI_6 NS_24 0 2.6990656075751079e-03
GC_6_25 b_6 NI_6 NS_25 0 -3.1433186425744572e-04
GC_6_26 b_6 NI_6 NS_26 0 -5.7769934798053858e-04
GC_6_27 b_6 NI_6 NS_27 0 -7.8696011499414573e-05
GC_6_28 b_6 NI_6 NS_28 0 -5.9334511719464733e-04
GC_6_29 b_6 NI_6 NS_29 0 -5.5416432522469229e-05
GC_6_30 b_6 NI_6 NS_30 0 1.9006831710440331e-04
GC_6_31 b_6 NI_6 NS_31 0 -9.2353677418877098e-05
GC_6_32 b_6 NI_6 NS_32 0 -8.7763296914338717e-05
GC_6_33 b_6 NI_6 NS_33 0 -7.7298069571654702e-05
GC_6_34 b_6 NI_6 NS_34 0 1.6349400313504522e-05
GC_6_35 b_6 NI_6 NS_35 0 6.5680347723196016e-05
GC_6_36 b_6 NI_6 NS_36 0 9.3310720197581733e-05
GC_6_37 b_6 NI_6 NS_37 0 -3.2476954394847924e-06
GC_6_38 b_6 NI_6 NS_38 0 -4.9509382717010810e-05
GC_6_39 b_6 NI_6 NS_39 0 -1.6742674685083045e-02
GC_6_40 b_6 NI_6 NS_40 0 -1.1938103742974620e-03
GC_6_41 b_6 NI_6 NS_41 0 6.4193301467349671e-04
GC_6_42 b_6 NI_6 NS_42 0 1.0394557259842689e-02
GC_6_43 b_6 NI_6 NS_43 0 -1.8237313571587631e-04
GC_6_44 b_6 NI_6 NS_44 0 2.2338028858786829e-05
GC_6_45 b_6 NI_6 NS_45 0 -4.1233282467569859e-05
GC_6_46 b_6 NI_6 NS_46 0 -1.4491918415844490e-05
GC_6_47 b_6 NI_6 NS_47 0 7.5915637400747376e-03
GC_6_48 b_6 NI_6 NS_48 0 7.4925562265614797e-03
GC_6_49 b_6 NI_6 NS_49 0 -2.9456115115578813e-05
GC_6_50 b_6 NI_6 NS_50 0 -2.2041753072573654e-06
GC_6_51 b_6 NI_6 NS_51 0 1.2167638135467167e-02
GC_6_52 b_6 NI_6 NS_52 0 -6.7260502262053816e-03
GC_6_53 b_6 NI_6 NS_53 0 -1.4499779181971472e-05
GC_6_54 b_6 NI_6 NS_54 0 1.2139489923852980e-05
GC_6_55 b_6 NI_6 NS_55 0 -2.2658371222055654e-05
GC_6_56 b_6 NI_6 NS_56 0 2.7670783827257258e-05
GC_6_57 b_6 NI_6 NS_57 0 5.6745343886767339e-06
GC_6_58 b_6 NI_6 NS_58 0 -2.9482457932476233e-06
GC_6_59 b_6 NI_6 NS_59 0 -1.2771761996347416e-05
GC_6_60 b_6 NI_6 NS_60 0 5.7272711877218923e-06
GC_6_61 b_6 NI_6 NS_61 0 -2.6452067773032237e-03
GC_6_62 b_6 NI_6 NS_62 0 3.9280406411299519e-03
GC_6_63 b_6 NI_6 NS_63 0 -1.1065164351958192e-04
GC_6_64 b_6 NI_6 NS_64 0 -8.0410195949890957e-04
GC_6_65 b_6 NI_6 NS_65 0 5.5547188456075515e-05
GC_6_66 b_6 NI_6 NS_66 0 -6.7263728795029394e-04
GC_6_67 b_6 NI_6 NS_67 0 -9.8895826249692615e-05
GC_6_68 b_6 NI_6 NS_68 0 1.2941657934378866e-04
GC_6_69 b_6 NI_6 NS_69 0 1.1513733522762177e-07
GC_6_70 b_6 NI_6 NS_70 0 -1.2995266343533173e-04
GC_6_71 b_6 NI_6 NS_71 0 -2.6014740141683634e-05
GC_6_72 b_6 NI_6 NS_72 0 -4.9425610736452481e-05
GC_6_73 b_6 NI_6 NS_73 0 1.2024054937647527e-05
GC_6_74 b_6 NI_6 NS_74 0 1.1972756381725557e-04
GC_6_75 b_6 NI_6 NS_75 0 4.5968798144789580e-06
GC_6_76 b_6 NI_6 NS_76 0 1.2806538886517006e-05
GC_6_77 b_6 NI_6 NS_77 0 -2.8443030229653634e-02
GC_6_78 b_6 NI_6 NS_78 0 1.4955325134402466e-03
GC_6_79 b_6 NI_6 NS_79 0 1.8247423708271621e-02
GC_6_80 b_6 NI_6 NS_80 0 5.3006359554845332e-03
GC_6_81 b_6 NI_6 NS_81 0 -4.5241668868645796e-05
GC_6_82 b_6 NI_6 NS_82 0 -2.7701767758547889e-04
GC_6_83 b_6 NI_6 NS_83 0 -3.9819765217001397e-05
GC_6_84 b_6 NI_6 NS_84 0 -2.6277233327688660e-06
GC_6_85 b_6 NI_6 NS_85 0 -7.1105909292300236e-03
GC_6_86 b_6 NI_6 NS_86 0 -1.1193699371304587e-02
GC_6_87 b_6 NI_6 NS_87 0 3.5139295641854737e-05
GC_6_88 b_6 NI_6 NS_88 0 1.6783429538419835e-06
GC_6_89 b_6 NI_6 NS_89 0 7.2413193891493277e-03
GC_6_90 b_6 NI_6 NS_90 0 -1.6741226091366287e-02
GC_6_91 b_6 NI_6 NS_91 0 -1.3405821588005844e-05
GC_6_92 b_6 NI_6 NS_92 0 2.0244596221327022e-06
GC_6_93 b_6 NI_6 NS_93 0 -1.5958425830094140e-05
GC_6_94 b_6 NI_6 NS_94 0 2.4840191377958053e-05
GC_6_95 b_6 NI_6 NS_95 0 1.9780828912749309e-05
GC_6_96 b_6 NI_6 NS_96 0 -1.0051588007276941e-05
GC_6_97 b_6 NI_6 NS_97 0 -7.0408773299358986e-06
GC_6_98 b_6 NI_6 NS_98 0 3.3239385818868089e-06
GC_6_99 b_6 NI_6 NS_99 0 -2.9706391025445698e-03
GC_6_100 b_6 NI_6 NS_100 0 1.8891379781008015e-03
GC_6_101 b_6 NI_6 NS_101 0 -2.5724740705391813e-04
GC_6_102 b_6 NI_6 NS_102 0 -4.5693238048794894e-04
GC_6_103 b_6 NI_6 NS_103 0 1.0923702697356215e-04
GC_6_104 b_6 NI_6 NS_104 0 -3.1934098702567087e-04
GC_6_105 b_6 NI_6 NS_105 0 -1.7160862918471313e-05
GC_6_106 b_6 NI_6 NS_106 0 1.0940888473132502e-04
GC_6_107 b_6 NI_6 NS_107 0 -1.6799826805548945e-05
GC_6_108 b_6 NI_6 NS_108 0 -1.6651536305036188e-05
GC_6_109 b_6 NI_6 NS_109 0 -2.6024370646772450e-05
GC_6_110 b_6 NI_6 NS_110 0 1.0673482640120225e-05
GC_6_111 b_6 NI_6 NS_111 0 6.7045706990544646e-05
GC_6_112 b_6 NI_6 NS_112 0 1.1878577288783087e-04
GC_6_113 b_6 NI_6 NS_113 0 3.5666404675524048e-05
GC_6_114 b_6 NI_6 NS_114 0 -7.8247845939503629e-06
GC_6_115 b_6 NI_6 NS_115 0 -1.2535064614446315e-02
GC_6_116 b_6 NI_6 NS_116 0 -1.4706200566388548e-03
GC_6_117 b_6 NI_6 NS_117 0 7.0061417083972771e-03
GC_6_118 b_6 NI_6 NS_118 0 2.7492837838096293e-02
GC_6_119 b_6 NI_6 NS_119 0 -1.6242382644635726e-04
GC_6_120 b_6 NI_6 NS_120 0 1.8916067541734682e-04
GC_6_121 b_6 NI_6 NS_121 0 -4.6484831708750337e-05
GC_6_122 b_6 NI_6 NS_122 0 8.3396306875866938e-06
GC_6_123 b_6 NI_6 NS_123 0 7.3644823016085232e-03
GC_6_124 b_6 NI_6 NS_124 0 1.0677175420320633e-02
GC_6_125 b_6 NI_6 NS_125 0 -3.0034911493637716e-05
GC_6_126 b_6 NI_6 NS_126 0 -2.0695126903528899e-06
GC_6_127 b_6 NI_6 NS_127 0 1.6169355974683705e-02
GC_6_128 b_6 NI_6 NS_128 0 -1.6385293973133777e-02
GC_6_129 b_6 NI_6 NS_129 0 -4.0273889922263768e-06
GC_6_130 b_6 NI_6 NS_130 0 1.3209526169688926e-05
GC_6_131 b_6 NI_6 NS_131 0 -2.0938410382263143e-05
GC_6_132 b_6 NI_6 NS_132 0 3.0007510323593079e-05
GC_6_133 b_6 NI_6 NS_133 0 1.5415329297651159e-05
GC_6_134 b_6 NI_6 NS_134 0 -3.3136707913854019e-06
GC_6_135 b_6 NI_6 NS_135 0 -1.2480173427360174e-05
GC_6_136 b_6 NI_6 NS_136 0 7.0579616439376450e-06
GC_6_137 b_6 NI_6 NS_137 0 -4.4794478254405641e-03
GC_6_138 b_6 NI_6 NS_138 0 2.4824909097018091e-03
GC_6_139 b_6 NI_6 NS_139 0 2.3590161818358890e-05
GC_6_140 b_6 NI_6 NS_140 0 -7.3605060328711550e-04
GC_6_141 b_6 NI_6 NS_141 0 3.2318228897186812e-04
GC_6_142 b_6 NI_6 NS_142 0 -4.2596740350556828e-04
GC_6_143 b_6 NI_6 NS_143 0 -7.6483272272492170e-05
GC_6_144 b_6 NI_6 NS_144 0 6.3435809244885910e-05
GC_6_145 b_6 NI_6 NS_145 0 6.4449089480138030e-06
GC_6_146 b_6 NI_6 NS_146 0 -3.1301388544875430e-05
GC_6_147 b_6 NI_6 NS_147 0 -1.9256637646027549e-05
GC_6_148 b_6 NI_6 NS_148 0 -9.9539770090668951e-06
GC_6_149 b_6 NI_6 NS_149 0 3.1383555308585167e-05
GC_6_150 b_6 NI_6 NS_150 0 9.2401336950679393e-05
GC_6_151 b_6 NI_6 NS_151 0 6.8905533651532561e-06
GC_6_152 b_6 NI_6 NS_152 0 1.2903108470830523e-05
GC_6_153 b_6 NI_6 NS_153 0 -2.1745834046004400e-02
GC_6_154 b_6 NI_6 NS_154 0 2.3989590655086874e-03
GC_6_155 b_6 NI_6 NS_155 0 3.8825843998651036e-02
GC_6_156 b_6 NI_6 NS_156 0 -5.8368559665246964e-03
GC_6_157 b_6 NI_6 NS_157 0 9.1005624035676001e-04
GC_6_158 b_6 NI_6 NS_158 0 5.6567779879795192e-05
GC_6_159 b_6 NI_6 NS_159 0 4.1684809742348629e-05
GC_6_160 b_6 NI_6 NS_160 0 -7.4955169525318750e-06
GC_6_161 b_6 NI_6 NS_161 0 3.6784426181686196e-02
GC_6_162 b_6 NI_6 NS_162 0 2.6844130346292905e-02
GC_6_163 b_6 NI_6 NS_163 0 2.9071436407629110e-05
GC_6_164 b_6 NI_6 NS_164 0 2.8921787919690581e-06
GC_6_165 b_6 NI_6 NS_165 0 -4.2909198152744139e-02
GC_6_166 b_6 NI_6 NS_166 0 2.1736354639412252e-02
GC_6_167 b_6 NI_6 NS_167 0 2.5196998414086705e-06
GC_6_168 b_6 NI_6 NS_168 0 1.0165348077836269e-05
GC_6_169 b_6 NI_6 NS_169 0 -9.0816122680975926e-07
GC_6_170 b_6 NI_6 NS_170 0 4.2851384694635271e-05
GC_6_171 b_6 NI_6 NS_171 0 1.4274262834426277e-07
GC_6_172 b_6 NI_6 NS_172 0 2.4290094309533522e-06
GC_6_173 b_6 NI_6 NS_173 0 7.4781608597825887e-09
GC_6_174 b_6 NI_6 NS_174 0 1.3773641616609153e-06
GC_6_175 b_6 NI_6 NS_175 0 -1.4315060264607055e-03
GC_6_176 b_6 NI_6 NS_176 0 4.2304523236850111e-03
GC_6_177 b_6 NI_6 NS_177 0 -4.5169519781934321e-04
GC_6_178 b_6 NI_6 NS_178 0 -4.4265543301014117e-04
GC_6_179 b_6 NI_6 NS_179 0 2.0190827442126113e-05
GC_6_180 b_6 NI_6 NS_180 0 -4.7709261777012822e-04
GC_6_181 b_6 NI_6 NS_181 0 -1.5234987500326455e-05
GC_6_182 b_6 NI_6 NS_182 0 1.7022630015282929e-04
GC_6_183 b_6 NI_6 NS_183 0 1.0710109813856949e-04
GC_6_184 b_6 NI_6 NS_184 0 1.2874252169460537e-05
GC_6_185 b_6 NI_6 NS_185 0 2.8948883795527483e-05
GC_6_186 b_6 NI_6 NS_186 0 -1.3241395338769503e-06
GC_6_187 b_6 NI_6 NS_187 0 2.0427696541343778e-04
GC_6_188 b_6 NI_6 NS_188 0 1.6541943896672602e-04
GC_6_189 b_6 NI_6 NS_189 0 1.0472500281365230e-04
GC_6_190 b_6 NI_6 NS_190 0 -7.7255590259628303e-05
GC_6_191 b_6 NI_6 NS_191 0 1.0994077786447423e-01
GC_6_192 b_6 NI_6 NS_192 0 -1.7455538146149275e-03
GC_6_193 b_6 NI_6 NS_193 0 1.5519177910829799e-02
GC_6_194 b_6 NI_6 NS_194 0 -5.6898240288479361e-02
GC_6_195 b_6 NI_6 NS_195 0 2.7536936671218023e-04
GC_6_196 b_6 NI_6 NS_196 0 -5.1701592008524715e-04
GC_6_197 b_6 NI_6 NS_197 0 4.1652644769935855e-05
GC_6_198 b_6 NI_6 NS_198 0 -6.8937446673382493e-05
GC_6_199 b_6 NI_6 NS_199 0 -1.7131915854760048e-02
GC_6_200 b_6 NI_6 NS_200 0 -1.8515945255155606e-03
GC_6_201 b_6 NI_6 NS_201 0 -1.3956468696667150e-05
GC_6_202 b_6 NI_6 NS_202 0 5.0221502200863603e-06
GC_6_203 b_6 NI_6 NS_203 0 -3.2526568309791226e-02
GC_6_204 b_6 NI_6 NS_204 0 1.6751006412242374e-02
GC_6_205 b_6 NI_6 NS_205 0 2.2423342302425366e-05
GC_6_206 b_6 NI_6 NS_206 0 -9.1029074500068392e-06
GC_6_207 b_6 NI_6 NS_207 0 7.2019102792375683e-06
GC_6_208 b_6 NI_6 NS_208 0 1.3673000962794939e-05
GC_6_209 b_6 NI_6 NS_209 0 5.8328899969460352e-06
GC_6_210 b_6 NI_6 NS_210 0 2.1875740713032747e-06
GC_6_211 b_6 NI_6 NS_211 0 1.1718536295253341e-06
GC_6_212 b_6 NI_6 NS_212 0 3.7787206987476339e-06
GC_6_213 b_6 NI_6 NS_213 0 -1.5401848153993156e-03
GC_6_214 b_6 NI_6 NS_214 0 4.1986615084338968e-03
GC_6_215 b_6 NI_6 NS_215 0 -2.8321992524984248e-04
GC_6_216 b_6 NI_6 NS_216 0 -3.7393824938184556e-04
GC_6_217 b_6 NI_6 NS_217 0 8.2277785809938697e-05
GC_6_218 b_6 NI_6 NS_218 0 -3.8230067520412039e-04
GC_6_219 b_6 NI_6 NS_219 0 -1.3980552672837969e-05
GC_6_220 b_6 NI_6 NS_220 0 1.2787294197505513e-04
GC_6_221 b_6 NI_6 NS_221 0 -2.4459991788184200e-05
GC_6_222 b_6 NI_6 NS_222 0 9.4118724338116867e-05
GC_6_223 b_6 NI_6 NS_223 0 9.9844994967619177e-06
GC_6_224 b_6 NI_6 NS_224 0 4.9041229197334953e-05
GC_6_225 b_6 NI_6 NS_225 0 1.5545181174459103e-04
GC_6_226 b_6 NI_6 NS_226 0 1.9072904449153868e-04
GC_6_227 b_6 NI_6 NS_227 0 1.0158206665301236e-04
GC_6_228 b_6 NI_6 NS_228 0 -2.2589185519967071e-05
GC_6_229 b_6 NI_6 NS_229 0 -4.7632657306742937e-03
GC_6_230 b_6 NI_6 NS_230 0 1.1838539911753793e-03
GC_6_231 b_6 NI_6 NS_231 0 -8.5305977930474272e-03
GC_6_232 b_6 NI_6 NS_232 0 -7.7284585353482975e-03
GC_6_233 b_6 NI_6 NS_233 0 -8.4684168395311927e-04
GC_6_234 b_6 NI_6 NS_234 0 7.5699160590785117e-04
GC_6_235 b_6 NI_6 NS_235 0 -6.4647184136860862e-05
GC_6_236 b_6 NI_6 NS_236 0 7.5006038547921657e-05
GC_6_237 b_6 NI_6 NS_237 0 -1.2298634047262504e-02
GC_6_238 b_6 NI_6 NS_238 0 -1.9887203737037489e-02
GC_6_239 b_6 NI_6 NS_239 0 -1.3677590782015585e-06
GC_6_240 b_6 NI_6 NS_240 0 -4.4368549678184122e-06
GC_6_241 b_6 NI_6 NS_241 0 1.3302945581129740e-02
GC_6_242 b_6 NI_6 NS_242 0 -1.5602803572070723e-02
GC_6_243 b_6 NI_6 NS_243 0 -3.6834928307845389e-05
GC_6_244 b_6 NI_6 NS_244 0 1.9926553206573709e-05
GC_6_245 b_6 NI_6 NS_245 0 -2.4867960648707335e-05
GC_6_246 b_6 NI_6 NS_246 0 3.4766566862742271e-05
GC_6_247 b_6 NI_6 NS_247 0 -1.8572325110472487e-05
GC_6_248 b_6 NI_6 NS_248 0 -6.5354527762376022e-06
GC_6_249 b_6 NI_6 NS_249 0 -6.5315417342349465e-08
GC_6_250 b_6 NI_6 NS_250 0 -3.5490755835153510e-06
GC_6_251 b_6 NI_6 NS_251 0 -3.1051608283568927e-03
GC_6_252 b_6 NI_6 NS_252 0 8.3221145296858440e-03
GC_6_253 b_6 NI_6 NS_253 0 -5.6527848020128228e-04
GC_6_254 b_6 NI_6 NS_254 0 -4.8607027766236051e-04
GC_6_255 b_6 NI_6 NS_255 0 2.5484804925910825e-04
GC_6_256 b_6 NI_6 NS_256 0 -5.0304004532042228e-04
GC_6_257 b_6 NI_6 NS_257 0 -2.8974802158225725e-06
GC_6_258 b_6 NI_6 NS_258 0 1.4068398074249817e-06
GC_6_259 b_6 NI_6 NS_259 0 5.7684704585646729e-05
GC_6_260 b_6 NI_6 NS_260 0 2.6390552606096882e-06
GC_6_261 b_6 NI_6 NS_261 0 1.0043004959814347e-05
GC_6_262 b_6 NI_6 NS_262 0 9.8196423512503278e-06
GC_6_263 b_6 NI_6 NS_263 0 6.5296925776613986e-05
GC_6_264 b_6 NI_6 NS_264 0 -4.0288371820707745e-05
GC_6_265 b_6 NI_6 NS_265 0 -9.9263695421574281e-06
GC_6_266 b_6 NI_6 NS_266 0 4.7257457385976639e-05
GC_6_267 b_6 NI_6 NS_267 0 2.9573265372323004e-02
GC_6_268 b_6 NI_6 NS_268 0 -1.4830406805773091e-03
GC_6_269 b_6 NI_6 NS_269 0 -1.2646239670250392e-02
GC_6_270 b_6 NI_6 NS_270 0 -6.0727356500991734e-03
GC_6_271 b_6 NI_6 NS_271 0 -3.1108993126685023e-05
GC_6_272 b_6 NI_6 NS_272 0 8.2220541461455488e-05
GC_6_273 b_6 NI_6 NS_273 0 -2.7396171835854671e-05
GC_6_274 b_6 NI_6 NS_274 0 3.6324090574262785e-06
GC_6_275 b_6 NI_6 NS_275 0 -4.4080161259694161e-05
GC_6_276 b_6 NI_6 NS_276 0 6.8137819574874553e-03
GC_6_277 b_6 NI_6 NS_277 0 -1.0403977004889512e-05
GC_6_278 b_6 NI_6 NS_278 0 3.1435323065702799e-06
GC_6_279 b_6 NI_6 NS_279 0 2.6202222640735477e-04
GC_6_280 b_6 NI_6 NS_280 0 -2.0575938581500492e-03
GC_6_281 b_6 NI_6 NS_281 0 -2.6268763252759796e-06
GC_6_282 b_6 NI_6 NS_282 0 9.4009084822871909e-06
GC_6_283 b_6 NI_6 NS_283 0 -1.4027405044686212e-05
GC_6_284 b_6 NI_6 NS_284 0 2.1783417539410715e-05
GC_6_285 b_6 NI_6 NS_285 0 -6.7500488409395686e-06
GC_6_286 b_6 NI_6 NS_286 0 -3.2851299791145545e-06
GC_6_287 b_6 NI_6 NS_287 0 -1.9503603921165499e-06
GC_6_288 b_6 NI_6 NS_288 0 1.5638322922314446e-06
GC_6_289 b_6 NI_6 NS_289 0 -2.8256108555331713e-03
GC_6_290 b_6 NI_6 NS_290 0 6.3954168080005711e-03
GC_6_291 b_6 NI_6 NS_291 0 -3.3374213518554640e-04
GC_6_292 b_6 NI_6 NS_292 0 -4.0864189890217834e-04
GC_6_293 b_6 NI_6 NS_293 0 2.9717058866606769e-04
GC_6_294 b_6 NI_6 NS_294 0 -3.2384159449768660e-04
GC_6_295 b_6 NI_6 NS_295 0 8.1266289352747392e-07
GC_6_296 b_6 NI_6 NS_296 0 2.5926503611537796e-05
GC_6_297 b_6 NI_6 NS_297 0 2.8552509586982133e-05
GC_6_298 b_6 NI_6 NS_298 0 5.5689693252509735e-05
GC_6_299 b_6 NI_6 NS_299 0 -7.3161748597333670e-06
GC_6_300 b_6 NI_6 NS_300 0 2.6861154563946500e-05
GC_6_301 b_6 NI_6 NS_301 0 6.4896431114341719e-05
GC_6_302 b_6 NI_6 NS_302 0 1.9837264967500716e-05
GC_6_303 b_6 NI_6 NS_303 0 -2.5470615851828096e-05
GC_6_304 b_6 NI_6 NS_304 0 3.6591043502717720e-05
GC_6_305 b_6 NI_6 NS_305 0 1.9369909629872239e-02
GC_6_306 b_6 NI_6 NS_306 0 1.3407412022835689e-03
GC_6_307 b_6 NI_6 NS_307 0 -1.1044775996933166e-02
GC_6_308 b_6 NI_6 NS_308 0 1.4728923974422884e-03
GC_6_309 b_6 NI_6 NS_309 0 -1.1275844141838515e-05
GC_6_310 b_6 NI_6 NS_310 0 6.0770032318208404e-04
GC_6_311 b_6 NI_6 NS_311 0 8.5155895502543125e-05
GC_6_312 b_6 NI_6 NS_312 0 3.9725735957245731e-05
GC_6_313 b_6 NI_6 NS_313 0 -7.2712313392968983e-03
GC_6_314 b_6 NI_6 NS_314 0 -4.6381228628405323e-03
GC_6_315 b_6 NI_6 NS_315 0 1.5243695786292264e-05
GC_6_316 b_6 NI_6 NS_316 0 2.7639549077002876e-06
GC_6_317 b_6 NI_6 NS_317 0 9.1275239220895664e-03
GC_6_318 b_6 NI_6 NS_318 0 -2.0116831025425433e-03
GC_6_319 b_6 NI_6 NS_319 0 1.9256185416612392e-05
GC_6_320 b_6 NI_6 NS_320 0 5.2898244886827429e-06
GC_6_321 b_6 NI_6 NS_321 0 -7.3249648691590445e-06
GC_6_322 b_6 NI_6 NS_322 0 3.9500945248384934e-05
GC_6_323 b_6 NI_6 NS_323 0 -2.2515948247121324e-05
GC_6_324 b_6 NI_6 NS_324 0 2.3587783336450142e-06
GC_6_325 b_6 NI_6 NS_325 0 1.0456075804579020e-05
GC_6_326 b_6 NI_6 NS_326 0 9.3929438819339596e-07
GC_6_327 b_6 NI_6 NS_327 0 -3.7796322598851496e-03
GC_6_328 b_6 NI_6 NS_328 0 2.2710433461240859e-03
GC_6_329 b_6 NI_6 NS_329 0 -1.6970497799358931e-04
GC_6_330 b_6 NI_6 NS_330 0 -3.9401925323042595e-04
GC_6_331 b_6 NI_6 NS_331 0 3.5638377145190392e-04
GC_6_332 b_6 NI_6 NS_332 0 -1.0417228147177746e-04
GC_6_333 b_6 NI_6 NS_333 0 2.1208569320225164e-05
GC_6_334 b_6 NI_6 NS_334 0 3.6309526965525646e-05
GC_6_335 b_6 NI_6 NS_335 0 -3.7965170420297923e-05
GC_6_336 b_6 NI_6 NS_336 0 2.2866307674457229e-05
GC_6_337 b_6 NI_6 NS_337 0 2.4354863670587275e-05
GC_6_338 b_6 NI_6 NS_338 0 3.1140607950157735e-05
GC_6_339 b_6 NI_6 NS_339 0 1.0021656663905051e-05
GC_6_340 b_6 NI_6 NS_340 0 1.0974691213020169e-04
GC_6_341 b_6 NI_6 NS_341 0 4.5625954127870879e-05
GC_6_342 b_6 NI_6 NS_342 0 2.0910946290219847e-05
GC_6_343 b_6 NI_6 NS_343 0 -8.9008808012522034e-03
GC_6_344 b_6 NI_6 NS_344 0 -1.3474895493992716e-03
GC_6_345 b_6 NI_6 NS_345 0 -2.0239223181490102e-03
GC_6_346 b_6 NI_6 NS_346 0 5.2287504723692365e-03
GC_6_347 b_6 NI_6 NS_347 0 -1.3293310109261858e-04
GC_6_348 b_6 NI_6 NS_348 0 2.0824799143282120e-04
GC_6_349 b_6 NI_6 NS_349 0 1.3275388490901689e-05
GC_6_350 b_6 NI_6 NS_350 0 3.3543679200831970e-05
GC_6_351 b_6 NI_6 NS_351 0 5.4760874488108211e-03
GC_6_352 b_6 NI_6 NS_352 0 2.7344701917840757e-03
GC_6_353 b_6 NI_6 NS_353 0 -1.4215157487167172e-05
GC_6_354 b_6 NI_6 NS_354 0 -1.6308133605897898e-06
GC_6_355 b_6 NI_6 NS_355 0 1.0116172779217275e-02
GC_6_356 b_6 NI_6 NS_356 0 -2.6917829508136698e-03
GC_6_357 b_6 NI_6 NS_357 0 1.3808184062339493e-05
GC_6_358 b_6 NI_6 NS_358 0 3.4374978849480493e-06
GC_6_359 b_6 NI_6 NS_359 0 -1.3984658688510413e-05
GC_6_360 b_6 NI_6 NS_360 0 3.4101812882519303e-05
GC_6_361 b_6 NI_6 NS_361 0 -1.2076039100346454e-05
GC_6_362 b_6 NI_6 NS_362 0 1.4372412453849523e-06
GC_6_363 b_6 NI_6 NS_363 0 9.1382312730643502e-06
GC_6_364 b_6 NI_6 NS_364 0 -6.7045380129544535e-08
GC_6_365 b_6 NI_6 NS_365 0 -3.3305839540494304e-03
GC_6_366 b_6 NI_6 NS_366 0 1.8528990606476010e-03
GC_6_367 b_6 NI_6 NS_367 0 4.9296604309937715e-06
GC_6_368 b_6 NI_6 NS_368 0 -4.6465916805445845e-04
GC_6_369 b_6 NI_6 NS_369 0 2.6858814370679988e-04
GC_6_370 b_6 NI_6 NS_370 0 -1.0414749630121421e-04
GC_6_371 b_6 NI_6 NS_371 0 4.8024677708898284e-05
GC_6_372 b_6 NI_6 NS_372 0 2.2857005649919665e-05
GC_6_373 b_6 NI_6 NS_373 0 7.0158416807869337e-06
GC_6_374 b_6 NI_6 NS_374 0 8.6173697951948342e-06
GC_6_375 b_6 NI_6 NS_375 0 1.8426448747428837e-05
GC_6_376 b_6 NI_6 NS_376 0 -1.1066141628106752e-06
GC_6_377 b_6 NI_6 NS_377 0 7.2414831215975758e-05
GC_6_378 b_6 NI_6 NS_378 0 -2.6824817425046697e-05
GC_6_379 b_6 NI_6 NS_379 0 9.9526931271987942e-07
GC_6_380 b_6 NI_6 NS_380 0 -4.1646978266789801e-05
GC_6_381 b_6 NI_6 NS_381 0 1.3114822262731397e-02
GC_6_382 b_6 NI_6 NS_382 0 1.1287923020912032e-03
GC_6_383 b_6 NI_6 NS_383 0 -1.0788723994419148e-02
GC_6_384 b_6 NI_6 NS_384 0 2.9521823125523952e-03
GC_6_385 b_6 NI_6 NS_385 0 2.9915111186120606e-04
GC_6_386 b_6 NI_6 NS_386 0 5.1595063720602237e-05
GC_6_387 b_6 NI_6 NS_387 0 8.4650006481452335e-05
GC_6_388 b_6 NI_6 NS_388 0 -1.4000916287810981e-05
GC_6_389 b_6 NI_6 NS_389 0 -2.0500065196476930e-03
GC_6_390 b_6 NI_6 NS_390 0 5.4371887755825365e-03
GC_6_391 b_6 NI_6 NS_391 0 1.8062075895192225e-05
GC_6_392 b_6 NI_6 NS_392 0 3.7088548662153396e-06
GC_6_393 b_6 NI_6 NS_393 0 5.7156272317106394e-03
GC_6_394 b_6 NI_6 NS_394 0 1.4786652268326795e-03
GC_6_395 b_6 NI_6 NS_395 0 3.4123296497911372e-05
GC_6_396 b_6 NI_6 NS_396 0 -2.7369729762554623e-07
GC_6_397 b_6 NI_6 NS_397 0 1.5640866446113549e-05
GC_6_398 b_6 NI_6 NS_398 0 1.1835072281932096e-05
GC_6_399 b_6 NI_6 NS_399 0 -2.3477141850726409e-05
GC_6_400 b_6 NI_6 NS_400 0 5.6195406368427391e-06
GC_6_401 b_6 NI_6 NS_401 0 8.5408221840995819e-06
GC_6_402 b_6 NI_6 NS_402 0 2.0225199225223345e-06
GC_6_403 b_6 NI_6 NS_403 0 -1.5488780184866743e-03
GC_6_404 b_6 NI_6 NS_404 0 4.1444040954818423e-04
GC_6_405 b_6 NI_6 NS_405 0 -1.3079521279808255e-04
GC_6_406 b_6 NI_6 NS_406 0 -5.4859077004818657e-05
GC_6_407 b_6 NI_6 NS_407 0 4.1675144403812705e-04
GC_6_408 b_6 NI_6 NS_408 0 2.3956983153773285e-04
GC_6_409 b_6 NI_6 NS_409 0 1.1903815705454928e-04
GC_6_410 b_6 NI_6 NS_410 0 -7.5516102275430041e-05
GC_6_411 b_6 NI_6 NS_411 0 -7.8642594342417767e-05
GC_6_412 b_6 NI_6 NS_412 0 -8.6887226570406744e-06
GC_6_413 b_6 NI_6 NS_413 0 4.2193945460612430e-05
GC_6_414 b_6 NI_6 NS_414 0 2.8009008894201596e-06
GC_6_415 b_6 NI_6 NS_415 0 -8.2703259167231185e-05
GC_6_416 b_6 NI_6 NS_416 0 -1.4121230860155231e-05
GC_6_417 b_6 NI_6 NS_417 0 -4.6013314241779921e-07
GC_6_418 b_6 NI_6 NS_418 0 -8.3682007542153606e-07
GC_6_419 b_6 NI_6 NS_419 0 -1.4088239326185917e-02
GC_6_420 b_6 NI_6 NS_420 0 -1.0866960669580082e-03
GC_6_421 b_6 NI_6 NS_421 0 1.3249442864496186e-03
GC_6_422 b_6 NI_6 NS_422 0 6.5898049814732754e-03
GC_6_423 b_6 NI_6 NS_423 0 1.1234248528794288e-04
GC_6_424 b_6 NI_6 NS_424 0 -6.0400334273695054e-06
GC_6_425 b_6 NI_6 NS_425 0 3.1672228217890750e-05
GC_6_426 b_6 NI_6 NS_426 0 2.9922279440085992e-05
GC_6_427 b_6 NI_6 NS_427 0 4.1149083185229316e-03
GC_6_428 b_6 NI_6 NS_428 0 -2.8040841273188660e-03
GC_6_429 b_6 NI_6 NS_429 0 -1.4314235365058203e-05
GC_6_430 b_6 NI_6 NS_430 0 -3.3588002410298285e-06
GC_6_431 b_6 NI_6 NS_431 0 8.5415946498472797e-03
GC_6_432 b_6 NI_6 NS_432 0 -4.8280732772959479e-03
GC_6_433 b_6 NI_6 NS_433 0 2.7116332238298046e-05
GC_6_434 b_6 NI_6 NS_434 0 7.1724483729699051e-06
GC_6_435 b_6 NI_6 NS_435 0 2.5055900516646149e-06
GC_6_436 b_6 NI_6 NS_436 0 2.2520618958433174e-05
GC_6_437 b_6 NI_6 NS_437 0 -1.7152523453575313e-05
GC_6_438 b_6 NI_6 NS_438 0 3.5290025261798042e-07
GC_6_439 b_6 NI_6 NS_439 0 6.5611811125495906e-06
GC_6_440 b_6 NI_6 NS_440 0 8.9861627068691186e-07
GC_6_441 b_6 NI_6 NS_441 0 -2.2232126197347987e-03
GC_6_442 b_6 NI_6 NS_442 0 1.7052796350615475e-03
GC_6_443 b_6 NI_6 NS_443 0 -2.2113546143513527e-06
GC_6_444 b_6 NI_6 NS_444 0 -3.1733486024637393e-04
GC_6_445 b_6 NI_6 NS_445 0 3.2575365247305965e-04
GC_6_446 b_6 NI_6 NS_446 0 1.2930465623372072e-04
GC_6_447 b_6 NI_6 NS_447 0 1.0804770674744857e-04
GC_6_448 b_6 NI_6 NS_448 0 -1.4473104946667723e-05
GC_6_449 b_6 NI_6 NS_449 0 -5.1592111448075151e-05
GC_6_450 b_6 NI_6 NS_450 0 -3.5809389137294981e-05
GC_6_451 b_6 NI_6 NS_451 0 2.7366968295980925e-05
GC_6_452 b_6 NI_6 NS_452 0 8.9972442812585297e-06
GC_6_453 b_6 NI_6 NS_453 0 -4.2073849390425144e-05
GC_6_454 b_6 NI_6 NS_454 0 -7.9946235798332259e-05
GC_6_455 b_6 NI_6 NS_455 0 -1.4389390620000891e-06
GC_6_456 b_6 NI_6 NS_456 0 -1.2323660978436695e-05
GD_6_1 b_6 NI_6 NA_1 0 -2.7828143504066158e-03
GD_6_2 b_6 NI_6 NA_2 0 2.3091107714769718e-04
GD_6_3 b_6 NI_6 NA_3 0 9.4849778154454667e-03
GD_6_4 b_6 NI_6 NA_4 0 -9.2659617208638665e-03
GD_6_5 b_6 NI_6 NA_5 0 -2.3084971838870136e-02
GD_6_6 b_6 NI_6 NA_6 0 -1.3701910501188355e-01
GD_6_7 b_6 NI_6 NA_7 0 2.0712623491270864e-02
GD_6_8 b_6 NI_6 NA_8 0 -5.9230083529004289e-03
GD_6_9 b_6 NI_6 NA_9 0 -7.2428147893526815e-03
GD_6_10 b_6 NI_6 NA_10 0 -1.6041207598697745e-04
GD_6_11 b_6 NI_6 NA_11 0 -5.6239217663542149e-03
GD_6_12 b_6 NI_6 NA_12 0 1.9761339788354447e-03
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 -1.4591039430947786e-02
GC_7_2 b_7 NI_7 NS_2 0 -9.7658055059331541e-04
GC_7_3 b_7 NI_7 NS_3 0 2.8852077840686502e-03
GC_7_4 b_7 NI_7 NS_4 0 1.0660650208638290e-02
GC_7_5 b_7 NI_7 NS_5 0 2.8906286199022543e-04
GC_7_6 b_7 NI_7 NS_6 0 -3.1790785783180367e-04
GC_7_7 b_7 NI_7 NS_7 0 5.7953693887811940e-05
GC_7_8 b_7 NI_7 NS_8 0 -8.9831698024520998e-06
GC_7_9 b_7 NI_7 NS_9 0 4.5969255258397172e-03
GC_7_10 b_7 NI_7 NS_10 0 -1.0911750089335076e-03
GC_7_11 b_7 NI_7 NS_11 0 -1.6371457080036895e-05
GC_7_12 b_7 NI_7 NS_12 0 3.5436117171179700e-06
GC_7_13 b_7 NI_7 NS_13 0 8.0994824451304358e-03
GC_7_14 b_7 NI_7 NS_14 0 -7.9715055066193075e-03
GC_7_15 b_7 NI_7 NS_15 0 -1.0754307088694789e-05
GC_7_16 b_7 NI_7 NS_16 0 2.8772909836960188e-06
GC_7_17 b_7 NI_7 NS_17 0 -1.7133823683918201e-05
GC_7_18 b_7 NI_7 NS_18 0 2.9860727726392600e-05
GC_7_19 b_7 NI_7 NS_19 0 3.7297693335812393e-05
GC_7_20 b_7 NI_7 NS_20 0 1.4573826510669856e-05
GC_7_21 b_7 NI_7 NS_21 0 2.3374286200376675e-06
GC_7_22 b_7 NI_7 NS_22 0 1.1095279742526186e-05
GC_7_23 b_7 NI_7 NS_23 0 2.6661279764482102e-04
GC_7_24 b_7 NI_7 NS_24 0 2.8025820877883123e-03
GC_7_25 b_7 NI_7 NS_25 0 -4.8458544112522315e-04
GC_7_26 b_7 NI_7 NS_26 0 -4.4663349170896596e-04
GC_7_27 b_7 NI_7 NS_27 0 -2.4748500617255577e-04
GC_7_28 b_7 NI_7 NS_28 0 -3.9011007671388252e-04
GC_7_29 b_7 NI_7 NS_29 0 -8.7726526472649798e-05
GC_7_30 b_7 NI_7 NS_30 0 3.5207544355866531e-04
GC_7_31 b_7 NI_7 NS_31 0 -2.8765151892729456e-05
GC_7_32 b_7 NI_7 NS_32 0 4.6273676925668970e-05
GC_7_33 b_7 NI_7 NS_33 0 1.2080954023670143e-05
GC_7_34 b_7 NI_7 NS_34 0 4.9149062650753473e-06
GC_7_35 b_7 NI_7 NS_35 0 -1.5958296707894682e-05
GC_7_36 b_7 NI_7 NS_36 0 8.6851713570332243e-05
GC_7_37 b_7 NI_7 NS_37 0 7.4550254093045947e-06
GC_7_38 b_7 NI_7 NS_38 0 -1.1848243012372821e-05
GC_7_39 b_7 NI_7 NS_39 0 9.5797274579637794e-03
GC_7_40 b_7 NI_7 NS_40 0 1.1362921366473502e-03
GC_7_41 b_7 NI_7 NS_41 0 -9.1222180329395934e-03
GC_7_42 b_7 NI_7 NS_42 0 5.8762687952091629e-03
GC_7_43 b_7 NI_7 NS_43 0 5.8317837863963239e-05
GC_7_44 b_7 NI_7 NS_44 0 6.7266213265939633e-05
GC_7_45 b_7 NI_7 NS_45 0 4.8866783032008899e-06
GC_7_46 b_7 NI_7 NS_46 0 -6.6602267616272374e-05
GC_7_47 b_7 NI_7 NS_47 0 -1.1382751734380883e-03
GC_7_48 b_7 NI_7 NS_48 0 6.6170703984179732e-03
GC_7_49 b_7 NI_7 NS_49 0 2.1092226113789361e-05
GC_7_50 b_7 NI_7 NS_50 0 7.7623620990658194e-07
GC_7_51 b_7 NI_7 NS_51 0 7.6360837826575422e-03
GC_7_52 b_7 NI_7 NS_52 0 -9.9560691936120176e-04
GC_7_53 b_7 NI_7 NS_53 0 1.3548836878607561e-05
GC_7_54 b_7 NI_7 NS_54 0 -1.8040040167328438e-05
GC_7_55 b_7 NI_7 NS_55 0 -6.0788735013486996e-06
GC_7_56 b_7 NI_7 NS_56 0 4.8589471192660978e-05
GC_7_57 b_7 NI_7 NS_57 0 1.0144241917143393e-05
GC_7_58 b_7 NI_7 NS_58 0 5.0180591204634060e-06
GC_7_59 b_7 NI_7 NS_59 0 6.2466646547757566e-06
GC_7_60 b_7 NI_7 NS_60 0 1.8153591569081980e-05
GC_7_61 b_7 NI_7 NS_61 0 -1.3092383322332770e-03
GC_7_62 b_7 NI_7 NS_62 0 2.3539068145778316e-03
GC_7_63 b_7 NI_7 NS_63 0 -1.6270977768932502e-04
GC_7_64 b_7 NI_7 NS_64 0 -6.2410769037255724e-04
GC_7_65 b_7 NI_7 NS_65 0 -4.0199953765321203e-05
GC_7_66 b_7 NI_7 NS_66 0 -4.2849867239029798e-04
GC_7_67 b_7 NI_7 NS_67 0 -8.5911551812560866e-05
GC_7_68 b_7 NI_7 NS_68 0 2.5324798329465464e-04
GC_7_69 b_7 NI_7 NS_69 0 -5.2747960491702451e-05
GC_7_70 b_7 NI_7 NS_70 0 2.7785313317617427e-06
GC_7_71 b_7 NI_7 NS_71 0 1.1869414351614081e-05
GC_7_72 b_7 NI_7 NS_72 0 8.1578857610943846e-06
GC_7_73 b_7 NI_7 NS_73 0 1.7327993700788851e-05
GC_7_74 b_7 NI_7 NS_74 0 6.5323147182124532e-05
GC_7_75 b_7 NI_7 NS_75 0 -1.3441361462984516e-05
GC_7_76 b_7 NI_7 NS_76 0 -2.4890730809086451e-05
GC_7_77 b_7 NI_7 NS_77 0 -1.4948248463461532e-02
GC_7_78 b_7 NI_7 NS_78 0 -1.3192706259983721e-03
GC_7_79 b_7 NI_7 NS_79 0 7.3863156286757339e-03
GC_7_80 b_7 NI_7 NS_80 0 1.1632345733802153e-02
GC_7_81 b_7 NI_7 NS_81 0 2.7340086753372187e-04
GC_7_82 b_7 NI_7 NS_82 0 4.0314973163680707e-04
GC_7_83 b_7 NI_7 NS_83 0 1.1059660825202290e-04
GC_7_84 b_7 NI_7 NS_84 0 4.2664613690145614e-05
GC_7_85 b_7 NI_7 NS_85 0 6.4063133492150755e-03
GC_7_86 b_7 NI_7 NS_86 0 3.6843272687977773e-03
GC_7_87 b_7 NI_7 NS_87 0 -1.5916833485211738e-05
GC_7_88 b_7 NI_7 NS_88 0 4.5528166410618609e-06
GC_7_89 b_7 NI_7 NS_89 0 9.7027095875884071e-03
GC_7_90 b_7 NI_7 NS_90 0 -8.5819826864380992e-03
GC_7_91 b_7 NI_7 NS_91 0 4.8954498937616184e-06
GC_7_92 b_7 NI_7 NS_92 0 3.5544329503547179e-05
GC_7_93 b_7 NI_7 NS_93 0 -1.5892109857427178e-05
GC_7_94 b_7 NI_7 NS_94 0 3.3464421294615727e-05
GC_7_95 b_7 NI_7 NS_95 0 3.6536315671004294e-05
GC_7_96 b_7 NI_7 NS_96 0 1.9463680783131911e-05
GC_7_97 b_7 NI_7 NS_97 0 2.2067272916012307e-06
GC_7_98 b_7 NI_7 NS_98 0 8.5370131434613556e-06
GC_7_99 b_7 NI_7 NS_99 0 -2.3718724775950032e-03
GC_7_100 b_7 NI_7 NS_100 0 2.7403022259772760e-03
GC_7_101 b_7 NI_7 NS_101 0 -4.5188584012324404e-04
GC_7_102 b_7 NI_7 NS_102 0 -4.1350773574039089e-04
GC_7_103 b_7 NI_7 NS_103 0 1.8327707241117807e-04
GC_7_104 b_7 NI_7 NS_104 0 -1.5941117763938441e-04
GC_7_105 b_7 NI_7 NS_105 0 2.1629174278441815e-05
GC_7_106 b_7 NI_7 NS_106 0 5.3189974798504938e-05
GC_7_107 b_7 NI_7 NS_107 0 9.8539765683223957e-06
GC_7_108 b_7 NI_7 NS_108 0 1.0981194963503939e-05
GC_7_109 b_7 NI_7 NS_109 0 2.1315752472903131e-06
GC_7_110 b_7 NI_7 NS_110 0 8.8401964699353915e-06
GC_7_111 b_7 NI_7 NS_111 0 4.7644035834303908e-05
GC_7_112 b_7 NI_7 NS_112 0 1.4610071661018845e-05
GC_7_113 b_7 NI_7 NS_113 0 7.0912135132987860e-06
GC_7_114 b_7 NI_7 NS_114 0 1.0019406203357358e-05
GC_7_115 b_7 NI_7 NS_115 0 1.9130790054337075e-02
GC_7_116 b_7 NI_7 NS_116 0 1.3328304558758147e-03
GC_7_117 b_7 NI_7 NS_117 0 -1.3764188946800097e-02
GC_7_118 b_7 NI_7 NS_118 0 6.4266401100535869e-03
GC_7_119 b_7 NI_7 NS_119 0 -3.0886927886213946e-04
GC_7_120 b_7 NI_7 NS_120 0 -7.8657093872683202e-05
GC_7_121 b_7 NI_7 NS_121 0 -1.5352813033027091e-05
GC_7_122 b_7 NI_7 NS_122 0 4.3631719422521753e-06
GC_7_123 b_7 NI_7 NS_123 0 -4.6961120787134556e-03
GC_7_124 b_7 NI_7 NS_124 0 -9.2008026549397271e-04
GC_7_125 b_7 NI_7 NS_125 0 1.8350372279492548e-05
GC_7_126 b_7 NI_7 NS_126 0 -1.1970604601772826e-06
GC_7_127 b_7 NI_7 NS_127 0 1.1931349163793814e-02
GC_7_128 b_7 NI_7 NS_128 0 9.1694644316643169e-04
GC_7_129 b_7 NI_7 NS_129 0 -5.8835638951700917e-06
GC_7_130 b_7 NI_7 NS_130 0 -1.2518223761967510e-05
GC_7_131 b_7 NI_7 NS_131 0 -5.3811163082872876e-06
GC_7_132 b_7 NI_7 NS_132 0 4.8502883470920306e-05
GC_7_133 b_7 NI_7 NS_133 0 1.9598194137975120e-05
GC_7_134 b_7 NI_7 NS_134 0 1.8926840081342172e-05
GC_7_135 b_7 NI_7 NS_135 0 6.6642187629042862e-06
GC_7_136 b_7 NI_7 NS_136 0 1.6179146985696948e-05
GC_7_137 b_7 NI_7 NS_137 0 -3.7345778026363938e-03
GC_7_138 b_7 NI_7 NS_138 0 1.7252066923856442e-03
GC_7_139 b_7 NI_7 NS_139 0 -1.0799806946569069e-04
GC_7_140 b_7 NI_7 NS_140 0 -6.4700217226983786e-04
GC_7_141 b_7 NI_7 NS_141 0 3.6372371820284137e-04
GC_7_142 b_7 NI_7 NS_142 0 -1.9917321978647694e-04
GC_7_143 b_7 NI_7 NS_143 0 -1.4366335878128976e-05
GC_7_144 b_7 NI_7 NS_144 0 3.8401983400048019e-05
GC_7_145 b_7 NI_7 NS_145 0 4.2523504481251161e-06
GC_7_146 b_7 NI_7 NS_146 0 3.7460609464263346e-06
GC_7_147 b_7 NI_7 NS_147 0 1.6991829423063963e-06
GC_7_148 b_7 NI_7 NS_148 0 1.2188882030769355e-05
GC_7_149 b_7 NI_7 NS_149 0 5.0773657789247703e-05
GC_7_150 b_7 NI_7 NS_150 0 1.6473765599626359e-05
GC_7_151 b_7 NI_7 NS_151 0 1.9250852681075274e-05
GC_7_152 b_7 NI_7 NS_152 0 -5.1454964696018956e-06
GC_7_153 b_7 NI_7 NS_153 0 2.6551105985365208e-02
GC_7_154 b_7 NI_7 NS_154 0 -1.4757388752052831e-03
GC_7_155 b_7 NI_7 NS_155 0 -6.1712372211028856e-03
GC_7_156 b_7 NI_7 NS_156 0 1.9720502815638256e-02
GC_7_157 b_7 NI_7 NS_157 0 -1.4235066297553159e-04
GC_7_158 b_7 NI_7 NS_158 0 1.0296618906411737e-03
GC_7_159 b_7 NI_7 NS_159 0 1.2377269919520544e-04
GC_7_160 b_7 NI_7 NS_160 0 6.8551102934550682e-05
GC_7_161 b_7 NI_7 NS_161 0 2.4205618401173705e-03
GC_7_162 b_7 NI_7 NS_162 0 6.0127969695976833e-03
GC_7_163 b_7 NI_7 NS_163 0 -9.5948552136531567e-06
GC_7_164 b_7 NI_7 NS_164 0 1.4383156852727286e-06
GC_7_165 b_7 NI_7 NS_165 0 1.6850290464837020e-02
GC_7_166 b_7 NI_7 NS_166 0 -1.2033678085478549e-02
GC_7_167 b_7 NI_7 NS_167 0 5.6735604419411063e-06
GC_7_168 b_7 NI_7 NS_168 0 5.8072186278396912e-05
GC_7_169 b_7 NI_7 NS_169 0 -2.5090032761234943e-05
GC_7_170 b_7 NI_7 NS_170 0 4.1323735968120821e-05
GC_7_171 b_7 NI_7 NS_171 0 -2.2207425061440676e-06
GC_7_172 b_7 NI_7 NS_172 0 -1.1920829753393022e-05
GC_7_173 b_7 NI_7 NS_173 0 -2.8888927125489576e-06
GC_7_174 b_7 NI_7 NS_174 0 -3.8367325322392859e-06
GC_7_175 b_7 NI_7 NS_175 0 -3.6730193222489532e-03
GC_7_176 b_7 NI_7 NS_176 0 8.2082606429911120e-03
GC_7_177 b_7 NI_7 NS_177 0 -7.3826905641672204e-04
GC_7_178 b_7 NI_7 NS_178 0 -5.4546509215744094e-04
GC_7_179 b_7 NI_7 NS_179 0 2.4652091005311340e-04
GC_7_180 b_7 NI_7 NS_180 0 -5.9443277937992192e-04
GC_7_181 b_7 NI_7 NS_181 0 -6.5436579030617211e-05
GC_7_182 b_7 NI_7 NS_182 0 1.1342642287878412e-05
GC_7_183 b_7 NI_7 NS_183 0 7.0676516732097656e-06
GC_7_184 b_7 NI_7 NS_184 0 -6.3151290720065011e-05
GC_7_185 b_7 NI_7 NS_185 0 2.8910893455744494e-05
GC_7_186 b_7 NI_7 NS_186 0 1.0863495146474084e-05
GC_7_187 b_7 NI_7 NS_187 0 3.0543311263083358e-05
GC_7_188 b_7 NI_7 NS_188 0 -4.8050873840168312e-05
GC_7_189 b_7 NI_7 NS_189 0 2.5507774239867824e-05
GC_7_190 b_7 NI_7 NS_190 0 3.9155712735015328e-05
GC_7_191 b_7 NI_7 NS_191 0 -4.7631775280434522e-03
GC_7_192 b_7 NI_7 NS_192 0 1.1838527108322951e-03
GC_7_193 b_7 NI_7 NS_193 0 -8.5306096678109469e-03
GC_7_194 b_7 NI_7 NS_194 0 -7.7284702072623239e-03
GC_7_195 b_7 NI_7 NS_195 0 -8.4684306955726989e-04
GC_7_196 b_7 NI_7 NS_196 0 7.5699168186039209e-04
GC_7_197 b_7 NI_7 NS_197 0 -6.4647416638296691e-05
GC_7_198 b_7 NI_7 NS_198 0 7.5006208940088355e-05
GC_7_199 b_7 NI_7 NS_199 0 -1.2298649327006110e-02
GC_7_200 b_7 NI_7 NS_200 0 -1.9887235737960095e-02
GC_7_201 b_7 NI_7 NS_201 0 -1.3677627369834707e-06
GC_7_202 b_7 NI_7 NS_202 0 -4.4368919178793024e-06
GC_7_203 b_7 NI_7 NS_203 0 1.3302923062922332e-02
GC_7_204 b_7 NI_7 NS_204 0 -1.5602780948391012e-02
GC_7_205 b_7 NI_7 NS_205 0 -3.6835016269748985e-05
GC_7_206 b_7 NI_7 NS_206 0 1.9926615380469904e-05
GC_7_207 b_7 NI_7 NS_207 0 -2.4868024843674796e-05
GC_7_208 b_7 NI_7 NS_208 0 3.4766611965720549e-05
GC_7_209 b_7 NI_7 NS_209 0 -1.8572373067132617e-05
GC_7_210 b_7 NI_7 NS_210 0 -6.5354434205385161e-06
GC_7_211 b_7 NI_7 NS_211 0 -6.5333652653461291e-08
GC_7_212 b_7 NI_7 NS_212 0 -3.5490892559510678e-06
GC_7_213 b_7 NI_7 NS_213 0 -3.1051564136441493e-03
GC_7_214 b_7 NI_7 NS_214 0 8.3221024995597508e-03
GC_7_215 b_7 NI_7 NS_215 0 -5.6527908221618006e-04
GC_7_216 b_7 NI_7 NS_216 0 -4.8606855280435490e-04
GC_7_217 b_7 NI_7 NS_217 0 2.5484804353981228e-04
GC_7_218 b_7 NI_7 NS_218 0 -5.0303752134977641e-04
GC_7_219 b_7 NI_7 NS_219 0 -2.8968904336502982e-06
GC_7_220 b_7 NI_7 NS_220 0 1.4068026191536544e-06
GC_7_221 b_7 NI_7 NS_221 0 5.7684659925864360e-05
GC_7_222 b_7 NI_7 NS_222 0 2.6389919285437939e-06
GC_7_223 b_7 NI_7 NS_223 0 1.0043142474308335e-05
GC_7_224 b_7 NI_7 NS_224 0 9.8196625003422260e-06
GC_7_225 b_7 NI_7 NS_225 0 6.5297140272336520e-05
GC_7_226 b_7 NI_7 NS_226 0 -4.0288196248727031e-05
GC_7_227 b_7 NI_7 NS_227 0 -9.9263422815182915e-06
GC_7_228 b_7 NI_7 NS_228 0 4.7257362947114134e-05
GC_7_229 b_7 NI_7 NS_229 0 8.8864262917655562e-02
GC_7_230 b_7 NI_7 NS_230 0 -1.7530432331854396e-03
GC_7_231 b_7 NI_7 NS_231 0 3.1152633229823892e-02
GC_7_232 b_7 NI_7 NS_232 0 -6.5484423834928918e-02
GC_7_233 b_7 NI_7 NS_233 0 -2.0158652669699417e-03
GC_7_234 b_7 NI_7 NS_234 0 -9.2769904698071525e-04
GC_7_235 b_7 NI_7 NS_235 0 -1.2361255740749808e-04
GC_7_236 b_7 NI_7 NS_236 0 -1.4261529413341033e-04
GC_7_237 b_7 NI_7 NS_237 0 -1.8366655226886502e-02
GC_7_238 b_7 NI_7 NS_238 0 -2.5716199671641329e-03
GC_7_239 b_7 NI_7 NS_239 0 -8.8955126443926941e-06
GC_7_240 b_7 NI_7 NS_240 0 4.2895321213183871e-06
GC_7_241 b_7 NI_7 NS_241 0 -4.6306452437342854e-02
GC_7_242 b_7 NI_7 NS_242 0 1.5118897994905806e-02
GC_7_243 b_7 NI_7 NS_243 0 -1.2750072033946203e-05
GC_7_244 b_7 NI_7 NS_244 0 -2.7099678049894707e-05
GC_7_245 b_7 NI_7 NS_245 0 -2.7183611477657222e-05
GC_7_246 b_7 NI_7 NS_246 0 -7.2516720931285981e-06
GC_7_247 b_7 NI_7 NS_247 0 7.1951319209412021e-08
GC_7_248 b_7 NI_7 NS_248 0 -3.7091730096453347e-05
GC_7_249 b_7 NI_7 NS_249 0 6.0051425000614293e-06
GC_7_250 b_7 NI_7 NS_250 0 -4.4763100492533469e-06
GC_7_251 b_7 NI_7 NS_251 0 -3.8598957349035507e-03
GC_7_252 b_7 NI_7 NS_252 0 4.8042659896723183e-03
GC_7_253 b_7 NI_7 NS_253 0 -5.8487957541046110e-04
GC_7_254 b_7 NI_7 NS_254 0 -3.2873687539825111e-04
GC_7_255 b_7 NI_7 NS_255 0 6.7797201617499840e-04
GC_7_256 b_7 NI_7 NS_256 0 -2.6476651013763926e-04
GC_7_257 b_7 NI_7 NS_257 0 6.4631576203966591e-05
GC_7_258 b_7 NI_7 NS_258 0 -3.0495536721723425e-04
GC_7_259 b_7 NI_7 NS_259 0 3.3370345978627137e-05
GC_7_260 b_7 NI_7 NS_260 0 -4.2874658252011854e-05
GC_7_261 b_7 NI_7 NS_261 0 -8.1813859278192549e-06
GC_7_262 b_7 NI_7 NS_262 0 8.1207602683916737e-06
GC_7_263 b_7 NI_7 NS_263 0 8.8962016744524651e-05
GC_7_264 b_7 NI_7 NS_264 0 -1.0571154774563148e-04
GC_7_265 b_7 NI_7 NS_265 0 4.5581128198220034e-05
GC_7_266 b_7 NI_7 NS_266 0 -4.0515143953035243e-05
GC_7_267 b_7 NI_7 NS_267 0 -2.6430119578274222e-02
GC_7_268 b_7 NI_7 NS_268 0 2.4154987827270805e-03
GC_7_269 b_7 NI_7 NS_269 0 4.1150524923219516e-02
GC_7_270 b_7 NI_7 NS_270 0 -7.7543965496153213e-03
GC_7_271 b_7 NI_7 NS_271 0 1.0291563980953193e-03
GC_7_272 b_7 NI_7 NS_272 0 3.0168894227148413e-04
GC_7_273 b_7 NI_7 NS_273 0 4.5884367525802784e-05
GC_7_274 b_7 NI_7 NS_274 0 -1.3705144700619561e-05
GC_7_275 b_7 NI_7 NS_275 0 3.7196820684468238e-02
GC_7_276 b_7 NI_7 NS_276 0 2.7481997496672007e-02
GC_7_277 b_7 NI_7 NS_277 0 2.8533926488436510e-05
GC_7_278 b_7 NI_7 NS_278 0 4.6184842469034984e-06
GC_7_279 b_7 NI_7 NS_279 0 -4.3148591878010130e-02
GC_7_280 b_7 NI_7 NS_280 0 2.2190135177862190e-02
GC_7_281 b_7 NI_7 NS_281 0 -7.6624553387217560e-07
GC_7_282 b_7 NI_7 NS_282 0 7.6915193712260664e-06
GC_7_283 b_7 NI_7 NS_283 0 5.3192602542421422e-07
GC_7_284 b_7 NI_7 NS_284 0 4.0564227641654015e-05
GC_7_285 b_7 NI_7 NS_285 0 -1.0410026990439835e-06
GC_7_286 b_7 NI_7 NS_286 0 -3.8972574626282825e-07
GC_7_287 b_7 NI_7 NS_287 0 1.1729931944756063e-07
GC_7_288 b_7 NI_7 NS_288 0 2.9844960375661491e-06
GC_7_289 b_7 NI_7 NS_289 0 -2.2472423045811129e-03
GC_7_290 b_7 NI_7 NS_290 0 3.3713556451761997e-03
GC_7_291 b_7 NI_7 NS_291 0 -4.2146298376553518e-04
GC_7_292 b_7 NI_7 NS_292 0 -1.8690559108323535e-04
GC_7_293 b_7 NI_7 NS_293 0 5.2627333709595885e-04
GC_7_294 b_7 NI_7 NS_294 0 4.2976169505283090e-05
GC_7_295 b_7 NI_7 NS_295 0 1.7611771453992397e-04
GC_7_296 b_7 NI_7 NS_296 0 -1.8447987448907036e-04
GC_7_297 b_7 NI_7 NS_297 0 7.5066435463922194e-05
GC_7_298 b_7 NI_7 NS_298 0 4.3977239132004162e-07
GC_7_299 b_7 NI_7 NS_299 0 -1.9816480754228630e-05
GC_7_300 b_7 NI_7 NS_300 0 2.8226058644121006e-05
GC_7_301 b_7 NI_7 NS_301 0 1.1324750055692437e-04
GC_7_302 b_7 NI_7 NS_302 0 -1.7512319675041322e-05
GC_7_303 b_7 NI_7 NS_303 0 6.3627870804952688e-05
GC_7_304 b_7 NI_7 NS_304 0 6.4845977258961063e-07
GC_7_305 b_7 NI_7 NS_305 0 -3.5973135004546707e-03
GC_7_306 b_7 NI_7 NS_306 0 -1.5461170934167041e-03
GC_7_307 b_7 NI_7 NS_307 0 -4.0555754377170873e-04
GC_7_308 b_7 NI_7 NS_308 0 5.9781059927271115e-03
GC_7_309 b_7 NI_7 NS_309 0 -1.4785748110485201e-03
GC_7_310 b_7 NI_7 NS_310 0 6.6776307075113925e-04
GC_7_311 b_7 NI_7 NS_311 0 -1.2692302933926683e-04
GC_7_312 b_7 NI_7 NS_312 0 2.9240992121099045e-05
GC_7_313 b_7 NI_7 NS_313 0 5.8380001641576470e-03
GC_7_314 b_7 NI_7 NS_314 0 1.1797739180318966e-02
GC_7_315 b_7 NI_7 NS_315 0 -2.2053616890083741e-05
GC_7_316 b_7 NI_7 NS_316 0 -7.1737839726005046e-06
GC_7_317 b_7 NI_7 NS_317 0 7.2099260200182416e-03
GC_7_318 b_7 NI_7 NS_318 0 -4.8472698763394320e-03
GC_7_319 b_7 NI_7 NS_319 0 -4.4848069223519898e-06
GC_7_320 b_7 NI_7 NS_320 0 -1.8274552566518402e-05
GC_7_321 b_7 NI_7 NS_321 0 -3.0872363932118875e-05
GC_7_322 b_7 NI_7 NS_322 0 4.7704070318466628e-05
GC_7_323 b_7 NI_7 NS_323 0 -3.3950246621169286e-05
GC_7_324 b_7 NI_7 NS_324 0 -5.2531708927601013e-05
GC_7_325 b_7 NI_7 NS_325 0 5.8095559559312941e-07
GC_7_326 b_7 NI_7 NS_326 0 -8.6792155007734145e-06
GC_7_327 b_7 NI_7 NS_327 0 -6.2436608171816416e-03
GC_7_328 b_7 NI_7 NS_328 0 1.2505413559934227e-03
GC_7_329 b_7 NI_7 NS_329 0 -2.9965405941675494e-04
GC_7_330 b_7 NI_7 NS_330 0 -3.8477792089532646e-04
GC_7_331 b_7 NI_7 NS_331 0 7.3897865234763636e-04
GC_7_332 b_7 NI_7 NS_332 0 2.7342933888444753e-05
GC_7_333 b_7 NI_7 NS_333 0 1.0899059650745573e-04
GC_7_334 b_7 NI_7 NS_334 0 -2.0159197696929449e-04
GC_7_335 b_7 NI_7 NS_335 0 6.5132763698716004e-06
GC_7_336 b_7 NI_7 NS_336 0 1.3315921514798726e-05
GC_7_337 b_7 NI_7 NS_337 0 -7.3989115692679347e-06
GC_7_338 b_7 NI_7 NS_338 0 2.3588150579731818e-05
GC_7_339 b_7 NI_7 NS_339 0 4.2783588773214238e-05
GC_7_340 b_7 NI_7 NS_340 0 3.3554394174611093e-06
GC_7_341 b_7 NI_7 NS_341 0 1.3081324307719082e-06
GC_7_342 b_7 NI_7 NS_342 0 9.6873980238220759e-06
GC_7_343 b_7 NI_7 NS_343 0 -2.4113817247040772e-02
GC_7_344 b_7 NI_7 NS_344 0 1.4730211553154917e-03
GC_7_345 b_7 NI_7 NS_345 0 1.4876817916475927e-02
GC_7_346 b_7 NI_7 NS_346 0 -2.3952720409711843e-03
GC_7_347 b_7 NI_7 NS_347 0 2.1084974370652362e-04
GC_7_348 b_7 NI_7 NS_348 0 2.1039126610700778e-05
GC_7_349 b_7 NI_7 NS_349 0 -2.3638661479953965e-05
GC_7_350 b_7 NI_7 NS_350 0 -5.1599070517634763e-06
GC_7_351 b_7 NI_7 NS_351 0 -8.0049530024044226e-03
GC_7_352 b_7 NI_7 NS_352 0 -1.2244925263476231e-02
GC_7_353 b_7 NI_7 NS_353 0 2.1888237836829523e-05
GC_7_354 b_7 NI_7 NS_354 0 6.3136533822527791e-06
GC_7_355 b_7 NI_7 NS_355 0 6.1156492879061121e-03
GC_7_356 b_7 NI_7 NS_356 0 -1.0678155870730099e-02
GC_7_357 b_7 NI_7 NS_357 0 -1.7101529303466072e-05
GC_7_358 b_7 NI_7 NS_358 0 -1.4847967548003028e-05
GC_7_359 b_7 NI_7 NS_359 0 -1.1403050423411634e-05
GC_7_360 b_7 NI_7 NS_360 0 4.8083309300717525e-05
GC_7_361 b_7 NI_7 NS_361 0 -1.8697623490148234e-05
GC_7_362 b_7 NI_7 NS_362 0 -2.1123706015564250e-05
GC_7_363 b_7 NI_7 NS_363 0 -6.0549883035682931e-07
GC_7_364 b_7 NI_7 NS_364 0 -6.8985296096225186e-06
GC_7_365 b_7 NI_7 NS_365 0 -4.2965371767886024e-03
GC_7_366 b_7 NI_7 NS_366 0 2.0134995314502802e-04
GC_7_367 b_7 NI_7 NS_367 0 -1.1511792763744222e-04
GC_7_368 b_7 NI_7 NS_368 0 -3.8955377435816667e-04
GC_7_369 b_7 NI_7 NS_369 0 4.4755695699804098e-04
GC_7_370 b_7 NI_7 NS_370 0 1.3354620333600465e-04
GC_7_371 b_7 NI_7 NS_371 0 1.7123512341871594e-04
GC_7_372 b_7 NI_7 NS_372 0 -1.2651890647244159e-04
GC_7_373 b_7 NI_7 NS_373 0 -1.6677576387093165e-05
GC_7_374 b_7 NI_7 NS_374 0 -8.2956715193798373e-06
GC_7_375 b_7 NI_7 NS_375 0 1.1422010803998404e-06
GC_7_376 b_7 NI_7 NS_376 0 6.7673954026321532e-06
GC_7_377 b_7 NI_7 NS_377 0 -1.1927060004964602e-06
GC_7_378 b_7 NI_7 NS_378 0 1.3996909095899032e-05
GC_7_379 b_7 NI_7 NS_379 0 3.0390360728356069e-05
GC_7_380 b_7 NI_7 NS_380 0 2.0363703722965163e-05
GC_7_381 b_7 NI_7 NS_381 0 -2.2063659944416017e-02
GC_7_382 b_7 NI_7 NS_382 0 -1.2404848703736428e-03
GC_7_383 b_7 NI_7 NS_383 0 9.0931973609006105e-03
GC_7_384 b_7 NI_7 NS_384 0 1.2497506561516710e-02
GC_7_385 b_7 NI_7 NS_385 0 6.5547088058883624e-04
GC_7_386 b_7 NI_7 NS_386 0 3.4687437035050406e-04
GC_7_387 b_7 NI_7 NS_387 0 -2.9912577744171773e-05
GC_7_388 b_7 NI_7 NS_388 0 3.8600164073962338e-06
GC_7_389 b_7 NI_7 NS_389 0 7.9879132492787931e-03
GC_7_390 b_7 NI_7 NS_390 0 6.9055013271336931e-03
GC_7_391 b_7 NI_7 NS_391 0 -2.2590324570722992e-05
GC_7_392 b_7 NI_7 NS_392 0 -5.6416831868798651e-06
GC_7_393 b_7 NI_7 NS_393 0 1.1053183017919112e-02
GC_7_394 b_7 NI_7 NS_394 0 -8.4975036314022690e-03
GC_7_395 b_7 NI_7 NS_395 0 2.0541792535917077e-05
GC_7_396 b_7 NI_7 NS_396 0 -4.9643565216708112e-05
GC_7_397 b_7 NI_7 NS_397 0 1.4412621487735023e-05
GC_7_398 b_7 NI_7 NS_398 0 4.8043992079186082e-05
GC_7_399 b_7 NI_7 NS_399 0 -4.6872944550867745e-05
GC_7_400 b_7 NI_7 NS_400 0 -3.9804246599222589e-05
GC_7_401 b_7 NI_7 NS_401 0 -3.0368104409710014e-06
GC_7_402 b_7 NI_7 NS_402 0 -5.5034364662922954e-06
GC_7_403 b_7 NI_7 NS_403 0 -3.5805352107349982e-03
GC_7_404 b_7 NI_7 NS_404 0 1.8314261858467526e-03
GC_7_405 b_7 NI_7 NS_405 0 -3.7094745397184232e-04
GC_7_406 b_7 NI_7 NS_406 0 -3.7654846238487801e-05
GC_7_407 b_7 NI_7 NS_407 0 8.8293593077682264e-04
GC_7_408 b_7 NI_7 NS_408 0 1.4453612870839733e-04
GC_7_409 b_7 NI_7 NS_409 0 1.0048099936950826e-04
GC_7_410 b_7 NI_7 NS_410 0 -4.0978111609649473e-04
GC_7_411 b_7 NI_7 NS_411 0 -5.3902229136908476e-05
GC_7_412 b_7 NI_7 NS_412 0 5.7204949883061926e-05
GC_7_413 b_7 NI_7 NS_413 0 -2.0528972068436257e-05
GC_7_414 b_7 NI_7 NS_414 0 1.2983139143910704e-05
GC_7_415 b_7 NI_7 NS_415 0 -4.3693801778395904e-05
GC_7_416 b_7 NI_7 NS_416 0 3.5040803794382619e-05
GC_7_417 b_7 NI_7 NS_417 0 -5.0896163221564445e-06
GC_7_418 b_7 NI_7 NS_418 0 1.4065395877779359e-08
GC_7_419 b_7 NI_7 NS_419 0 2.5101600701566959e-02
GC_7_420 b_7 NI_7 NS_420 0 1.2306792507807238e-03
GC_7_421 b_7 NI_7 NS_421 0 -1.5318726835486620e-02
GC_7_422 b_7 NI_7 NS_422 0 1.2333990014425946e-03
GC_7_423 b_7 NI_7 NS_423 0 4.0036534898762219e-04
GC_7_424 b_7 NI_7 NS_424 0 -2.5192064561226844e-04
GC_7_425 b_7 NI_7 NS_425 0 -1.1137216305158501e-05
GC_7_426 b_7 NI_7 NS_426 0 -1.9943676154290536e-05
GC_7_427 b_7 NI_7 NS_427 0 -8.2920104843385110e-03
GC_7_428 b_7 NI_7 NS_428 0 -7.8176457287028461e-03
GC_7_429 b_7 NI_7 NS_429 0 2.0757398919958137e-05
GC_7_430 b_7 NI_7 NS_430 0 6.5884437285511361e-06
GC_7_431 b_7 NI_7 NS_431 0 9.6915207014852730e-03
GC_7_432 b_7 NI_7 NS_432 0 1.5047245657696933e-03
GC_7_433 b_7 NI_7 NS_433 0 -3.6979050380963488e-06
GC_7_434 b_7 NI_7 NS_434 0 -4.2165211781882023e-05
GC_7_435 b_7 NI_7 NS_435 0 9.1468708630295745e-06
GC_7_436 b_7 NI_7 NS_436 0 5.0465035246189457e-05
GC_7_437 b_7 NI_7 NS_437 0 -2.3246744563939462e-05
GC_7_438 b_7 NI_7 NS_438 0 -2.5611693693045768e-05
GC_7_439 b_7 NI_7 NS_439 0 -1.4746513884070386e-06
GC_7_440 b_7 NI_7 NS_440 0 -4.7835129953357569e-06
GC_7_441 b_7 NI_7 NS_441 0 -4.4927216494639894e-03
GC_7_442 b_7 NI_7 NS_442 0 5.5513105877920605e-04
GC_7_443 b_7 NI_7 NS_443 0 -1.2390154984313494e-04
GC_7_444 b_7 NI_7 NS_444 0 -2.8585112831755829e-04
GC_7_445 b_7 NI_7 NS_445 0 7.4983181754985969e-04
GC_7_446 b_7 NI_7 NS_446 0 3.7004261922730962e-04
GC_7_447 b_7 NI_7 NS_447 0 2.6737625307316870e-04
GC_7_448 b_7 NI_7 NS_448 0 -3.1089052016405286e-04
GC_7_449 b_7 NI_7 NS_449 0 -7.3772211173709485e-05
GC_7_450 b_7 NI_7 NS_450 0 9.0525509306995044e-06
GC_7_451 b_7 NI_7 NS_451 0 -1.6263136282165976e-05
GC_7_452 b_7 NI_7 NS_452 0 1.7046765708274505e-06
GC_7_453 b_7 NI_7 NS_453 0 -6.9786045833731584e-05
GC_7_454 b_7 NI_7 NS_454 0 1.7597504523417348e-05
GC_7_455 b_7 NI_7 NS_455 0 -4.2029240995787246e-06
GC_7_456 b_7 NI_7 NS_456 0 3.9083091467222365e-06
GD_7_1 b_7 NI_7 NA_1 0 -2.5259757570995456e-03
GD_7_2 b_7 NI_7 NA_2 0 -6.3704701671097709e-03
GD_7_3 b_7 NI_7 NA_3 0 -9.2750432992688807e-03
GD_7_4 b_7 NI_7 NA_4 0 -8.9592395435854084e-03
GD_7_5 b_7 NI_7 NA_5 0 -3.4465806932342760e-02
GD_7_6 b_7 NI_7 NA_6 0 2.0712576101638753e-02
GD_7_7 b_7 NI_7 NA_7 0 -8.0922755250270817e-02
GD_7_8 b_7 NI_7 NA_8 0 -2.1049626403373187e-02
GD_7_9 b_7 NI_7 NA_9 0 7.1528125093672521e-03
GD_7_10 b_7 NI_7 NA_10 0 1.1951586823095705e-02
GD_7_11 b_7 NI_7 NA_11 0 -6.5418334461556068e-03
GD_7_12 b_7 NI_7 NA_12 0 -7.8439671122404412e-03
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 7.8588000288786937e-03
GC_8_2 b_8 NI_8 NS_2 0 1.1231922144294840e-03
GC_8_3 b_8 NI_8 NS_3 0 -8.2820768904528740e-03
GC_8_4 b_8 NI_8 NS_4 0 7.9316652815912530e-03
GC_8_5 b_8 NI_8 NS_5 0 -3.4436464601069504e-05
GC_8_6 b_8 NI_8 NS_6 0 -2.6131778744015877e-04
GC_8_7 b_8 NI_8 NS_7 0 3.8415778429252966e-05
GC_8_8 b_8 NI_8 NS_8 0 -1.9608479105329055e-05
GC_8_9 b_8 NI_8 NS_9 0 -1.1514677090752267e-03
GC_8_10 b_8 NI_8 NS_10 0 6.1453857588627467e-03
GC_8_11 b_8 NI_8 NS_11 0 2.7449146874490862e-05
GC_8_12 b_8 NI_8 NS_12 0 -1.0349987711489159e-06
GC_8_13 b_8 NI_8 NS_13 0 7.4352770063286786e-03
GC_8_14 b_8 NI_8 NS_14 0 -2.8375799472765998e-03
GC_8_15 b_8 NI_8 NS_15 0 7.3955670456024892e-07
GC_8_16 b_8 NI_8 NS_16 0 -7.0808109089295189e-06
GC_8_17 b_8 NI_8 NS_17 0 -1.1393056333389523e-05
GC_8_18 b_8 NI_8 NS_18 0 1.0295582253533218e-05
GC_8_19 b_8 NI_8 NS_19 0 2.1144149664126777e-05
GC_8_20 b_8 NI_8 NS_20 0 6.8775960121361872e-06
GC_8_21 b_8 NI_8 NS_21 0 -1.7141208164293109e-05
GC_8_22 b_8 NI_8 NS_22 0 9.5060663785102206e-06
GC_8_23 b_8 NI_8 NS_23 0 -5.1229178302076195e-04
GC_8_24 b_8 NI_8 NS_24 0 2.3450323446358320e-03
GC_8_25 b_8 NI_8 NS_25 0 -2.2840220833152296e-04
GC_8_26 b_8 NI_8 NS_26 0 -4.3184760874949549e-04
GC_8_27 b_8 NI_8 NS_27 0 -4.1612137967063501e-05
GC_8_28 b_8 NI_8 NS_28 0 -3.8982279836094664e-04
GC_8_29 b_8 NI_8 NS_29 0 -1.7938570056191390e-04
GC_8_30 b_8 NI_8 NS_30 0 2.4931402442780515e-04
GC_8_31 b_8 NI_8 NS_31 0 -6.5061200442651456e-05
GC_8_32 b_8 NI_8 NS_32 0 -1.7574791957100171e-05
GC_8_33 b_8 NI_8 NS_33 0 1.4895950101112089e-05
GC_8_34 b_8 NI_8 NS_34 0 1.0951563586983982e-05
GC_8_35 b_8 NI_8 NS_35 0 -3.9192373033960824e-05
GC_8_36 b_8 NI_8 NS_36 0 6.8776219945739946e-05
GC_8_37 b_8 NI_8 NS_37 0 1.3677043023185759e-05
GC_8_38 b_8 NI_8 NS_38 0 -1.2745177252819924e-05
GC_8_39 b_8 NI_8 NS_39 0 -1.9134362644894865e-02
GC_8_40 b_8 NI_8 NS_40 0 -1.0287209278749961e-03
GC_8_41 b_8 NI_8 NS_41 0 3.5560044033521271e-03
GC_8_42 b_8 NI_8 NS_42 0 8.3936622486899398e-03
GC_8_43 b_8 NI_8 NS_43 0 2.4696250363082820e-05
GC_8_44 b_8 NI_8 NS_44 0 -9.1459538476170520e-05
GC_8_45 b_8 NI_8 NS_45 0 -4.5822750417312331e-05
GC_8_46 b_8 NI_8 NS_46 0 1.8035158084167162e-05
GC_8_47 b_8 NI_8 NS_47 0 4.9834073875528817e-03
GC_8_48 b_8 NI_8 NS_48 0 -1.0725628902769685e-03
GC_8_49 b_8 NI_8 NS_49 0 -2.0578175068814621e-05
GC_8_50 b_8 NI_8 NS_50 0 2.5749348500155169e-06
GC_8_51 b_8 NI_8 NS_51 0 9.3384410248491794e-03
GC_8_52 b_8 NI_8 NS_52 0 -7.4118648758797505e-03
GC_8_53 b_8 NI_8 NS_53 0 9.0332022518739258e-07
GC_8_54 b_8 NI_8 NS_54 0 2.6095644444398158e-05
GC_8_55 b_8 NI_8 NS_55 0 -1.5577253491193212e-05
GC_8_56 b_8 NI_8 NS_56 0 2.6682652818221125e-05
GC_8_57 b_8 NI_8 NS_57 0 4.6316653135743823e-06
GC_8_58 b_8 NI_8 NS_58 0 1.1817104459644428e-07
GC_8_59 b_8 NI_8 NS_59 0 -2.7670382488710180e-05
GC_8_60 b_8 NI_8 NS_60 0 1.5730610033737863e-05
GC_8_61 b_8 NI_8 NS_61 0 -1.7663299645196370e-03
GC_8_62 b_8 NI_8 NS_62 0 3.2729635629340859e-03
GC_8_63 b_8 NI_8 NS_63 0 -1.9692330688164281e-05
GC_8_64 b_8 NI_8 NS_64 0 -5.6525883000338017e-04
GC_8_65 b_8 NI_8 NS_65 0 1.3175728919236451e-04
GC_8_66 b_8 NI_8 NS_66 0 -4.6464254822218870e-04
GC_8_67 b_8 NI_8 NS_67 0 -1.6935430692580859e-04
GC_8_68 b_8 NI_8 NS_68 0 1.6192602519558548e-04
GC_8_69 b_8 NI_8 NS_69 0 -3.0382759317478527e-05
GC_8_70 b_8 NI_8 NS_70 0 -5.4079139476874523e-05
GC_8_71 b_8 NI_8 NS_71 0 7.2710182407532685e-06
GC_8_72 b_8 NI_8 NS_72 0 4.8473519793037493e-06
GC_8_73 b_8 NI_8 NS_73 0 -9.8035972644828044e-06
GC_8_74 b_8 NI_8 NS_74 0 5.4741363155495601e-05
GC_8_75 b_8 NI_8 NS_75 0 -1.3758539791658053e-06
GC_8_76 b_8 NI_8 NS_76 0 -2.8254307464332939e-05
GC_8_77 b_8 NI_8 NS_77 0 7.3101835112056529e-03
GC_8_78 b_8 NI_8 NS_78 0 1.3556891546286712e-03
GC_8_79 b_8 NI_8 NS_79 0 -6.4264511280333206e-03
GC_8_80 b_8 NI_8 NS_80 0 2.9716196593923896e-03
GC_8_81 b_8 NI_8 NS_81 0 1.1174861511909687e-04
GC_8_82 b_8 NI_8 NS_82 0 5.3071251233338421e-05
GC_8_83 b_8 NI_8 NS_83 0 4.3955713662675676e-05
GC_8_84 b_8 NI_8 NS_84 0 1.5663266758180485e-05
GC_8_85 b_8 NI_8 NS_85 0 -5.9821136283822610e-03
GC_8_86 b_8 NI_8 NS_86 0 -3.4130180138898817e-03
GC_8_87 b_8 NI_8 NS_87 0 2.3284955101653639e-05
GC_8_88 b_8 NI_8 NS_88 0 -2.9307736660153736e-06
GC_8_89 b_8 NI_8 NS_89 0 9.0967655268249861e-03
GC_8_90 b_8 NI_8 NS_90 0 -4.9040823807714792e-03
GC_8_91 b_8 NI_8 NS_91 0 -4.2593950068529259e-06
GC_8_92 b_8 NI_8 NS_92 0 -6.9905538011086718e-06
GC_8_93 b_8 NI_8 NS_93 0 -1.2409624478089027e-05
GC_8_94 b_8 NI_8 NS_94 0 2.4964429735507514e-05
GC_8_95 b_8 NI_8 NS_95 0 1.6655919325570886e-05
GC_8_96 b_8 NI_8 NS_96 0 1.0331494841896193e-05
GC_8_97 b_8 NI_8 NS_97 0 -1.4970434225169068e-05
GC_8_98 b_8 NI_8 NS_98 0 8.5887983976173513e-06
GC_8_99 b_8 NI_8 NS_99 0 -2.9815286025429437e-03
GC_8_100 b_8 NI_8 NS_100 0 2.3381584965287546e-03
GC_8_101 b_8 NI_8 NS_101 0 -2.4070282055448948e-04
GC_8_102 b_8 NI_8 NS_102 0 -4.0204341911355483e-04
GC_8_103 b_8 NI_8 NS_103 0 2.3789438915000106e-04
GC_8_104 b_8 NI_8 NS_104 0 -8.6089137382537985e-05
GC_8_105 b_8 NI_8 NS_105 0 8.8884754347398292e-06
GC_8_106 b_8 NI_8 NS_106 0 5.1377114100196989e-05
GC_8_107 b_8 NI_8 NS_107 0 -6.7248433831970596e-06
GC_8_108 b_8 NI_8 NS_108 0 6.5462505152147674e-06
GC_8_109 b_8 NI_8 NS_109 0 2.0543238312191801e-06
GC_8_110 b_8 NI_8 NS_110 0 1.1084961639383054e-05
GC_8_111 b_8 NI_8 NS_111 0 4.1186746661218593e-05
GC_8_112 b_8 NI_8 NS_112 0 4.8813998553325050e-05
GC_8_113 b_8 NI_8 NS_113 0 2.7087346652772202e-06
GC_8_114 b_8 NI_8 NS_114 0 8.0925177797437968e-06
GC_8_115 b_8 NI_8 NS_115 0 -5.0893612613850967e-04
GC_8_116 b_8 NI_8 NS_116 0 -1.3150662623033717e-03
GC_8_117 b_8 NI_8 NS_117 0 -7.4776836713396190e-03
GC_8_118 b_8 NI_8 NS_118 0 8.3598885178417237e-03
GC_8_119 b_8 NI_8 NS_119 0 -3.8133435673700691e-05
GC_8_120 b_8 NI_8 NS_120 0 -1.0974056418991172e-04
GC_8_121 b_8 NI_8 NS_121 0 -7.0939415659858386e-05
GC_8_122 b_8 NI_8 NS_122 0 2.3385597289418907e-05
GC_8_123 b_8 NI_8 NS_123 0 5.1211511531292532e-03
GC_8_124 b_8 NI_8 NS_124 0 2.8105855286699815e-03
GC_8_125 b_8 NI_8 NS_125 0 -2.0552488980242408e-05
GC_8_126 b_8 NI_8 NS_126 0 3.4759209509511308e-06
GC_8_127 b_8 NI_8 NS_127 0 1.3221075214391996e-02
GC_8_128 b_8 NI_8 NS_128 0 -1.5087094666463717e-03
GC_8_129 b_8 NI_8 NS_129 0 7.1089052131673034e-06
GC_8_130 b_8 NI_8 NS_130 0 2.1873766811152582e-05
GC_8_131 b_8 NI_8 NS_131 0 -1.8966019485989927e-05
GC_8_132 b_8 NI_8 NS_132 0 2.6956899612527810e-05
GC_8_133 b_8 NI_8 NS_133 0 7.8610290273619060e-06
GC_8_134 b_8 NI_8 NS_134 0 6.4805483493355233e-06
GC_8_135 b_8 NI_8 NS_135 0 -2.6456425778527157e-05
GC_8_136 b_8 NI_8 NS_136 0 1.7036490860116436e-05
GC_8_137 b_8 NI_8 NS_137 0 -4.3093171803429472e-03
GC_8_138 b_8 NI_8 NS_138 0 1.8529421028523978e-03
GC_8_139 b_8 NI_8 NS_139 0 5.7634782086147171e-05
GC_8_140 b_8 NI_8 NS_140 0 -5.4673613287662673e-04
GC_8_141 b_8 NI_8 NS_141 0 4.2509239786602009e-04
GC_8_142 b_8 NI_8 NS_142 0 -1.1110466476065567e-04
GC_8_143 b_8 NI_8 NS_143 0 -2.5198730024227441e-05
GC_8_144 b_8 NI_8 NS_144 0 1.6541176019398553e-05
GC_8_145 b_8 NI_8 NS_145 0 -2.0511442418888074e-06
GC_8_146 b_8 NI_8 NS_146 0 3.3909093262095477e-06
GC_8_147 b_8 NI_8 NS_147 0 -5.3559873280116897e-06
GC_8_148 b_8 NI_8 NS_148 0 3.9828627185612331e-06
GC_8_149 b_8 NI_8 NS_149 0 4.4739474978270880e-05
GC_8_150 b_8 NI_8 NS_150 0 4.1455044588949126e-05
GC_8_151 b_8 NI_8 NS_151 0 1.4547153849628127e-05
GC_8_152 b_8 NI_8 NS_152 0 3.0054691807065033e-06
GC_8_153 b_8 NI_8 NS_153 0 -2.4968812220719492e-03
GC_8_154 b_8 NI_8 NS_154 0 1.1659568370898223e-03
GC_8_155 b_8 NI_8 NS_155 0 1.4957083777879163e-03
GC_8_156 b_8 NI_8 NS_156 0 -6.3561230572526601e-03
GC_8_157 b_8 NI_8 NS_157 0 -5.5637035661352143e-05
GC_8_158 b_8 NI_8 NS_158 0 7.7035146985619124e-04
GC_8_159 b_8 NI_8 NS_159 0 3.6593702921272038e-05
GC_8_160 b_8 NI_8 NS_160 0 9.7289965761496270e-05
GC_8_161 b_8 NI_8 NS_161 0 -1.2769254916876522e-02
GC_8_162 b_8 NI_8 NS_162 0 -1.9886414107110912e-02
GC_8_163 b_8 NI_8 NS_163 0 -7.7314411583063185e-07
GC_8_164 b_8 NI_8 NS_164 0 -4.9343868086894477e-06
GC_8_165 b_8 NI_8 NS_165 0 7.6753409303586236e-03
GC_8_166 b_8 NI_8 NS_166 0 -1.7877285429264814e-02
GC_8_167 b_8 NI_8 NS_167 0 -1.7263036440540588e-05
GC_8_168 b_8 NI_8 NS_168 0 8.4619820579784366e-06
GC_8_169 b_8 NI_8 NS_169 0 -2.0330060093519994e-05
GC_8_170 b_8 NI_8 NS_170 0 4.7619491856742888e-05
GC_8_171 b_8 NI_8 NS_171 0 -6.0874961126016848e-06
GC_8_172 b_8 NI_8 NS_172 0 -3.4049012524784488e-06
GC_8_173 b_8 NI_8 NS_173 0 3.9523565425445907e-07
GC_8_174 b_8 NI_8 NS_174 0 -5.6836590220427050e-06
GC_8_175 b_8 NI_8 NS_175 0 -3.8285971216547444e-03
GC_8_176 b_8 NI_8 NS_176 0 8.7866558284996395e-03
GC_8_177 b_8 NI_8 NS_177 0 -5.2098441261411643e-04
GC_8_178 b_8 NI_8 NS_178 0 -5.8846879211546640e-04
GC_8_179 b_8 NI_8 NS_179 0 3.7056573192875502e-04
GC_8_180 b_8 NI_8 NS_180 0 -5.3886326461690998e-04
GC_8_181 b_8 NI_8 NS_181 0 -7.1652826442721737e-05
GC_8_182 b_8 NI_8 NS_182 0 -1.4464696549362869e-05
GC_8_183 b_8 NI_8 NS_183 0 6.0196205312946926e-05
GC_8_184 b_8 NI_8 NS_184 0 -2.0499744792191697e-05
GC_8_185 b_8 NI_8 NS_185 0 1.4083566917590647e-05
GC_8_186 b_8 NI_8 NS_186 0 2.2907078739473003e-05
GC_8_187 b_8 NI_8 NS_187 0 5.9660611732491392e-05
GC_8_188 b_8 NI_8 NS_188 0 -2.4588717818683568e-05
GC_8_189 b_8 NI_8 NS_189 0 -1.2183550304362696e-06
GC_8_190 b_8 NI_8 NS_190 0 4.4775909793180460e-05
GC_8_191 b_8 NI_8 NS_191 0 2.9573452492089401e-02
GC_8_192 b_8 NI_8 NS_192 0 -1.4830417326759586e-03
GC_8_193 b_8 NI_8 NS_193 0 -1.2646361476794496e-02
GC_8_194 b_8 NI_8 NS_194 0 -6.0727707501738917e-03
GC_8_195 b_8 NI_8 NS_195 0 -3.1105797549848654e-05
GC_8_196 b_8 NI_8 NS_196 0 8.2220534885231629e-05
GC_8_197 b_8 NI_8 NS_197 0 -2.7395587181923589e-05
GC_8_198 b_8 NI_8 NS_198 0 3.6323587237261178e-06
GC_8_199 b_8 NI_8 NS_199 0 -4.4100564696039774e-05
GC_8_200 b_8 NI_8 NS_200 0 6.8137491509456241e-03
GC_8_201 b_8 NI_8 NS_201 0 -1.0403993557755315e-05
GC_8_202 b_8 NI_8 NS_202 0 3.1435212014762258e-06
GC_8_203 b_8 NI_8 NS_203 0 2.6204689550149147e-04
GC_8_204 b_8 NI_8 NS_204 0 -2.0575200576341160e-03
GC_8_205 b_8 NI_8 NS_205 0 -2.6266620744576270e-06
GC_8_206 b_8 NI_8 NS_206 0 9.4009480776909814e-06
GC_8_207 b_8 NI_8 NS_207 0 -1.4027249819578200e-05
GC_8_208 b_8 NI_8 NS_208 0 2.1783472189045532e-05
GC_8_209 b_8 NI_8 NS_209 0 -6.7499816981529471e-06
GC_8_210 b_8 NI_8 NS_210 0 -3.2850486753576677e-06
GC_8_211 b_8 NI_8 NS_211 0 -1.9503719021686099e-06
GC_8_212 b_8 NI_8 NS_212 0 1.5638797245032633e-06
GC_8_213 b_8 NI_8 NS_213 0 -2.8256319588491350e-03
GC_8_214 b_8 NI_8 NS_214 0 6.3954058637100660e-03
GC_8_215 b_8 NI_8 NS_215 0 -3.3373888449924466e-04
GC_8_216 b_8 NI_8 NS_216 0 -4.0864123423146978e-04
GC_8_217 b_8 NI_8 NS_217 0 2.9717446074543582e-04
GC_8_218 b_8 NI_8 NS_218 0 -3.2384175975272233e-04
GC_8_219 b_8 NI_8 NS_219 0 8.1259255737615088e-07
GC_8_220 b_8 NI_8 NS_220 0 2.5925674912882502e-05
GC_8_221 b_8 NI_8 NS_221 0 2.8552417556957551e-05
GC_8_222 b_8 NI_8 NS_222 0 5.5689733412113933e-05
GC_8_223 b_8 NI_8 NS_223 0 -7.3161193262340345e-06
GC_8_224 b_8 NI_8 NS_224 0 2.6860984851663201e-05
GC_8_225 b_8 NI_8 NS_225 0 6.4896685221899861e-05
GC_8_226 b_8 NI_8 NS_226 0 1.9837000436813265e-05
GC_8_227 b_8 NI_8 NS_227 0 -2.5470736448887223e-05
GC_8_228 b_8 NI_8 NS_228 0 3.6590995087997876e-05
GC_8_229 b_8 NI_8 NS_229 0 -2.6430329890764610e-02
GC_8_230 b_8 NI_8 NS_230 0 2.4155009219326844e-03
GC_8_231 b_8 NI_8 NS_231 0 4.1150593760105277e-02
GC_8_232 b_8 NI_8 NS_232 0 -7.7543366216423909e-03
GC_8_233 b_8 NI_8 NS_233 0 1.0291547649831196e-03
GC_8_234 b_8 NI_8 NS_234 0 3.0168849805186282e-04
GC_8_235 b_8 NI_8 NS_235 0 4.5884142861453736e-05
GC_8_236 b_8 NI_8 NS_236 0 -1.3704892734004157e-05
GC_8_237 b_8 NI_8 NS_237 0 3.7196858398950906e-02
GC_8_238 b_8 NI_8 NS_238 0 2.7482066029435159e-02
GC_8_239 b_8 NI_8 NS_239 0 2.8533979851086780e-05
GC_8_240 b_8 NI_8 NS_240 0 4.6185702174119663e-06
GC_8_241 b_8 NI_8 NS_241 0 -4.3148541346375240e-02
GC_8_242 b_8 NI_8 NS_242 0 2.2190063296667881e-02
GC_8_243 b_8 NI_8 NS_243 0 -7.6623487340396499e-07
GC_8_244 b_8 NI_8 NS_244 0 7.6916005080952437e-06
GC_8_245 b_8 NI_8 NS_245 0 5.3196599027701083e-07
GC_8_246 b_8 NI_8 NS_246 0 4.0564258067870750e-05
GC_8_247 b_8 NI_8 NS_247 0 -1.0409664787617497e-06
GC_8_248 b_8 NI_8 NS_248 0 -3.8970530785700447e-07
GC_8_249 b_8 NI_8 NS_249 0 1.1731080121854274e-07
GC_8_250 b_8 NI_8 NS_250 0 2.9845212521654217e-06
GC_8_251 b_8 NI_8 NS_251 0 -2.2472534250058433e-03
GC_8_252 b_8 NI_8 NS_252 0 3.3713861984286712e-03
GC_8_253 b_8 NI_8 NS_253 0 -4.2146102229600129e-04
GC_8_254 b_8 NI_8 NS_254 0 -1.8690925447174898e-04
GC_8_255 b_8 NI_8 NS_255 0 5.2627434684961714e-04
GC_8_256 b_8 NI_8 NS_256 0 4.2969898035290135e-05
GC_8_257 b_8 NI_8 NS_257 0 1.7611621216866705e-04
GC_8_258 b_8 NI_8 NS_258 0 -1.8448007587048559e-04
GC_8_259 b_8 NI_8 NS_259 0 7.5066519492227138e-05
GC_8_260 b_8 NI_8 NS_260 0 4.4000002607025435e-07
GC_8_261 b_8 NI_8 NS_261 0 -1.9816873127485929e-05
GC_8_262 b_8 NI_8 NS_262 0 2.8225889624476552e-05
GC_8_263 b_8 NI_8 NS_263 0 1.1324706029788932e-04
GC_8_264 b_8 NI_8 NS_264 0 -1.7512934643589226e-05
GC_8_265 b_8 NI_8 NS_265 0 6.3627719420243043e-05
GC_8_266 b_8 NI_8 NS_266 0 6.4869250413955847e-07
GC_8_267 b_8 NI_8 NS_267 0 1.1682166450804650e-01
GC_8_268 b_8 NI_8 NS_268 0 -1.7616266930335297e-03
GC_8_269 b_8 NI_8 NS_269 0 1.0922005887119125e-02
GC_8_270 b_8 NI_8 NS_270 0 -5.9833124517292197e-02
GC_8_271 b_8 NI_8 NS_271 0 7.4039555529890210e-05
GC_8_272 b_8 NI_8 NS_272 0 -5.9476320904995909e-04
GC_8_273 b_8 NI_8 NS_273 0 5.4986538597033358e-05
GC_8_274 b_8 NI_8 NS_274 0 -6.7845406627100465e-05
GC_8_275 b_8 NI_8 NS_275 0 -1.8452082943804883e-02
GC_8_276 b_8 NI_8 NS_276 0 -3.7316232717870415e-03
GC_8_277 b_8 NI_8 NS_277 0 -1.4376171095803010e-05
GC_8_278 b_8 NI_8 NS_278 0 3.6054998099803132e-06
GC_8_279 b_8 NI_8 NS_279 0 -3.0100417633255761e-02
GC_8_280 b_8 NI_8 NS_280 0 1.9743304603094737e-02
GC_8_281 b_8 NI_8 NS_281 0 3.3781054893545121e-05
GC_8_282 b_8 NI_8 NS_282 0 -1.0107365614994272e-05
GC_8_283 b_8 NI_8 NS_283 0 9.9305370058900829e-06
GC_8_284 b_8 NI_8 NS_284 0 4.8870763835163646e-06
GC_8_285 b_8 NI_8 NS_285 0 1.1039558460300069e-05
GC_8_286 b_8 NI_8 NS_286 0 -5.7288362746882212e-06
GC_8_287 b_8 NI_8 NS_287 0 2.2314560599368257e-07
GC_8_288 b_8 NI_8 NS_288 0 8.9200671143893780e-06
GC_8_289 b_8 NI_8 NS_289 0 -4.3612994674114324e-03
GC_8_290 b_8 NI_8 NS_290 0 3.8052976081828236e-03
GC_8_291 b_8 NI_8 NS_291 0 -1.7276762807969046e-04
GC_8_292 b_8 NI_8 NS_292 0 -2.9302330470647040e-04
GC_8_293 b_8 NI_8 NS_293 0 6.0389075466311232e-04
GC_8_294 b_8 NI_8 NS_294 0 1.7374642995075137e-04
GC_8_295 b_8 NI_8 NS_295 0 2.3379901148804552e-04
GC_8_296 b_8 NI_8 NS_296 0 -1.1472256044216965e-04
GC_8_297 b_8 NI_8 NS_297 0 3.2417886433877552e-05
GC_8_298 b_8 NI_8 NS_298 0 5.3872765219700202e-05
GC_8_299 b_8 NI_8 NS_299 0 -8.6289151015557037e-06
GC_8_300 b_8 NI_8 NS_300 0 1.0657387771644543e-05
GC_8_301 b_8 NI_8 NS_301 0 1.3305451140500202e-04
GC_8_302 b_8 NI_8 NS_302 0 6.2809568287655596e-05
GC_8_303 b_8 NI_8 NS_303 0 4.8967696114973702e-05
GC_8_304 b_8 NI_8 NS_304 0 2.2306020018149647e-05
GC_8_305 b_8 NI_8 NS_305 0 -2.5747213379074822e-02
GC_8_306 b_8 NI_8 NS_306 0 1.4965428367406074e-03
GC_8_307 b_8 NI_8 NS_307 0 1.5316510189651460e-02
GC_8_308 b_8 NI_8 NS_308 0 3.2312651584604263e-03
GC_8_309 b_8 NI_8 NS_309 0 -4.4279029139443131e-05
GC_8_310 b_8 NI_8 NS_310 0 3.5380712334446410e-05
GC_8_311 b_8 NI_8 NS_311 0 -5.4393398026999202e-06
GC_8_312 b_8 NI_8 NS_312 0 -1.3016320764415001e-05
GC_8_313 b_8 NI_8 NS_313 0 -7.0734574377485735e-03
GC_8_314 b_8 NI_8 NS_314 0 -1.0892133453368050e-02
GC_8_315 b_8 NI_8 NS_315 0 2.5449632785282621e-05
GC_8_316 b_8 NI_8 NS_316 0 1.0189853687520895e-05
GC_8_317 b_8 NI_8 NS_317 0 9.5300076516754463e-03
GC_8_318 b_8 NI_8 NS_318 0 -1.3617274588679357e-02
GC_8_319 b_8 NI_8 NS_319 0 -2.2052044427182055e-06
GC_8_320 b_8 NI_8 NS_320 0 5.8092054007672716e-06
GC_8_321 b_8 NI_8 NS_321 0 -1.1424147189214219e-05
GC_8_322 b_8 NI_8 NS_322 0 3.9426820382556401e-05
GC_8_323 b_8 NI_8 NS_323 0 -1.0480641076646154e-05
GC_8_324 b_8 NI_8 NS_324 0 -2.2687840171352904e-05
GC_8_325 b_8 NI_8 NS_325 0 1.8238871256883022e-05
GC_8_326 b_8 NI_8 NS_326 0 -2.9463978215647549e-06
GC_8_327 b_8 NI_8 NS_327 0 -5.1151007530429414e-03
GC_8_328 b_8 NI_8 NS_328 0 8.2621791085545516e-04
GC_8_329 b_8 NI_8 NS_329 0 -1.6163107454145214e-04
GC_8_330 b_8 NI_8 NS_330 0 -3.1633006893380861e-04
GC_8_331 b_8 NI_8 NS_331 0 6.0852111889602020e-04
GC_8_332 b_8 NI_8 NS_332 0 2.1537823018098653e-04
GC_8_333 b_8 NI_8 NS_333 0 1.6376614984907169e-04
GC_8_334 b_8 NI_8 NS_334 0 -1.1783953836951381e-04
GC_8_335 b_8 NI_8 NS_335 0 -1.3253833765780750e-05
GC_8_336 b_8 NI_8 NS_336 0 1.1335378105575963e-05
GC_8_337 b_8 NI_8 NS_337 0 -1.8347763510256801e-05
GC_8_338 b_8 NI_8 NS_338 0 9.8702340024981514e-06
GC_8_339 b_8 NI_8 NS_339 0 3.7851420729887182e-05
GC_8_340 b_8 NI_8 NS_340 0 3.3543610657218423e-05
GC_8_341 b_8 NI_8 NS_341 0 -3.5980668227272342e-06
GC_8_342 b_8 NI_8 NS_342 0 6.3681324060339424e-06
GC_8_343 b_8 NI_8 NS_343 0 -1.5982575393725554e-02
GC_8_344 b_8 NI_8 NS_344 0 -1.5163477925050333e-03
GC_8_345 b_8 NI_8 NS_345 0 1.0314742800452432e-02
GC_8_346 b_8 NI_8 NS_346 0 2.2248737834155173e-02
GC_8_347 b_8 NI_8 NS_347 0 -2.6378405080704502e-04
GC_8_348 b_8 NI_8 NS_348 0 4.3028376808757450e-04
GC_8_349 b_8 NI_8 NS_349 0 -1.3837731871376411e-05
GC_8_350 b_8 NI_8 NS_350 0 3.8170344073895171e-05
GC_8_351 b_8 NI_8 NS_351 0 6.8934973873173650e-03
GC_8_352 b_8 NI_8 NS_352 0 9.4223723104126574e-03
GC_8_353 b_8 NI_8 NS_353 0 -2.2150590461911566e-05
GC_8_354 b_8 NI_8 NS_354 0 -9.3857844636299131e-06
GC_8_355 b_8 NI_8 NS_355 0 1.2955492626767600e-02
GC_8_356 b_8 NI_8 NS_356 0 -1.4354712241189381e-02
GC_8_357 b_8 NI_8 NS_357 0 4.9111385388435823e-06
GC_8_358 b_8 NI_8 NS_358 0 1.2586769693765095e-05
GC_8_359 b_8 NI_8 NS_359 0 -1.7380033963321392e-05
GC_8_360 b_8 NI_8 NS_360 0 3.1536607213563099e-05
GC_8_361 b_8 NI_8 NS_361 0 -7.0170438318977441e-06
GC_8_362 b_8 NI_8 NS_362 0 -1.4031556072566027e-05
GC_8_363 b_8 NI_8 NS_363 0 1.7502692615673181e-05
GC_8_364 b_8 NI_8 NS_364 0 -3.1218177692031184e-06
GC_8_365 b_8 NI_8 NS_365 0 -4.3699029535698500e-03
GC_8_366 b_8 NI_8 NS_366 0 5.4981967886625098e-04
GC_8_367 b_8 NI_8 NS_367 0 -1.7784136674074632e-06
GC_8_368 b_8 NI_8 NS_368 0 -3.8108286816283576e-04
GC_8_369 b_8 NI_8 NS_369 0 4.0701006708126244e-04
GC_8_370 b_8 NI_8 NS_370 0 1.6191009681837054e-04
GC_8_371 b_8 NI_8 NS_371 0 1.7798919805811240e-04
GC_8_372 b_8 NI_8 NS_372 0 -5.8431438129054612e-05
GC_8_373 b_8 NI_8 NS_373 0 -8.3320149059618518e-06
GC_8_374 b_8 NI_8 NS_374 0 -1.8244211428170002e-05
GC_8_375 b_8 NI_8 NS_375 0 4.3794128966736336e-06
GC_8_376 b_8 NI_8 NS_376 0 -3.4524980505818874e-06
GC_8_377 b_8 NI_8 NS_377 0 4.7232566251657871e-06
GC_8_378 b_8 NI_8 NS_378 0 2.2794910311728148e-06
GC_8_379 b_8 NI_8 NS_379 0 9.3957677778344759e-06
GC_8_380 b_8 NI_8 NS_380 0 2.8025186589905643e-05
GC_8_381 b_8 NI_8 NS_381 0 2.8297154795743438e-02
GC_8_382 b_8 NI_8 NS_382 0 1.2246467983558689e-03
GC_8_383 b_8 NI_8 NS_383 0 -1.6132337420508278e-02
GC_8_384 b_8 NI_8 NS_384 0 4.6064867323175147e-03
GC_8_385 b_8 NI_8 NS_385 0 -1.8478216740815790e-04
GC_8_386 b_8 NI_8 NS_386 0 2.2349568838709984e-05
GC_8_387 b_8 NI_8 NS_387 0 -3.0699506901544379e-05
GC_8_388 b_8 NI_8 NS_388 0 -2.3502102580789786e-05
GC_8_389 b_8 NI_8 NS_389 0 -6.7574240948204377e-03
GC_8_390 b_8 NI_8 NS_390 0 -5.1973173953047099e-03
GC_8_391 b_8 NI_8 NS_391 0 2.4010533293720503e-05
GC_8_392 b_8 NI_8 NS_392 0 8.4647330984192373e-06
GC_8_393 b_8 NI_8 NS_393 0 9.5680607181625604e-03
GC_8_394 b_8 NI_8 NS_394 0 3.5539559523425045e-03
GC_8_395 b_8 NI_8 NS_395 0 7.1087483862184915e-06
GC_8_396 b_8 NI_8 NS_396 0 2.2745072323852721e-05
GC_8_397 b_8 NI_8 NS_397 0 1.2237726089310596e-05
GC_8_398 b_8 NI_8 NS_398 0 1.0377902862393515e-05
GC_8_399 b_8 NI_8 NS_399 0 -1.3763294106940889e-05
GC_8_400 b_8 NI_8 NS_400 0 -2.4632484855183445e-05
GC_8_401 b_8 NI_8 NS_401 0 1.4186591373960014e-05
GC_8_402 b_8 NI_8 NS_402 0 -2.1387179134397884e-06
GC_8_403 b_8 NI_8 NS_403 0 -3.4617925165965329e-03
GC_8_404 b_8 NI_8 NS_404 0 -3.5295011324543157e-04
GC_8_405 b_8 NI_8 NS_405 0 -1.8078946594143186e-04
GC_8_406 b_8 NI_8 NS_406 0 -4.3805294607143753e-05
GC_8_407 b_8 NI_8 NS_407 0 7.3200114904677408e-04
GC_8_408 b_8 NI_8 NS_408 0 4.4593049467913450e-04
GC_8_409 b_8 NI_8 NS_409 0 2.5334491170446238e-04
GC_8_410 b_8 NI_8 NS_410 0 -2.9257227275923859e-04
GC_8_411 b_8 NI_8 NS_411 0 -8.4269998886085380e-05
GC_8_412 b_8 NI_8 NS_412 0 -2.4066527969983921e-05
GC_8_413 b_8 NI_8 NS_413 0 -1.2715345111585833e-05
GC_8_414 b_8 NI_8 NS_414 0 -5.0281232220395564e-06
GC_8_415 b_8 NI_8 NS_415 0 -4.7195189734775557e-05
GC_8_416 b_8 NI_8 NS_416 0 1.9038928760654751e-05
GC_8_417 b_8 NI_8 NS_417 0 -1.7447400822591291e-07
GC_8_418 b_8 NI_8 NS_418 0 -8.9067774978087589e-06
GC_8_419 b_8 NI_8 NS_419 0 -1.2024433379659185e-02
GC_8_420 b_8 NI_8 NS_420 0 -1.2442109045579207e-03
GC_8_421 b_8 NI_8 NS_421 0 -1.0347567126437588e-03
GC_8_422 b_8 NI_8 NS_422 0 6.3022529176531292e-03
GC_8_423 b_8 NI_8 NS_423 0 -1.0767891859427630e-04
GC_8_424 b_8 NI_8 NS_424 0 1.3149046397893633e-04
GC_8_425 b_8 NI_8 NS_425 0 -1.7619034737817181e-05
GC_8_426 b_8 NI_8 NS_426 0 2.5005051235902252e-05
GC_8_427 b_8 NI_8 NS_427 0 6.4245074773071507e-03
GC_8_428 b_8 NI_8 NS_428 0 5.3972795590063426e-03
GC_8_429 b_8 NI_8 NS_429 0 -2.0900525773201872e-05
GC_8_430 b_8 NI_8 NS_430 0 -9.3292573121341445e-06
GC_8_431 b_8 NI_8 NS_431 0 1.0828321284358686e-02
GC_8_432 b_8 NI_8 NS_432 0 -2.3432928089228426e-03
GC_8_433 b_8 NI_8 NS_433 0 1.4900248939487674e-06
GC_8_434 b_8 NI_8 NS_434 0 2.6190485214042985e-05
GC_8_435 b_8 NI_8 NS_435 0 -2.0215352034863811e-06
GC_8_436 b_8 NI_8 NS_436 0 1.9913358433729285e-05
GC_8_437 b_8 NI_8 NS_437 0 -9.8157715280737369e-06
GC_8_438 b_8 NI_8 NS_438 0 -1.7651170899028115e-05
GC_8_439 b_8 NI_8 NS_439 0 1.2915118200176349e-05
GC_8_440 b_8 NI_8 NS_440 0 -1.9935660814462444e-06
GC_8_441 b_8 NI_8 NS_441 0 -3.7951734444448821e-03
GC_8_442 b_8 NI_8 NS_442 0 7.3353535760163960e-04
GC_8_443 b_8 NI_8 NS_443 0 -5.4173872003808263e-05
GC_8_444 b_8 NI_8 NS_444 0 -2.7771820885448279e-04
GC_8_445 b_8 NI_8 NS_445 0 5.5434420268272023e-04
GC_8_446 b_8 NI_8 NS_446 0 4.3605653007613103e-04
GC_8_447 b_8 NI_8 NS_447 0 3.1508650867247579e-04
GC_8_448 b_8 NI_8 NS_448 0 -1.6637727118000783e-04
GC_8_449 b_8 NI_8 NS_449 0 -5.4558664553268218e-05
GC_8_450 b_8 NI_8 NS_450 0 -6.1811172781022720e-05
GC_8_451 b_8 NI_8 NS_451 0 -5.2605692122670523e-06
GC_8_452 b_8 NI_8 NS_452 0 -2.0217799158825165e-05
GC_8_453 b_8 NI_8 NS_453 0 -6.2970224657927734e-05
GC_8_454 b_8 NI_8 NS_454 0 -3.4757401194867292e-05
GC_8_455 b_8 NI_8 NS_455 0 -7.8834052236581859e-06
GC_8_456 b_8 NI_8 NS_456 0 -7.1414417023166478e-07
GD_8_1 b_8 NI_8 NA_1 0 -5.6748397637676768e-03
GD_8_2 b_8 NI_8 NA_2 0 3.0898138514031258e-03
GD_8_3 b_8 NI_8 NA_3 0 -2.1882992235460839e-03
GD_8_4 b_8 NI_8 NA_4 0 -4.7772950745000268e-03
GD_8_5 b_8 NI_8 NA_5 0 1.0065895716837824e-02
GD_8_6 b_8 NI_8 NA_6 0 -5.9230547200081205e-03
GD_8_7 b_8 NI_8 NA_7 0 -2.1049566512056674e-02
GD_8_8 b_8 NI_8 NA_8 0 -1.3750158455180100e-01
GD_8_9 b_8 NI_8 NA_9 0 9.2424307347686776e-03
GD_8_10 b_8 NI_8 NA_10 0 -5.7611603571999046e-03
GD_8_11 b_8 NI_8 NA_11 0 -1.1769257409425761e-02
GD_8_12 b_8 NI_8 NA_12 0 1.9486947452406419e-04
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 1.1317846909168554e-02
GC_9_2 b_9 NI_9 NS_2 0 -7.4996209223750221e-04
GC_9_3 b_9 NI_9 NS_3 0 -1.1349914246277234e-02
GC_9_4 b_9 NI_9 NS_4 0 6.3516953002048116e-03
GC_9_5 b_9 NI_9 NS_5 0 4.2981285794357508e-04
GC_9_6 b_9 NI_9 NS_6 0 -6.0569243150607860e-04
GC_9_7 b_9 NI_9 NS_7 0 1.5495008814622911e-04
GC_9_8 b_9 NI_9 NS_8 0 -1.5851044536326918e-04
GC_9_9 b_9 NI_9 NS_9 0 7.1863970781915092e-04
GC_9_10 b_9 NI_9 NS_10 0 -4.9678857769805415e-03
GC_9_11 b_9 NI_9 NS_11 0 -1.9006975440549182e-05
GC_9_12 b_9 NI_9 NS_12 0 3.9729465420012817e-05
GC_9_13 b_9 NI_9 NS_13 0 7.1329700573697155e-03
GC_9_14 b_9 NI_9 NS_14 0 1.0861145264091634e-03
GC_9_15 b_9 NI_9 NS_15 0 -2.6156627482817244e-05
GC_9_16 b_9 NI_9 NS_16 0 1.0729414119782133e-05
GC_9_17 b_9 NI_9 NS_17 0 -2.8017541769606065e-05
GC_9_18 b_9 NI_9 NS_18 0 3.9785805505329395e-05
GC_9_19 b_9 NI_9 NS_19 0 1.3432539216401369e-04
GC_9_20 b_9 NI_9 NS_20 0 -1.0815765844283430e-06
GC_9_21 b_9 NI_9 NS_21 0 4.4661571027535008e-05
GC_9_22 b_9 NI_9 NS_22 0 3.4175002446302435e-05
GC_9_23 b_9 NI_9 NS_23 0 -1.1001500825620436e-03
GC_9_24 b_9 NI_9 NS_24 0 1.2466326469056765e-03
GC_9_25 b_9 NI_9 NS_25 0 -1.4387290870435560e-04
GC_9_26 b_9 NI_9 NS_26 0 -5.6899670426060556e-04
GC_9_27 b_9 NI_9 NS_27 0 9.2176364879940559e-05
GC_9_28 b_9 NI_9 NS_28 0 -3.2726725055553239e-04
GC_9_29 b_9 NI_9 NS_29 0 -1.3793730350241561e-04
GC_9_30 b_9 NI_9 NS_30 0 2.1575653114539657e-04
GC_9_31 b_9 NI_9 NS_31 0 -2.8127144537810374e-05
GC_9_32 b_9 NI_9 NS_32 0 -6.3699364599758006e-05
GC_9_33 b_9 NI_9 NS_33 0 -2.8324406061405524e-05
GC_9_34 b_9 NI_9 NS_34 0 3.5070483877531103e-05
GC_9_35 b_9 NI_9 NS_35 0 -3.5357340706684911e-06
GC_9_36 b_9 NI_9 NS_36 0 7.1642899279759182e-05
GC_9_37 b_9 NI_9 NS_37 0 1.7217129568183952e-05
GC_9_38 b_9 NI_9 NS_38 0 -2.3061900515346572e-05
GC_9_39 b_9 NI_9 NS_39 0 -6.7356598241214280e-03
GC_9_40 b_9 NI_9 NS_40 0 8.2734071811470331e-04
GC_9_41 b_9 NI_9 NS_41 0 1.0004116334779818e-03
GC_9_42 b_9 NI_9 NS_42 0 -9.2292258028096995e-03
GC_9_43 b_9 NI_9 NS_43 0 -3.7290995368841931e-06
GC_9_44 b_9 NI_9 NS_44 0 8.0043085120871428e-04
GC_9_45 b_9 NI_9 NS_45 0 3.8383281640492193e-05
GC_9_46 b_9 NI_9 NS_46 0 1.3981021004995969e-04
GC_9_47 b_9 NI_9 NS_47 0 2.1076518538504239e-05
GC_9_48 b_9 NI_9 NS_48 0 7.0555444534625214e-03
GC_9_49 b_9 NI_9 NS_49 0 2.2150435451787994e-05
GC_9_50 b_9 NI_9 NS_50 0 -3.1865290876123054e-05
GC_9_51 b_9 NI_9 NS_51 0 2.8332225129098089e-04
GC_9_52 b_9 NI_9 NS_52 0 3.7445680827114494e-03
GC_9_53 b_9 NI_9 NS_53 0 4.8671932700318945e-05
GC_9_54 b_9 NI_9 NS_54 0 6.0519247532071576e-05
GC_9_55 b_9 NI_9 NS_55 0 -1.5301196958295103e-05
GC_9_56 b_9 NI_9 NS_56 0 8.8606400887231070e-05
GC_9_57 b_9 NI_9 NS_57 0 1.8994450202642704e-05
GC_9_58 b_9 NI_9 NS_58 0 2.0650509051951945e-05
GC_9_59 b_9 NI_9 NS_59 0 7.3548899092420572e-05
GC_9_60 b_9 NI_9 NS_60 0 5.0569615428426661e-05
GC_9_61 b_9 NI_9 NS_61 0 -1.5520368945437929e-03
GC_9_62 b_9 NI_9 NS_62 0 9.3328118619805261e-05
GC_9_63 b_9 NI_9 NS_63 0 2.2341433470965356e-04
GC_9_64 b_9 NI_9 NS_64 0 -5.9917130291025299e-04
GC_9_65 b_9 NI_9 NS_65 0 1.8599127156008493e-04
GC_9_66 b_9 NI_9 NS_66 0 -2.9580204084492966e-04
GC_9_67 b_9 NI_9 NS_67 0 -1.2185274036026872e-04
GC_9_68 b_9 NI_9 NS_68 0 1.6010891160465513e-04
GC_9_69 b_9 NI_9 NS_69 0 2.5411546232834217e-05
GC_9_70 b_9 NI_9 NS_70 0 -6.7811011127050214e-05
GC_9_71 b_9 NI_9 NS_71 0 -2.6913042009196982e-05
GC_9_72 b_9 NI_9 NS_72 0 6.8254596859998787e-06
GC_9_73 b_9 NI_9 NS_73 0 -3.1762904185281503e-05
GC_9_74 b_9 NI_9 NS_74 0 6.7560569555513372e-05
GC_9_75 b_9 NI_9 NS_75 0 5.8021985107358573e-06
GC_9_76 b_9 NI_9 NS_76 0 6.4614343203871718e-07
GC_9_77 b_9 NI_9 NS_77 0 4.2067826467191496e-03
GC_9_78 b_9 NI_9 NS_78 0 -1.1129306658367050e-03
GC_9_79 b_9 NI_9 NS_79 0 -8.5750357551100942e-03
GC_9_80 b_9 NI_9 NS_80 0 5.7767702739952922e-03
GC_9_81 b_9 NI_9 NS_81 0 6.9631235485622626e-04
GC_9_82 b_9 NI_9 NS_82 0 -2.2695997482215883e-04
GC_9_83 b_9 NI_9 NS_83 0 1.9031227212822121e-04
GC_9_84 b_9 NI_9 NS_84 0 -1.4908480119933448e-04
GC_9_85 b_9 NI_9 NS_85 0 2.5814904204589846e-03
GC_9_86 b_9 NI_9 NS_86 0 -4.7567008128469737e-03
GC_9_87 b_9 NI_9 NS_87 0 -2.0078536995327253e-05
GC_9_88 b_9 NI_9 NS_88 0 3.9966635048464217e-05
GC_9_89 b_9 NI_9 NS_89 0 8.5037714248666681e-03
GC_9_90 b_9 NI_9 NS_90 0 2.2810105944712387e-03
GC_9_91 b_9 NI_9 NS_91 0 -4.9935997119355270e-06
GC_9_92 b_9 NI_9 NS_92 0 -6.8607536271045349e-06
GC_9_93 b_9 NI_9 NS_93 0 -2.8732385516456630e-05
GC_9_94 b_9 NI_9 NS_94 0 4.8234664563478642e-05
GC_9_95 b_9 NI_9 NS_95 0 1.4192795760467343e-04
GC_9_96 b_9 NI_9 NS_96 0 1.0455911537463721e-05
GC_9_97 b_9 NI_9 NS_97 0 4.1046190970473911e-05
GC_9_98 b_9 NI_9 NS_98 0 2.4656107968712888e-05
GC_9_99 b_9 NI_9 NS_99 0 -2.1812850937461842e-03
GC_9_100 b_9 NI_9 NS_100 0 -3.9477110509401756e-04
GC_9_101 b_9 NI_9 NS_101 0 -1.6432132904675329e-04
GC_9_102 b_9 NI_9 NS_102 0 -4.2855348306879333e-04
GC_9_103 b_9 NI_9 NS_103 0 2.7431652131619619e-04
GC_9_104 b_9 NI_9 NS_104 0 1.6460290356926316e-05
GC_9_105 b_9 NI_9 NS_105 0 3.1324875752324771e-06
GC_9_106 b_9 NI_9 NS_106 0 4.9385224734606252e-05
GC_9_107 b_9 NI_9 NS_107 0 -9.3997448024606568e-06
GC_9_108 b_9 NI_9 NS_108 0 -1.9125069423998065e-05
GC_9_109 b_9 NI_9 NS_109 0 -1.6169992414524030e-05
GC_9_110 b_9 NI_9 NS_110 0 2.0283494595593792e-05
GC_9_111 b_9 NI_9 NS_111 0 -4.4479276537857836e-06
GC_9_112 b_9 NI_9 NS_112 0 6.6246393070713337e-05
GC_9_113 b_9 NI_9 NS_113 0 1.9521411808189205e-05
GC_9_114 b_9 NI_9 NS_114 0 8.2199544208150993e-06
GC_9_115 b_9 NI_9 NS_115 0 7.1472111691862359e-03
GC_9_116 b_9 NI_9 NS_116 0 1.1225186416300270e-03
GC_9_117 b_9 NI_9 NS_117 0 -5.9685641258190886e-03
GC_9_118 b_9 NI_9 NS_118 0 -5.5599305444885812e-03
GC_9_119 b_9 NI_9 NS_119 0 3.1555540495829292e-05
GC_9_120 b_9 NI_9 NS_120 0 5.9865771796870657e-04
GC_9_121 b_9 NI_9 NS_121 0 9.9759916442992218e-05
GC_9_122 b_9 NI_9 NS_122 0 1.6334922023101295e-04
GC_9_123 b_9 NI_9 NS_123 0 -1.7806241626158405e-03
GC_9_124 b_9 NI_9 NS_124 0 5.9238109280109041e-03
GC_9_125 b_9 NI_9 NS_125 0 2.3591994635792472e-05
GC_9_126 b_9 NI_9 NS_126 0 -3.1794465650556350e-05
GC_9_127 b_9 NI_9 NS_127 0 3.0199844776659956e-03
GC_9_128 b_9 NI_9 NS_128 0 6.4399034581179666e-03
GC_9_129 b_9 NI_9 NS_129 0 5.2755109251917821e-05
GC_9_130 b_9 NI_9 NS_130 0 3.7785179183352527e-05
GC_9_131 b_9 NI_9 NS_131 0 -9.9972118822922724e-06
GC_9_132 b_9 NI_9 NS_132 0 8.0791505042817144e-05
GC_9_133 b_9 NI_9 NS_133 0 7.8379289181548868e-05
GC_9_134 b_9 NI_9 NS_134 0 4.6936552188083872e-05
GC_9_135 b_9 NI_9 NS_135 0 7.5986283828544557e-05
GC_9_136 b_9 NI_9 NS_136 0 4.3037380953136219e-05
GC_9_137 b_9 NI_9 NS_137 0 -2.5617243920460888e-03
GC_9_138 b_9 NI_9 NS_138 0 -1.1726537634188985e-03
GC_9_139 b_9 NI_9 NS_139 0 2.3700120237656448e-04
GC_9_140 b_9 NI_9 NS_140 0 -5.3062445546570892e-04
GC_9_141 b_9 NI_9 NS_141 0 4.1876523776095565e-04
GC_9_142 b_9 NI_9 NS_142 0 1.5535967855127863e-05
GC_9_143 b_9 NI_9 NS_143 0 -2.5761325501375171e-05
GC_9_144 b_9 NI_9 NS_144 0 2.0424502628397802e-05
GC_9_145 b_9 NI_9 NS_145 0 4.6496898283326888e-06
GC_9_146 b_9 NI_9 NS_146 0 -2.3589861617407522e-05
GC_9_147 b_9 NI_9 NS_147 0 -2.3101843972903341e-05
GC_9_148 b_9 NI_9 NS_148 0 7.3311779801843317e-06
GC_9_149 b_9 NI_9 NS_149 0 -1.2044537963404091e-05
GC_9_150 b_9 NI_9 NS_150 0 4.6556792854740533e-05
GC_9_151 b_9 NI_9 NS_151 0 7.2529010180875736e-06
GC_9_152 b_9 NI_9 NS_152 0 7.5927115370154787e-06
GC_9_153 b_9 NI_9 NS_153 0 -1.8458570578173916e-02
GC_9_154 b_9 NI_9 NS_154 0 -1.2992302062736607e-03
GC_9_155 b_9 NI_9 NS_155 0 6.6807679844281828e-03
GC_9_156 b_9 NI_9 NS_156 0 1.1259901687325139e-02
GC_9_157 b_9 NI_9 NS_157 0 6.4840587871553513e-04
GC_9_158 b_9 NI_9 NS_158 0 7.7943032507661212e-04
GC_9_159 b_9 NI_9 NS_159 0 2.0724747859150378e-04
GC_9_160 b_9 NI_9 NS_160 0 -8.8605641203122807e-05
GC_9_161 b_9 NI_9 NS_161 0 6.8035709786535481e-03
GC_9_162 b_9 NI_9 NS_162 0 4.2614827044972622e-03
GC_9_163 b_9 NI_9 NS_163 0 -1.0369154422193501e-05
GC_9_164 b_9 NI_9 NS_164 0 5.9754201010277255e-07
GC_9_165 b_9 NI_9 NS_165 0 1.2412887755124950e-02
GC_9_166 b_9 NI_9 NS_166 0 -9.3231865013479170e-03
GC_9_167 b_9 NI_9 NS_167 0 5.0526679156251888e-06
GC_9_168 b_9 NI_9 NS_168 0 -1.1262527017345053e-05
GC_9_169 b_9 NI_9 NS_169 0 -3.8782744082103667e-05
GC_9_170 b_9 NI_9 NS_170 0 6.8361256916129692e-05
GC_9_171 b_9 NI_9 NS_171 0 -5.0518868627619856e-06
GC_9_172 b_9 NI_9 NS_172 0 -3.5392426408159015e-05
GC_9_173 b_9 NI_9 NS_173 0 -1.0250114836097576e-05
GC_9_174 b_9 NI_9 NS_174 0 -7.7961387274425920e-07
GC_9_175 b_9 NI_9 NS_175 0 -3.9060152856283149e-03
GC_9_176 b_9 NI_9 NS_176 0 3.3805389120997015e-03
GC_9_177 b_9 NI_9 NS_177 0 -3.3049530117038284e-04
GC_9_178 b_9 NI_9 NS_178 0 -5.6535378714512371e-04
GC_9_179 b_9 NI_9 NS_179 0 4.1296670869508072e-04
GC_9_180 b_9 NI_9 NS_180 0 -2.7804546597949120e-04
GC_9_181 b_9 NI_9 NS_181 0 -4.7327208213053721e-05
GC_9_182 b_9 NI_9 NS_182 0 1.8362586347399990e-05
GC_9_183 b_9 NI_9 NS_183 0 3.0442468559524016e-05
GC_9_184 b_9 NI_9 NS_184 0 2.3584987270137939e-05
GC_9_185 b_9 NI_9 NS_185 0 9.3130662535285868e-06
GC_9_186 b_9 NI_9 NS_186 0 -8.5491721310445514e-06
GC_9_187 b_9 NI_9 NS_187 0 2.5839611868826467e-05
GC_9_188 b_9 NI_9 NS_188 0 1.0007697354826691e-04
GC_9_189 b_9 NI_9 NS_189 0 6.1105615013979650e-05
GC_9_190 b_9 NI_9 NS_190 0 3.5028443535479024e-06
GC_9_191 b_9 NI_9 NS_191 0 1.9370008079876429e-02
GC_9_192 b_9 NI_9 NS_192 0 1.3407414668932672e-03
GC_9_193 b_9 NI_9 NS_193 0 -1.1044871577328049e-02
GC_9_194 b_9 NI_9 NS_194 0 1.4728989695773137e-03
GC_9_195 b_9 NI_9 NS_195 0 -1.1271923567607490e-05
GC_9_196 b_9 NI_9 NS_196 0 6.0769933292453902e-04
GC_9_197 b_9 NI_9 NS_197 0 8.5156505779864126e-05
GC_9_198 b_9 NI_9 NS_198 0 3.9725213477171023e-05
GC_9_199 b_9 NI_9 NS_199 0 -7.2712345802166799e-03
GC_9_200 b_9 NI_9 NS_200 0 -4.6381214841478618e-03
GC_9_201 b_9 NI_9 NS_201 0 1.5243686596368601e-05
GC_9_202 b_9 NI_9 NS_202 0 2.7639759709437234e-06
GC_9_203 b_9 NI_9 NS_203 0 9.1275708751375612e-03
GC_9_204 b_9 NI_9 NS_204 0 -2.0116506356940597e-03
GC_9_205 b_9 NI_9 NS_205 0 1.9256385896365345e-05
GC_9_206 b_9 NI_9 NS_206 0 5.2896859990754580e-06
GC_9_207 b_9 NI_9 NS_207 0 -7.3248183816056737e-06
GC_9_208 b_9 NI_9 NS_208 0 3.9500880507983919e-05
GC_9_209 b_9 NI_9 NS_209 0 -2.2515852979356737e-05
GC_9_210 b_9 NI_9 NS_210 0 2.3587931829221904e-06
GC_9_211 b_9 NI_9 NS_211 0 1.0456095974342807e-05
GC_9_212 b_9 NI_9 NS_212 0 9.3933019081355003e-07
GC_9_213 b_9 NI_9 NS_213 0 -3.7796532470370158e-03
GC_9_214 b_9 NI_9 NS_214 0 2.2710480241147266e-03
GC_9_215 b_9 NI_9 NS_215 0 -1.6970201057722387e-04
GC_9_216 b_9 NI_9 NS_216 0 -3.9402012322136120e-04
GC_9_217 b_9 NI_9 NS_217 0 3.5638748653454860e-04
GC_9_218 b_9 NI_9 NS_218 0 -1.0417493368696448e-04
GC_9_219 b_9 NI_9 NS_219 0 2.1207830011539976e-05
GC_9_220 b_9 NI_9 NS_220 0 3.6308683577401984e-05
GC_9_221 b_9 NI_9 NS_221 0 -3.7965160385089195e-05
GC_9_222 b_9 NI_9 NS_222 0 2.2866453998489001e-05
GC_9_223 b_9 NI_9 NS_223 0 2.4354667566221720e-05
GC_9_224 b_9 NI_9 NS_224 0 3.1140423487043586e-05
GC_9_225 b_9 NI_9 NS_225 0 1.0021621536003254e-05
GC_9_226 b_9 NI_9 NS_226 0 1.0974635683771028e-04
GC_9_227 b_9 NI_9 NS_227 0 4.5625773606299996e-05
GC_9_228 b_9 NI_9 NS_228 0 2.0911045641551760e-05
GC_9_229 b_9 NI_9 NS_229 0 -3.5977709462462907e-03
GC_9_230 b_9 NI_9 NS_230 0 -1.5461173173129980e-03
GC_9_231 b_9 NI_9 NS_231 0 -4.0516485870699197e-04
GC_9_232 b_9 NI_9 NS_232 0 5.9781605552543648e-03
GC_9_233 b_9 NI_9 NS_233 0 -1.4785880317639822e-03
GC_9_234 b_9 NI_9 NS_234 0 6.6776346815027845e-04
GC_9_235 b_9 NI_9 NS_235 0 -1.2692552700586628e-04
GC_9_236 b_9 NI_9 NS_236 0 2.9241847670888462e-05
GC_9_237 b_9 NI_9 NS_237 0 5.8380267635876615e-03
GC_9_238 b_9 NI_9 NS_238 0 1.1797757476155473e-02
GC_9_239 b_9 NI_9 NS_239 0 -2.2053576729776790e-05
GC_9_240 b_9 NI_9 NS_240 0 -7.1738644701531505e-06
GC_9_241 b_9 NI_9 NS_241 0 7.2097659349842176e-03
GC_9_242 b_9 NI_9 NS_242 0 -4.8474732482815600e-03
GC_9_243 b_9 NI_9 NS_243 0 -4.4856586051763419e-06
GC_9_244 b_9 NI_9 NS_244 0 -1.8274377433869869e-05
GC_9_245 b_9 NI_9 NS_245 0 -3.0872943530322502e-05
GC_9_246 b_9 NI_9 NS_246 0 4.7704093681313354e-05
GC_9_247 b_9 NI_9 NS_247 0 -3.3950532858020239e-05
GC_9_248 b_9 NI_9 NS_248 0 -5.2531876338285056e-05
GC_9_249 b_9 NI_9 NS_249 0 5.8096170953312290e-07
GC_9_250 b_9 NI_9 NS_250 0 -8.6793507933413432e-06
GC_9_251 b_9 NI_9 NS_251 0 -6.2435638071343278e-03
GC_9_252 b_9 NI_9 NS_252 0 1.2505554317875311e-03
GC_9_253 b_9 NI_9 NS_253 0 -2.9966899900690764e-04
GC_9_254 b_9 NI_9 NS_254 0 -3.8477894442332335e-04
GC_9_255 b_9 NI_9 NS_255 0 7.3896027545717214e-04
GC_9_256 b_9 NI_9 NS_256 0 2.7349328783128630e-05
GC_9_257 b_9 NI_9 NS_257 0 1.0899243380228496e-04
GC_9_258 b_9 NI_9 NS_258 0 -2.0158806936307149e-04
GC_9_259 b_9 NI_9 NS_259 0 6.5136392619110667e-06
GC_9_260 b_9 NI_9 NS_260 0 1.3315515239115227e-05
GC_9_261 b_9 NI_9 NS_261 0 -7.3988222451200766e-06
GC_9_262 b_9 NI_9 NS_262 0 2.3589107798274814e-05
GC_9_263 b_9 NI_9 NS_263 0 4.2782929663923133e-05
GC_9_264 b_9 NI_9 NS_264 0 3.3571612379238611e-06
GC_9_265 b_9 NI_9 NS_265 0 1.3087777777090761e-06
GC_9_266 b_9 NI_9 NS_266 0 9.6873893269206259e-06
GC_9_267 b_9 NI_9 NS_267 0 -2.5745354540253479e-02
GC_9_268 b_9 NI_9 NS_268 0 1.4965376926811475e-03
GC_9_269 b_9 NI_9 NS_269 0 1.5315578048357852e-02
GC_9_270 b_9 NI_9 NS_270 0 3.2312461848881505e-03
GC_9_271 b_9 NI_9 NS_271 0 -4.4270981279000691e-05
GC_9_272 b_9 NI_9 NS_272 0 3.5369900752481731e-05
GC_9_273 b_9 NI_9 NS_273 0 -5.4379372455174740e-06
GC_9_274 b_9 NI_9 NS_274 0 -1.3017535263879351e-05
GC_9_275 b_9 NI_9 NS_275 0 -7.0736360678231901e-03
GC_9_276 b_9 NI_9 NS_276 0 -1.0892381103453797e-02
GC_9_277 b_9 NI_9 NS_277 0 2.5449279997197973e-05
GC_9_278 b_9 NI_9 NS_278 0 1.0189729737277478e-05
GC_9_279 b_9 NI_9 NS_279 0 9.5301436641444803e-03
GC_9_280 b_9 NI_9 NS_280 0 -1.3616712848149439e-02
GC_9_281 b_9 NI_9 NS_281 0 -2.2046047045552154e-06
GC_9_282 b_9 NI_9 NS_282 0 5.8090006668073752e-06
GC_9_283 b_9 NI_9 NS_283 0 -1.1423730996034475e-05
GC_9_284 b_9 NI_9 NS_284 0 3.9426785195992757e-05
GC_9_285 b_9 NI_9 NS_285 0 -1.0480500437734298e-05
GC_9_286 b_9 NI_9 NS_286 0 -2.2687676885996928e-05
GC_9_287 b_9 NI_9 NS_287 0 1.8238792981375619e-05
GC_9_288 b_9 NI_9 NS_288 0 -2.9463018871039155e-06
GC_9_289 b_9 NI_9 NS_289 0 -5.1152167972296839e-03
GC_9_290 b_9 NI_9 NS_290 0 8.2609025226963089e-04
GC_9_291 b_9 NI_9 NS_291 0 -1.6161617382377455e-04
GC_9_292 b_9 NI_9 NS_292 0 -3.1631441119582960e-04
GC_9_293 b_9 NI_9 NS_293 0 6.0854893106374009e-04
GC_9_294 b_9 NI_9 NS_294 0 2.1539245663147548e-04
GC_9_295 b_9 NI_9 NS_295 0 1.6376869698170950e-04
GC_9_296 b_9 NI_9 NS_296 0 -1.1784623911383725e-04
GC_9_297 b_9 NI_9 NS_297 0 -1.3254416909790467e-05
GC_9_298 b_9 NI_9 NS_298 0 1.1335205198773640e-05
GC_9_299 b_9 NI_9 NS_299 0 -1.8346957020651098e-05
GC_9_300 b_9 NI_9 NS_300 0 9.8695836189060627e-06
GC_9_301 b_9 NI_9 NS_301 0 3.7853865648077903e-05
GC_9_302 b_9 NI_9 NS_302 0 3.3542233740124151e-05
GC_9_303 b_9 NI_9 NS_303 0 -3.5988201737895024e-06
GC_9_304 b_9 NI_9 NS_304 0 6.3676203424591225e-06
GC_9_305 b_9 NI_9 NS_305 0 3.3615911392428269e-02
GC_9_306 b_9 NI_9 NS_306 0 -1.8239320146785981e-03
GC_9_307 b_9 NI_9 NS_307 0 5.3940324068789618e-02
GC_9_308 b_9 NI_9 NS_308 0 -6.8253605372553358e-02
GC_9_309 b_9 NI_9 NS_309 0 -2.6863291885298990e-03
GC_9_310 b_9 NI_9 NS_310 0 -1.0631900225639317e-03
GC_9_311 b_9 NI_9 NS_311 0 -4.6008082633728427e-04
GC_9_312 b_9 NI_9 NS_312 0 1.1650505655785578e-04
GC_9_313 b_9 NI_9 NS_313 0 -8.9905474291296483e-03
GC_9_314 b_9 NI_9 NS_314 0 1.6549385490036383e-02
GC_9_315 b_9 NI_9 NS_315 0 -4.0162814944679759e-05
GC_9_316 b_9 NI_9 NS_316 0 -9.5760859653042007e-05
GC_9_317 b_9 NI_9 NS_317 0 -4.1561918444982970e-02
GC_9_318 b_9 NI_9 NS_318 0 8.4174136174726532e-03
GC_9_319 b_9 NI_9 NS_319 0 -7.8097199005751136e-05
GC_9_320 b_9 NI_9 NS_320 0 -3.7565354332188621e-05
GC_9_321 b_9 NI_9 NS_321 0 -7.6367681399253085e-05
GC_9_322 b_9 NI_9 NS_322 0 8.7336607431034920e-05
GC_9_323 b_9 NI_9 NS_323 0 -1.9183451748169873e-04
GC_9_324 b_9 NI_9 NS_324 0 -9.5236596667179187e-05
GC_9_325 b_9 NI_9 NS_325 0 -3.7648588992257272e-05
GC_9_326 b_9 NI_9 NS_326 0 -3.8268280200710054e-05
GC_9_327 b_9 NI_9 NS_327 0 -8.0752411485829258e-03
GC_9_328 b_9 NI_9 NS_328 0 3.8247640451628795e-03
GC_9_329 b_9 NI_9 NS_329 0 -2.6106628219185708e-04
GC_9_330 b_9 NI_9 NS_330 0 -4.7138674605787478e-04
GC_9_331 b_9 NI_9 NS_331 0 6.6426048994132434e-04
GC_9_332 b_9 NI_9 NS_332 0 8.2066035082568019e-05
GC_9_333 b_9 NI_9 NS_333 0 8.4327715952289148e-05
GC_9_334 b_9 NI_9 NS_334 0 -1.3649504059648712e-04
GC_9_335 b_9 NI_9 NS_335 0 -1.0317793012824025e-05
GC_9_336 b_9 NI_9 NS_336 0 8.6081399959687983e-06
GC_9_337 b_9 NI_9 NS_337 0 2.2066249970220835e-05
GC_9_338 b_9 NI_9 NS_338 0 -1.9013679249819626e-06
GC_9_339 b_9 NI_9 NS_339 0 -6.2137459788323175e-06
GC_9_340 b_9 NI_9 NS_340 0 2.3091889141764406e-05
GC_9_341 b_9 NI_9 NS_341 0 4.4029298004566510e-06
GC_9_342 b_9 NI_9 NS_342 0 1.7298660109007575e-05
GC_9_343 b_9 NI_9 NS_343 0 3.8119423149045102e-02
GC_9_344 b_9 NI_9 NS_344 0 2.2971178845214522e-03
GC_9_345 b_9 NI_9 NS_345 0 1.2353684121591803e-02
GC_9_346 b_9 NI_9 NS_346 0 -1.9939009732102601e-02
GC_9_347 b_9 NI_9 NS_347 0 1.5278508017496320e-03
GC_9_348 b_9 NI_9 NS_348 0 3.5031091715703395e-05
GC_9_349 b_9 NI_9 NS_349 0 4.1315897875601011e-05
GC_9_350 b_9 NI_9 NS_350 0 -7.0089271326092332e-06
GC_9_351 b_9 NI_9 NS_351 0 2.3295484863662359e-02
GC_9_352 b_9 NI_9 NS_352 0 1.8086309135933831e-03
GC_9_353 b_9 NI_9 NS_353 0 4.3610970443957944e-05
GC_9_354 b_9 NI_9 NS_354 0 9.1844388480353555e-05
GC_9_355 b_9 NI_9 NS_355 0 -4.3234578638930272e-02
GC_9_356 b_9 NI_9 NS_356 0 4.1033419292500428e-02
GC_9_357 b_9 NI_9 NS_357 0 -2.6657138388584630e-06
GC_9_358 b_9 NI_9 NS_358 0 -5.2305756345326379e-06
GC_9_359 b_9 NI_9 NS_359 0 -1.6873158405456550e-05
GC_9_360 b_9 NI_9 NS_360 0 7.9286578063751054e-05
GC_9_361 b_9 NI_9 NS_361 0 -8.9759983804186898e-05
GC_9_362 b_9 NI_9 NS_362 0 -2.6595067042051891e-05
GC_9_363 b_9 NI_9 NS_363 0 -3.2770294385636900e-05
GC_9_364 b_9 NI_9 NS_364 0 -2.7262810870137458e-05
GC_9_365 b_9 NI_9 NS_365 0 -4.6019021892612574e-03
GC_9_366 b_9 NI_9 NS_366 0 -1.7320656985325715e-03
GC_9_367 b_9 NI_9 NS_367 0 1.1156467732135068e-04
GC_9_368 b_9 NI_9 NS_368 0 -1.9781066761801006e-04
GC_9_369 b_9 NI_9 NS_369 0 3.5639383954378989e-04
GC_9_370 b_9 NI_9 NS_370 0 3.7496818599918463e-04
GC_9_371 b_9 NI_9 NS_371 0 1.7010908206913211e-04
GC_9_372 b_9 NI_9 NS_372 0 -3.0864861384420831e-05
GC_9_373 b_9 NI_9 NS_373 0 2.7422255109372638e-05
GC_9_374 b_9 NI_9 NS_374 0 3.4740371452733563e-07
GC_9_375 b_9 NI_9 NS_375 0 1.9365782872248011e-05
GC_9_376 b_9 NI_9 NS_376 0 1.6928810604587076e-05
GC_9_377 b_9 NI_9 NS_377 0 1.2643494950441816e-05
GC_9_378 b_9 NI_9 NS_378 0 4.9589104720033801e-05
GC_9_379 b_9 NI_9 NS_379 0 2.9057004280682399e-05
GC_9_380 b_9 NI_9 NS_380 0 -9.9991786833282200e-06
GC_9_381 b_9 NI_9 NS_381 0 -2.9758681962329933e-02
GC_9_382 b_9 NI_9 NS_382 0 -1.3212972475662955e-03
GC_9_383 b_9 NI_9 NS_383 0 1.8973426635920384e-02
GC_9_384 b_9 NI_9 NS_384 0 2.6527168163548592e-02
GC_9_385 b_9 NI_9 NS_385 0 -5.4241342184880876e-04
GC_9_386 b_9 NI_9 NS_386 0 9.5578595217108298e-04
GC_9_387 b_9 NI_9 NS_387 0 -2.6747221338567934e-04
GC_9_388 b_9 NI_9 NS_388 0 3.1348149335912141e-04
GC_9_389 b_9 NI_9 NS_389 0 1.3303980754570524e-02
GC_9_390 b_9 NI_9 NS_390 0 2.7451555401063293e-02
GC_9_391 b_9 NI_9 NS_391 0 -3.8837905278745543e-05
GC_9_392 b_9 NI_9 NS_392 0 -9.5372219309270662e-05
GC_9_393 b_9 NI_9 NS_393 0 2.1886915822181968e-02
GC_9_394 b_9 NI_9 NS_394 0 -2.2631570258835651e-02
GC_9_395 b_9 NI_9 NS_395 0 -5.0525371153022285e-05
GC_9_396 b_9 NI_9 NS_396 0 3.9152150965229183e-05
GC_9_397 b_9 NI_9 NS_397 0 2.1200187170393960e-06
GC_9_398 b_9 NI_9 NS_398 0 8.5625207000171122e-05
GC_9_399 b_9 NI_9 NS_399 0 -2.2649302449206121e-04
GC_9_400 b_9 NI_9 NS_400 0 -5.8352245949547796e-05
GC_9_401 b_9 NI_9 NS_401 0 -3.5799778335783432e-05
GC_9_402 b_9 NI_9 NS_402 0 -2.8441041298384344e-05
GC_9_403 b_9 NI_9 NS_403 0 -6.6681135069017782e-03
GC_9_404 b_9 NI_9 NS_404 0 7.8488431533054424e-03
GC_9_405 b_9 NI_9 NS_405 0 -5.0473766259451918e-04
GC_9_406 b_9 NI_9 NS_406 0 -2.2428286242269662e-04
GC_9_407 b_9 NI_9 NS_407 0 7.8076199286783953e-04
GC_9_408 b_9 NI_9 NS_408 0 9.5966782919948472e-05
GC_9_409 b_9 NI_9 NS_409 0 1.2484169720081143e-04
GC_9_410 b_9 NI_9 NS_410 0 -3.0756743818986229e-04
GC_9_411 b_9 NI_9 NS_411 0 8.9479459476694239e-06
GC_9_412 b_9 NI_9 NS_412 0 -6.8018145398816293e-06
GC_9_413 b_9 NI_9 NS_413 0 4.1386917219501204e-05
GC_9_414 b_9 NI_9 NS_414 0 -4.5503052693097296e-05
GC_9_415 b_9 NI_9 NS_415 0 -3.7154907226333802e-06
GC_9_416 b_9 NI_9 NS_416 0 -4.9683592176823018e-05
GC_9_417 b_9 NI_9 NS_417 0 -1.6767613467668368e-05
GC_9_418 b_9 NI_9 NS_418 0 -6.4755703468880777e-06
GC_9_419 b_9 NI_9 NS_419 0 6.1541202250942811e-02
GC_9_420 b_9 NI_9 NS_420 0 9.5437186245519014e-04
GC_9_421 b_9 NI_9 NS_421 0 -2.6950858120779055e-02
GC_9_422 b_9 NI_9 NS_422 0 -1.2663222532447806e-02
GC_9_423 b_9 NI_9 NS_423 0 4.7137588335846185e-04
GC_9_424 b_9 NI_9 NS_424 0 1.3870783261366000e-04
GC_9_425 b_9 NI_9 NS_425 0 -4.6727010236436558e-05
GC_9_426 b_9 NI_9 NS_426 0 5.6056417463444103e-05
GC_9_427 b_9 NI_9 NS_427 0 -2.4925378287592326e-02
GC_9_428 b_9 NI_9 NS_428 0 -4.3043023868461011e-02
GC_9_429 b_9 NI_9 NS_429 0 1.5386758560291591e-05
GC_9_430 b_9 NI_9 NS_430 0 8.4355514080787218e-05
GC_9_431 b_9 NI_9 NS_431 0 9.2900882340972261e-03
GC_9_432 b_9 NI_9 NS_432 0 -9.2114384340989675e-04
GC_9_433 b_9 NI_9 NS_433 0 -5.7921462395721772e-05
GC_9_434 b_9 NI_9 NS_434 0 1.7622754724637924e-05
GC_9_435 b_9 NI_9 NS_435 0 1.6763970859317871e-06
GC_9_436 b_9 NI_9 NS_436 0 7.8001716865188373e-05
GC_9_437 b_9 NI_9 NS_437 0 -1.2523407726074438e-04
GC_9_438 b_9 NI_9 NS_438 0 -5.0911600599733481e-05
GC_9_439 b_9 NI_9 NS_439 0 -2.6961110551043744e-05
GC_9_440 b_9 NI_9 NS_440 0 -2.7879677141066555e-05
GC_9_441 b_9 NI_9 NS_441 0 -7.0543733042151046e-03
GC_9_442 b_9 NI_9 NS_442 0 3.8062549984276156e-03
GC_9_443 b_9 NI_9 NS_443 0 -7.9301365822698975e-05
GC_9_444 b_9 NI_9 NS_444 0 -3.1437330186147983e-04
GC_9_445 b_9 NI_9 NS_445 0 6.5690676114676895e-04
GC_9_446 b_9 NI_9 NS_446 0 3.8222619464051941e-04
GC_9_447 b_9 NI_9 NS_447 0 2.4397648307596814e-04
GC_9_448 b_9 NI_9 NS_448 0 -1.9371650450460647e-04
GC_9_449 b_9 NI_9 NS_449 0 2.0415190854114966e-05
GC_9_450 b_9 NI_9 NS_450 0 4.4957149995675729e-06
GC_9_451 b_9 NI_9 NS_451 0 4.9454484405663989e-05
GC_9_452 b_9 NI_9 NS_452 0 -9.7842609570475814e-06
GC_9_453 b_9 NI_9 NS_453 0 9.4871109340513576e-06
GC_9_454 b_9 NI_9 NS_454 0 -3.3875678798557717e-05
GC_9_455 b_9 NI_9 NS_455 0 -2.5459732210032395e-06
GC_9_456 b_9 NI_9 NS_456 0 -1.1194190447181381e-05
GD_9_1 b_9 NI_9 NA_1 0 -6.0496872185284139e-03
GD_9_2 b_9 NI_9 NA_2 0 5.6987302099214820e-03
GD_9_3 b_9 NI_9 NA_3 0 -5.1206598920046174e-03
GD_9_4 b_9 NI_9 NA_4 0 -1.8005639314467015e-03
GD_9_5 b_9 NI_9 NA_5 0 -7.3345395710348186e-03
GD_9_6 b_9 NI_9 NA_6 0 -7.2428412570775275e-03
GD_9_7 b_9 NI_9 NA_7 0 7.1529226489252104e-03
GD_9_8 b_9 NI_9 NA_8 0 9.2416185279420304e-03
GD_9_9 b_9 NI_9 NA_9 0 -5.7718379124423069e-02
GD_9_10 b_9 NI_9 NA_10 0 -3.7437997018895212e-02
GD_9_11 b_9 NI_9 NA_11 0 -1.9098073043337330e-02
GD_9_12 b_9 NI_9 NA_12 0 -1.0314169785713761e-02
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 9.4379903484938764e-03
GC_10_2 b_10 NI_10 NS_2 0 7.6168694393267478e-04
GC_10_3 b_10 NI_10 NS_3 0 -7.2022367026068701e-03
GC_10_4 b_10 NI_10 NS_4 0 9.2347499530668947e-04
GC_10_5 b_10 NI_10 NS_5 0 8.7782947869176426e-05
GC_10_6 b_10 NI_10 NS_6 0 -1.4229333300813508e-04
GC_10_7 b_10 NI_10 NS_7 0 6.1952230574390980e-05
GC_10_8 b_10 NI_10 NS_8 0 -4.5140297071354825e-05
GC_10_9 b_10 NI_10 NS_9 0 -1.0155001352133064e-03
GC_10_10 b_10 NI_10 NS_10 0 5.0973698583507889e-03
GC_10_11 b_10 NI_10 NS_11 0 2.2250675801794268e-05
GC_10_12 b_10 NI_10 NS_12 0 -3.3073358398619051e-05
GC_10_13 b_10 NI_10 NS_13 0 2.4284135883846526e-03
GC_10_14 b_10 NI_10 NS_14 0 2.4954487484093110e-03
GC_10_15 b_10 NI_10 NS_15 0 -1.1169595720511763e-05
GC_10_16 b_10 NI_10 NS_16 0 2.0638223923911895e-05
GC_10_17 b_10 NI_10 NS_17 0 -2.9919615079133713e-05
GC_10_18 b_10 NI_10 NS_18 0 3.3750456097066169e-05
GC_10_19 b_10 NI_10 NS_19 0 6.9109567876441528e-05
GC_10_20 b_10 NI_10 NS_20 0 -8.2387412109726782e-06
GC_10_21 b_10 NI_10 NS_21 0 3.7904532781263533e-05
GC_10_22 b_10 NI_10 NS_22 0 3.0649349528501178e-05
GC_10_23 b_10 NI_10 NS_23 0 -5.5284349563609143e-04
GC_10_24 b_10 NI_10 NS_24 0 6.0960219288546020e-04
GC_10_25 b_10 NI_10 NS_25 0 7.5290367564529695e-05
GC_10_26 b_10 NI_10 NS_26 0 -5.9360258726339214e-04
GC_10_27 b_10 NI_10 NS_27 0 -1.1403398323497179e-05
GC_10_28 b_10 NI_10 NS_28 0 -3.1205388655161989e-04
GC_10_29 b_10 NI_10 NS_29 0 -1.4002843941390410e-04
GC_10_30 b_10 NI_10 NS_30 0 1.5161295240105689e-04
GC_10_31 b_10 NI_10 NS_31 0 -1.5366726402107859e-05
GC_10_32 b_10 NI_10 NS_32 0 3.9513789107584104e-06
GC_10_33 b_10 NI_10 NS_33 0 -1.2901270150809404e-05
GC_10_34 b_10 NI_10 NS_34 0 5.9710716822454871e-05
GC_10_35 b_10 NI_10 NS_35 0 1.0584336325094494e-05
GC_10_36 b_10 NI_10 NS_36 0 -1.4312742408808855e-05
GC_10_37 b_10 NI_10 NS_37 0 -1.3643712998194805e-05
GC_10_38 b_10 NI_10 NS_38 0 9.2996541632320967e-07
GC_10_39 b_10 NI_10 NS_39 0 7.7921969089085738e-03
GC_10_40 b_10 NI_10 NS_40 0 -8.1321745016285391e-04
GC_10_41 b_10 NI_10 NS_41 0 -7.5104897507362340e-03
GC_10_42 b_10 NI_10 NS_42 0 -4.0556804053710699e-03
GC_10_43 b_10 NI_10 NS_43 0 1.0926551063463790e-04
GC_10_44 b_10 NI_10 NS_44 0 2.0190808178968203e-04
GC_10_45 b_10 NI_10 NS_45 0 3.4348656593414286e-05
GC_10_46 b_10 NI_10 NS_46 0 9.5203085717516611e-05
GC_10_47 b_10 NI_10 NS_47 0 -2.0547264048763591e-04
GC_10_48 b_10 NI_10 NS_48 0 -6.8745847269247665e-03
GC_10_49 b_10 NI_10 NS_49 0 -2.3831848667020335e-05
GC_10_50 b_10 NI_10 NS_50 0 2.8334788256346724e-05
GC_10_51 b_10 NI_10 NS_51 0 3.9174173761262745e-03
GC_10_52 b_10 NI_10 NS_52 0 5.0602341298025058e-03
GC_10_53 b_10 NI_10 NS_53 0 5.7307072016445859e-05
GC_10_54 b_10 NI_10 NS_54 0 5.4375054285860746e-05
GC_10_55 b_10 NI_10 NS_55 0 -1.4927843388986412e-05
GC_10_56 b_10 NI_10 NS_56 0 6.5501137991632452e-05
GC_10_57 b_10 NI_10 NS_57 0 1.3431857238267234e-05
GC_10_58 b_10 NI_10 NS_58 0 1.5206213385899240e-05
GC_10_59 b_10 NI_10 NS_59 0 6.0601845909927559e-05
GC_10_60 b_10 NI_10 NS_60 0 4.6012871445150076e-05
GC_10_61 b_10 NI_10 NS_61 0 -2.2717875896521322e-03
GC_10_62 b_10 NI_10 NS_62 0 3.9767776404575243e-04
GC_10_63 b_10 NI_10 NS_63 0 3.8241501678092310e-04
GC_10_64 b_10 NI_10 NS_64 0 -6.7399758626471415e-04
GC_10_65 b_10 NI_10 NS_65 0 1.6608438916437444e-04
GC_10_66 b_10 NI_10 NS_66 0 -3.6132682948697821e-04
GC_10_67 b_10 NI_10 NS_67 0 -1.2799367628360596e-04
GC_10_68 b_10 NI_10 NS_68 0 9.4649733690508068e-05
GC_10_69 b_10 NI_10 NS_69 0 -2.1317674709613808e-05
GC_10_70 b_10 NI_10 NS_70 0 -7.8121854076295340e-06
GC_10_71 b_10 NI_10 NS_71 0 -4.4546552899888745e-05
GC_10_72 b_10 NI_10 NS_72 0 1.0524004674583242e-05
GC_10_73 b_10 NI_10 NS_73 0 3.0892384518069330e-05
GC_10_74 b_10 NI_10 NS_74 0 -2.8808519947237921e-06
GC_10_75 b_10 NI_10 NS_75 0 7.5764294526146051e-06
GC_10_76 b_10 NI_10 NS_76 0 1.6179605440116628e-06
GC_10_77 b_10 NI_10 NS_77 0 1.3481314461212876e-02
GC_10_78 b_10 NI_10 NS_78 0 1.1270839926274801e-03
GC_10_79 b_10 NI_10 NS_79 0 -9.5721183869524676e-03
GC_10_80 b_10 NI_10 NS_80 0 1.2007839633793095e-03
GC_10_81 b_10 NI_10 NS_81 0 2.3592254125013131e-04
GC_10_82 b_10 NI_10 NS_82 0 -2.1851889153327498e-04
GC_10_83 b_10 NI_10 NS_83 0 6.7386324266736274e-05
GC_10_84 b_10 NI_10 NS_84 0 -6.1486903451215424e-05
GC_10_85 b_10 NI_10 NS_85 0 -2.0750373229901234e-03
GC_10_86 b_10 NI_10 NS_86 0 5.6028578657436757e-03
GC_10_87 b_10 NI_10 NS_87 0 2.3440936349190155e-05
GC_10_88 b_10 NI_10 NS_88 0 -3.3427826397956492e-05
GC_10_89 b_10 NI_10 NS_89 0 3.6181762005694012e-03
GC_10_90 b_10 NI_10 NS_90 0 4.4649809987568493e-03
GC_10_91 b_10 NI_10 NS_91 0 -1.7556471519911999e-05
GC_10_92 b_10 NI_10 NS_92 0 -9.8179535378387229e-06
GC_10_93 b_10 NI_10 NS_93 0 -2.2334745323429076e-05
GC_10_94 b_10 NI_10 NS_94 0 4.2470999405369936e-05
GC_10_95 b_10 NI_10 NS_95 0 7.6370032637165637e-05
GC_10_96 b_10 NI_10 NS_96 0 -2.4913480113564247e-06
GC_10_97 b_10 NI_10 NS_97 0 3.5651919786888616e-05
GC_10_98 b_10 NI_10 NS_98 0 2.3031348336486263e-05
GC_10_99 b_10 NI_10 NS_99 0 -1.3671874192019032e-03
GC_10_100 b_10 NI_10 NS_100 0 -7.7234369625365108e-04
GC_10_101 b_10 NI_10 NS_101 0 4.7757957389924680e-05
GC_10_102 b_10 NI_10 NS_102 0 -4.3130279378351857e-04
GC_10_103 b_10 NI_10 NS_103 0 1.3790379773758612e-04
GC_10_104 b_10 NI_10 NS_104 0 2.0909340420989686e-05
GC_10_105 b_10 NI_10 NS_105 0 2.5085832592425018e-05
GC_10_106 b_10 NI_10 NS_106 0 4.9385458652437667e-05
GC_10_107 b_10 NI_10 NS_107 0 -6.1958848193347164e-06
GC_10_108 b_10 NI_10 NS_108 0 -3.0096494140338460e-06
GC_10_109 b_10 NI_10 NS_109 0 -1.0205732802798304e-05
GC_10_110 b_10 NI_10 NS_110 0 2.1584069982005138e-05
GC_10_111 b_10 NI_10 NS_111 0 2.8935838892203092e-05
GC_10_112 b_10 NI_10 NS_112 0 3.0488833967802398e-06
GC_10_113 b_10 NI_10 NS_113 0 4.7198941896832179e-06
GC_10_114 b_10 NI_10 NS_114 0 -9.0580250550141212e-06
GC_10_115 b_10 NI_10 NS_115 0 9.8335405310515933e-03
GC_10_116 b_10 NI_10 NS_116 0 -1.1184866204153505e-03
GC_10_117 b_10 NI_10 NS_117 0 -8.9641725997885897e-03
GC_10_118 b_10 NI_10 NS_118 0 -2.7022998601686585e-03
GC_10_119 b_10 NI_10 NS_119 0 1.4215151153032404e-04
GC_10_120 b_10 NI_10 NS_120 0 1.7288164290281085e-04
GC_10_121 b_10 NI_10 NS_121 0 4.9934378841612073e-05
GC_10_122 b_10 NI_10 NS_122 0 9.8026904304897078e-05
GC_10_123 b_10 NI_10 NS_123 0 8.0739659815351320e-04
GC_10_124 b_10 NI_10 NS_124 0 -6.7270701221655424e-03
GC_10_125 b_10 NI_10 NS_125 0 -2.5664887807669964e-05
GC_10_126 b_10 NI_10 NS_126 0 2.8406616156355259e-05
GC_10_127 b_10 NI_10 NS_127 0 4.4520168973041369e-03
GC_10_128 b_10 NI_10 NS_128 0 6.7708519599191932e-03
GC_10_129 b_10 NI_10 NS_129 0 5.8580162283204681e-05
GC_10_130 b_10 NI_10 NS_130 0 2.6941983612918479e-05
GC_10_131 b_10 NI_10 NS_131 0 -1.7983212555279232e-05
GC_10_132 b_10 NI_10 NS_132 0 5.9731475074863496e-05
GC_10_133 b_10 NI_10 NS_133 0 4.6612495938382389e-05
GC_10_134 b_10 NI_10 NS_134 0 2.1553275315607320e-05
GC_10_135 b_10 NI_10 NS_135 0 6.5181206767107625e-05
GC_10_136 b_10 NI_10 NS_136 0 4.0000004012528492e-05
GC_10_137 b_10 NI_10 NS_137 0 -2.5410209426888850e-03
GC_10_138 b_10 NI_10 NS_138 0 -8.8530435054689116e-04
GC_10_139 b_10 NI_10 NS_139 0 3.9370779001252906e-04
GC_10_140 b_10 NI_10 NS_140 0 -5.3416742642412528e-04
GC_10_141 b_10 NI_10 NS_141 0 3.0598776752266632e-04
GC_10_142 b_10 NI_10 NS_142 0 -6.9971218195091726e-05
GC_10_143 b_10 NI_10 NS_143 0 -1.5587634291218238e-05
GC_10_144 b_10 NI_10 NS_144 0 1.8616194975057651e-05
GC_10_145 b_10 NI_10 NS_145 0 -1.0442446808739100e-05
GC_10_146 b_10 NI_10 NS_146 0 -8.9639404652769531e-06
GC_10_147 b_10 NI_10 NS_147 0 -2.0186797858370707e-05
GC_10_148 b_10 NI_10 NS_148 0 5.7592249150796708e-06
GC_10_149 b_10 NI_10 NS_149 0 2.4797665937652780e-05
GC_10_150 b_10 NI_10 NS_150 0 -3.3063946650519344e-06
GC_10_151 b_10 NI_10 NS_151 0 4.5254632177187744e-06
GC_10_152 b_10 NI_10 NS_152 0 6.8548261321419156e-06
GC_10_153 b_10 NI_10 NS_153 0 1.0944170740129827e-02
GC_10_154 b_10 NI_10 NS_154 0 1.3496456981999070e-03
GC_10_155 b_10 NI_10 NS_155 0 -1.2355658574303676e-02
GC_10_156 b_10 NI_10 NS_156 0 2.0266962996839662e-03
GC_10_157 b_10 NI_10 NS_157 0 3.0286033960542241e-04
GC_10_158 b_10 NI_10 NS_158 0 -5.5942401945680367e-05
GC_10_159 b_10 NI_10 NS_159 0 7.4864323896525560e-05
GC_10_160 b_10 NI_10 NS_160 0 -6.3940496968093672e-05
GC_10_161 b_10 NI_10 NS_161 0 -4.2789482767755741e-03
GC_10_162 b_10 NI_10 NS_162 0 -5.6119776758759878e-04
GC_10_163 b_10 NI_10 NS_163 0 1.3780875058243109e-05
GC_10_164 b_10 NI_10 NS_164 0 2.2699881228296596e-06
GC_10_165 b_10 NI_10 NS_165 0 1.1409463318914456e-02
GC_10_166 b_10 NI_10 NS_166 0 1.6019415398492729e-03
GC_10_167 b_10 NI_10 NS_167 0 -2.1548363144454436e-05
GC_10_168 b_10 NI_10 NS_168 0 -3.1646781906316395e-05
GC_10_169 b_10 NI_10 NS_169 0 -1.7189195469216145e-05
GC_10_170 b_10 NI_10 NS_170 0 5.5921558996780222e-05
GC_10_171 b_10 NI_10 NS_171 0 1.1204098210629585e-06
GC_10_172 b_10 NI_10 NS_172 0 -1.8508564807027557e-05
GC_10_173 b_10 NI_10 NS_173 0 -7.9308527843013070e-06
GC_10_174 b_10 NI_10 NS_174 0 -5.7425691802748489e-07
GC_10_175 b_10 NI_10 NS_175 0 -3.7107580507947458e-03
GC_10_176 b_10 NI_10 NS_176 0 1.3307979249318289e-03
GC_10_177 b_10 NI_10 NS_177 0 5.5028435902109891e-06
GC_10_178 b_10 NI_10 NS_178 0 -6.2287303750332610e-04
GC_10_179 b_10 NI_10 NS_179 0 3.2648864059855353e-04
GC_10_180 b_10 NI_10 NS_180 0 -1.7113665473680528e-04
GC_10_181 b_10 NI_10 NS_181 0 1.8901080766294166e-05
GC_10_182 b_10 NI_10 NS_182 0 -8.2982848668053146e-06
GC_10_183 b_10 NI_10 NS_183 0 8.1963119548269902e-06
GC_10_184 b_10 NI_10 NS_184 0 -1.1917951488226548e-05
GC_10_185 b_10 NI_10 NS_185 0 -2.2657084303827808e-05
GC_10_186 b_10 NI_10 NS_186 0 -1.3419710363475165e-05
GC_10_187 b_10 NI_10 NS_187 0 6.4454940719837616e-05
GC_10_188 b_10 NI_10 NS_188 0 -5.1900177604833111e-05
GC_10_189 b_10 NI_10 NS_189 0 -1.9762567331051415e-05
GC_10_190 b_10 NI_10 NS_190 0 -4.2241836157926336e-05
GC_10_191 b_10 NI_10 NS_191 0 -8.9009039068153276e-03
GC_10_192 b_10 NI_10 NS_192 0 -1.3474891042239588e-03
GC_10_193 b_10 NI_10 NS_193 0 -2.0239400735629757e-03
GC_10_194 b_10 NI_10 NS_194 0 5.2287519009650311e-03
GC_10_195 b_10 NI_10 NS_195 0 -1.3293117749463266e-04
GC_10_196 b_10 NI_10 NS_196 0 2.0824785929209451e-04
GC_10_197 b_10 NI_10 NS_197 0 1.3275692557363985e-05
GC_10_198 b_10 NI_10 NS_198 0 3.3543471568744571e-05
GC_10_199 b_10 NI_10 NS_199 0 5.4760933835810858e-03
GC_10_200 b_10 NI_10 NS_200 0 2.7344827144192689e-03
GC_10_201 b_10 NI_10 NS_201 0 -1.4215150657641639e-05
GC_10_202 b_10 NI_10 NS_202 0 -1.6307927714006435e-06
GC_10_203 b_10 NI_10 NS_203 0 1.0116194408685657e-02
GC_10_204 b_10 NI_10 NS_204 0 -2.6917852764692172e-03
GC_10_205 b_10 NI_10 NS_205 0 1.3808286754993898e-05
GC_10_206 b_10 NI_10 NS_206 0 3.4374378633866931e-06
GC_10_207 b_10 NI_10 NS_207 0 -1.3984584939155149e-05
GC_10_208 b_10 NI_10 NS_208 0 3.4101781242089735e-05
GC_10_209 b_10 NI_10 NS_209 0 -1.2075990167911117e-05
GC_10_210 b_10 NI_10 NS_210 0 1.4372460949201602e-06
GC_10_211 b_10 NI_10 NS_211 0 9.1382436911932601e-06
GC_10_212 b_10 NI_10 NS_212 0 -6.7027722001587201e-08
GC_10_213 b_10 NI_10 NS_213 0 -3.3305916708277010e-03
GC_10_214 b_10 NI_10 NS_214 0 1.8529063419789938e-03
GC_10_215 b_10 NI_10 NS_215 0 4.9308852511701567e-06
GC_10_216 b_10 NI_10 NS_216 0 -4.6466034185078643e-04
GC_10_217 b_10 NI_10 NS_217 0 2.6858897064058256e-04
GC_10_218 b_10 NI_10 NS_218 0 -1.0414960723172922e-04
GC_10_219 b_10 NI_10 NS_219 0 4.8024189839655124e-05
GC_10_220 b_10 NI_10 NS_220 0 2.2856870451952514e-05
GC_10_221 b_10 NI_10 NS_221 0 7.0158643934500438e-06
GC_10_222 b_10 NI_10 NS_222 0 8.6174287116913664e-06
GC_10_223 b_10 NI_10 NS_223 0 1.8426341764534190e-05
GC_10_224 b_10 NI_10 NS_224 0 -1.1066626827999448e-06
GC_10_225 b_10 NI_10 NS_225 0 7.2414717976304862e-05
GC_10_226 b_10 NI_10 NS_226 0 -2.6825032757170435e-05
GC_10_227 b_10 NI_10 NS_227 0 9.9520967550548455e-07
GC_10_228 b_10 NI_10 NS_228 0 -4.1646903874745335e-05
GC_10_229 b_10 NI_10 NS_229 0 -2.4112243421142803e-02
GC_10_230 b_10 NI_10 NS_230 0 1.4730135136552499e-03
GC_10_231 b_10 NI_10 NS_231 0 1.4876220840276143e-02
GC_10_232 b_10 NI_10 NS_232 0 -2.3953699740304562e-03
GC_10_233 b_10 NI_10 NS_233 0 2.1084605692689131e-04
GC_10_234 b_10 NI_10 NS_234 0 2.1031897943993997e-05
GC_10_235 b_10 NI_10 NS_235 0 -2.3639261700425282e-05
GC_10_236 b_10 NI_10 NS_236 0 -5.1595780335728009e-06
GC_10_237 b_10 NI_10 NS_237 0 -8.0051480608333593e-03
GC_10_238 b_10 NI_10 NS_238 0 -1.2245231716655369e-02
GC_10_239 b_10 NI_10 NS_239 0 2.1887848468152405e-05
GC_10_240 b_10 NI_10 NS_240 0 6.3133388693476109e-06
GC_10_241 b_10 NI_10 NS_241 0 6.1155468229604675e-03
GC_10_242 b_10 NI_10 NS_242 0 -1.0677698665093514e-02
GC_10_243 b_10 NI_10 NS_243 0 -1.7101627140765224e-05
GC_10_244 b_10 NI_10 NS_244 0 -1.4847722855170524e-05
GC_10_245 b_10 NI_10 NS_245 0 -1.1403084944160053e-05
GC_10_246 b_10 NI_10 NS_246 0 4.8083516853010681e-05
GC_10_247 b_10 NI_10 NS_247 0 -1.8697713599127601e-05
GC_10_248 b_10 NI_10 NS_248 0 -2.1123609439320645e-05
GC_10_249 b_10 NI_10 NS_249 0 -6.0556988818997383e-07
GC_10_250 b_10 NI_10 NS_250 0 -6.8985572094447156e-06
GC_10_251 b_10 NI_10 NS_251 0 -4.2965421981393456e-03
GC_10_252 b_10 NI_10 NS_252 0 2.0119180889228042e-04
GC_10_253 b_10 NI_10 NS_253 0 -1.1512098237070457e-04
GC_10_254 b_10 NI_10 NS_254 0 -3.8953460584192440e-04
GC_10_255 b_10 NI_10 NS_255 0 4.4756393971484061e-04
GC_10_256 b_10 NI_10 NS_256 0 1.3357744451760880e-04
GC_10_257 b_10 NI_10 NS_257 0 1.7124256750736117e-04
GC_10_258 b_10 NI_10 NS_258 0 -1.2652129182092638e-04
GC_10_259 b_10 NI_10 NS_259 0 -1.6678129363065428e-05
GC_10_260 b_10 NI_10 NS_260 0 -8.2963750411584869e-06
GC_10_261 b_10 NI_10 NS_261 0 1.1437716997777356e-06
GC_10_262 b_10 NI_10 NS_262 0 6.7674329462041710e-06
GC_10_263 b_10 NI_10 NS_263 0 -1.1895340877261689e-06
GC_10_264 b_10 NI_10 NS_264 0 1.3998226370687503e-05
GC_10_265 b_10 NI_10 NS_265 0 3.0390325374904444e-05
GC_10_266 b_10 NI_10 NS_266 0 2.0362526871568657e-05
GC_10_267 b_10 NI_10 NS_267 0 -1.5982046220309663e-02
GC_10_268 b_10 NI_10 NS_268 0 -1.5163490837181044e-03
GC_10_269 b_10 NI_10 NS_269 0 1.0314462558101882e-02
GC_10_270 b_10 NI_10 NS_270 0 2.2248713364982950e-02
GC_10_271 b_10 NI_10 NS_271 0 -2.6378094819725869e-04
GC_10_272 b_10 NI_10 NS_272 0 4.3028149633284063e-04
GC_10_273 b_10 NI_10 NS_273 0 -1.3837196025189993e-05
GC_10_274 b_10 NI_10 NS_274 0 3.8170119986278707e-05
GC_10_275 b_10 NI_10 NS_275 0 6.8934481583097429e-03
GC_10_276 b_10 NI_10 NS_276 0 9.4223067075043208e-03
GC_10_277 b_10 NI_10 NS_277 0 -2.2150683662866841e-05
GC_10_278 b_10 NI_10 NS_278 0 -9.3857991455956528e-06
GC_10_279 b_10 NI_10 NS_279 0 1.2955541139946869e-02
GC_10_280 b_10 NI_10 NS_280 0 -1.4354532997746626e-02
GC_10_281 b_10 NI_10 NS_281 0 4.9113415316699182e-06
GC_10_282 b_10 NI_10 NS_282 0 1.2586786758519486e-05
GC_10_283 b_10 NI_10 NS_283 0 -1.7379887332537018e-05
GC_10_284 b_10 NI_10 NS_284 0 3.1536670455491510e-05
GC_10_285 b_10 NI_10 NS_285 0 -7.0169962877865841e-06
GC_10_286 b_10 NI_10 NS_286 0 -1.4031457987323992e-05
GC_10_287 b_10 NI_10 NS_287 0 1.7502657514875347e-05
GC_10_288 b_10 NI_10 NS_288 0 -3.1217753180603299e-06
GC_10_289 b_10 NI_10 NS_289 0 -4.3699462740916005e-03
GC_10_290 b_10 NI_10 NS_290 0 5.4977835055190663e-04
GC_10_291 b_10 NI_10 NS_291 0 -1.7725634798774787e-06
GC_10_292 b_10 NI_10 NS_292 0 -3.8107774520761709e-04
GC_10_293 b_10 NI_10 NS_293 0 4.0701999869383141e-04
GC_10_294 b_10 NI_10 NS_294 0 1.6191437326907102e-04
GC_10_295 b_10 NI_10 NS_295 0 1.7799000932638897e-04
GC_10_296 b_10 NI_10 NS_296 0 -5.8433726125533116e-05
GC_10_297 b_10 NI_10 NS_297 0 -8.3323528612178273e-06
GC_10_298 b_10 NI_10 NS_298 0 -1.8244213094078600e-05
GC_10_299 b_10 NI_10 NS_299 0 4.3798197544120547e-06
GC_10_300 b_10 NI_10 NS_300 0 -3.4529297897865611e-06
GC_10_301 b_10 NI_10 NS_301 0 4.7242518180958716e-06
GC_10_302 b_10 NI_10 NS_302 0 2.2791047102450693e-06
GC_10_303 b_10 NI_10 NS_303 0 9.3955146002553513e-06
GC_10_304 b_10 NI_10 NS_304 0 2.8024907074551126e-05
GC_10_305 b_10 NI_10 NS_305 0 3.8120006653767774e-02
GC_10_306 b_10 NI_10 NS_306 0 2.2971138896204363e-03
GC_10_307 b_10 NI_10 NS_307 0 1.2353267202868459e-02
GC_10_308 b_10 NI_10 NS_308 0 -1.9939162004279736e-02
GC_10_309 b_10 NI_10 NS_309 0 1.5278723613196248e-03
GC_10_310 b_10 NI_10 NS_310 0 3.5029179274735491e-05
GC_10_311 b_10 NI_10 NS_311 0 4.1319094132670505e-05
GC_10_312 b_10 NI_10 NS_312 0 -7.0118540408861886e-06
GC_10_313 b_10 NI_10 NS_313 0 2.3295403345166835e-02
GC_10_314 b_10 NI_10 NS_314 0 1.8084948937525020e-03
GC_10_315 b_10 NI_10 NS_315 0 4.3610870537124921e-05
GC_10_316 b_10 NI_10 NS_316 0 9.1844256953310731e-05
GC_10_317 b_10 NI_10 NS_317 0 -4.3234548618815614e-02
GC_10_318 b_10 NI_10 NS_318 0 4.1033638144166655e-02
GC_10_319 b_10 NI_10 NS_319 0 -2.6648980577572929e-06
GC_10_320 b_10 NI_10 NS_320 0 -5.2314745046151768e-06
GC_10_321 b_10 NI_10 NS_321 0 -1.6872682655160079e-05
GC_10_322 b_10 NI_10 NS_322 0 7.9286109576271464e-05
GC_10_323 b_10 NI_10 NS_323 0 -8.9759691428086991e-05
GC_10_324 b_10 NI_10 NS_324 0 -2.6595141804483044e-05
GC_10_325 b_10 NI_10 NS_325 0 -3.2770221591688805e-05
GC_10_326 b_10 NI_10 NS_326 0 -2.7262748503146014e-05
GC_10_327 b_10 NI_10 NS_327 0 -4.6019315417753521e-03
GC_10_328 b_10 NI_10 NS_328 0 -1.7321018277720803e-03
GC_10_329 b_10 NI_10 NS_329 0 1.1156783938872234e-04
GC_10_330 b_10 NI_10 NS_330 0 -1.9780919370238924e-04
GC_10_331 b_10 NI_10 NS_331 0 3.5639726874750423e-04
GC_10_332 b_10 NI_10 NS_332 0 3.7497160376676476e-04
GC_10_333 b_10 NI_10 NS_333 0 1.7011003156755376e-04
GC_10_334 b_10 NI_10 NS_334 0 -3.0865486276652642e-05
GC_10_335 b_10 NI_10 NS_335 0 2.7422085587741399e-05
GC_10_336 b_10 NI_10 NS_336 0 3.4724031384383386e-07
GC_10_337 b_10 NI_10 NS_337 0 1.9366190458186600e-05
GC_10_338 b_10 NI_10 NS_338 0 1.6928785234428384e-05
GC_10_339 b_10 NI_10 NS_339 0 1.2644096038730807e-05
GC_10_340 b_10 NI_10 NS_340 0 4.9589356588088941e-05
GC_10_341 b_10 NI_10 NS_341 0 2.9057018593954362e-05
GC_10_342 b_10 NI_10 NS_342 0 -9.9994199386400228e-06
GC_10_343 b_10 NI_10 NS_343 0 4.8618403262691012e-02
GC_10_344 b_10 NI_10 NS_344 0 -1.7609209191877999e-03
GC_10_345 b_10 NI_10 NS_345 0 4.6135578503255628e-02
GC_10_346 b_10 NI_10 NS_346 0 -5.4327626944676743e-02
GC_10_347 b_10 NI_10 NS_347 0 -4.5044019406316184e-04
GC_10_348 b_10 NI_10 NS_348 0 3.7491840703232388e-04
GC_10_349 b_10 NI_10 NS_349 0 -1.1571225458418209e-05
GC_10_350 b_10 NI_10 NS_350 0 1.1061801350388812e-04
GC_10_351 b_10 NI_10 NS_351 0 -6.6945599549177023e-03
GC_10_352 b_10 NI_10 NS_352 0 1.7899868822433419e-02
GC_10_353 b_10 NI_10 NS_353 0 -2.5611566228420524e-05
GC_10_354 b_10 NI_10 NS_354 0 -8.1050342601411940e-05
GC_10_355 b_10 NI_10 NS_355 0 -3.0042620181318182e-02
GC_10_356 b_10 NI_10 NS_356 0 7.6797497113262414e-03
GC_10_357 b_10 NI_10 NS_357 0 -1.8546140584491211e-05
GC_10_358 b_10 NI_10 NS_358 0 2.7916012970268470e-05
GC_10_359 b_10 NI_10 NS_359 0 -4.4632211923040384e-05
GC_10_360 b_10 NI_10 NS_360 0 7.5621735727828215e-05
GC_10_361 b_10 NI_10 NS_361 0 -6.2162162490957164e-05
GC_10_362 b_10 NI_10 NS_362 0 -1.3658335187300115e-05
GC_10_363 b_10 NI_10 NS_363 0 -2.7426795827615103e-05
GC_10_364 b_10 NI_10 NS_364 0 -3.3539239217590905e-05
GC_10_365 b_10 NI_10 NS_365 0 -3.5293194866156566e-03
GC_10_366 b_10 NI_10 NS_366 0 2.2912129794367777e-03
GC_10_367 b_10 NI_10 NS_367 0 1.4935355430018606e-04
GC_10_368 b_10 NI_10 NS_368 0 -3.5226812611956318e-04
GC_10_369 b_10 NI_10 NS_369 0 3.1764363581102887e-04
GC_10_370 b_10 NI_10 NS_370 0 6.2974560019346879e-05
GC_10_371 b_10 NI_10 NS_371 0 1.2930670251606603e-04
GC_10_372 b_10 NI_10 NS_372 0 -5.2313805772889139e-05
GC_10_373 b_10 NI_10 NS_373 0 1.2043747627155808e-05
GC_10_374 b_10 NI_10 NS_374 0 9.0755021418639666e-06
GC_10_375 b_10 NI_10 NS_375 0 7.1403598975567657e-06
GC_10_376 b_10 NI_10 NS_376 0 -2.1102327897015260e-05
GC_10_377 b_10 NI_10 NS_377 0 -4.2651012133835756e-06
GC_10_378 b_10 NI_10 NS_378 0 -4.2365021629586419e-05
GC_10_379 b_10 NI_10 NS_379 0 -2.5740792854628425e-05
GC_10_380 b_10 NI_10 NS_380 0 -3.3902956563772624e-06
GC_10_381 b_10 NI_10 NS_381 0 5.7049805530080412e-02
GC_10_382 b_10 NI_10 NS_382 0 9.2459103948133150e-04
GC_10_383 b_10 NI_10 NS_383 0 -3.4891474033354131e-02
GC_10_384 b_10 NI_10 NS_384 0 -1.4433131859337230e-02
GC_10_385 b_10 NI_10 NS_385 0 -6.2029530685235200e-04
GC_10_386 b_10 NI_10 NS_386 0 2.6308391115533369e-04
GC_10_387 b_10 NI_10 NS_387 0 -1.3720883005254440e-04
GC_10_388 b_10 NI_10 NS_388 0 1.2168603009896299e-04
GC_10_389 b_10 NI_10 NS_389 0 -2.4467120521553646e-02
GC_10_390 b_10 NI_10 NS_390 0 -4.3613909873158961e-02
GC_10_391 b_10 NI_10 NS_391 0 1.5965592363683892e-05
GC_10_392 b_10 NI_10 NS_392 0 8.3164444572729940e-05
GC_10_393 b_10 NI_10 NS_393 0 1.3305732156688716e-02
GC_10_394 b_10 NI_10 NS_394 0 -2.1369016957191938e-04
GC_10_395 b_10 NI_10 NS_395 0 -2.5929284441616845e-05
GC_10_396 b_10 NI_10 NS_396 0 5.0407167693001589e-05
GC_10_397 b_10 NI_10 NS_397 0 -5.8767281978336969e-06
GC_10_398 b_10 NI_10 NS_398 0 3.9648046323389993e-05
GC_10_399 b_10 NI_10 NS_399 0 -1.1890108408902688e-04
GC_10_400 b_10 NI_10 NS_400 0 -2.7602376799180241e-05
GC_10_401 b_10 NI_10 NS_401 0 -2.4374109266254137e-05
GC_10_402 b_10 NI_10 NS_402 0 -2.5382640210774570e-05
GC_10_403 b_10 NI_10 NS_403 0 -5.4409749353955088e-03
GC_10_404 b_10 NI_10 NS_404 0 4.1782945557269245e-03
GC_10_405 b_10 NI_10 NS_405 0 -1.5878093538416522e-04
GC_10_406 b_10 NI_10 NS_406 0 -2.5094067076768186e-04
GC_10_407 b_10 NI_10 NS_407 0 6.2372590304789221e-04
GC_10_408 b_10 NI_10 NS_408 0 2.1594250633765553e-04
GC_10_409 b_10 NI_10 NS_409 0 1.8537009019696868e-04
GC_10_410 b_10 NI_10 NS_410 0 -2.3875302199764947e-04
GC_10_411 b_10 NI_10 NS_411 0 3.4179840332053541e-05
GC_10_412 b_10 NI_10 NS_412 0 1.3039545485477453e-05
GC_10_413 b_10 NI_10 NS_413 0 3.2311118834437607e-05
GC_10_414 b_10 NI_10 NS_414 0 -3.5399657659314476e-05
GC_10_415 b_10 NI_10 NS_415 0 -7.1059500383841714e-06
GC_10_416 b_10 NI_10 NS_416 0 1.8975202538938102e-05
GC_10_417 b_10 NI_10 NS_417 0 -3.8058795023185931e-06
GC_10_418 b_10 NI_10 NS_418 0 -5.9631428859058883e-06
GC_10_419 b_10 NI_10 NS_419 0 -3.9907462552120146e-03
GC_10_420 b_10 NI_10 NS_420 0 -1.4032328031731911e-03
GC_10_421 b_10 NI_10 NS_421 0 1.2077943006268302e-03
GC_10_422 b_10 NI_10 NS_422 0 -3.5921095464235106e-03
GC_10_423 b_10 NI_10 NS_423 0 -4.1901655624453912e-04
GC_10_424 b_10 NI_10 NS_424 0 5.7189086426440931e-04
GC_10_425 b_10 NI_10 NS_425 0 -5.6536612121570353e-05
GC_10_426 b_10 NI_10 NS_426 0 1.0476005672297238e-04
GC_10_427 b_10 NI_10 NS_427 0 7.7236945158374913e-03
GC_10_428 b_10 NI_10 NS_428 0 2.3103097487258056e-02
GC_10_429 b_10 NI_10 NS_429 0 -2.6971168581682481e-05
GC_10_430 b_10 NI_10 NS_430 0 -8.4231210674609716e-05
GC_10_431 b_10 NI_10 NS_431 0 4.9533168271373206e-03
GC_10_432 b_10 NI_10 NS_432 0 -3.6202481250936515e-03
GC_10_433 b_10 NI_10 NS_433 0 -4.2869874335046379e-05
GC_10_434 b_10 NI_10 NS_434 0 5.8576309458925962e-05
GC_10_435 b_10 NI_10 NS_435 0 -2.6275634749957401e-05
GC_10_436 b_10 NI_10 NS_436 0 5.8114226528874556e-05
GC_10_437 b_10 NI_10 NS_437 0 -8.0537850511464294e-05
GC_10_438 b_10 NI_10 NS_438 0 -2.7887353272553584e-05
GC_10_439 b_10 NI_10 NS_439 0 -2.1091488772656007e-05
GC_10_440 b_10 NI_10 NS_440 0 -3.1106294827211774e-05
GC_10_441 b_10 NI_10 NS_441 0 -5.5316221982171570e-03
GC_10_442 b_10 NI_10 NS_442 0 3.7852963150724370e-03
GC_10_443 b_10 NI_10 NS_443 0 7.4445149685532303e-05
GC_10_444 b_10 NI_10 NS_444 0 -3.2468976442515839e-04
GC_10_445 b_10 NI_10 NS_445 0 5.1446924293904034e-04
GC_10_446 b_10 NI_10 NS_446 0 2.6685035426966775e-04
GC_10_447 b_10 NI_10 NS_447 0 2.4742019067437666e-04
GC_10_448 b_10 NI_10 NS_448 0 -1.4105279881308132e-04
GC_10_449 b_10 NI_10 NS_449 0 1.7317911586527770e-05
GC_10_450 b_10 NI_10 NS_450 0 3.3421662533460864e-05
GC_10_451 b_10 NI_10 NS_451 0 4.1579282264894099e-05
GC_10_452 b_10 NI_10 NS_452 0 -2.5194919010954322e-05
GC_10_453 b_10 NI_10 NS_453 0 -1.6418360978852971e-05
GC_10_454 b_10 NI_10 NS_454 0 -1.2561232004454082e-05
GC_10_455 b_10 NI_10 NS_455 0 -1.0595204124503212e-05
GC_10_456 b_10 NI_10 NS_456 0 -1.1811286991780449e-05
GD_10_1 b_10 NI_10 NA_1 0 -3.2465259657341481e-03
GD_10_2 b_10 NI_10 NA_2 0 -8.2354181119865340e-04
GD_10_3 b_10 NI_10 NA_3 0 -5.0829437010726890e-03
GD_10_4 b_10 NI_10 NA_4 0 -2.8725085569522696e-03
GD_10_5 b_10 NI_10 NA_5 0 -3.1499964760540356e-03
GD_10_6 b_10 NI_10 NA_6 0 -1.6038739131278573e-04
GD_10_7 b_10 NI_10 NA_7 0 1.1950900823398225e-02
GD_10_8 b_10 NI_10 NA_8 0 -5.7613799841656609e-03
GD_10_9 b_10 NI_10 NA_9 0 -3.7438033902145895e-02
GD_10_10 b_10 NI_10 NA_10 0 -1.2004894330214973e-01
GD_10_11 b_10 NI_10 NA_11 0 1.7503028800809936e-03
GD_10_12 b_10 NI_10 NA_12 0 1.4508872502093674e-03
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 8.5420431837792514e-03
GC_11_2 b_11 NI_11 NS_2 0 -4.9689565496506582e-04
GC_11_3 b_11 NI_11 NS_3 0 -6.6709328344836802e-03
GC_11_4 b_11 NI_11 NS_4 0 3.0245579775209476e-03
GC_11_5 b_11 NI_11 NS_5 0 4.1888015309182059e-05
GC_11_6 b_11 NI_11 NS_6 0 -2.6210771300021910e-05
GC_11_7 b_11 NI_11 NS_7 0 1.7916199006957933e-04
GC_11_8 b_11 NI_11 NS_8 0 -1.6276130920364097e-04
GC_11_9 b_11 NI_11 NS_9 0 -1.1767274335482790e-04
GC_11_10 b_11 NI_11 NS_10 0 -4.2758630039716828e-03
GC_11_11 b_11 NI_11 NS_11 0 -1.6650485302682404e-05
GC_11_12 b_11 NI_11 NS_12 0 3.6525995883256354e-05
GC_11_13 b_11 NI_11 NS_13 0 2.4608797864107430e-03
GC_11_14 b_11 NI_11 NS_14 0 7.9712518572635084e-04
GC_11_15 b_11 NI_11 NS_15 0 -4.0240806327151764e-06
GC_11_16 b_11 NI_11 NS_16 0 1.0939352581962854e-05
GC_11_17 b_11 NI_11 NS_17 0 1.0195247565800430e-05
GC_11_18 b_11 NI_11 NS_18 0 2.1819429176216493e-05
GC_11_19 b_11 NI_11 NS_19 0 1.3691770930120763e-04
GC_11_20 b_11 NI_11 NS_20 0 -1.9802490680622586e-05
GC_11_21 b_11 NI_11 NS_21 0 3.3573887954335791e-05
GC_11_22 b_11 NI_11 NS_22 0 2.3801839166632560e-05
GC_11_23 b_11 NI_11 NS_23 0 2.5634391886516806e-04
GC_11_24 b_11 NI_11 NS_24 0 1.1311513672013051e-04
GC_11_25 b_11 NI_11 NS_25 0 -2.0051802624497213e-04
GC_11_26 b_11 NI_11 NS_26 0 -2.4647199272213974e-04
GC_11_27 b_11 NI_11 NS_27 0 2.8763145924846129e-05
GC_11_28 b_11 NI_11 NS_28 0 6.7721919230652003e-05
GC_11_29 b_11 NI_11 NS_29 0 -9.6072866483684036e-05
GC_11_30 b_11 NI_11 NS_30 0 2.0919730836595888e-04
GC_11_31 b_11 NI_11 NS_31 0 8.5562393209248200e-06
GC_11_32 b_11 NI_11 NS_32 0 -7.2599892198543981e-05
GC_11_33 b_11 NI_11 NS_33 0 1.7602015256688587e-06
GC_11_34 b_11 NI_11 NS_34 0 7.5003885766292711e-05
GC_11_35 b_11 NI_11 NS_35 0 -2.2612257548687217e-05
GC_11_36 b_11 NI_11 NS_36 0 -1.9114406176336275e-05
GC_11_37 b_11 NI_11 NS_37 0 1.0465233138159147e-05
GC_11_38 b_11 NI_11 NS_38 0 6.6405199964782080e-06
GC_11_39 b_11 NI_11 NS_39 0 -6.0891852958693043e-03
GC_11_40 b_11 NI_11 NS_40 0 5.1284650432848150e-04
GC_11_41 b_11 NI_11 NS_41 0 2.0297472888782899e-03
GC_11_42 b_11 NI_11 NS_42 0 -7.2133118646992038e-03
GC_11_43 b_11 NI_11 NS_43 0 1.6451874685510198e-05
GC_11_44 b_11 NI_11 NS_44 0 3.8607096380780746e-04
GC_11_45 b_11 NI_11 NS_45 0 6.7671084316645437e-06
GC_11_46 b_11 NI_11 NS_46 0 1.6247958468643191e-04
GC_11_47 b_11 NI_11 NS_47 0 -6.3360781915316460e-05
GC_11_48 b_11 NI_11 NS_48 0 4.4581844958769502e-03
GC_11_49 b_11 NI_11 NS_49 0 1.8118273775085381e-05
GC_11_50 b_11 NI_11 NS_50 0 -3.1341300750460272e-05
GC_11_51 b_11 NI_11 NS_51 0 -1.8164054216542973e-03
GC_11_52 b_11 NI_11 NS_52 0 2.2732239350762747e-03
GC_11_53 b_11 NI_11 NS_53 0 1.5959970783231875e-05
GC_11_54 b_11 NI_11 NS_54 0 6.2604114563906659e-05
GC_11_55 b_11 NI_11 NS_55 0 2.2756973179480537e-05
GC_11_56 b_11 NI_11 NS_56 0 3.8454738855284607e-05
GC_11_57 b_11 NI_11 NS_57 0 1.5255492898900992e-05
GC_11_58 b_11 NI_11 NS_58 0 1.1679475479847519e-05
GC_11_59 b_11 NI_11 NS_59 0 5.7222165834358814e-05
GC_11_60 b_11 NI_11 NS_60 0 3.4478820538945022e-05
GC_11_61 b_11 NI_11 NS_61 0 -2.1949110433376305e-04
GC_11_62 b_11 NI_11 NS_62 0 -4.2445101749880151e-04
GC_11_63 b_11 NI_11 NS_63 0 7.1380895382932739e-05
GC_11_64 b_11 NI_11 NS_64 0 -3.0009868893515388e-04
GC_11_65 b_11 NI_11 NS_65 0 1.0856493515135171e-04
GC_11_66 b_11 NI_11 NS_66 0 -1.0592213910149152e-05
GC_11_67 b_11 NI_11 NS_67 0 -7.5738159593269046e-05
GC_11_68 b_11 NI_11 NS_68 0 1.5424535578477061e-04
GC_11_69 b_11 NI_11 NS_69 0 5.0741647705658734e-05
GC_11_70 b_11 NI_11 NS_70 0 -3.6179205698019870e-05
GC_11_71 b_11 NI_11 NS_71 0 -5.7671907870550490e-05
GC_11_72 b_11 NI_11 NS_72 0 4.0656278711928189e-05
GC_11_73 b_11 NI_11 NS_73 0 -2.2724737390586107e-05
GC_11_74 b_11 NI_11 NS_74 0 -4.9982570680484243e-05
GC_11_75 b_11 NI_11 NS_75 0 3.6063728521047501e-06
GC_11_76 b_11 NI_11 NS_76 0 3.9597413920792075e-06
GC_11_77 b_11 NI_11 NS_77 0 1.7525362303539183e-02
GC_11_78 b_11 NI_11 NS_78 0 -8.1893421755909303e-04
GC_11_79 b_11 NI_11 NS_79 0 -1.4206764830202967e-02
GC_11_80 b_11 NI_11 NS_80 0 2.3391777555343777e-03
GC_11_81 b_11 NI_11 NS_81 0 7.4477688474910574e-04
GC_11_82 b_11 NI_11 NS_82 0 -3.6149539531685963e-04
GC_11_83 b_11 NI_11 NS_83 0 1.8738094276051474e-04
GC_11_84 b_11 NI_11 NS_84 0 -2.1661004444174599e-04
GC_11_85 b_11 NI_11 NS_85 0 -6.6974409716547109e-04
GC_11_86 b_11 NI_11 NS_86 0 -7.4150412276779423e-03
GC_11_87 b_11 NI_11 NS_87 0 -1.8566598256101503e-05
GC_11_88 b_11 NI_11 NS_88 0 3.7166812781215435e-05
GC_11_89 b_11 NI_11 NS_89 0 4.6432890730919371e-03
GC_11_90 b_11 NI_11 NS_90 0 4.4301367098203140e-03
GC_11_91 b_11 NI_11 NS_91 0 2.2013975945596037e-05
GC_11_92 b_11 NI_11 NS_92 0 -4.2412613220417553e-05
GC_11_93 b_11 NI_11 NS_93 0 9.7578187939158288e-06
GC_11_94 b_11 NI_11 NS_94 0 3.8359227730863962e-05
GC_11_95 b_11 NI_11 NS_95 0 1.4627977345489632e-04
GC_11_96 b_11 NI_11 NS_96 0 -6.4987142821654993e-06
GC_11_97 b_11 NI_11 NS_97 0 3.0306541983693589e-05
GC_11_98 b_11 NI_11 NS_98 0 1.7091779988808225e-05
GC_11_99 b_11 NI_11 NS_99 0 -8.3197623757195235e-04
GC_11_100 b_11 NI_11 NS_100 0 -6.9564568981070319e-04
GC_11_101 b_11 NI_11 NS_101 0 -2.3649265687185908e-04
GC_11_102 b_11 NI_11 NS_102 0 -1.4542255679426014e-04
GC_11_103 b_11 NI_11 NS_103 0 2.9862197228757922e-04
GC_11_104 b_11 NI_11 NS_104 0 3.2664965089344064e-04
GC_11_105 b_11 NI_11 NS_105 0 7.2063762540506695e-05
GC_11_106 b_11 NI_11 NS_106 0 -3.4202924107805993e-05
GC_11_107 b_11 NI_11 NS_107 0 -2.0604201750674301e-05
GC_11_108 b_11 NI_11 NS_108 0 -2.6419099489580971e-05
GC_11_109 b_11 NI_11 NS_109 0 -8.1635789630065121e-06
GC_11_110 b_11 NI_11 NS_110 0 3.0365222612408889e-05
GC_11_111 b_11 NI_11 NS_111 0 -4.2276543837686215e-05
GC_11_112 b_11 NI_11 NS_112 0 -1.6526256016336749e-05
GC_11_113 b_11 NI_11 NS_113 0 1.1538916547362811e-06
GC_11_114 b_11 NI_11 NS_114 0 2.4982027479547950e-06
GC_11_115 b_11 NI_11 NS_115 0 3.3126596613846627e-03
GC_11_116 b_11 NI_11 NS_116 0 7.6895886125138405e-04
GC_11_117 b_11 NI_11 NS_117 0 -4.0804260636653133e-03
GC_11_118 b_11 NI_11 NS_118 0 -4.7421802485423051e-03
GC_11_119 b_11 NI_11 NS_119 0 1.2052527085649286e-04
GC_11_120 b_11 NI_11 NS_120 0 4.2767875907711239e-04
GC_11_121 b_11 NI_11 NS_121 0 7.2140352954886289e-05
GC_11_122 b_11 NI_11 NS_122 0 1.5686266901200540e-04
GC_11_123 b_11 NI_11 NS_123 0 -7.2547632277717735e-04
GC_11_124 b_11 NI_11 NS_124 0 5.5616549360361757e-03
GC_11_125 b_11 NI_11 NS_125 0 1.9791492922850782e-05
GC_11_126 b_11 NI_11 NS_126 0 -3.1303820290398339e-05
GC_11_127 b_11 NI_11 NS_127 0 1.0265401594665893e-03
GC_11_128 b_11 NI_11 NS_128 0 4.0272104390693250e-03
GC_11_129 b_11 NI_11 NS_129 0 4.0325297025798445e-05
GC_11_130 b_11 NI_11 NS_130 0 6.4029924599100672e-05
GC_11_131 b_11 NI_11 NS_131 0 2.0007415655734661e-05
GC_11_132 b_11 NI_11 NS_132 0 3.5171261858122946e-05
GC_11_133 b_11 NI_11 NS_133 0 8.1185149988564567e-05
GC_11_134 b_11 NI_11 NS_134 0 3.3200219430358155e-05
GC_11_135 b_11 NI_11 NS_135 0 5.8665200647834321e-05
GC_11_136 b_11 NI_11 NS_136 0 2.8730280284445550e-05
GC_11_137 b_11 NI_11 NS_137 0 -1.1141920502589168e-03
GC_11_138 b_11 NI_11 NS_138 0 -6.3143431710119724e-04
GC_11_139 b_11 NI_11 NS_139 0 7.1121968156985441e-06
GC_11_140 b_11 NI_11 NS_140 0 -2.8415371547900296e-04
GC_11_141 b_11 NI_11 NS_141 0 3.5994522869320134e-04
GC_11_142 b_11 NI_11 NS_142 0 2.2121729450357274e-04
GC_11_143 b_11 NI_11 NS_143 0 4.4364872261815712e-05
GC_11_144 b_11 NI_11 NS_144 0 -3.9892057308413064e-05
GC_11_145 b_11 NI_11 NS_145 0 -1.1723750058447194e-05
GC_11_146 b_11 NI_11 NS_146 0 -2.6256859215662192e-05
GC_11_147 b_11 NI_11 NS_147 0 -3.0778161146104479e-05
GC_11_148 b_11 NI_11 NS_148 0 1.5045823068562403e-05
GC_11_149 b_11 NI_11 NS_149 0 -3.4281893598740826e-05
GC_11_150 b_11 NI_11 NS_150 0 -3.5248847782545268e-05
GC_11_151 b_11 NI_11 NS_151 0 -1.7825968454980562e-06
GC_11_152 b_11 NI_11 NS_152 0 2.4531358641748597e-06
GC_11_153 b_11 NI_11 NS_153 0 -1.2243432774686921e-02
GC_11_154 b_11 NI_11 NS_154 0 -1.0230968460256660e-03
GC_11_155 b_11 NI_11 NS_155 0 -5.2688289784614184e-04
GC_11_156 b_11 NI_11 NS_156 0 7.4680601639112382e-03
GC_11_157 b_11 NI_11 NS_157 0 1.0116748945626355e-03
GC_11_158 b_11 NI_11 NS_158 0 -7.4477932689710443e-05
GC_11_159 b_11 NI_11 NS_159 0 1.4568491338366252e-04
GC_11_160 b_11 NI_11 NS_160 0 -1.9821039552117185e-04
GC_11_161 b_11 NI_11 NS_161 0 3.9935582346728778e-03
GC_11_162 b_11 NI_11 NS_162 0 -2.3501744492664327e-03
GC_11_163 b_11 NI_11 NS_163 0 -1.1344459634711998e-05
GC_11_164 b_11 NI_11 NS_164 0 -2.1422769433543885e-06
GC_11_165 b_11 NI_11 NS_165 0 8.1840014622498163e-03
GC_11_166 b_11 NI_11 NS_166 0 -5.2425608440929078e-03
GC_11_167 b_11 NI_11 NS_167 0 2.9233158852827346e-05
GC_11_168 b_11 NI_11 NS_168 0 -7.8957702806176222e-05
GC_11_169 b_11 NI_11 NS_169 0 3.9330266992239816e-06
GC_11_170 b_11 NI_11 NS_170 0 5.2531833338573226e-05
GC_11_171 b_11 NI_11 NS_171 0 -1.3963020794233089e-05
GC_11_172 b_11 NI_11 NS_172 0 -3.7407667576585411e-05
GC_11_173 b_11 NI_11 NS_173 0 -8.1075950892301587e-06
GC_11_174 b_11 NI_11 NS_174 0 -3.9234399312245435e-07
GC_11_175 b_11 NI_11 NS_175 0 -1.0696844035196478e-03
GC_11_176 b_11 NI_11 NS_176 0 1.6545896083485518e-03
GC_11_177 b_11 NI_11 NS_177 0 -3.1129565434633071e-04
GC_11_178 b_11 NI_11 NS_178 0 -1.3497352017881239e-04
GC_11_179 b_11 NI_11 NS_179 0 4.6296712715869059e-04
GC_11_180 b_11 NI_11 NS_180 0 8.7032084946215551e-05
GC_11_181 b_11 NI_11 NS_181 0 8.1031649819519555e-06
GC_11_182 b_11 NI_11 NS_182 0 -1.2224610267076385e-04
GC_11_183 b_11 NI_11 NS_183 0 -1.0120762403129076e-05
GC_11_184 b_11 NI_11 NS_184 0 5.3253370814242539e-05
GC_11_185 b_11 NI_11 NS_185 0 -2.8254819143599052e-05
GC_11_186 b_11 NI_11 NS_186 0 -1.6647624459342361e-05
GC_11_187 b_11 NI_11 NS_187 0 -1.0520166346544245e-04
GC_11_188 b_11 NI_11 NS_188 0 -2.4069902982602841e-06
GC_11_189 b_11 NI_11 NS_189 0 -2.8863550039254355e-06
GC_11_190 b_11 NI_11 NS_190 0 1.4300268014075762e-05
GC_11_191 b_11 NI_11 NS_191 0 1.3114856444320096e-02
GC_11_192 b_11 NI_11 NS_192 0 1.1287921871285104e-03
GC_11_193 b_11 NI_11 NS_193 0 -1.0788738729235747e-02
GC_11_194 b_11 NI_11 NS_194 0 2.9521786035010995e-03
GC_11_195 b_11 NI_11 NS_195 0 2.9915102791764269e-04
GC_11_196 b_11 NI_11 NS_196 0 5.1595076986915273e-05
GC_11_197 b_11 NI_11 NS_197 0 8.4650006558517643e-05
GC_11_198 b_11 NI_11 NS_198 0 -1.4000869427872668e-05
GC_11_199 b_11 NI_11 NS_199 0 -2.0500101926737950e-03
GC_11_200 b_11 NI_11 NS_200 0 5.4371834794486977e-03
GC_11_201 b_11 NI_11 NS_201 0 1.8062068985590932e-05
GC_11_202 b_11 NI_11 NS_202 0 3.7088510021526249e-06
GC_11_203 b_11 NI_11 NS_203 0 5.7156278871774687e-03
GC_11_204 b_11 NI_11 NS_204 0 1.4786778216009362e-03
GC_11_205 b_11 NI_11 NS_205 0 3.4123297156194431e-05
GC_11_206 b_11 NI_11 NS_206 0 -2.7367596253348879e-07
GC_11_207 b_11 NI_11 NS_207 0 1.5640866245024478e-05
GC_11_208 b_11 NI_11 NS_208 0 1.1835090364461678e-05
GC_11_209 b_11 NI_11 NS_209 0 -2.3477147428090500e-05
GC_11_210 b_11 NI_11 NS_210 0 5.6195528008901743e-06
GC_11_211 b_11 NI_11 NS_211 0 8.5408159137197197e-06
GC_11_212 b_11 NI_11 NS_212 0 2.0225222035646312e-06
GC_11_213 b_11 NI_11 NS_213 0 -1.5488808633677435e-03
GC_11_214 b_11 NI_11 NS_214 0 4.1443659195217918e-04
GC_11_215 b_11 NI_11 NS_215 0 -1.3079482927369710e-04
GC_11_216 b_11 NI_11 NS_216 0 -5.4858474997280199e-05
GC_11_217 b_11 NI_11 NS_217 0 4.1675239723779371e-04
GC_11_218 b_11 NI_11 NS_218 0 2.3957042027785219e-04
GC_11_219 b_11 NI_11 NS_219 0 1.1903826655270087e-04
GC_11_220 b_11 NI_11 NS_220 0 -7.5516366903426993e-05
GC_11_221 b_11 NI_11 NS_221 0 -7.8642619061494175e-05
GC_11_222 b_11 NI_11 NS_222 0 -8.6887067834865197e-06
GC_11_223 b_11 NI_11 NS_223 0 4.2193956511448782e-05
GC_11_224 b_11 NI_11 NS_224 0 2.8008480703952345e-06
GC_11_225 b_11 NI_11 NS_225 0 -8.2703156371833773e-05
GC_11_226 b_11 NI_11 NS_226 0 -1.4121307633726938e-05
GC_11_227 b_11 NI_11 NS_227 0 -4.6017501060223501e-07
GC_11_228 b_11 NI_11 NS_228 0 -8.3683952462201037e-07
GC_11_229 b_11 NI_11 NS_229 0 -2.2063229378628986e-02
GC_11_230 b_11 NI_11 NS_230 0 -1.2404852964999977e-03
GC_11_231 b_11 NI_11 NS_231 0 9.0929508719168536e-03
GC_11_232 b_11 NI_11 NS_232 0 1.2497558860945040e-02
GC_11_233 b_11 NI_11 NS_233 0 6.5547352832035367e-04
GC_11_234 b_11 NI_11 NS_234 0 3.4687006714260364e-04
GC_11_235 b_11 NI_11 NS_235 0 -2.9912152876675814e-05
GC_11_236 b_11 NI_11 NS_236 0 3.8593595422283616e-06
GC_11_237 b_11 NI_11 NS_237 0 7.9878843901873137e-03
GC_11_238 b_11 NI_11 NS_238 0 6.9054687179096255e-03
GC_11_239 b_11 NI_11 NS_239 0 -2.2590374667124456e-05
GC_11_240 b_11 NI_11 NS_240 0 -5.6416706621680126e-06
GC_11_241 b_11 NI_11 NS_241 0 1.1053267339791938e-02
GC_11_242 b_11 NI_11 NS_242 0 -8.4973923246830785e-03
GC_11_243 b_11 NI_11 NS_243 0 2.0542000162352375e-05
GC_11_244 b_11 NI_11 NS_244 0 -4.9643739044583268e-05
GC_11_245 b_11 NI_11 NS_245 0 1.4412777535290286e-05
GC_11_246 b_11 NI_11 NS_246 0 4.8043892583669744e-05
GC_11_247 b_11 NI_11 NS_247 0 -4.6872858290059584e-05
GC_11_248 b_11 NI_11 NS_248 0 -3.9804231913452411e-05
GC_11_249 b_11 NI_11 NS_249 0 -3.0368042457981146e-06
GC_11_250 b_11 NI_11 NS_250 0 -5.5033948731942925e-06
GC_11_251 b_11 NI_11 NS_251 0 -3.5805773166813501e-03
GC_11_252 b_11 NI_11 NS_252 0 1.8314129807043907e-03
GC_11_253 b_11 NI_11 NS_253 0 -3.7094216759325712e-04
GC_11_254 b_11 NI_11 NS_254 0 -3.7653035760137121e-05
GC_11_255 b_11 NI_11 NS_255 0 8.8294476670418732e-04
GC_11_256 b_11 NI_11 NS_256 0 1.4453598956108940e-04
GC_11_257 b_11 NI_11 NS_257 0 1.0048072975890485e-04
GC_11_258 b_11 NI_11 NS_258 0 -4.0978329630046668e-04
GC_11_259 b_11 NI_11 NS_259 0 -5.3902400866281962e-05
GC_11_260 b_11 NI_11 NS_260 0 5.7205110140767192e-05
GC_11_261 b_11 NI_11 NS_261 0 -2.0528967647485662e-05
GC_11_262 b_11 NI_11 NS_262 0 1.2982711468007774e-05
GC_11_263 b_11 NI_11 NS_263 0 -4.3693364824250030e-05
GC_11_264 b_11 NI_11 NS_264 0 3.5039981113676949e-05
GC_11_265 b_11 NI_11 NS_265 0 -5.0899314481643429e-06
GC_11_266 b_11 NI_11 NS_266 0 1.4045253616946629e-08
GC_11_267 b_11 NI_11 NS_267 0 2.8297173310085019e-02
GC_11_268 b_11 NI_11 NS_268 0 1.2246464029386319e-03
GC_11_269 b_11 NI_11 NS_269 0 -1.6132322407377355e-02
GC_11_270 b_11 NI_11 NS_270 0 4.6064719487240750e-03
GC_11_271 b_11 NI_11 NS_271 0 -1.8478349238667237e-04
GC_11_272 b_11 NI_11 NS_272 0 2.2350023366089958e-05
GC_11_273 b_11 NI_11 NS_273 0 -3.0699696909636315e-05
GC_11_274 b_11 NI_11 NS_274 0 -2.3501896501964950e-05
GC_11_275 b_11 NI_11 NS_275 0 -6.7574310849061779e-03
GC_11_276 b_11 NI_11 NS_276 0 -5.1973307776146003e-03
GC_11_277 b_11 NI_11 NS_277 0 2.4010518317242742e-05
GC_11_278 b_11 NI_11 NS_278 0 8.4647095462183932e-06
GC_11_279 b_11 NI_11 NS_279 0 9.5680349106861094e-03
GC_11_280 b_11 NI_11 NS_280 0 3.5539638562877267e-03
GC_11_281 b_11 NI_11 NS_281 0 7.1086763883097732e-06
GC_11_282 b_11 NI_11 NS_282 0 2.2745131365106848e-05
GC_11_283 b_11 NI_11 NS_283 0 1.2237669091177928e-05
GC_11_284 b_11 NI_11 NS_284 0 1.0377937578020044e-05
GC_11_285 b_11 NI_11 NS_285 0 -1.3763336448629433e-05
GC_11_286 b_11 NI_11 NS_286 0 -2.4632483289900633e-05
GC_11_287 b_11 NI_11 NS_287 0 1.4186578687330027e-05
GC_11_288 b_11 NI_11 NS_288 0 -2.1387317662892086e-06
GC_11_289 b_11 NI_11 NS_289 0 -3.4617839640117272e-03
GC_11_290 b_11 NI_11 NS_290 0 -3.5295960105517939e-04
GC_11_291 b_11 NI_11 NS_291 0 -1.8079087103754467e-04
GC_11_292 b_11 NI_11 NS_292 0 -4.3804089303866842e-05
GC_11_293 b_11 NI_11 NS_293 0 7.3199983272278883e-04
GC_11_294 b_11 NI_11 NS_294 0 4.4593318676220290e-04
GC_11_295 b_11 NI_11 NS_295 0 2.5334563905114889e-04
GC_11_296 b_11 NI_11 NS_296 0 -2.9257201342546278e-04
GC_11_297 b_11 NI_11 NS_297 0 -8.4270049136394082e-05
GC_11_298 b_11 NI_11 NS_298 0 -2.4066599994600728e-05
GC_11_299 b_11 NI_11 NS_299 0 -1.2715183653510639e-05
GC_11_300 b_11 NI_11 NS_300 0 -5.0280919033906111e-06
GC_11_301 b_11 NI_11 NS_301 0 -4.7194961268532305e-05
GC_11_302 b_11 NI_11 NS_302 0 1.9039237232810966e-05
GC_11_303 b_11 NI_11 NS_303 0 -1.7441535283474903e-07
GC_11_304 b_11 NI_11 NS_304 0 -8.9069053975575698e-06
GC_11_305 b_11 NI_11 NS_305 0 -2.9758686994037664e-02
GC_11_306 b_11 NI_11 NS_306 0 -1.3212972999271306e-03
GC_11_307 b_11 NI_11 NS_307 0 1.8973454099461957e-02
GC_11_308 b_11 NI_11 NS_308 0 2.6527160896856524e-02
GC_11_309 b_11 NI_11 NS_309 0 -5.4241460335888647e-04
GC_11_310 b_11 NI_11 NS_310 0 9.5578596284331258e-04
GC_11_311 b_11 NI_11 NS_311 0 -2.6747247108127110e-04
GC_11_312 b_11 NI_11 NS_312 0 3.1348153485449582e-04
GC_11_313 b_11 NI_11 NS_313 0 1.3303976698581754e-02
GC_11_314 b_11 NI_11 NS_314 0 2.7451548727576037e-02
GC_11_315 b_11 NI_11 NS_315 0 -3.8837928196611817e-05
GC_11_316 b_11 NI_11 NS_316 0 -9.5372240676790300e-05
GC_11_317 b_11 NI_11 NS_317 0 2.1886886830289453e-02
GC_11_318 b_11 NI_11 NS_318 0 -2.2631573862302405e-02
GC_11_319 b_11 NI_11 NS_319 0 -5.0525476161445574e-05
GC_11_320 b_11 NI_11 NS_320 0 3.9152150457078525e-05
GC_11_321 b_11 NI_11 NS_321 0 2.1199397131008649e-06
GC_11_322 b_11 NI_11 NS_322 0 8.5625200610919675e-05
GC_11_323 b_11 NI_11 NS_323 0 -2.2649306888483593e-04
GC_11_324 b_11 NI_11 NS_324 0 -5.8352278748121529e-05
GC_11_325 b_11 NI_11 NS_325 0 -3.5799782575350721e-05
GC_11_326 b_11 NI_11 NS_326 0 -2.8441069964313928e-05
GC_11_327 b_11 NI_11 NS_327 0 -6.6681002619813261e-03
GC_11_328 b_11 NI_11 NS_328 0 7.8488365759612974e-03
GC_11_329 b_11 NI_11 NS_329 0 -5.0473947264516230e-04
GC_11_330 b_11 NI_11 NS_330 0 -2.2428200475591207e-04
GC_11_331 b_11 NI_11 NS_331 0 7.8075953692517642e-04
GC_11_332 b_11 NI_11 NS_332 0 9.5968416066302762e-05
GC_11_333 b_11 NI_11 NS_333 0 1.2484201203428257e-04
GC_11_334 b_11 NI_11 NS_334 0 -3.0756669888434775e-04
GC_11_335 b_11 NI_11 NS_335 0 8.9479246938943914e-06
GC_11_336 b_11 NI_11 NS_336 0 -6.8019709971402551e-06
GC_11_337 b_11 NI_11 NS_337 0 4.1387139876546132e-05
GC_11_338 b_11 NI_11 NS_338 0 -4.5502875869675838e-05
GC_11_339 b_11 NI_11 NS_339 0 -3.7154871645335171e-06
GC_11_340 b_11 NI_11 NS_340 0 -4.9682904267592117e-05
GC_11_341 b_11 NI_11 NS_341 0 -1.6767404744238353e-05
GC_11_342 b_11 NI_11 NS_342 0 -6.4757179785663409e-06
GC_11_343 b_11 NI_11 NS_343 0 5.7049334366697423e-02
GC_11_344 b_11 NI_11 NS_344 0 9.2458667546044433e-04
GC_11_345 b_11 NI_11 NS_345 0 -3.4891118115797634e-02
GC_11_346 b_11 NI_11 NS_346 0 -1.4434479294245361e-02
GC_11_347 b_11 NI_11 NS_347 0 -6.2028509819578997e-04
GC_11_348 b_11 NI_11 NS_348 0 2.6315366158804961e-04
GC_11_349 b_11 NI_11 NS_349 0 -1.3720226006819309e-04
GC_11_350 b_11 NI_11 NS_350 0 1.2169639549909166e-04
GC_11_351 b_11 NI_11 NS_351 0 -2.4467227914756737e-02
GC_11_352 b_11 NI_11 NS_352 0 -4.3614096720367930e-02
GC_11_353 b_11 NI_11 NS_353 0 1.5965248284230578e-05
GC_11_354 b_11 NI_11 NS_354 0 8.3164201595976869e-05
GC_11_355 b_11 NI_11 NS_355 0 1.3305170308541010e-02
GC_11_356 b_11 NI_11 NS_356 0 -2.1310553191137530e-04
GC_11_357 b_11 NI_11 NS_357 0 -2.5927784724858720e-05
GC_11_358 b_11 NI_11 NS_358 0 5.0410634161256108e-05
GC_11_359 b_11 NI_11 NS_359 0 -5.8761442150335742e-06
GC_11_360 b_11 NI_11 NS_360 0 3.9650498084956317e-05
GC_11_361 b_11 NI_11 NS_361 0 -1.1890160423336639e-04
GC_11_362 b_11 NI_11 NS_362 0 -2.7600973257612936e-05
GC_11_363 b_11 NI_11 NS_363 0 -2.4374749935815833e-05
GC_11_364 b_11 NI_11 NS_364 0 -2.5382462477963791e-05
GC_11_365 b_11 NI_11 NS_365 0 -5.4410008621515191e-03
GC_11_366 b_11 NI_11 NS_366 0 4.1779973124300568e-03
GC_11_367 b_11 NI_11 NS_367 0 -1.5876734011551814e-04
GC_11_368 b_11 NI_11 NS_368 0 -2.5089711230726855e-04
GC_11_369 b_11 NI_11 NS_369 0 6.2375804344798271e-04
GC_11_370 b_11 NI_11 NS_370 0 2.1598650365279459e-04
GC_11_371 b_11 NI_11 NS_371 0 1.8537918445404262e-04
GC_11_372 b_11 NI_11 NS_372 0 -2.3876091100791491e-04
GC_11_373 b_11 NI_11 NS_373 0 3.4178604654706713e-05
GC_11_374 b_11 NI_11 NS_374 0 1.3038952980007208e-05
GC_11_375 b_11 NI_11 NS_375 0 3.2313415911120940e-05
GC_11_376 b_11 NI_11 NS_376 0 -3.5400564416623729e-05
GC_11_377 b_11 NI_11 NS_377 0 -7.1009824621884441e-06
GC_11_378 b_11 NI_11 NS_378 0 1.8975510006222506e-05
GC_11_379 b_11 NI_11 NS_379 0 -3.8064296291005859e-06
GC_11_380 b_11 NI_11 NS_380 0 -5.9647414025911526e-06
GC_11_381 b_11 NI_11 NS_381 0 3.8286173448358642e-02
GC_11_382 b_11 NI_11 NS_382 0 -1.3309973624776889e-03
GC_11_383 b_11 NI_11 NS_383 0 6.1900653263971123e-02
GC_11_384 b_11 NI_11 NS_384 0 -6.4202552868157556e-02
GC_11_385 b_11 NI_11 NS_385 0 -3.2415295004883716e-03
GC_11_386 b_11 NI_11 NS_386 0 -9.1959309900846106e-04
GC_11_387 b_11 NI_11 NS_387 0 -4.7155107535035081e-04
GC_11_388 b_11 NI_11 NS_388 0 2.6540388252082036e-04
GC_11_389 b_11 NI_11 NS_389 0 -1.1397807938122945e-02
GC_11_390 b_11 NI_11 NS_390 0 1.6821755050486015e-02
GC_11_391 b_11 NI_11 NS_391 0 -3.6016276661829929e-05
GC_11_392 b_11 NI_11 NS_392 0 -9.0266375601688470e-05
GC_11_393 b_11 NI_11 NS_393 0 -5.0764418314765768e-02
GC_11_394 b_11 NI_11 NS_394 0 9.0817216836928700e-04
GC_11_395 b_11 NI_11 NS_395 0 -1.2165976354201439e-04
GC_11_396 b_11 NI_11 NS_396 0 6.7618745686309347e-05
GC_11_397 b_11 NI_11 NS_397 0 2.2585910586083706e-05
GC_11_398 b_11 NI_11 NS_398 0 -5.1825724620381355e-06
GC_11_399 b_11 NI_11 NS_399 0 -2.3807806114253780e-04
GC_11_400 b_11 NI_11 NS_400 0 -4.6289812722526048e-05
GC_11_401 b_11 NI_11 NS_401 0 -2.4204043251134825e-05
GC_11_402 b_11 NI_11 NS_402 0 -1.9328395888998225e-05
GC_11_403 b_11 NI_11 NS_403 0 -4.7034602251975035e-03
GC_11_404 b_11 NI_11 NS_404 0 5.7772967818827620e-03
GC_11_405 b_11 NI_11 NS_405 0 -4.3215011077842269e-04
GC_11_406 b_11 NI_11 NS_406 0 2.7890337098331720e-05
GC_11_407 b_11 NI_11 NS_407 0 1.0353915511806036e-03
GC_11_408 b_11 NI_11 NS_408 0 5.4720082942092110e-05
GC_11_409 b_11 NI_11 NS_409 0 9.0552880573762897e-05
GC_11_410 b_11 NI_11 NS_410 0 -4.8846080529011825e-04
GC_11_411 b_11 NI_11 NS_411 0 1.2429564265412465e-04
GC_11_412 b_11 NI_11 NS_412 0 -5.4213025294888374e-05
GC_11_413 b_11 NI_11 NS_413 0 6.0125016523340616e-05
GC_11_414 b_11 NI_11 NS_414 0 -7.9557303331191556e-05
GC_11_415 b_11 NI_11 NS_415 0 7.8831357355413982e-05
GC_11_416 b_11 NI_11 NS_416 0 -3.1635641199367456e-06
GC_11_417 b_11 NI_11 NS_417 0 -1.2216753409198436e-05
GC_11_418 b_11 NI_11 NS_418 0 -1.3554710853422533e-05
GC_11_419 b_11 NI_11 NS_419 0 1.9324373648156312e-02
GC_11_420 b_11 NI_11 NS_420 0 1.8259620081006261e-03
GC_11_421 b_11 NI_11 NS_421 0 2.4610410480565930e-02
GC_11_422 b_11 NI_11 NS_422 0 -1.6224651574562422e-02
GC_11_423 b_11 NI_11 NS_423 0 1.2917168901901033e-03
GC_11_424 b_11 NI_11 NS_424 0 6.9502506043464524e-05
GC_11_425 b_11 NI_11 NS_425 0 1.4149587769442107e-05
GC_11_426 b_11 NI_11 NS_426 0 3.4006069791268352e-05
GC_11_427 b_11 NI_11 NS_427 0 2.6070945074820391e-02
GC_11_428 b_11 NI_11 NS_428 0 2.4077603128284781e-03
GC_11_429 b_11 NI_11 NS_429 0 4.0640875540198221e-05
GC_11_430 b_11 NI_11 NS_430 0 8.6258653861871832e-05
GC_11_431 b_11 NI_11 NS_431 0 -4.5704222947255409e-02
GC_11_432 b_11 NI_11 NS_432 0 3.2071097015620963e-02
GC_11_433 b_11 NI_11 NS_433 0 -3.9747579253640223e-05
GC_11_434 b_11 NI_11 NS_434 0 8.1760321655267203e-05
GC_11_435 b_11 NI_11 NS_435 0 5.0752801873980368e-05
GC_11_436 b_11 NI_11 NS_436 0 1.6309091262461509e-05
GC_11_437 b_11 NI_11 NS_437 0 -1.2946889790428124e-04
GC_11_438 b_11 NI_11 NS_438 0 -3.4899506157469947e-05
GC_11_439 b_11 NI_11 NS_439 0 -2.0618630734140787e-05
GC_11_440 b_11 NI_11 NS_440 0 -1.5588245023491003e-05
GC_11_441 b_11 NI_11 NS_441 0 -4.0752602899988858e-03
GC_11_442 b_11 NI_11 NS_442 0 3.0867286752573095e-04
GC_11_443 b_11 NI_11 NS_443 0 -1.2734754794673476e-04
GC_11_444 b_11 NI_11 NS_444 0 6.9394274904934123e-05
GC_11_445 b_11 NI_11 NS_445 0 8.2501101247835088e-04
GC_11_446 b_11 NI_11 NS_446 0 6.2737999790004348e-04
GC_11_447 b_11 NI_11 NS_447 0 3.2408905210367712e-04
GC_11_448 b_11 NI_11 NS_448 0 -3.6391678140871984e-04
GC_11_449 b_11 NI_11 NS_449 0 1.4130506387190415e-04
GC_11_450 b_11 NI_11 NS_450 0 1.9597992956074212e-05
GC_11_451 b_11 NI_11 NS_451 0 8.5959879890491829e-05
GC_11_452 b_11 NI_11 NS_452 0 -8.1241377704726684e-06
GC_11_453 b_11 NI_11 NS_453 0 3.7362849658474951e-05
GC_11_454 b_11 NI_11 NS_454 0 7.7182121489254685e-05
GC_11_455 b_11 NI_11 NS_455 0 1.2980536820677831e-05
GC_11_456 b_11 NI_11 NS_456 0 -1.2819386219481447e-05
GD_11_1 b_11 NI_11 NA_1 0 -3.5471377605590338e-03
GD_11_2 b_11 NI_11 NA_2 0 5.6421795812681749e-03
GD_11_3 b_11 NI_11 NA_3 0 -5.8234354061276923e-03
GD_11_4 b_11 NI_11 NA_4 0 3.3123519438670821e-04
GD_11_5 b_11 NI_11 NA_5 0 -4.7349378475581623e-04
GD_11_6 b_11 NI_11 NA_6 0 -5.6239373596878141e-03
GD_11_7 b_11 NI_11 NA_7 0 -6.5420482390400447e-03
GD_11_8 b_11 NI_11 NA_8 0 -1.1769265684899829e-02
GD_11_9 b_11 NI_11 NA_9 0 -1.9098073287263952e-02
GD_11_10 b_11 NI_11 NA_10 0 1.7510448623952767e-03
GD_11_11 b_11 NI_11 NA_11 0 -6.4455764844236194e-02
GD_11_12 b_11 NI_11 NA_12 0 -3.3054978222160282e-02
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 -1.2388825442102504e-03
GC_12_2 b_12 NI_12 NS_2 0 5.1570788076757792e-04
GC_12_3 b_12 NI_12 NS_3 0 -6.5344504657048293e-04
GC_12_4 b_12 NI_12 NS_4 0 -9.2584737458167898e-04
GC_12_5 b_12 NI_12 NS_5 0 -9.1862827878091678e-05
GC_12_6 b_12 NI_12 NS_6 0 2.2352062221736203e-04
GC_12_7 b_12 NI_12 NS_7 0 7.3111050249512164e-05
GC_12_8 b_12 NI_12 NS_8 0 -1.0500400947839343e-05
GC_12_9 b_12 NI_12 NS_9 0 2.7464067920455515e-05
GC_12_10 b_12 NI_12 NS_10 0 4.5900457558491611e-03
GC_12_11 b_12 NI_12 NS_11 0 1.9614338149760619e-05
GC_12_12 b_12 NI_12 NS_12 0 -3.2331325345561492e-05
GC_12_13 b_12 NI_12 NS_13 0 4.1682719671909266e-04
GC_12_14 b_12 NI_12 NS_14 0 2.0359940910366484e-04
GC_12_15 b_12 NI_12 NS_15 0 5.9368040964213770e-06
GC_12_16 b_12 NI_12 NS_16 0 3.3468406794044595e-05
GC_12_17 b_12 NI_12 NS_17 0 -5.4465320740411660e-07
GC_12_18 b_12 NI_12 NS_18 0 3.3307329034361184e-05
GC_12_19 b_12 NI_12 NS_19 0 8.3237859594566808e-05
GC_12_20 b_12 NI_12 NS_20 0 1.5054112595105116e-07
GC_12_21 b_12 NI_12 NS_21 0 2.7190039265534389e-05
GC_12_22 b_12 NI_12 NS_22 0 2.6244528753374182e-05
GC_12_23 b_12 NI_12 NS_23 0 -2.5004210648727400e-05
GC_12_24 b_12 NI_12 NS_24 0 4.9807781378454429e-04
GC_12_25 b_12 NI_12 NS_25 0 9.8187095191162583e-05
GC_12_26 b_12 NI_12 NS_26 0 -4.7654015516249636e-04
GC_12_27 b_12 NI_12 NS_27 0 -1.0710130519884615e-05
GC_12_28 b_12 NI_12 NS_28 0 -1.2070446451163193e-04
GC_12_29 b_12 NI_12 NS_29 0 -1.9293923169937498e-04
GC_12_30 b_12 NI_12 NS_30 0 1.7760741312731920e-04
GC_12_31 b_12 NI_12 NS_31 0 3.9441100685244725e-05
GC_12_32 b_12 NI_12 NS_32 0 -4.2471890637876249e-05
GC_12_33 b_12 NI_12 NS_33 0 -4.4345430973438804e-05
GC_12_34 b_12 NI_12 NS_34 0 6.7680670416849317e-05
GC_12_35 b_12 NI_12 NS_35 0 7.0036031387887396e-06
GC_12_36 b_12 NI_12 NS_36 0 -4.1817284445404211e-05
GC_12_37 b_12 NI_12 NS_37 0 -1.3573455891045298e-06
GC_12_38 b_12 NI_12 NS_38 0 1.1220228347569958e-05
GC_12_39 b_12 NI_12 NS_39 0 6.3440273537645284e-03
GC_12_40 b_12 NI_12 NS_40 0 -5.5836212371708732e-04
GC_12_41 b_12 NI_12 NS_41 0 -5.2521354059643175e-03
GC_12_42 b_12 NI_12 NS_42 0 -4.4858919985252448e-03
GC_12_43 b_12 NI_12 NS_43 0 8.0084189599060696e-05
GC_12_44 b_12 NI_12 NS_44 0 8.9793323054880697e-05
GC_12_45 b_12 NI_12 NS_45 0 -5.5760985825788784e-06
GC_12_46 b_12 NI_12 NS_46 0 1.2806696076042624e-04
GC_12_47 b_12 NI_12 NS_47 0 -7.8554938379383924e-04
GC_12_48 b_12 NI_12 NS_48 0 -5.9315644706753158e-03
GC_12_49 b_12 NI_12 NS_49 0 -2.0761648140112290e-05
GC_12_50 b_12 NI_12 NS_50 0 2.6683462969164912e-05
GC_12_51 b_12 NI_12 NS_51 0 1.9552677789372260e-03
GC_12_52 b_12 NI_12 NS_52 0 4.1918097444532130e-03
GC_12_53 b_12 NI_12 NS_53 0 3.8972368019414821e-05
GC_12_54 b_12 NI_12 NS_54 0 5.5701498248370561e-05
GC_12_55 b_12 NI_12 NS_55 0 1.2633154222321443e-05
GC_12_56 b_12 NI_12 NS_56 0 4.0861843182636973e-05
GC_12_57 b_12 NI_12 NS_57 0 1.1063479671776688e-05
GC_12_58 b_12 NI_12 NS_58 0 8.6024590067058689e-06
GC_12_59 b_12 NI_12 NS_59 0 4.6828889300880019e-05
GC_12_60 b_12 NI_12 NS_60 0 3.9094896278237631e-05
GC_12_61 b_12 NI_12 NS_61 0 -1.8761098161632211e-03
GC_12_62 b_12 NI_12 NS_62 0 1.1360974652175114e-04
GC_12_63 b_12 NI_12 NS_63 0 4.4578299979821452e-04
GC_12_64 b_12 NI_12 NS_64 0 -5.3001939029482235e-04
GC_12_65 b_12 NI_12 NS_65 0 2.3017874819296455e-04
GC_12_66 b_12 NI_12 NS_66 0 -2.2603696905037471e-04
GC_12_67 b_12 NI_12 NS_67 0 -1.6770901069250465e-04
GC_12_68 b_12 NI_12 NS_68 0 9.9079444074836058e-05
GC_12_69 b_12 NI_12 NS_69 0 4.4992851025052334e-05
GC_12_70 b_12 NI_12 NS_70 0 3.5276150125949222e-06
GC_12_71 b_12 NI_12 NS_71 0 -7.5820287950918470e-05
GC_12_72 b_12 NI_12 NS_72 0 -7.5058192899285440e-06
GC_12_73 b_12 NI_12 NS_73 0 2.5241059467078368e-05
GC_12_74 b_12 NI_12 NS_74 0 -7.2477178280915330e-05
GC_12_75 b_12 NI_12 NS_75 0 -2.9014235024573518e-06
GC_12_76 b_12 NI_12 NS_76 0 9.9041220864345716e-06
GC_12_77 b_12 NI_12 NS_77 0 7.3339076078213286e-03
GC_12_78 b_12 NI_12 NS_78 0 8.2243797316050571e-04
GC_12_79 b_12 NI_12 NS_79 0 -7.3854185849669025e-03
GC_12_80 b_12 NI_12 NS_80 0 1.6955081630884354e-03
GC_12_81 b_12 NI_12 NS_81 0 1.4765753779779221e-04
GC_12_82 b_12 NI_12 NS_82 0 -9.3134357725069964e-05
GC_12_83 b_12 NI_12 NS_83 0 6.8656691191737148e-05
GC_12_84 b_12 NI_12 NS_84 0 -6.8102414599616323e-05
GC_12_85 b_12 NI_12 NS_85 0 -3.6468616493767395e-04
GC_12_86 b_12 NI_12 NS_86 0 6.6707434395170380e-03
GC_12_87 b_12 NI_12 NS_87 0 2.0794162488936908e-05
GC_12_88 b_12 NI_12 NS_88 0 -3.2738976778469039e-05
GC_12_89 b_12 NI_12 NS_89 0 3.6219187070852502e-03
GC_12_90 b_12 NI_12 NS_90 0 2.6309995188893058e-03
GC_12_91 b_12 NI_12 NS_91 0 4.4586128149690108e-06
GC_12_92 b_12 NI_12 NS_92 0 -2.3074162712801853e-05
GC_12_93 b_12 NI_12 NS_93 0 -2.4885310129145392e-06
GC_12_94 b_12 NI_12 NS_94 0 4.5350771888842988e-05
GC_12_95 b_12 NI_12 NS_95 0 8.7426867667210256e-05
GC_12_96 b_12 NI_12 NS_96 0 6.9923347943043929e-06
GC_12_97 b_12 NI_12 NS_97 0 2.5887691573404132e-05
GC_12_98 b_12 NI_12 NS_98 0 1.9262437901660157e-05
GC_12_99 b_12 NI_12 NS_99 0 -1.2001189261312869e-03
GC_12_100 b_12 NI_12 NS_100 0 -2.2059248448488440e-04
GC_12_101 b_12 NI_12 NS_101 0 1.5451284741028968e-05
GC_12_102 b_12 NI_12 NS_102 0 -3.6371149544032631e-04
GC_12_103 b_12 NI_12 NS_103 0 1.9751339640343351e-04
GC_12_104 b_12 NI_12 NS_104 0 2.3879432312760192e-04
GC_12_105 b_12 NI_12 NS_105 0 6.3161983642696714e-05
GC_12_106 b_12 NI_12 NS_106 0 7.5036777713908563e-06
GC_12_107 b_12 NI_12 NS_107 0 -5.0935582554959460e-06
GC_12_108 b_12 NI_12 NS_108 0 -2.8261363163849652e-05
GC_12_109 b_12 NI_12 NS_109 0 -2.3421881886198583e-05
GC_12_110 b_12 NI_12 NS_110 0 1.8312295358042118e-05
GC_12_111 b_12 NI_12 NS_111 0 -1.4242374161090816e-05
GC_12_112 b_12 NI_12 NS_112 0 -4.4664993607254028e-05
GC_12_113 b_12 NI_12 NS_113 0 -2.1349428600753784e-06
GC_12_114 b_12 NI_12 NS_114 0 -1.4680901807195112e-06
GC_12_115 b_12 NI_12 NS_115 0 1.7604529112116150e-02
GC_12_116 b_12 NI_12 NS_116 0 -8.5633039341564564e-04
GC_12_117 b_12 NI_12 NS_117 0 -1.2299201138022959e-02
GC_12_118 b_12 NI_12 NS_118 0 -4.1211416403004004e-03
GC_12_119 b_12 NI_12 NS_119 0 2.8176342796296057e-04
GC_12_120 b_12 NI_12 NS_120 0 3.6191572332329330e-06
GC_12_121 b_12 NI_12 NS_121 0 4.2441040353210352e-05
GC_12_122 b_12 NI_12 NS_122 0 8.1711269724230395e-05
GC_12_123 b_12 NI_12 NS_123 0 -1.4405612172868579e-03
GC_12_124 b_12 NI_12 NS_124 0 -8.7482261617895761e-03
GC_12_125 b_12 NI_12 NS_125 0 -2.3899052769040151e-05
GC_12_126 b_12 NI_12 NS_126 0 2.6164878620311938e-05
GC_12_127 b_12 NI_12 NS_127 0 3.3222373240285484e-03
GC_12_128 b_12 NI_12 NS_128 0 7.6830806418595240e-03
GC_12_129 b_12 NI_12 NS_129 0 5.0517525227131519e-05
GC_12_130 b_12 NI_12 NS_130 0 3.7503006546175213e-05
GC_12_131 b_12 NI_12 NS_131 0 5.7796531238281520e-06
GC_12_132 b_12 NI_12 NS_132 0 3.3711642636119574e-05
GC_12_133 b_12 NI_12 NS_133 0 4.9011858228137959e-05
GC_12_134 b_12 NI_12 NS_134 0 2.3614323501646825e-05
GC_12_135 b_12 NI_12 NS_135 0 5.0475002051129334e-05
GC_12_136 b_12 NI_12 NS_136 0 3.4328931840794889e-05
GC_12_137 b_12 NI_12 NS_137 0 -2.4659121598534441e-03
GC_12_138 b_12 NI_12 NS_138 0 -9.0314061139446780e-04
GC_12_139 b_12 NI_12 NS_139 0 3.9476870359991882e-04
GC_12_140 b_12 NI_12 NS_140 0 -4.2264640429812860e-04
GC_12_141 b_12 NI_12 NS_141 0 3.9089060941585206e-04
GC_12_142 b_12 NI_12 NS_142 0 1.3971483575583117e-04
GC_12_143 b_12 NI_12 NS_143 0 2.7987828693065576e-05
GC_12_144 b_12 NI_12 NS_144 0 -2.7292050403953945e-05
GC_12_145 b_12 NI_12 NS_145 0 -1.9097269766530833e-06
GC_12_146 b_12 NI_12 NS_146 0 -2.3373105906829697e-05
GC_12_147 b_12 NI_12 NS_147 0 -3.4922820252420641e-05
GC_12_148 b_12 NI_12 NS_148 0 -1.2539740367185492e-05
GC_12_149 b_12 NI_12 NS_149 0 1.0813188431810437e-06
GC_12_150 b_12 NI_12 NS_150 0 -6.3106493668506927e-05
GC_12_151 b_12 NI_12 NS_151 0 -1.0039034769220428e-05
GC_12_152 b_12 NI_12 NS_152 0 1.9683122489054912e-06
GC_12_153 b_12 NI_12 NS_153 0 2.4018996698136980e-02
GC_12_154 b_12 NI_12 NS_154 0 1.1010201447625397e-03
GC_12_155 b_12 NI_12 NS_155 0 -1.9027009242466607e-02
GC_12_156 b_12 NI_12 NS_156 0 7.3243253322235026e-03
GC_12_157 b_12 NI_12 NS_157 0 3.8569117359880516e-04
GC_12_158 b_12 NI_12 NS_158 0 -5.4604650668031230e-04
GC_12_159 b_12 NI_12 NS_159 0 5.4856257518595211e-05
GC_12_160 b_12 NI_12 NS_160 0 -1.2298823757739819e-04
GC_12_161 b_12 NI_12 NS_161 0 -2.3024327170735105e-03
GC_12_162 b_12 NI_12 NS_162 0 4.9587851438758638e-03
GC_12_163 b_12 NI_12 NS_163 0 1.3957685499604118e-05
GC_12_164 b_12 NI_12 NS_164 0 3.3806055890689592e-06
GC_12_165 b_12 NI_12 NS_165 0 1.0233691946064549e-02
GC_12_166 b_12 NI_12 NS_166 0 3.6585802624339620e-03
GC_12_167 b_12 NI_12 NS_167 0 5.4704750943985096e-06
GC_12_168 b_12 NI_12 NS_168 0 -7.3520369880879669e-05
GC_12_169 b_12 NI_12 NS_169 0 2.3386192790466898e-06
GC_12_170 b_12 NI_12 NS_170 0 5.4777985307491346e-05
GC_12_171 b_12 NI_12 NS_171 0 -1.5233820805677375e-06
GC_12_172 b_12 NI_12 NS_172 0 -2.2211119628799266e-05
GC_12_173 b_12 NI_12 NS_173 0 -7.1498490860936472e-06
GC_12_174 b_12 NI_12 NS_174 0 -1.1892699893730989e-07
GC_12_175 b_12 NI_12 NS_175 0 -2.9512127474892237e-03
GC_12_176 b_12 NI_12 NS_176 0 9.2747166149726335e-04
GC_12_177 b_12 NI_12 NS_177 0 4.8664963677192475e-05
GC_12_178 b_12 NI_12 NS_178 0 -4.2792125847203267e-04
GC_12_179 b_12 NI_12 NS_179 0 4.7332972900830325e-04
GC_12_180 b_12 NI_12 NS_180 0 1.3517346545459307e-04
GC_12_181 b_12 NI_12 NS_181 0 7.2379933189993873e-05
GC_12_182 b_12 NI_12 NS_182 0 -9.4996586345582097e-05
GC_12_183 b_12 NI_12 NS_183 0 -3.6983196776517167e-05
GC_12_184 b_12 NI_12 NS_184 0 2.9796093852031758e-05
GC_12_185 b_12 NI_12 NS_185 0 -1.3266341366905431e-05
GC_12_186 b_12 NI_12 NS_186 0 -3.7228765631737632e-05
GC_12_187 b_12 NI_12 NS_187 0 -4.8364519770384895e-05
GC_12_188 b_12 NI_12 NS_188 0 -6.2144760198920923e-05
GC_12_189 b_12 NI_12 NS_189 0 -1.4212830254186757e-05
GC_12_190 b_12 NI_12 NS_190 0 -1.2309937077662281e-05
GC_12_191 b_12 NI_12 NS_191 0 -1.4088304669649186e-02
GC_12_192 b_12 NI_12 NS_192 0 -1.0866958898526958e-03
GC_12_193 b_12 NI_12 NS_193 0 1.3249853507821124e-03
GC_12_194 b_12 NI_12 NS_194 0 6.5898160568060443e-03
GC_12_195 b_12 NI_12 NS_195 0 1.1234161350507224e-04
GC_12_196 b_12 NI_12 NS_196 0 -6.0400192500942730e-06
GC_12_197 b_12 NI_12 NS_197 0 3.1672087146299499e-05
GC_12_198 b_12 NI_12 NS_198 0 2.9922287482082545e-05
GC_12_199 b_12 NI_12 NS_199 0 4.1149147959997079e-03
GC_12_200 b_12 NI_12 NS_200 0 -2.8040753210849191e-03
GC_12_201 b_12 NI_12 NS_201 0 -1.4314224980518962e-05
GC_12_202 b_12 NI_12 NS_202 0 -3.3587957084119994e-06
GC_12_203 b_12 NI_12 NS_203 0 8.5415851608764016e-03
GC_12_204 b_12 NI_12 NS_204 0 -4.8281004028392551e-03
GC_12_205 b_12 NI_12 NS_205 0 2.7116288948781598e-05
GC_12_206 b_12 NI_12 NS_206 0 7.1724243176393610e-06
GC_12_207 b_12 NI_12 NS_207 0 2.5055564330296788e-06
GC_12_208 b_12 NI_12 NS_208 0 2.2520586271314222e-05
GC_12_209 b_12 NI_12 NS_209 0 -1.7152534686315369e-05
GC_12_210 b_12 NI_12 NS_210 0 3.5286659907732887e-07
GC_12_211 b_12 NI_12 NS_211 0 6.5611895269879101e-06
GC_12_212 b_12 NI_12 NS_212 0 8.9860183051808890e-07
GC_12_213 b_12 NI_12 NS_213 0 -2.2232034335620218e-03
GC_12_214 b_12 NI_12 NS_214 0 1.7052843549858186e-03
GC_12_215 b_12 NI_12 NS_215 0 -2.2128331011658456e-06
GC_12_216 b_12 NI_12 NS_216 0 -3.1733554249632789e-04
GC_12_217 b_12 NI_12 NS_217 0 3.2575136928568693e-04
GC_12_218 b_12 NI_12 NS_218 0 1.2930472088864498e-04
GC_12_219 b_12 NI_12 NS_219 0 1.0804781745927847e-04
GC_12_220 b_12 NI_12 NS_220 0 -1.4472565870555564e-05
GC_12_221 b_12 NI_12 NS_221 0 -5.1592080369773523e-05
GC_12_222 b_12 NI_12 NS_222 0 -3.5809430872382297e-05
GC_12_223 b_12 NI_12 NS_223 0 2.7366979860232018e-05
GC_12_224 b_12 NI_12 NS_224 0 8.9973384497699922e-06
GC_12_225 b_12 NI_12 NS_225 0 -4.2073923759820138e-05
GC_12_226 b_12 NI_12 NS_226 0 -7.9946031758876206e-05
GC_12_227 b_12 NI_12 NS_227 0 -1.4388678165732527e-06
GC_12_228 b_12 NI_12 NS_228 0 -1.2323670389603531e-05
GC_12_229 b_12 NI_12 NS_229 0 2.5101940825261036e-02
GC_12_230 b_12 NI_12 NS_230 0 1.2306803088253640e-03
GC_12_231 b_12 NI_12 NS_231 0 -1.5319010348000289e-02
GC_12_232 b_12 NI_12 NS_232 0 1.2334705487002913e-03
GC_12_233 b_12 NI_12 NS_233 0 4.0037202462424039e-04
GC_12_234 b_12 NI_12 NS_234 0 -2.5192403282558112e-04
GC_12_235 b_12 NI_12 NS_235 0 -1.1135957935176143e-05
GC_12_236 b_12 NI_12 NS_236 0 -1.9944508875750319e-05
GC_12_237 b_12 NI_12 NS_237 0 -8.2920145035604818e-03
GC_12_238 b_12 NI_12 NS_238 0 -7.8176301452083270e-03
GC_12_239 b_12 NI_12 NS_239 0 2.0757395355752152e-05
GC_12_240 b_12 NI_12 NS_240 0 6.5885413460309340e-06
GC_12_241 b_12 NI_12 NS_241 0 9.6916873840354953e-03
GC_12_242 b_12 NI_12 NS_242 0 1.5048201768907189e-03
GC_12_243 b_12 NI_12 NS_243 0 -3.6974035772841365e-06
GC_12_244 b_12 NI_12 NS_244 0 -4.2165414133699021e-05
GC_12_245 b_12 NI_12 NS_245 0 9.1472481130520652e-06
GC_12_246 b_12 NI_12 NS_246 0 5.0464975181949823e-05
GC_12_247 b_12 NI_12 NS_247 0 -2.3246503880317829e-05
GC_12_248 b_12 NI_12 NS_248 0 -2.5611586815583026e-05
GC_12_249 b_12 NI_12 NS_249 0 -1.4746173154437371e-06
GC_12_250 b_12 NI_12 NS_250 0 -4.7833955845162427e-06
GC_12_251 b_12 NI_12 NS_251 0 -4.4927979944853948e-03
GC_12_252 b_12 NI_12 NS_252 0 5.5514703034557238e-04
GC_12_253 b_12 NI_12 NS_253 0 -1.2389013769969004e-04
GC_12_254 b_12 NI_12 NS_254 0 -2.8585289622000870e-04
GC_12_255 b_12 NI_12 NS_255 0 7.4984684787331158e-04
GC_12_256 b_12 NI_12 NS_256 0 3.7003287543925962e-04
GC_12_257 b_12 NI_12 NS_257 0 2.6737328466704433e-04
GC_12_258 b_12 NI_12 NS_258 0 -3.1089398838066455e-04
GC_12_259 b_12 NI_12 NS_259 0 -7.3772187443221451e-05
GC_12_260 b_12 NI_12 NS_260 0 9.0530301402097635e-06
GC_12_261 b_12 NI_12 NS_261 0 -1.6263784106878825e-05
GC_12_262 b_12 NI_12 NS_262 0 1.7040621495946332e-06
GC_12_263 b_12 NI_12 NS_263 0 -6.9786365033808626e-05
GC_12_264 b_12 NI_12 NS_264 0 1.7595481546145244e-05
GC_12_265 b_12 NI_12 NS_265 0 -4.2035135348020037e-06
GC_12_266 b_12 NI_12 NS_266 0 3.9087288441553234e-06
GC_12_267 b_12 NI_12 NS_267 0 -1.2024290963616036e-02
GC_12_268 b_12 NI_12 NS_268 0 -1.2442110538276882e-03
GC_12_269 b_12 NI_12 NS_269 0 -1.0348783870395126e-03
GC_12_270 b_12 NI_12 NS_270 0 6.3022320988442388e-03
GC_12_271 b_12 NI_12 NS_271 0 -1.0767414905710969e-04
GC_12_272 b_12 NI_12 NS_272 0 1.3149005157559791e-04
GC_12_273 b_12 NI_12 NS_273 0 -1.7618238300344924e-05
GC_12_274 b_12 NI_12 NS_274 0 2.5004625560831346e-05
GC_12_275 b_12 NI_12 NS_275 0 6.4244963775913749e-03
GC_12_276 b_12 NI_12 NS_276 0 5.3972674569762302e-03
GC_12_277 b_12 NI_12 NS_277 0 -2.0900543873148605e-05
GC_12_278 b_12 NI_12 NS_278 0 -9.3292487436721408e-06
GC_12_279 b_12 NI_12 NS_279 0 1.0828363347881459e-02
GC_12_280 b_12 NI_12 NS_280 0 -2.3432337652792594e-03
GC_12_281 b_12 NI_12 NS_281 0 1.4902858605314354e-06
GC_12_282 b_12 NI_12 NS_282 0 2.6190389987764821e-05
GC_12_283 b_12 NI_12 NS_283 0 -2.0213523454190823e-06
GC_12_284 b_12 NI_12 NS_284 0 1.9913327460180961e-05
GC_12_285 b_12 NI_12 NS_285 0 -9.8156709909186419e-06
GC_12_286 b_12 NI_12 NS_286 0 -1.7651127931715003e-05
GC_12_287 b_12 NI_12 NS_287 0 1.2915127865872281e-05
GC_12_288 b_12 NI_12 NS_288 0 -1.9935220034297260e-06
GC_12_289 b_12 NI_12 NS_289 0 -3.7951979825777654e-03
GC_12_290 b_12 NI_12 NS_290 0 7.3353217299771409e-04
GC_12_291 b_12 NI_12 NS_291 0 -5.4170219611830990e-05
GC_12_292 b_12 NI_12 NS_292 0 -2.7771829004707142e-04
GC_12_293 b_12 NI_12 NS_293 0 5.5434861326842462e-04
GC_12_294 b_12 NI_12 NS_294 0 4.3605478596231157e-04
GC_12_295 b_12 NI_12 NS_295 0 3.1508600448481970e-04
GC_12_296 b_12 NI_12 NS_296 0 -1.6637823169661904e-04
GC_12_297 b_12 NI_12 NS_297 0 -5.4558732120559403e-05
GC_12_298 b_12 NI_12 NS_298 0 -6.1811073174402852e-05
GC_12_299 b_12 NI_12 NS_299 0 -5.2606163843478750e-06
GC_12_300 b_12 NI_12 NS_300 0 -2.0218009465938109e-05
GC_12_301 b_12 NI_12 NS_301 0 -6.2970124835074612e-05
GC_12_302 b_12 NI_12 NS_302 0 -3.4757842676726541e-05
GC_12_303 b_12 NI_12 NS_303 0 -7.8835567455566365e-06
GC_12_304 b_12 NI_12 NS_304 0 -7.1411293831639518e-07
GC_12_305 b_12 NI_12 NS_305 0 6.1549451467470942e-02
GC_12_306 b_12 NI_12 NS_306 0 9.5435913655154069e-04
GC_12_307 b_12 NI_12 NS_307 0 -2.6956996408427733e-02
GC_12_308 b_12 NI_12 NS_308 0 -1.2662677667600127e-02
GC_12_309 b_12 NI_12 NS_309 0 4.7154061418605445e-04
GC_12_310 b_12 NI_12 NS_310 0 1.3859687425550179e-04
GC_12_311 b_12 NI_12 NS_311 0 -4.6704500522467127e-05
GC_12_312 b_12 NI_12 NS_312 0 5.6032126540921393e-05
GC_12_313 b_12 NI_12 NS_313 0 -2.4925961546799148e-02
GC_12_314 b_12 NI_12 NS_314 0 -4.3043716941874449e-02
GC_12_315 b_12 NI_12 NS_315 0 1.5385858092046948e-05
GC_12_316 b_12 NI_12 NS_316 0 8.4355774166293057e-05
GC_12_317 b_12 NI_12 NS_317 0 9.2923077572863375e-03
GC_12_318 b_12 NI_12 NS_318 0 -9.1890547795164498e-04
GC_12_319 b_12 NI_12 NS_319 0 -5.7912398526722552e-05
GC_12_320 b_12 NI_12 NS_320 0 1.7616921711044991e-05
GC_12_321 b_12 NI_12 NS_321 0 1.6834984640431453e-06
GC_12_322 b_12 NI_12 NS_322 0 7.7999056826739789e-05
GC_12_323 b_12 NI_12 NS_323 0 -1.2522934373937949e-04
GC_12_324 b_12 NI_12 NS_324 0 -5.0910373111965625e-05
GC_12_325 b_12 NI_12 NS_325 0 -2.6960201685462587e-05
GC_12_326 b_12 NI_12 NS_326 0 -2.7877580355378020e-05
GC_12_327 b_12 NI_12 NS_327 0 -7.0552791417224847e-03
GC_12_328 b_12 NI_12 NS_328 0 3.8063648158357137e-03
GC_12_329 b_12 NI_12 NS_329 0 -7.9176714967057565e-05
GC_12_330 b_12 NI_12 NS_330 0 -3.1444028502902429e-04
GC_12_331 b_12 NI_12 NS_331 0 6.5701089771306976e-04
GC_12_332 b_12 NI_12 NS_332 0 3.8212016663924608e-04
GC_12_333 b_12 NI_12 NS_333 0 2.4395151486950126e-04
GC_12_334 b_12 NI_12 NS_334 0 -1.9373666579693705e-04
GC_12_335 b_12 NI_12 NS_335 0 2.0414292333049289e-05
GC_12_336 b_12 NI_12 NS_336 0 4.4982600911834046e-06
GC_12_337 b_12 NI_12 NS_337 0 4.9452132932785473e-05
GC_12_338 b_12 NI_12 NS_338 0 -9.7884512090600308e-06
GC_12_339 b_12 NI_12 NS_339 0 9.4846921821963336e-06
GC_12_340 b_12 NI_12 NS_340 0 -3.3887524023719954e-05
GC_12_341 b_12 NI_12 NS_341 0 -2.5490564892210598e-06
GC_12_342 b_12 NI_12 NS_342 0 -1.1191832878186759e-05
GC_12_343 b_12 NI_12 NS_343 0 -3.9916585068793123e-03
GC_12_344 b_12 NI_12 NS_344 0 -1.4032278192640131e-03
GC_12_345 b_12 NI_12 NS_345 0 1.2082218267701953e-03
GC_12_346 b_12 NI_12 NS_346 0 -3.5917479803100707e-03
GC_12_347 b_12 NI_12 NS_347 0 -4.1902446852482434e-04
GC_12_348 b_12 NI_12 NS_348 0 5.7188056653865017e-04
GC_12_349 b_12 NI_12 NS_349 0 -5.6538884009705925e-05
GC_12_350 b_12 NI_12 NS_350 0 1.0475821578036266e-04
GC_12_351 b_12 NI_12 NS_351 0 7.7238301850074765e-03
GC_12_352 b_12 NI_12 NS_352 0 2.3103306775711829e-02
GC_12_353 b_12 NI_12 NS_353 0 -2.6970885334208828e-05
GC_12_354 b_12 NI_12 NS_354 0 -8.4231024255522721e-05
GC_12_355 b_12 NI_12 NS_355 0 4.9534010180389493e-03
GC_12_356 b_12 NI_12 NS_356 0 -3.6206886090693426e-03
GC_12_357 b_12 NI_12 NS_357 0 -4.2870548797579085e-05
GC_12_358 b_12 NI_12 NS_358 0 5.8575512772678242e-05
GC_12_359 b_12 NI_12 NS_359 0 -2.6276023128607194e-05
GC_12_360 b_12 NI_12 NS_360 0 5.8113573800104901e-05
GC_12_361 b_12 NI_12 NS_361 0 -8.0537824774178972e-05
GC_12_362 b_12 NI_12 NS_362 0 -2.7887847570776732e-05
GC_12_363 b_12 NI_12 NS_363 0 -2.1091288334360743e-05
GC_12_364 b_12 NI_12 NS_364 0 -3.1106430432040301e-05
GC_12_365 b_12 NI_12 NS_365 0 -5.5315695579933408e-03
GC_12_366 b_12 NI_12 NS_366 0 3.7854277310765553e-03
GC_12_367 b_12 NI_12 NS_367 0 7.4435053720349988e-05
GC_12_368 b_12 NI_12 NS_368 0 -3.2470451702593811e-04
GC_12_369 b_12 NI_12 NS_369 0 5.1445409462628621e-04
GC_12_370 b_12 NI_12 NS_370 0 2.6683517591263124e-04
GC_12_371 b_12 NI_12 NS_371 0 2.4741697273722907e-04
GC_12_372 b_12 NI_12 NS_372 0 -1.4104963968017067e-04
GC_12_373 b_12 NI_12 NS_373 0 1.7318431456874249e-05
GC_12_374 b_12 NI_12 NS_374 0 3.3422048819287838e-05
GC_12_375 b_12 NI_12 NS_375 0 4.1578134612994011e-05
GC_12_376 b_12 NI_12 NS_376 0 -2.5194692290109258e-05
GC_12_377 b_12 NI_12 NS_377 0 -1.6420324710283742e-05
GC_12_378 b_12 NI_12 NS_378 0 -1.2561684208362316e-05
GC_12_379 b_12 NI_12 NS_379 0 -1.0595135737760303e-05
GC_12_380 b_12 NI_12 NS_380 0 -1.1810554843928240e-05
GC_12_381 b_12 NI_12 NS_381 0 1.9324914772620161e-02
GC_12_382 b_12 NI_12 NS_382 0 1.8259581239176840e-03
GC_12_383 b_12 NI_12 NS_383 0 2.4610014218715982e-02
GC_12_384 b_12 NI_12 NS_384 0 -1.6224792397864018e-02
GC_12_385 b_12 NI_12 NS_385 0 1.2917387942377237e-03
GC_12_386 b_12 NI_12 NS_386 0 6.9499816279832796e-05
GC_12_387 b_12 NI_12 NS_387 0 1.4152682802604328e-05
GC_12_388 b_12 NI_12 NS_388 0 3.4002850615308249e-05
GC_12_389 b_12 NI_12 NS_389 0 2.6070867504164236e-02
GC_12_390 b_12 NI_12 NS_390 0 2.4076294161360216e-03
GC_12_391 b_12 NI_12 NS_391 0 4.0640778335563702e-05
GC_12_392 b_12 NI_12 NS_392 0 8.6258519797654843e-05
GC_12_393 b_12 NI_12 NS_393 0 -4.5704197166866946e-02
GC_12_394 b_12 NI_12 NS_394 0 3.2071294129808810e-02
GC_12_395 b_12 NI_12 NS_395 0 -3.9746822267682283e-05
GC_12_396 b_12 NI_12 NS_396 0 8.1759322601852744e-05
GC_12_397 b_12 NI_12 NS_397 0 5.0753236232348428e-05
GC_12_398 b_12 NI_12 NS_398 0 1.6308559567710754e-05
GC_12_399 b_12 NI_12 NS_399 0 -1.2946861140450015e-04
GC_12_400 b_12 NI_12 NS_400 0 -3.4899623416817219e-05
GC_12_401 b_12 NI_12 NS_401 0 -2.0618545807178833e-05
GC_12_402 b_12 NI_12 NS_402 0 -1.5588196153313841e-05
GC_12_403 b_12 NI_12 NS_403 0 -4.0752824822775638e-03
GC_12_404 b_12 NI_12 NS_404 0 3.0864237097900427e-04
GC_12_405 b_12 NI_12 NS_405 0 -1.2734555558199060e-04
GC_12_406 b_12 NI_12 NS_406 0 6.9394917361303057e-05
GC_12_407 b_12 NI_12 NS_407 0 8.2501262153308126e-04
GC_12_408 b_12 NI_12 NS_408 0 6.2738303929307717e-04
GC_12_409 b_12 NI_12 NS_409 0 3.2408995017440466e-04
GC_12_410 b_12 NI_12 NS_410 0 -3.6391699203389653e-04
GC_12_411 b_12 NI_12 NS_411 0 1.4130494843646817e-04
GC_12_412 b_12 NI_12 NS_412 0 1.9597813940017679e-05
GC_12_413 b_12 NI_12 NS_413 0 8.5960245584447117e-05
GC_12_414 b_12 NI_12 NS_414 0 -8.1240769707845320e-06
GC_12_415 b_12 NI_12 NS_415 0 3.7363303006013260e-05
GC_12_416 b_12 NI_12 NS_416 0 7.7182493250622659e-05
GC_12_417 b_12 NI_12 NS_417 0 1.2980610408085520e-05
GC_12_418 b_12 NI_12 NS_418 0 -1.2819596620948699e-05
GC_12_419 b_12 NI_12 NS_419 0 5.3135767835832931e-02
GC_12_420 b_12 NI_12 NS_420 0 -1.3729443511873722e-03
GC_12_421 b_12 NI_12 NS_421 0 4.7404299234929642e-02
GC_12_422 b_12 NI_12 NS_422 0 -5.7877658332268725e-02
GC_12_423 b_12 NI_12 NS_423 0 -9.1869523162396781e-04
GC_12_424 b_12 NI_12 NS_424 0 1.5787934982705541e-04
GC_12_425 b_12 NI_12 NS_425 0 -8.8526087329860939e-05
GC_12_426 b_12 NI_12 NS_426 0 1.0837687541784398e-04
GC_12_427 b_12 NI_12 NS_427 0 -1.0387345511389210e-02
GC_12_428 b_12 NI_12 NS_428 0 1.4918761185154564e-02
GC_12_429 b_12 NI_12 NS_429 0 -2.4057386879081404e-05
GC_12_430 b_12 NI_12 NS_430 0 -7.8548462980428728e-05
GC_12_431 b_12 NI_12 NS_431 0 -3.1560782781964808e-02
GC_12_432 b_12 NI_12 NS_432 0 4.8383278051938828e-03
GC_12_433 b_12 NI_12 NS_433 0 -8.0460533701025863e-05
GC_12_434 b_12 NI_12 NS_434 0 1.0420417377853900e-04
GC_12_435 b_12 NI_12 NS_435 0 5.3551215992539158e-06
GC_12_436 b_12 NI_12 NS_436 0 3.1411642922183388e-05
GC_12_437 b_12 NI_12 NS_437 0 -9.0109998802105206e-05
GC_12_438 b_12 NI_12 NS_438 0 -3.8765404488954239e-05
GC_12_439 b_12 NI_12 NS_439 0 -1.6414935739687740e-05
GC_12_440 b_12 NI_12 NS_440 0 -2.5460862599559124e-05
GC_12_441 b_12 NI_12 NS_441 0 -5.6806829920272002e-03
GC_12_442 b_12 NI_12 NS_442 0 3.3226943144100182e-03
GC_12_443 b_12 NI_12 NS_443 0 8.8009377890074332e-06
GC_12_444 b_12 NI_12 NS_444 0 -2.0378112899052271e-04
GC_12_445 b_12 NI_12 NS_445 0 7.4352201691413702e-04
GC_12_446 b_12 NI_12 NS_446 0 5.9674241151683584e-04
GC_12_447 b_12 NI_12 NS_447 0 4.2413489842206775e-04
GC_12_448 b_12 NI_12 NS_448 0 -2.6297856694334007e-04
GC_12_449 b_12 NI_12 NS_449 0 8.2983135877598725e-05
GC_12_450 b_12 NI_12 NS_450 0 9.8516678845932134e-05
GC_12_451 b_12 NI_12 NS_451 0 8.7320007672957766e-05
GC_12_452 b_12 NI_12 NS_452 0 8.9209413373004594e-06
GC_12_453 b_12 NI_12 NS_453 0 1.6387352154161776e-05
GC_12_454 b_12 NI_12 NS_454 0 4.8391450927281000e-05
GC_12_455 b_12 NI_12 NS_455 0 2.7586089354142148e-06
GC_12_456 b_12 NI_12 NS_456 0 -1.2518199609393377e-05
GD_12_1 b_12 NI_12 NA_1 0 1.1841352763398796e-03
GD_12_2 b_12 NI_12 NA_2 0 2.7985605476178423e-04
GD_12_3 b_12 NI_12 NA_3 0 -2.6553130234307043e-03
GD_12_4 b_12 NI_12 NA_4 0 -3.7050037427891320e-03
GD_12_5 b_12 NI_12 NA_5 0 -1.0633092857226828e-02
GD_12_6 b_12 NI_12 NA_6 0 1.9761535138168728e-03
GD_12_7 b_12 NI_12 NA_7 0 -7.8441362722564134e-03
GD_12_8 b_12 NI_12 NA_8 0 1.9484509102620680e-04
GD_12_9 b_12 NI_12 NA_9 0 -1.0316605182123047e-02
GD_12_10 b_12 NI_12 NA_10 0 1.4511168839527399e-03
GD_12_11 b_12 NI_12 NA_11 0 -3.3054995099955499e-02
GD_12_12 b_12 NI_12 NA_12 0 -1.1846587620059205e-01
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 3.4413071814985372e+00
GS_1_1 0 NS_1 NA_1 0 1.0694336352474016e+00
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 3.0797075048869470e+01
GS_2_1 0 NS_2 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 3/4
CS_3 NS_3 0 9.9999999999999998e-13
CS_4 NS_4 0 9.9999999999999998e-13
RS_3 NS_3 0 8.9335977936087705e+00
RS_4 NS_4 0 8.9335977936087705e+00
GL_3 0 NS_3 NS_4 0 2.2441700641819512e-01
GL_4 0 NS_4 NS_3 0 -2.2441700641819512e-01
GS_3_1 0 NS_3 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 5.9158463852536897e+01
RS_6 NS_6 0 5.9158463852536897e+01
GL_5 0 NS_5 NS_6 0 2.6680991281534006e-01
GL_6 0 NS_6 NS_5 0 -2.6680991281534006e-01
GS_5_1 0 NS_5 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 9.2065834236318878e+01
RS_8 NS_8 0 9.2065834236318864e+01
GL_7 0 NS_7 NS_8 0 2.4567219632280338e-01
GL_8 0 NS_8 NS_7 0 -2.4567219632280338e-01
GS_7_1 0 NS_7 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 1.4764174191595519e+01
RS_10 NS_10 0 1.4764174191595517e+01
GL_9 0 NS_9 NS_10 0 1.4400577194218670e-02
GL_10 0 NS_10 NS_9 0 -1.4400577194218670e-02
GS_9_1 0 NS_9 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 9.7834937041354195e+01
RS_12 NS_12 0 9.7834937041354195e+01
GL_11 0 NS_11 NS_12 0 6.3371310235267833e-02
GL_12 0 NS_12 NS_11 0 -6.3371310235267833e-02
GS_11_1 0 NS_11 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 1.4785099744646029e+01
RS_14 NS_14 0 1.4785099744646031e+01
GL_13 0 NS_13 NS_14 0 1.5607347485362127e-01
GL_14 0 NS_14 NS_13 0 -1.5607347485362127e-01
GS_13_1 0 NS_13 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 1.3466736941644649e+02
RS_16 NS_16 0 1.3466736941644649e+02
GL_15 0 NS_15 NS_16 0 2.3468192685328568e-01
GL_16 0 NS_16 NS_15 0 -2.3468192685328568e-01
GS_15_1 0 NS_15 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 1.5102368550954495e+02
RS_18 NS_18 0 1.5102368550954495e+02
GL_17 0 NS_17 NS_18 0 2.2562219216120838e-01
GL_18 0 NS_18 NS_17 0 -2.2562219216120838e-01
GS_17_1 0 NS_17 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 1.6979945400908466e+02
RS_20 NS_20 0 1.6979945400908468e+02
GL_19 0 NS_19 NS_20 0 2.1538055438627146e-01
GL_20 0 NS_20 NS_19 0 -2.1538055438627146e-01
GS_19_1 0 NS_19 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 2.2834543421620666e+02
RS_22 NS_22 0 2.2834543421620666e+02
GL_21 0 NS_21 NS_22 0 2.0391309107915187e-01
GL_22 0 NS_22 NS_21 0 -2.0391309107915187e-01
GS_21_1 0 NS_21 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 3.4087022095623759e+01
RS_24 NS_24 0 3.4087022095623759e+01
GL_23 0 NS_23 NS_24 0 1.5530350392230499e-01
GL_24 0 NS_24 NS_23 0 -1.5530350392230499e-01
GS_23_1 0 NS_23 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 7.5761470378414444e+01
RS_26 NS_26 0 7.5761470378414444e+01
GL_25 0 NS_25 NS_26 0 1.6902428843873585e-01
GL_26 0 NS_26 NS_25 0 -1.6902428843873585e-01
GS_25_1 0 NS_25 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 1.1061014882057984e+02
RS_28 NS_28 0 1.1061014882057984e+02
GL_27 0 NS_27 NS_28 0 1.5628591857280719e-01
GL_28 0 NS_28 NS_27 0 -1.5628591857280719e-01
GS_27_1 0 NS_27 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 1.9636019836512071e+02
RS_30 NS_30 0 1.9636019836512071e+02
GL_29 0 NS_29 NS_30 0 1.5213319862255134e-01
GL_30 0 NS_30 NS_29 0 -1.5213319862255134e-01
GS_29_1 0 NS_29 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 4.3243187986905582e+02
RS_32 NS_32 0 4.3243187986905582e+02
GL_31 0 NS_31 NS_32 0 1.3841574306468743e-01
GL_32 0 NS_32 NS_31 0 -1.3841574306468743e-01
GS_31_1 0 NS_31 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 3.6825571251433115e+02
RS_34 NS_34 0 3.6825571251433115e+02
GL_33 0 NS_33 NS_34 0 1.3950469341450047e-01
GL_34 0 NS_34 NS_33 0 -1.3950469341450047e-01
GS_33_1 0 NS_33 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 3.0711053107765838e+02
RS_36 NS_36 0 3.0711053107765838e+02
GL_35 0 NS_35 NS_36 0 1.4553496077846845e-01
GL_36 0 NS_36 NS_35 0 -1.4553496077846845e-01
GS_35_1 0 NS_35 NA_1 0 1.0694336352474016e+00
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 4.6727671488342185e+02
RS_38 NS_38 0 4.6727671488342185e+02
GL_37 0 NS_37 NS_38 0 1.4422859584763473e-01
GL_38 0 NS_38 NS_37 0 -1.4422859584763473e-01
GS_37_1 0 NS_37 NA_1 0 1.0694336352474016e+00
*
* Real pole n. 39
CS_39 NS_39 0 9.9999999999999998e-13
RS_39 NS_39 0 3.4413071814985372e+00
GS_39_2 0 NS_39 NA_2 0 1.0694336352474016e+00
*
* Real pole n. 40
CS_40 NS_40 0 9.9999999999999998e-13
RS_40 NS_40 0 3.0797075048869470e+01
GS_40_2 0 NS_40 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 8.9335977936087705e+00
RS_42 NS_42 0 8.9335977936087705e+00
GL_41 0 NS_41 NS_42 0 2.2441700641819512e-01
GL_42 0 NS_42 NS_41 0 -2.2441700641819512e-01
GS_41_2 0 NS_41 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 5.9158463852536897e+01
RS_44 NS_44 0 5.9158463852536897e+01
GL_43 0 NS_43 NS_44 0 2.6680991281534006e-01
GL_44 0 NS_44 NS_43 0 -2.6680991281534006e-01
GS_43_2 0 NS_43 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 45/46
CS_45 NS_45 0 9.9999999999999998e-13
CS_46 NS_46 0 9.9999999999999998e-13
RS_45 NS_45 0 9.2065834236318878e+01
RS_46 NS_46 0 9.2065834236318864e+01
GL_45 0 NS_45 NS_46 0 2.4567219632280338e-01
GL_46 0 NS_46 NS_45 0 -2.4567219632280338e-01
GS_45_2 0 NS_45 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 1.4764174191595519e+01
RS_48 NS_48 0 1.4764174191595517e+01
GL_47 0 NS_47 NS_48 0 1.4400577194218670e-02
GL_48 0 NS_48 NS_47 0 -1.4400577194218670e-02
GS_47_2 0 NS_47 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 9.7834937041354195e+01
RS_50 NS_50 0 9.7834937041354195e+01
GL_49 0 NS_49 NS_50 0 6.3371310235267833e-02
GL_50 0 NS_50 NS_49 0 -6.3371310235267833e-02
GS_49_2 0 NS_49 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 1.4785099744646029e+01
RS_52 NS_52 0 1.4785099744646031e+01
GL_51 0 NS_51 NS_52 0 1.5607347485362127e-01
GL_52 0 NS_52 NS_51 0 -1.5607347485362127e-01
GS_51_2 0 NS_51 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 1.3466736941644649e+02
RS_54 NS_54 0 1.3466736941644649e+02
GL_53 0 NS_53 NS_54 0 2.3468192685328568e-01
GL_54 0 NS_54 NS_53 0 -2.3468192685328568e-01
GS_53_2 0 NS_53 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 1.5102368550954495e+02
RS_56 NS_56 0 1.5102368550954495e+02
GL_55 0 NS_55 NS_56 0 2.2562219216120838e-01
GL_56 0 NS_56 NS_55 0 -2.2562219216120838e-01
GS_55_2 0 NS_55 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 1.6979945400908466e+02
RS_58 NS_58 0 1.6979945400908468e+02
GL_57 0 NS_57 NS_58 0 2.1538055438627146e-01
GL_58 0 NS_58 NS_57 0 -2.1538055438627146e-01
GS_57_2 0 NS_57 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 2.2834543421620666e+02
RS_60 NS_60 0 2.2834543421620666e+02
GL_59 0 NS_59 NS_60 0 2.0391309107915187e-01
GL_60 0 NS_60 NS_59 0 -2.0391309107915187e-01
GS_59_2 0 NS_59 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 3.4087022095623759e+01
RS_62 NS_62 0 3.4087022095623759e+01
GL_61 0 NS_61 NS_62 0 1.5530350392230499e-01
GL_62 0 NS_62 NS_61 0 -1.5530350392230499e-01
GS_61_2 0 NS_61 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 7.5761470378414444e+01
RS_64 NS_64 0 7.5761470378414444e+01
GL_63 0 NS_63 NS_64 0 1.6902428843873585e-01
GL_64 0 NS_64 NS_63 0 -1.6902428843873585e-01
GS_63_2 0 NS_63 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 1.1061014882057984e+02
RS_66 NS_66 0 1.1061014882057984e+02
GL_65 0 NS_65 NS_66 0 1.5628591857280719e-01
GL_66 0 NS_66 NS_65 0 -1.5628591857280719e-01
GS_65_2 0 NS_65 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 1.9636019836512071e+02
RS_68 NS_68 0 1.9636019836512071e+02
GL_67 0 NS_67 NS_68 0 1.5213319862255134e-01
GL_68 0 NS_68 NS_67 0 -1.5213319862255134e-01
GS_67_2 0 NS_67 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 4.3243187986905582e+02
RS_70 NS_70 0 4.3243187986905582e+02
GL_69 0 NS_69 NS_70 0 1.3841574306468743e-01
GL_70 0 NS_70 NS_69 0 -1.3841574306468743e-01
GS_69_2 0 NS_69 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 3.6825571251433115e+02
RS_72 NS_72 0 3.6825571251433115e+02
GL_71 0 NS_71 NS_72 0 1.3950469341450047e-01
GL_72 0 NS_72 NS_71 0 -1.3950469341450047e-01
GS_71_2 0 NS_71 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 3.0711053107765838e+02
RS_74 NS_74 0 3.0711053107765838e+02
GL_73 0 NS_73 NS_74 0 1.4553496077846845e-01
GL_74 0 NS_74 NS_73 0 -1.4553496077846845e-01
GS_73_2 0 NS_73 NA_2 0 1.0694336352474016e+00
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 4.6727671488342185e+02
RS_76 NS_76 0 4.6727671488342185e+02
GL_75 0 NS_75 NS_76 0 1.4422859584763473e-01
GL_76 0 NS_76 NS_75 0 -1.4422859584763473e-01
GS_75_2 0 NS_75 NA_2 0 1.0694336352474016e+00
*
* Real pole n. 77
CS_77 NS_77 0 9.9999999999999998e-13
RS_77 NS_77 0 3.4413071814985372e+00
GS_77_3 0 NS_77 NA_3 0 1.0694336352474016e+00
*
* Real pole n. 78
CS_78 NS_78 0 9.9999999999999998e-13
RS_78 NS_78 0 3.0797075048869470e+01
GS_78_3 0 NS_78 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 8.9335977936087705e+00
RS_80 NS_80 0 8.9335977936087705e+00
GL_79 0 NS_79 NS_80 0 2.2441700641819512e-01
GL_80 0 NS_80 NS_79 0 -2.2441700641819512e-01
GS_79_3 0 NS_79 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 5.9158463852536897e+01
RS_82 NS_82 0 5.9158463852536897e+01
GL_81 0 NS_81 NS_82 0 2.6680991281534006e-01
GL_82 0 NS_82 NS_81 0 -2.6680991281534006e-01
GS_81_3 0 NS_81 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 9.2065834236318878e+01
RS_84 NS_84 0 9.2065834236318864e+01
GL_83 0 NS_83 NS_84 0 2.4567219632280338e-01
GL_84 0 NS_84 NS_83 0 -2.4567219632280338e-01
GS_83_3 0 NS_83 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 1.4764174191595519e+01
RS_86 NS_86 0 1.4764174191595517e+01
GL_85 0 NS_85 NS_86 0 1.4400577194218670e-02
GL_86 0 NS_86 NS_85 0 -1.4400577194218670e-02
GS_85_3 0 NS_85 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 9.7834937041354195e+01
RS_88 NS_88 0 9.7834937041354195e+01
GL_87 0 NS_87 NS_88 0 6.3371310235267833e-02
GL_88 0 NS_88 NS_87 0 -6.3371310235267833e-02
GS_87_3 0 NS_87 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 89/90
CS_89 NS_89 0 9.9999999999999998e-13
CS_90 NS_90 0 9.9999999999999998e-13
RS_89 NS_89 0 1.4785099744646029e+01
RS_90 NS_90 0 1.4785099744646031e+01
GL_89 0 NS_89 NS_90 0 1.5607347485362127e-01
GL_90 0 NS_90 NS_89 0 -1.5607347485362127e-01
GS_89_3 0 NS_89 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 1.3466736941644649e+02
RS_92 NS_92 0 1.3466736941644649e+02
GL_91 0 NS_91 NS_92 0 2.3468192685328568e-01
GL_92 0 NS_92 NS_91 0 -2.3468192685328568e-01
GS_91_3 0 NS_91 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 1.5102368550954495e+02
RS_94 NS_94 0 1.5102368550954495e+02
GL_93 0 NS_93 NS_94 0 2.2562219216120838e-01
GL_94 0 NS_94 NS_93 0 -2.2562219216120838e-01
GS_93_3 0 NS_93 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 1.6979945400908466e+02
RS_96 NS_96 0 1.6979945400908468e+02
GL_95 0 NS_95 NS_96 0 2.1538055438627146e-01
GL_96 0 NS_96 NS_95 0 -2.1538055438627146e-01
GS_95_3 0 NS_95 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 2.2834543421620666e+02
RS_98 NS_98 0 2.2834543421620666e+02
GL_97 0 NS_97 NS_98 0 2.0391309107915187e-01
GL_98 0 NS_98 NS_97 0 -2.0391309107915187e-01
GS_97_3 0 NS_97 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 3.4087022095623759e+01
RS_100 NS_100 0 3.4087022095623759e+01
GL_99 0 NS_99 NS_100 0 1.5530350392230499e-01
GL_100 0 NS_100 NS_99 0 -1.5530350392230499e-01
GS_99_3 0 NS_99 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 7.5761470378414444e+01
RS_102 NS_102 0 7.5761470378414444e+01
GL_101 0 NS_101 NS_102 0 1.6902428843873585e-01
GL_102 0 NS_102 NS_101 0 -1.6902428843873585e-01
GS_101_3 0 NS_101 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 1.1061014882057984e+02
RS_104 NS_104 0 1.1061014882057984e+02
GL_103 0 NS_103 NS_104 0 1.5628591857280719e-01
GL_104 0 NS_104 NS_103 0 -1.5628591857280719e-01
GS_103_3 0 NS_103 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 1.9636019836512071e+02
RS_106 NS_106 0 1.9636019836512071e+02
GL_105 0 NS_105 NS_106 0 1.5213319862255134e-01
GL_106 0 NS_106 NS_105 0 -1.5213319862255134e-01
GS_105_3 0 NS_105 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 4.3243187986905582e+02
RS_108 NS_108 0 4.3243187986905582e+02
GL_107 0 NS_107 NS_108 0 1.3841574306468743e-01
GL_108 0 NS_108 NS_107 0 -1.3841574306468743e-01
GS_107_3 0 NS_107 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 3.6825571251433115e+02
RS_110 NS_110 0 3.6825571251433115e+02
GL_109 0 NS_109 NS_110 0 1.3950469341450047e-01
GL_110 0 NS_110 NS_109 0 -1.3950469341450047e-01
GS_109_3 0 NS_109 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 3.0711053107765838e+02
RS_112 NS_112 0 3.0711053107765838e+02
GL_111 0 NS_111 NS_112 0 1.4553496077846845e-01
GL_112 0 NS_112 NS_111 0 -1.4553496077846845e-01
GS_111_3 0 NS_111 NA_3 0 1.0694336352474016e+00
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 4.6727671488342185e+02
RS_114 NS_114 0 4.6727671488342185e+02
GL_113 0 NS_113 NS_114 0 1.4422859584763473e-01
GL_114 0 NS_114 NS_113 0 -1.4422859584763473e-01
GS_113_3 0 NS_113 NA_3 0 1.0694336352474016e+00
*
* Real pole n. 115
CS_115 NS_115 0 9.9999999999999998e-13
RS_115 NS_115 0 3.4413071814985372e+00
GS_115_4 0 NS_115 NA_4 0 1.0694336352474016e+00
*
* Real pole n. 116
CS_116 NS_116 0 9.9999999999999998e-13
RS_116 NS_116 0 3.0797075048869470e+01
GS_116_4 0 NS_116 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 8.9335977936087705e+00
RS_118 NS_118 0 8.9335977936087705e+00
GL_117 0 NS_117 NS_118 0 2.2441700641819512e-01
GL_118 0 NS_118 NS_117 0 -2.2441700641819512e-01
GS_117_4 0 NS_117 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 5.9158463852536897e+01
RS_120 NS_120 0 5.9158463852536897e+01
GL_119 0 NS_119 NS_120 0 2.6680991281534006e-01
GL_120 0 NS_120 NS_119 0 -2.6680991281534006e-01
GS_119_4 0 NS_119 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 9.2065834236318878e+01
RS_122 NS_122 0 9.2065834236318864e+01
GL_121 0 NS_121 NS_122 0 2.4567219632280338e-01
GL_122 0 NS_122 NS_121 0 -2.4567219632280338e-01
GS_121_4 0 NS_121 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 1.4764174191595519e+01
RS_124 NS_124 0 1.4764174191595517e+01
GL_123 0 NS_123 NS_124 0 1.4400577194218670e-02
GL_124 0 NS_124 NS_123 0 -1.4400577194218670e-02
GS_123_4 0 NS_123 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 9.7834937041354195e+01
RS_126 NS_126 0 9.7834937041354195e+01
GL_125 0 NS_125 NS_126 0 6.3371310235267833e-02
GL_126 0 NS_126 NS_125 0 -6.3371310235267833e-02
GS_125_4 0 NS_125 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 1.4785099744646029e+01
RS_128 NS_128 0 1.4785099744646031e+01
GL_127 0 NS_127 NS_128 0 1.5607347485362127e-01
GL_128 0 NS_128 NS_127 0 -1.5607347485362127e-01
GS_127_4 0 NS_127 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 1.3466736941644649e+02
RS_130 NS_130 0 1.3466736941644649e+02
GL_129 0 NS_129 NS_130 0 2.3468192685328568e-01
GL_130 0 NS_130 NS_129 0 -2.3468192685328568e-01
GS_129_4 0 NS_129 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 1.5102368550954495e+02
RS_132 NS_132 0 1.5102368550954495e+02
GL_131 0 NS_131 NS_132 0 2.2562219216120838e-01
GL_132 0 NS_132 NS_131 0 -2.2562219216120838e-01
GS_131_4 0 NS_131 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 133/134
CS_133 NS_133 0 9.9999999999999998e-13
CS_134 NS_134 0 9.9999999999999998e-13
RS_133 NS_133 0 1.6979945400908466e+02
RS_134 NS_134 0 1.6979945400908468e+02
GL_133 0 NS_133 NS_134 0 2.1538055438627146e-01
GL_134 0 NS_134 NS_133 0 -2.1538055438627146e-01
GS_133_4 0 NS_133 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 2.2834543421620666e+02
RS_136 NS_136 0 2.2834543421620666e+02
GL_135 0 NS_135 NS_136 0 2.0391309107915187e-01
GL_136 0 NS_136 NS_135 0 -2.0391309107915187e-01
GS_135_4 0 NS_135 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 3.4087022095623759e+01
RS_138 NS_138 0 3.4087022095623759e+01
GL_137 0 NS_137 NS_138 0 1.5530350392230499e-01
GL_138 0 NS_138 NS_137 0 -1.5530350392230499e-01
GS_137_4 0 NS_137 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 7.5761470378414444e+01
RS_140 NS_140 0 7.5761470378414444e+01
GL_139 0 NS_139 NS_140 0 1.6902428843873585e-01
GL_140 0 NS_140 NS_139 0 -1.6902428843873585e-01
GS_139_4 0 NS_139 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 1.1061014882057984e+02
RS_142 NS_142 0 1.1061014882057984e+02
GL_141 0 NS_141 NS_142 0 1.5628591857280719e-01
GL_142 0 NS_142 NS_141 0 -1.5628591857280719e-01
GS_141_4 0 NS_141 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 1.9636019836512071e+02
RS_144 NS_144 0 1.9636019836512071e+02
GL_143 0 NS_143 NS_144 0 1.5213319862255134e-01
GL_144 0 NS_144 NS_143 0 -1.5213319862255134e-01
GS_143_4 0 NS_143 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 4.3243187986905582e+02
RS_146 NS_146 0 4.3243187986905582e+02
GL_145 0 NS_145 NS_146 0 1.3841574306468743e-01
GL_146 0 NS_146 NS_145 0 -1.3841574306468743e-01
GS_145_4 0 NS_145 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 3.6825571251433115e+02
RS_148 NS_148 0 3.6825571251433115e+02
GL_147 0 NS_147 NS_148 0 1.3950469341450047e-01
GL_148 0 NS_148 NS_147 0 -1.3950469341450047e-01
GS_147_4 0 NS_147 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 3.0711053107765838e+02
RS_150 NS_150 0 3.0711053107765838e+02
GL_149 0 NS_149 NS_150 0 1.4553496077846845e-01
GL_150 0 NS_150 NS_149 0 -1.4553496077846845e-01
GS_149_4 0 NS_149 NA_4 0 1.0694336352474016e+00
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 4.6727671488342185e+02
RS_152 NS_152 0 4.6727671488342185e+02
GL_151 0 NS_151 NS_152 0 1.4422859584763473e-01
GL_152 0 NS_152 NS_151 0 -1.4422859584763473e-01
GS_151_4 0 NS_151 NA_4 0 1.0694336352474016e+00
*
* Real pole n. 153
CS_153 NS_153 0 9.9999999999999998e-13
RS_153 NS_153 0 3.4413071814985372e+00
GS_153_5 0 NS_153 NA_5 0 1.0694336352474016e+00
*
* Real pole n. 154
CS_154 NS_154 0 9.9999999999999998e-13
RS_154 NS_154 0 3.0797075048869470e+01
GS_154_5 0 NS_154 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 8.9335977936087705e+00
RS_156 NS_156 0 8.9335977936087705e+00
GL_155 0 NS_155 NS_156 0 2.2441700641819512e-01
GL_156 0 NS_156 NS_155 0 -2.2441700641819512e-01
GS_155_5 0 NS_155 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 5.9158463852536897e+01
RS_158 NS_158 0 5.9158463852536897e+01
GL_157 0 NS_157 NS_158 0 2.6680991281534006e-01
GL_158 0 NS_158 NS_157 0 -2.6680991281534006e-01
GS_157_5 0 NS_157 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 9.2065834236318878e+01
RS_160 NS_160 0 9.2065834236318864e+01
GL_159 0 NS_159 NS_160 0 2.4567219632280338e-01
GL_160 0 NS_160 NS_159 0 -2.4567219632280338e-01
GS_159_5 0 NS_159 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 1.4764174191595519e+01
RS_162 NS_162 0 1.4764174191595517e+01
GL_161 0 NS_161 NS_162 0 1.4400577194218670e-02
GL_162 0 NS_162 NS_161 0 -1.4400577194218670e-02
GS_161_5 0 NS_161 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 163/164
CS_163 NS_163 0 9.9999999999999998e-13
CS_164 NS_164 0 9.9999999999999998e-13
RS_163 NS_163 0 9.7834937041354195e+01
RS_164 NS_164 0 9.7834937041354195e+01
GL_163 0 NS_163 NS_164 0 6.3371310235267833e-02
GL_164 0 NS_164 NS_163 0 -6.3371310235267833e-02
GS_163_5 0 NS_163 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 1.4785099744646029e+01
RS_166 NS_166 0 1.4785099744646031e+01
GL_165 0 NS_165 NS_166 0 1.5607347485362127e-01
GL_166 0 NS_166 NS_165 0 -1.5607347485362127e-01
GS_165_5 0 NS_165 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 1.3466736941644649e+02
RS_168 NS_168 0 1.3466736941644649e+02
GL_167 0 NS_167 NS_168 0 2.3468192685328568e-01
GL_168 0 NS_168 NS_167 0 -2.3468192685328568e-01
GS_167_5 0 NS_167 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 1.5102368550954495e+02
RS_170 NS_170 0 1.5102368550954495e+02
GL_169 0 NS_169 NS_170 0 2.2562219216120838e-01
GL_170 0 NS_170 NS_169 0 -2.2562219216120838e-01
GS_169_5 0 NS_169 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 1.6979945400908466e+02
RS_172 NS_172 0 1.6979945400908468e+02
GL_171 0 NS_171 NS_172 0 2.1538055438627146e-01
GL_172 0 NS_172 NS_171 0 -2.1538055438627146e-01
GS_171_5 0 NS_171 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 2.2834543421620666e+02
RS_174 NS_174 0 2.2834543421620666e+02
GL_173 0 NS_173 NS_174 0 2.0391309107915187e-01
GL_174 0 NS_174 NS_173 0 -2.0391309107915187e-01
GS_173_5 0 NS_173 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 3.4087022095623759e+01
RS_176 NS_176 0 3.4087022095623759e+01
GL_175 0 NS_175 NS_176 0 1.5530350392230499e-01
GL_176 0 NS_176 NS_175 0 -1.5530350392230499e-01
GS_175_5 0 NS_175 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 177/178
CS_177 NS_177 0 9.9999999999999998e-13
CS_178 NS_178 0 9.9999999999999998e-13
RS_177 NS_177 0 7.5761470378414444e+01
RS_178 NS_178 0 7.5761470378414444e+01
GL_177 0 NS_177 NS_178 0 1.6902428843873585e-01
GL_178 0 NS_178 NS_177 0 -1.6902428843873585e-01
GS_177_5 0 NS_177 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 1.1061014882057984e+02
RS_180 NS_180 0 1.1061014882057984e+02
GL_179 0 NS_179 NS_180 0 1.5628591857280719e-01
GL_180 0 NS_180 NS_179 0 -1.5628591857280719e-01
GS_179_5 0 NS_179 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 181/182
CS_181 NS_181 0 9.9999999999999998e-13
CS_182 NS_182 0 9.9999999999999998e-13
RS_181 NS_181 0 1.9636019836512071e+02
RS_182 NS_182 0 1.9636019836512071e+02
GL_181 0 NS_181 NS_182 0 1.5213319862255134e-01
GL_182 0 NS_182 NS_181 0 -1.5213319862255134e-01
GS_181_5 0 NS_181 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 183/184
CS_183 NS_183 0 9.9999999999999998e-13
CS_184 NS_184 0 9.9999999999999998e-13
RS_183 NS_183 0 4.3243187986905582e+02
RS_184 NS_184 0 4.3243187986905582e+02
GL_183 0 NS_183 NS_184 0 1.3841574306468743e-01
GL_184 0 NS_184 NS_183 0 -1.3841574306468743e-01
GS_183_5 0 NS_183 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 3.6825571251433115e+02
RS_186 NS_186 0 3.6825571251433115e+02
GL_185 0 NS_185 NS_186 0 1.3950469341450047e-01
GL_186 0 NS_186 NS_185 0 -1.3950469341450047e-01
GS_185_5 0 NS_185 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 3.0711053107765838e+02
RS_188 NS_188 0 3.0711053107765838e+02
GL_187 0 NS_187 NS_188 0 1.4553496077846845e-01
GL_188 0 NS_188 NS_187 0 -1.4553496077846845e-01
GS_187_5 0 NS_187 NA_5 0 1.0694336352474016e+00
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 4.6727671488342185e+02
RS_190 NS_190 0 4.6727671488342185e+02
GL_189 0 NS_189 NS_190 0 1.4422859584763473e-01
GL_190 0 NS_190 NS_189 0 -1.4422859584763473e-01
GS_189_5 0 NS_189 NA_5 0 1.0694336352474016e+00
*
* Real pole n. 191
CS_191 NS_191 0 9.9999999999999998e-13
RS_191 NS_191 0 3.4413071814985372e+00
GS_191_6 0 NS_191 NA_6 0 1.0694336352474016e+00
*
* Real pole n. 192
CS_192 NS_192 0 9.9999999999999998e-13
RS_192 NS_192 0 3.0797075048869470e+01
GS_192_6 0 NS_192 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 8.9335977936087705e+00
RS_194 NS_194 0 8.9335977936087705e+00
GL_193 0 NS_193 NS_194 0 2.2441700641819512e-01
GL_194 0 NS_194 NS_193 0 -2.2441700641819512e-01
GS_193_6 0 NS_193 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 5.9158463852536897e+01
RS_196 NS_196 0 5.9158463852536897e+01
GL_195 0 NS_195 NS_196 0 2.6680991281534006e-01
GL_196 0 NS_196 NS_195 0 -2.6680991281534006e-01
GS_195_6 0 NS_195 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 9.2065834236318878e+01
RS_198 NS_198 0 9.2065834236318864e+01
GL_197 0 NS_197 NS_198 0 2.4567219632280338e-01
GL_198 0 NS_198 NS_197 0 -2.4567219632280338e-01
GS_197_6 0 NS_197 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 1.4764174191595519e+01
RS_200 NS_200 0 1.4764174191595517e+01
GL_199 0 NS_199 NS_200 0 1.4400577194218670e-02
GL_200 0 NS_200 NS_199 0 -1.4400577194218670e-02
GS_199_6 0 NS_199 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 201/202
CS_201 NS_201 0 9.9999999999999998e-13
CS_202 NS_202 0 9.9999999999999998e-13
RS_201 NS_201 0 9.7834937041354195e+01
RS_202 NS_202 0 9.7834937041354195e+01
GL_201 0 NS_201 NS_202 0 6.3371310235267833e-02
GL_202 0 NS_202 NS_201 0 -6.3371310235267833e-02
GS_201_6 0 NS_201 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 203/204
CS_203 NS_203 0 9.9999999999999998e-13
CS_204 NS_204 0 9.9999999999999998e-13
RS_203 NS_203 0 1.4785099744646029e+01
RS_204 NS_204 0 1.4785099744646031e+01
GL_203 0 NS_203 NS_204 0 1.5607347485362127e-01
GL_204 0 NS_204 NS_203 0 -1.5607347485362127e-01
GS_203_6 0 NS_203 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 1.3466736941644649e+02
RS_206 NS_206 0 1.3466736941644649e+02
GL_205 0 NS_205 NS_206 0 2.3468192685328568e-01
GL_206 0 NS_206 NS_205 0 -2.3468192685328568e-01
GS_205_6 0 NS_205 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 1.5102368550954495e+02
RS_208 NS_208 0 1.5102368550954495e+02
GL_207 0 NS_207 NS_208 0 2.2562219216120838e-01
GL_208 0 NS_208 NS_207 0 -2.2562219216120838e-01
GS_207_6 0 NS_207 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 1.6979945400908466e+02
RS_210 NS_210 0 1.6979945400908468e+02
GL_209 0 NS_209 NS_210 0 2.1538055438627146e-01
GL_210 0 NS_210 NS_209 0 -2.1538055438627146e-01
GS_209_6 0 NS_209 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 2.2834543421620666e+02
RS_212 NS_212 0 2.2834543421620666e+02
GL_211 0 NS_211 NS_212 0 2.0391309107915187e-01
GL_212 0 NS_212 NS_211 0 -2.0391309107915187e-01
GS_211_6 0 NS_211 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 3.4087022095623759e+01
RS_214 NS_214 0 3.4087022095623759e+01
GL_213 0 NS_213 NS_214 0 1.5530350392230499e-01
GL_214 0 NS_214 NS_213 0 -1.5530350392230499e-01
GS_213_6 0 NS_213 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 7.5761470378414444e+01
RS_216 NS_216 0 7.5761470378414444e+01
GL_215 0 NS_215 NS_216 0 1.6902428843873585e-01
GL_216 0 NS_216 NS_215 0 -1.6902428843873585e-01
GS_215_6 0 NS_215 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 1.1061014882057984e+02
RS_218 NS_218 0 1.1061014882057984e+02
GL_217 0 NS_217 NS_218 0 1.5628591857280719e-01
GL_218 0 NS_218 NS_217 0 -1.5628591857280719e-01
GS_217_6 0 NS_217 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 1.9636019836512071e+02
RS_220 NS_220 0 1.9636019836512071e+02
GL_219 0 NS_219 NS_220 0 1.5213319862255134e-01
GL_220 0 NS_220 NS_219 0 -1.5213319862255134e-01
GS_219_6 0 NS_219 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 221/222
CS_221 NS_221 0 9.9999999999999998e-13
CS_222 NS_222 0 9.9999999999999998e-13
RS_221 NS_221 0 4.3243187986905582e+02
RS_222 NS_222 0 4.3243187986905582e+02
GL_221 0 NS_221 NS_222 0 1.3841574306468743e-01
GL_222 0 NS_222 NS_221 0 -1.3841574306468743e-01
GS_221_6 0 NS_221 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 223/224
CS_223 NS_223 0 9.9999999999999998e-13
CS_224 NS_224 0 9.9999999999999998e-13
RS_223 NS_223 0 3.6825571251433115e+02
RS_224 NS_224 0 3.6825571251433115e+02
GL_223 0 NS_223 NS_224 0 1.3950469341450047e-01
GL_224 0 NS_224 NS_223 0 -1.3950469341450047e-01
GS_223_6 0 NS_223 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 225/226
CS_225 NS_225 0 9.9999999999999998e-13
CS_226 NS_226 0 9.9999999999999998e-13
RS_225 NS_225 0 3.0711053107765838e+02
RS_226 NS_226 0 3.0711053107765838e+02
GL_225 0 NS_225 NS_226 0 1.4553496077846845e-01
GL_226 0 NS_226 NS_225 0 -1.4553496077846845e-01
GS_225_6 0 NS_225 NA_6 0 1.0694336352474016e+00
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 4.6727671488342185e+02
RS_228 NS_228 0 4.6727671488342185e+02
GL_227 0 NS_227 NS_228 0 1.4422859584763473e-01
GL_228 0 NS_228 NS_227 0 -1.4422859584763473e-01
GS_227_6 0 NS_227 NA_6 0 1.0694336352474016e+00
*
* Real pole n. 229
CS_229 NS_229 0 9.9999999999999998e-13
RS_229 NS_229 0 3.4413071814985372e+00
GS_229_7 0 NS_229 NA_7 0 1.0694336352474016e+00
*
* Real pole n. 230
CS_230 NS_230 0 9.9999999999999998e-13
RS_230 NS_230 0 3.0797075048869470e+01
GS_230_7 0 NS_230 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 8.9335977936087705e+00
RS_232 NS_232 0 8.9335977936087705e+00
GL_231 0 NS_231 NS_232 0 2.2441700641819512e-01
GL_232 0 NS_232 NS_231 0 -2.2441700641819512e-01
GS_231_7 0 NS_231 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 5.9158463852536897e+01
RS_234 NS_234 0 5.9158463852536897e+01
GL_233 0 NS_233 NS_234 0 2.6680991281534006e-01
GL_234 0 NS_234 NS_233 0 -2.6680991281534006e-01
GS_233_7 0 NS_233 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 9.2065834236318878e+01
RS_236 NS_236 0 9.2065834236318864e+01
GL_235 0 NS_235 NS_236 0 2.4567219632280338e-01
GL_236 0 NS_236 NS_235 0 -2.4567219632280338e-01
GS_235_7 0 NS_235 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 1.4764174191595519e+01
RS_238 NS_238 0 1.4764174191595517e+01
GL_237 0 NS_237 NS_238 0 1.4400577194218670e-02
GL_238 0 NS_238 NS_237 0 -1.4400577194218670e-02
GS_237_7 0 NS_237 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 9.7834937041354195e+01
RS_240 NS_240 0 9.7834937041354195e+01
GL_239 0 NS_239 NS_240 0 6.3371310235267833e-02
GL_240 0 NS_240 NS_239 0 -6.3371310235267833e-02
GS_239_7 0 NS_239 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 241/242
CS_241 NS_241 0 9.9999999999999998e-13
CS_242 NS_242 0 9.9999999999999998e-13
RS_241 NS_241 0 1.4785099744646029e+01
RS_242 NS_242 0 1.4785099744646031e+01
GL_241 0 NS_241 NS_242 0 1.5607347485362127e-01
GL_242 0 NS_242 NS_241 0 -1.5607347485362127e-01
GS_241_7 0 NS_241 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 243/244
CS_243 NS_243 0 9.9999999999999998e-13
CS_244 NS_244 0 9.9999999999999998e-13
RS_243 NS_243 0 1.3466736941644649e+02
RS_244 NS_244 0 1.3466736941644649e+02
GL_243 0 NS_243 NS_244 0 2.3468192685328568e-01
GL_244 0 NS_244 NS_243 0 -2.3468192685328568e-01
GS_243_7 0 NS_243 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 245/246
CS_245 NS_245 0 9.9999999999999998e-13
CS_246 NS_246 0 9.9999999999999998e-13
RS_245 NS_245 0 1.5102368550954495e+02
RS_246 NS_246 0 1.5102368550954495e+02
GL_245 0 NS_245 NS_246 0 2.2562219216120838e-01
GL_246 0 NS_246 NS_245 0 -2.2562219216120838e-01
GS_245_7 0 NS_245 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 247/248
CS_247 NS_247 0 9.9999999999999998e-13
CS_248 NS_248 0 9.9999999999999998e-13
RS_247 NS_247 0 1.6979945400908466e+02
RS_248 NS_248 0 1.6979945400908468e+02
GL_247 0 NS_247 NS_248 0 2.1538055438627146e-01
GL_248 0 NS_248 NS_247 0 -2.1538055438627146e-01
GS_247_7 0 NS_247 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 249/250
CS_249 NS_249 0 9.9999999999999998e-13
CS_250 NS_250 0 9.9999999999999998e-13
RS_249 NS_249 0 2.2834543421620666e+02
RS_250 NS_250 0 2.2834543421620666e+02
GL_249 0 NS_249 NS_250 0 2.0391309107915187e-01
GL_250 0 NS_250 NS_249 0 -2.0391309107915187e-01
GS_249_7 0 NS_249 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 251/252
CS_251 NS_251 0 9.9999999999999998e-13
CS_252 NS_252 0 9.9999999999999998e-13
RS_251 NS_251 0 3.4087022095623759e+01
RS_252 NS_252 0 3.4087022095623759e+01
GL_251 0 NS_251 NS_252 0 1.5530350392230499e-01
GL_252 0 NS_252 NS_251 0 -1.5530350392230499e-01
GS_251_7 0 NS_251 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 253/254
CS_253 NS_253 0 9.9999999999999998e-13
CS_254 NS_254 0 9.9999999999999998e-13
RS_253 NS_253 0 7.5761470378414444e+01
RS_254 NS_254 0 7.5761470378414444e+01
GL_253 0 NS_253 NS_254 0 1.6902428843873585e-01
GL_254 0 NS_254 NS_253 0 -1.6902428843873585e-01
GS_253_7 0 NS_253 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 255/256
CS_255 NS_255 0 9.9999999999999998e-13
CS_256 NS_256 0 9.9999999999999998e-13
RS_255 NS_255 0 1.1061014882057984e+02
RS_256 NS_256 0 1.1061014882057984e+02
GL_255 0 NS_255 NS_256 0 1.5628591857280719e-01
GL_256 0 NS_256 NS_255 0 -1.5628591857280719e-01
GS_255_7 0 NS_255 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 257/258
CS_257 NS_257 0 9.9999999999999998e-13
CS_258 NS_258 0 9.9999999999999998e-13
RS_257 NS_257 0 1.9636019836512071e+02
RS_258 NS_258 0 1.9636019836512071e+02
GL_257 0 NS_257 NS_258 0 1.5213319862255134e-01
GL_258 0 NS_258 NS_257 0 -1.5213319862255134e-01
GS_257_7 0 NS_257 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 259/260
CS_259 NS_259 0 9.9999999999999998e-13
CS_260 NS_260 0 9.9999999999999998e-13
RS_259 NS_259 0 4.3243187986905582e+02
RS_260 NS_260 0 4.3243187986905582e+02
GL_259 0 NS_259 NS_260 0 1.3841574306468743e-01
GL_260 0 NS_260 NS_259 0 -1.3841574306468743e-01
GS_259_7 0 NS_259 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 261/262
CS_261 NS_261 0 9.9999999999999998e-13
CS_262 NS_262 0 9.9999999999999998e-13
RS_261 NS_261 0 3.6825571251433115e+02
RS_262 NS_262 0 3.6825571251433115e+02
GL_261 0 NS_261 NS_262 0 1.3950469341450047e-01
GL_262 0 NS_262 NS_261 0 -1.3950469341450047e-01
GS_261_7 0 NS_261 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 263/264
CS_263 NS_263 0 9.9999999999999998e-13
CS_264 NS_264 0 9.9999999999999998e-13
RS_263 NS_263 0 3.0711053107765838e+02
RS_264 NS_264 0 3.0711053107765838e+02
GL_263 0 NS_263 NS_264 0 1.4553496077846845e-01
GL_264 0 NS_264 NS_263 0 -1.4553496077846845e-01
GS_263_7 0 NS_263 NA_7 0 1.0694336352474016e+00
*
* Complex pair n. 265/266
CS_265 NS_265 0 9.9999999999999998e-13
CS_266 NS_266 0 9.9999999999999998e-13
RS_265 NS_265 0 4.6727671488342185e+02
RS_266 NS_266 0 4.6727671488342185e+02
GL_265 0 NS_265 NS_266 0 1.4422859584763473e-01
GL_266 0 NS_266 NS_265 0 -1.4422859584763473e-01
GS_265_7 0 NS_265 NA_7 0 1.0694336352474016e+00
*
* Real pole n. 267
CS_267 NS_267 0 9.9999999999999998e-13
RS_267 NS_267 0 3.4413071814985372e+00
GS_267_8 0 NS_267 NA_8 0 1.0694336352474016e+00
*
* Real pole n. 268
CS_268 NS_268 0 9.9999999999999998e-13
RS_268 NS_268 0 3.0797075048869470e+01
GS_268_8 0 NS_268 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 269/270
CS_269 NS_269 0 9.9999999999999998e-13
CS_270 NS_270 0 9.9999999999999998e-13
RS_269 NS_269 0 8.9335977936087705e+00
RS_270 NS_270 0 8.9335977936087705e+00
GL_269 0 NS_269 NS_270 0 2.2441700641819512e-01
GL_270 0 NS_270 NS_269 0 -2.2441700641819512e-01
GS_269_8 0 NS_269 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 271/272
CS_271 NS_271 0 9.9999999999999998e-13
CS_272 NS_272 0 9.9999999999999998e-13
RS_271 NS_271 0 5.9158463852536897e+01
RS_272 NS_272 0 5.9158463852536897e+01
GL_271 0 NS_271 NS_272 0 2.6680991281534006e-01
GL_272 0 NS_272 NS_271 0 -2.6680991281534006e-01
GS_271_8 0 NS_271 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 273/274
CS_273 NS_273 0 9.9999999999999998e-13
CS_274 NS_274 0 9.9999999999999998e-13
RS_273 NS_273 0 9.2065834236318878e+01
RS_274 NS_274 0 9.2065834236318864e+01
GL_273 0 NS_273 NS_274 0 2.4567219632280338e-01
GL_274 0 NS_274 NS_273 0 -2.4567219632280338e-01
GS_273_8 0 NS_273 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 275/276
CS_275 NS_275 0 9.9999999999999998e-13
CS_276 NS_276 0 9.9999999999999998e-13
RS_275 NS_275 0 1.4764174191595519e+01
RS_276 NS_276 0 1.4764174191595517e+01
GL_275 0 NS_275 NS_276 0 1.4400577194218670e-02
GL_276 0 NS_276 NS_275 0 -1.4400577194218670e-02
GS_275_8 0 NS_275 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 277/278
CS_277 NS_277 0 9.9999999999999998e-13
CS_278 NS_278 0 9.9999999999999998e-13
RS_277 NS_277 0 9.7834937041354195e+01
RS_278 NS_278 0 9.7834937041354195e+01
GL_277 0 NS_277 NS_278 0 6.3371310235267833e-02
GL_278 0 NS_278 NS_277 0 -6.3371310235267833e-02
GS_277_8 0 NS_277 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 279/280
CS_279 NS_279 0 9.9999999999999998e-13
CS_280 NS_280 0 9.9999999999999998e-13
RS_279 NS_279 0 1.4785099744646029e+01
RS_280 NS_280 0 1.4785099744646031e+01
GL_279 0 NS_279 NS_280 0 1.5607347485362127e-01
GL_280 0 NS_280 NS_279 0 -1.5607347485362127e-01
GS_279_8 0 NS_279 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 281/282
CS_281 NS_281 0 9.9999999999999998e-13
CS_282 NS_282 0 9.9999999999999998e-13
RS_281 NS_281 0 1.3466736941644649e+02
RS_282 NS_282 0 1.3466736941644649e+02
GL_281 0 NS_281 NS_282 0 2.3468192685328568e-01
GL_282 0 NS_282 NS_281 0 -2.3468192685328568e-01
GS_281_8 0 NS_281 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 283/284
CS_283 NS_283 0 9.9999999999999998e-13
CS_284 NS_284 0 9.9999999999999998e-13
RS_283 NS_283 0 1.5102368550954495e+02
RS_284 NS_284 0 1.5102368550954495e+02
GL_283 0 NS_283 NS_284 0 2.2562219216120838e-01
GL_284 0 NS_284 NS_283 0 -2.2562219216120838e-01
GS_283_8 0 NS_283 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 285/286
CS_285 NS_285 0 9.9999999999999998e-13
CS_286 NS_286 0 9.9999999999999998e-13
RS_285 NS_285 0 1.6979945400908466e+02
RS_286 NS_286 0 1.6979945400908468e+02
GL_285 0 NS_285 NS_286 0 2.1538055438627146e-01
GL_286 0 NS_286 NS_285 0 -2.1538055438627146e-01
GS_285_8 0 NS_285 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 287/288
CS_287 NS_287 0 9.9999999999999998e-13
CS_288 NS_288 0 9.9999999999999998e-13
RS_287 NS_287 0 2.2834543421620666e+02
RS_288 NS_288 0 2.2834543421620666e+02
GL_287 0 NS_287 NS_288 0 2.0391309107915187e-01
GL_288 0 NS_288 NS_287 0 -2.0391309107915187e-01
GS_287_8 0 NS_287 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 289/290
CS_289 NS_289 0 9.9999999999999998e-13
CS_290 NS_290 0 9.9999999999999998e-13
RS_289 NS_289 0 3.4087022095623759e+01
RS_290 NS_290 0 3.4087022095623759e+01
GL_289 0 NS_289 NS_290 0 1.5530350392230499e-01
GL_290 0 NS_290 NS_289 0 -1.5530350392230499e-01
GS_289_8 0 NS_289 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 291/292
CS_291 NS_291 0 9.9999999999999998e-13
CS_292 NS_292 0 9.9999999999999998e-13
RS_291 NS_291 0 7.5761470378414444e+01
RS_292 NS_292 0 7.5761470378414444e+01
GL_291 0 NS_291 NS_292 0 1.6902428843873585e-01
GL_292 0 NS_292 NS_291 0 -1.6902428843873585e-01
GS_291_8 0 NS_291 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 293/294
CS_293 NS_293 0 9.9999999999999998e-13
CS_294 NS_294 0 9.9999999999999998e-13
RS_293 NS_293 0 1.1061014882057984e+02
RS_294 NS_294 0 1.1061014882057984e+02
GL_293 0 NS_293 NS_294 0 1.5628591857280719e-01
GL_294 0 NS_294 NS_293 0 -1.5628591857280719e-01
GS_293_8 0 NS_293 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 295/296
CS_295 NS_295 0 9.9999999999999998e-13
CS_296 NS_296 0 9.9999999999999998e-13
RS_295 NS_295 0 1.9636019836512071e+02
RS_296 NS_296 0 1.9636019836512071e+02
GL_295 0 NS_295 NS_296 0 1.5213319862255134e-01
GL_296 0 NS_296 NS_295 0 -1.5213319862255134e-01
GS_295_8 0 NS_295 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 297/298
CS_297 NS_297 0 9.9999999999999998e-13
CS_298 NS_298 0 9.9999999999999998e-13
RS_297 NS_297 0 4.3243187986905582e+02
RS_298 NS_298 0 4.3243187986905582e+02
GL_297 0 NS_297 NS_298 0 1.3841574306468743e-01
GL_298 0 NS_298 NS_297 0 -1.3841574306468743e-01
GS_297_8 0 NS_297 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 299/300
CS_299 NS_299 0 9.9999999999999998e-13
CS_300 NS_300 0 9.9999999999999998e-13
RS_299 NS_299 0 3.6825571251433115e+02
RS_300 NS_300 0 3.6825571251433115e+02
GL_299 0 NS_299 NS_300 0 1.3950469341450047e-01
GL_300 0 NS_300 NS_299 0 -1.3950469341450047e-01
GS_299_8 0 NS_299 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 301/302
CS_301 NS_301 0 9.9999999999999998e-13
CS_302 NS_302 0 9.9999999999999998e-13
RS_301 NS_301 0 3.0711053107765838e+02
RS_302 NS_302 0 3.0711053107765838e+02
GL_301 0 NS_301 NS_302 0 1.4553496077846845e-01
GL_302 0 NS_302 NS_301 0 -1.4553496077846845e-01
GS_301_8 0 NS_301 NA_8 0 1.0694336352474016e+00
*
* Complex pair n. 303/304
CS_303 NS_303 0 9.9999999999999998e-13
CS_304 NS_304 0 9.9999999999999998e-13
RS_303 NS_303 0 4.6727671488342185e+02
RS_304 NS_304 0 4.6727671488342185e+02
GL_303 0 NS_303 NS_304 0 1.4422859584763473e-01
GL_304 0 NS_304 NS_303 0 -1.4422859584763473e-01
GS_303_8 0 NS_303 NA_8 0 1.0694336352474016e+00
*
* Real pole n. 305
CS_305 NS_305 0 9.9999999999999998e-13
RS_305 NS_305 0 3.4413071814985372e+00
GS_305_9 0 NS_305 NA_9 0 1.0694336352474016e+00
*
* Real pole n. 306
CS_306 NS_306 0 9.9999999999999998e-13
RS_306 NS_306 0 3.0797075048869470e+01
GS_306_9 0 NS_306 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 307/308
CS_307 NS_307 0 9.9999999999999998e-13
CS_308 NS_308 0 9.9999999999999998e-13
RS_307 NS_307 0 8.9335977936087705e+00
RS_308 NS_308 0 8.9335977936087705e+00
GL_307 0 NS_307 NS_308 0 2.2441700641819512e-01
GL_308 0 NS_308 NS_307 0 -2.2441700641819512e-01
GS_307_9 0 NS_307 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 309/310
CS_309 NS_309 0 9.9999999999999998e-13
CS_310 NS_310 0 9.9999999999999998e-13
RS_309 NS_309 0 5.9158463852536897e+01
RS_310 NS_310 0 5.9158463852536897e+01
GL_309 0 NS_309 NS_310 0 2.6680991281534006e-01
GL_310 0 NS_310 NS_309 0 -2.6680991281534006e-01
GS_309_9 0 NS_309 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 311/312
CS_311 NS_311 0 9.9999999999999998e-13
CS_312 NS_312 0 9.9999999999999998e-13
RS_311 NS_311 0 9.2065834236318878e+01
RS_312 NS_312 0 9.2065834236318864e+01
GL_311 0 NS_311 NS_312 0 2.4567219632280338e-01
GL_312 0 NS_312 NS_311 0 -2.4567219632280338e-01
GS_311_9 0 NS_311 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 313/314
CS_313 NS_313 0 9.9999999999999998e-13
CS_314 NS_314 0 9.9999999999999998e-13
RS_313 NS_313 0 1.4764174191595519e+01
RS_314 NS_314 0 1.4764174191595517e+01
GL_313 0 NS_313 NS_314 0 1.4400577194218670e-02
GL_314 0 NS_314 NS_313 0 -1.4400577194218670e-02
GS_313_9 0 NS_313 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 315/316
CS_315 NS_315 0 9.9999999999999998e-13
CS_316 NS_316 0 9.9999999999999998e-13
RS_315 NS_315 0 9.7834937041354195e+01
RS_316 NS_316 0 9.7834937041354195e+01
GL_315 0 NS_315 NS_316 0 6.3371310235267833e-02
GL_316 0 NS_316 NS_315 0 -6.3371310235267833e-02
GS_315_9 0 NS_315 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 317/318
CS_317 NS_317 0 9.9999999999999998e-13
CS_318 NS_318 0 9.9999999999999998e-13
RS_317 NS_317 0 1.4785099744646029e+01
RS_318 NS_318 0 1.4785099744646031e+01
GL_317 0 NS_317 NS_318 0 1.5607347485362127e-01
GL_318 0 NS_318 NS_317 0 -1.5607347485362127e-01
GS_317_9 0 NS_317 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 319/320
CS_319 NS_319 0 9.9999999999999998e-13
CS_320 NS_320 0 9.9999999999999998e-13
RS_319 NS_319 0 1.3466736941644649e+02
RS_320 NS_320 0 1.3466736941644649e+02
GL_319 0 NS_319 NS_320 0 2.3468192685328568e-01
GL_320 0 NS_320 NS_319 0 -2.3468192685328568e-01
GS_319_9 0 NS_319 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 321/322
CS_321 NS_321 0 9.9999999999999998e-13
CS_322 NS_322 0 9.9999999999999998e-13
RS_321 NS_321 0 1.5102368550954495e+02
RS_322 NS_322 0 1.5102368550954495e+02
GL_321 0 NS_321 NS_322 0 2.2562219216120838e-01
GL_322 0 NS_322 NS_321 0 -2.2562219216120838e-01
GS_321_9 0 NS_321 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 323/324
CS_323 NS_323 0 9.9999999999999998e-13
CS_324 NS_324 0 9.9999999999999998e-13
RS_323 NS_323 0 1.6979945400908466e+02
RS_324 NS_324 0 1.6979945400908468e+02
GL_323 0 NS_323 NS_324 0 2.1538055438627146e-01
GL_324 0 NS_324 NS_323 0 -2.1538055438627146e-01
GS_323_9 0 NS_323 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 325/326
CS_325 NS_325 0 9.9999999999999998e-13
CS_326 NS_326 0 9.9999999999999998e-13
RS_325 NS_325 0 2.2834543421620666e+02
RS_326 NS_326 0 2.2834543421620666e+02
GL_325 0 NS_325 NS_326 0 2.0391309107915187e-01
GL_326 0 NS_326 NS_325 0 -2.0391309107915187e-01
GS_325_9 0 NS_325 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 327/328
CS_327 NS_327 0 9.9999999999999998e-13
CS_328 NS_328 0 9.9999999999999998e-13
RS_327 NS_327 0 3.4087022095623759e+01
RS_328 NS_328 0 3.4087022095623759e+01
GL_327 0 NS_327 NS_328 0 1.5530350392230499e-01
GL_328 0 NS_328 NS_327 0 -1.5530350392230499e-01
GS_327_9 0 NS_327 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 329/330
CS_329 NS_329 0 9.9999999999999998e-13
CS_330 NS_330 0 9.9999999999999998e-13
RS_329 NS_329 0 7.5761470378414444e+01
RS_330 NS_330 0 7.5761470378414444e+01
GL_329 0 NS_329 NS_330 0 1.6902428843873585e-01
GL_330 0 NS_330 NS_329 0 -1.6902428843873585e-01
GS_329_9 0 NS_329 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 331/332
CS_331 NS_331 0 9.9999999999999998e-13
CS_332 NS_332 0 9.9999999999999998e-13
RS_331 NS_331 0 1.1061014882057984e+02
RS_332 NS_332 0 1.1061014882057984e+02
GL_331 0 NS_331 NS_332 0 1.5628591857280719e-01
GL_332 0 NS_332 NS_331 0 -1.5628591857280719e-01
GS_331_9 0 NS_331 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 333/334
CS_333 NS_333 0 9.9999999999999998e-13
CS_334 NS_334 0 9.9999999999999998e-13
RS_333 NS_333 0 1.9636019836512071e+02
RS_334 NS_334 0 1.9636019836512071e+02
GL_333 0 NS_333 NS_334 0 1.5213319862255134e-01
GL_334 0 NS_334 NS_333 0 -1.5213319862255134e-01
GS_333_9 0 NS_333 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 335/336
CS_335 NS_335 0 9.9999999999999998e-13
CS_336 NS_336 0 9.9999999999999998e-13
RS_335 NS_335 0 4.3243187986905582e+02
RS_336 NS_336 0 4.3243187986905582e+02
GL_335 0 NS_335 NS_336 0 1.3841574306468743e-01
GL_336 0 NS_336 NS_335 0 -1.3841574306468743e-01
GS_335_9 0 NS_335 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 337/338
CS_337 NS_337 0 9.9999999999999998e-13
CS_338 NS_338 0 9.9999999999999998e-13
RS_337 NS_337 0 3.6825571251433115e+02
RS_338 NS_338 0 3.6825571251433115e+02
GL_337 0 NS_337 NS_338 0 1.3950469341450047e-01
GL_338 0 NS_338 NS_337 0 -1.3950469341450047e-01
GS_337_9 0 NS_337 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 339/340
CS_339 NS_339 0 9.9999999999999998e-13
CS_340 NS_340 0 9.9999999999999998e-13
RS_339 NS_339 0 3.0711053107765838e+02
RS_340 NS_340 0 3.0711053107765838e+02
GL_339 0 NS_339 NS_340 0 1.4553496077846845e-01
GL_340 0 NS_340 NS_339 0 -1.4553496077846845e-01
GS_339_9 0 NS_339 NA_9 0 1.0694336352474016e+00
*
* Complex pair n. 341/342
CS_341 NS_341 0 9.9999999999999998e-13
CS_342 NS_342 0 9.9999999999999998e-13
RS_341 NS_341 0 4.6727671488342185e+02
RS_342 NS_342 0 4.6727671488342185e+02
GL_341 0 NS_341 NS_342 0 1.4422859584763473e-01
GL_342 0 NS_342 NS_341 0 -1.4422859584763473e-01
GS_341_9 0 NS_341 NA_9 0 1.0694336352474016e+00
*
* Real pole n. 343
CS_343 NS_343 0 9.9999999999999998e-13
RS_343 NS_343 0 3.4413071814985372e+00
GS_343_10 0 NS_343 NA_10 0 1.0694336352474016e+00
*
* Real pole n. 344
CS_344 NS_344 0 9.9999999999999998e-13
RS_344 NS_344 0 3.0797075048869470e+01
GS_344_10 0 NS_344 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 345/346
CS_345 NS_345 0 9.9999999999999998e-13
CS_346 NS_346 0 9.9999999999999998e-13
RS_345 NS_345 0 8.9335977936087705e+00
RS_346 NS_346 0 8.9335977936087705e+00
GL_345 0 NS_345 NS_346 0 2.2441700641819512e-01
GL_346 0 NS_346 NS_345 0 -2.2441700641819512e-01
GS_345_10 0 NS_345 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 347/348
CS_347 NS_347 0 9.9999999999999998e-13
CS_348 NS_348 0 9.9999999999999998e-13
RS_347 NS_347 0 5.9158463852536897e+01
RS_348 NS_348 0 5.9158463852536897e+01
GL_347 0 NS_347 NS_348 0 2.6680991281534006e-01
GL_348 0 NS_348 NS_347 0 -2.6680991281534006e-01
GS_347_10 0 NS_347 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 349/350
CS_349 NS_349 0 9.9999999999999998e-13
CS_350 NS_350 0 9.9999999999999998e-13
RS_349 NS_349 0 9.2065834236318878e+01
RS_350 NS_350 0 9.2065834236318864e+01
GL_349 0 NS_349 NS_350 0 2.4567219632280338e-01
GL_350 0 NS_350 NS_349 0 -2.4567219632280338e-01
GS_349_10 0 NS_349 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 351/352
CS_351 NS_351 0 9.9999999999999998e-13
CS_352 NS_352 0 9.9999999999999998e-13
RS_351 NS_351 0 1.4764174191595519e+01
RS_352 NS_352 0 1.4764174191595517e+01
GL_351 0 NS_351 NS_352 0 1.4400577194218670e-02
GL_352 0 NS_352 NS_351 0 -1.4400577194218670e-02
GS_351_10 0 NS_351 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 353/354
CS_353 NS_353 0 9.9999999999999998e-13
CS_354 NS_354 0 9.9999999999999998e-13
RS_353 NS_353 0 9.7834937041354195e+01
RS_354 NS_354 0 9.7834937041354195e+01
GL_353 0 NS_353 NS_354 0 6.3371310235267833e-02
GL_354 0 NS_354 NS_353 0 -6.3371310235267833e-02
GS_353_10 0 NS_353 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 355/356
CS_355 NS_355 0 9.9999999999999998e-13
CS_356 NS_356 0 9.9999999999999998e-13
RS_355 NS_355 0 1.4785099744646029e+01
RS_356 NS_356 0 1.4785099744646031e+01
GL_355 0 NS_355 NS_356 0 1.5607347485362127e-01
GL_356 0 NS_356 NS_355 0 -1.5607347485362127e-01
GS_355_10 0 NS_355 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 357/358
CS_357 NS_357 0 9.9999999999999998e-13
CS_358 NS_358 0 9.9999999999999998e-13
RS_357 NS_357 0 1.3466736941644649e+02
RS_358 NS_358 0 1.3466736941644649e+02
GL_357 0 NS_357 NS_358 0 2.3468192685328568e-01
GL_358 0 NS_358 NS_357 0 -2.3468192685328568e-01
GS_357_10 0 NS_357 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 359/360
CS_359 NS_359 0 9.9999999999999998e-13
CS_360 NS_360 0 9.9999999999999998e-13
RS_359 NS_359 0 1.5102368550954495e+02
RS_360 NS_360 0 1.5102368550954495e+02
GL_359 0 NS_359 NS_360 0 2.2562219216120838e-01
GL_360 0 NS_360 NS_359 0 -2.2562219216120838e-01
GS_359_10 0 NS_359 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 361/362
CS_361 NS_361 0 9.9999999999999998e-13
CS_362 NS_362 0 9.9999999999999998e-13
RS_361 NS_361 0 1.6979945400908466e+02
RS_362 NS_362 0 1.6979945400908468e+02
GL_361 0 NS_361 NS_362 0 2.1538055438627146e-01
GL_362 0 NS_362 NS_361 0 -2.1538055438627146e-01
GS_361_10 0 NS_361 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 363/364
CS_363 NS_363 0 9.9999999999999998e-13
CS_364 NS_364 0 9.9999999999999998e-13
RS_363 NS_363 0 2.2834543421620666e+02
RS_364 NS_364 0 2.2834543421620666e+02
GL_363 0 NS_363 NS_364 0 2.0391309107915187e-01
GL_364 0 NS_364 NS_363 0 -2.0391309107915187e-01
GS_363_10 0 NS_363 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 365/366
CS_365 NS_365 0 9.9999999999999998e-13
CS_366 NS_366 0 9.9999999999999998e-13
RS_365 NS_365 0 3.4087022095623759e+01
RS_366 NS_366 0 3.4087022095623759e+01
GL_365 0 NS_365 NS_366 0 1.5530350392230499e-01
GL_366 0 NS_366 NS_365 0 -1.5530350392230499e-01
GS_365_10 0 NS_365 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 367/368
CS_367 NS_367 0 9.9999999999999998e-13
CS_368 NS_368 0 9.9999999999999998e-13
RS_367 NS_367 0 7.5761470378414444e+01
RS_368 NS_368 0 7.5761470378414444e+01
GL_367 0 NS_367 NS_368 0 1.6902428843873585e-01
GL_368 0 NS_368 NS_367 0 -1.6902428843873585e-01
GS_367_10 0 NS_367 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 369/370
CS_369 NS_369 0 9.9999999999999998e-13
CS_370 NS_370 0 9.9999999999999998e-13
RS_369 NS_369 0 1.1061014882057984e+02
RS_370 NS_370 0 1.1061014882057984e+02
GL_369 0 NS_369 NS_370 0 1.5628591857280719e-01
GL_370 0 NS_370 NS_369 0 -1.5628591857280719e-01
GS_369_10 0 NS_369 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 371/372
CS_371 NS_371 0 9.9999999999999998e-13
CS_372 NS_372 0 9.9999999999999998e-13
RS_371 NS_371 0 1.9636019836512071e+02
RS_372 NS_372 0 1.9636019836512071e+02
GL_371 0 NS_371 NS_372 0 1.5213319862255134e-01
GL_372 0 NS_372 NS_371 0 -1.5213319862255134e-01
GS_371_10 0 NS_371 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 373/374
CS_373 NS_373 0 9.9999999999999998e-13
CS_374 NS_374 0 9.9999999999999998e-13
RS_373 NS_373 0 4.3243187986905582e+02
RS_374 NS_374 0 4.3243187986905582e+02
GL_373 0 NS_373 NS_374 0 1.3841574306468743e-01
GL_374 0 NS_374 NS_373 0 -1.3841574306468743e-01
GS_373_10 0 NS_373 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 375/376
CS_375 NS_375 0 9.9999999999999998e-13
CS_376 NS_376 0 9.9999999999999998e-13
RS_375 NS_375 0 3.6825571251433115e+02
RS_376 NS_376 0 3.6825571251433115e+02
GL_375 0 NS_375 NS_376 0 1.3950469341450047e-01
GL_376 0 NS_376 NS_375 0 -1.3950469341450047e-01
GS_375_10 0 NS_375 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 377/378
CS_377 NS_377 0 9.9999999999999998e-13
CS_378 NS_378 0 9.9999999999999998e-13
RS_377 NS_377 0 3.0711053107765838e+02
RS_378 NS_378 0 3.0711053107765838e+02
GL_377 0 NS_377 NS_378 0 1.4553496077846845e-01
GL_378 0 NS_378 NS_377 0 -1.4553496077846845e-01
GS_377_10 0 NS_377 NA_10 0 1.0694336352474016e+00
*
* Complex pair n. 379/380
CS_379 NS_379 0 9.9999999999999998e-13
CS_380 NS_380 0 9.9999999999999998e-13
RS_379 NS_379 0 4.6727671488342185e+02
RS_380 NS_380 0 4.6727671488342185e+02
GL_379 0 NS_379 NS_380 0 1.4422859584763473e-01
GL_380 0 NS_380 NS_379 0 -1.4422859584763473e-01
GS_379_10 0 NS_379 NA_10 0 1.0694336352474016e+00
*
* Real pole n. 381
CS_381 NS_381 0 9.9999999999999998e-13
RS_381 NS_381 0 3.4413071814985372e+00
GS_381_11 0 NS_381 NA_11 0 1.0694336352474016e+00
*
* Real pole n. 382
CS_382 NS_382 0 9.9999999999999998e-13
RS_382 NS_382 0 3.0797075048869470e+01
GS_382_11 0 NS_382 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 383/384
CS_383 NS_383 0 9.9999999999999998e-13
CS_384 NS_384 0 9.9999999999999998e-13
RS_383 NS_383 0 8.9335977936087705e+00
RS_384 NS_384 0 8.9335977936087705e+00
GL_383 0 NS_383 NS_384 0 2.2441700641819512e-01
GL_384 0 NS_384 NS_383 0 -2.2441700641819512e-01
GS_383_11 0 NS_383 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 385/386
CS_385 NS_385 0 9.9999999999999998e-13
CS_386 NS_386 0 9.9999999999999998e-13
RS_385 NS_385 0 5.9158463852536897e+01
RS_386 NS_386 0 5.9158463852536897e+01
GL_385 0 NS_385 NS_386 0 2.6680991281534006e-01
GL_386 0 NS_386 NS_385 0 -2.6680991281534006e-01
GS_385_11 0 NS_385 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 387/388
CS_387 NS_387 0 9.9999999999999998e-13
CS_388 NS_388 0 9.9999999999999998e-13
RS_387 NS_387 0 9.2065834236318878e+01
RS_388 NS_388 0 9.2065834236318864e+01
GL_387 0 NS_387 NS_388 0 2.4567219632280338e-01
GL_388 0 NS_388 NS_387 0 -2.4567219632280338e-01
GS_387_11 0 NS_387 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 389/390
CS_389 NS_389 0 9.9999999999999998e-13
CS_390 NS_390 0 9.9999999999999998e-13
RS_389 NS_389 0 1.4764174191595519e+01
RS_390 NS_390 0 1.4764174191595517e+01
GL_389 0 NS_389 NS_390 0 1.4400577194218670e-02
GL_390 0 NS_390 NS_389 0 -1.4400577194218670e-02
GS_389_11 0 NS_389 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 391/392
CS_391 NS_391 0 9.9999999999999998e-13
CS_392 NS_392 0 9.9999999999999998e-13
RS_391 NS_391 0 9.7834937041354195e+01
RS_392 NS_392 0 9.7834937041354195e+01
GL_391 0 NS_391 NS_392 0 6.3371310235267833e-02
GL_392 0 NS_392 NS_391 0 -6.3371310235267833e-02
GS_391_11 0 NS_391 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 393/394
CS_393 NS_393 0 9.9999999999999998e-13
CS_394 NS_394 0 9.9999999999999998e-13
RS_393 NS_393 0 1.4785099744646029e+01
RS_394 NS_394 0 1.4785099744646031e+01
GL_393 0 NS_393 NS_394 0 1.5607347485362127e-01
GL_394 0 NS_394 NS_393 0 -1.5607347485362127e-01
GS_393_11 0 NS_393 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 395/396
CS_395 NS_395 0 9.9999999999999998e-13
CS_396 NS_396 0 9.9999999999999998e-13
RS_395 NS_395 0 1.3466736941644649e+02
RS_396 NS_396 0 1.3466736941644649e+02
GL_395 0 NS_395 NS_396 0 2.3468192685328568e-01
GL_396 0 NS_396 NS_395 0 -2.3468192685328568e-01
GS_395_11 0 NS_395 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 397/398
CS_397 NS_397 0 9.9999999999999998e-13
CS_398 NS_398 0 9.9999999999999998e-13
RS_397 NS_397 0 1.5102368550954495e+02
RS_398 NS_398 0 1.5102368550954495e+02
GL_397 0 NS_397 NS_398 0 2.2562219216120838e-01
GL_398 0 NS_398 NS_397 0 -2.2562219216120838e-01
GS_397_11 0 NS_397 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 399/400
CS_399 NS_399 0 9.9999999999999998e-13
CS_400 NS_400 0 9.9999999999999998e-13
RS_399 NS_399 0 1.6979945400908466e+02
RS_400 NS_400 0 1.6979945400908468e+02
GL_399 0 NS_399 NS_400 0 2.1538055438627146e-01
GL_400 0 NS_400 NS_399 0 -2.1538055438627146e-01
GS_399_11 0 NS_399 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 401/402
CS_401 NS_401 0 9.9999999999999998e-13
CS_402 NS_402 0 9.9999999999999998e-13
RS_401 NS_401 0 2.2834543421620666e+02
RS_402 NS_402 0 2.2834543421620666e+02
GL_401 0 NS_401 NS_402 0 2.0391309107915187e-01
GL_402 0 NS_402 NS_401 0 -2.0391309107915187e-01
GS_401_11 0 NS_401 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 403/404
CS_403 NS_403 0 9.9999999999999998e-13
CS_404 NS_404 0 9.9999999999999998e-13
RS_403 NS_403 0 3.4087022095623759e+01
RS_404 NS_404 0 3.4087022095623759e+01
GL_403 0 NS_403 NS_404 0 1.5530350392230499e-01
GL_404 0 NS_404 NS_403 0 -1.5530350392230499e-01
GS_403_11 0 NS_403 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 405/406
CS_405 NS_405 0 9.9999999999999998e-13
CS_406 NS_406 0 9.9999999999999998e-13
RS_405 NS_405 0 7.5761470378414444e+01
RS_406 NS_406 0 7.5761470378414444e+01
GL_405 0 NS_405 NS_406 0 1.6902428843873585e-01
GL_406 0 NS_406 NS_405 0 -1.6902428843873585e-01
GS_405_11 0 NS_405 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 407/408
CS_407 NS_407 0 9.9999999999999998e-13
CS_408 NS_408 0 9.9999999999999998e-13
RS_407 NS_407 0 1.1061014882057984e+02
RS_408 NS_408 0 1.1061014882057984e+02
GL_407 0 NS_407 NS_408 0 1.5628591857280719e-01
GL_408 0 NS_408 NS_407 0 -1.5628591857280719e-01
GS_407_11 0 NS_407 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 409/410
CS_409 NS_409 0 9.9999999999999998e-13
CS_410 NS_410 0 9.9999999999999998e-13
RS_409 NS_409 0 1.9636019836512071e+02
RS_410 NS_410 0 1.9636019836512071e+02
GL_409 0 NS_409 NS_410 0 1.5213319862255134e-01
GL_410 0 NS_410 NS_409 0 -1.5213319862255134e-01
GS_409_11 0 NS_409 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 411/412
CS_411 NS_411 0 9.9999999999999998e-13
CS_412 NS_412 0 9.9999999999999998e-13
RS_411 NS_411 0 4.3243187986905582e+02
RS_412 NS_412 0 4.3243187986905582e+02
GL_411 0 NS_411 NS_412 0 1.3841574306468743e-01
GL_412 0 NS_412 NS_411 0 -1.3841574306468743e-01
GS_411_11 0 NS_411 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 413/414
CS_413 NS_413 0 9.9999999999999998e-13
CS_414 NS_414 0 9.9999999999999998e-13
RS_413 NS_413 0 3.6825571251433115e+02
RS_414 NS_414 0 3.6825571251433115e+02
GL_413 0 NS_413 NS_414 0 1.3950469341450047e-01
GL_414 0 NS_414 NS_413 0 -1.3950469341450047e-01
GS_413_11 0 NS_413 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 415/416
CS_415 NS_415 0 9.9999999999999998e-13
CS_416 NS_416 0 9.9999999999999998e-13
RS_415 NS_415 0 3.0711053107765838e+02
RS_416 NS_416 0 3.0711053107765838e+02
GL_415 0 NS_415 NS_416 0 1.4553496077846845e-01
GL_416 0 NS_416 NS_415 0 -1.4553496077846845e-01
GS_415_11 0 NS_415 NA_11 0 1.0694336352474016e+00
*
* Complex pair n. 417/418
CS_417 NS_417 0 9.9999999999999998e-13
CS_418 NS_418 0 9.9999999999999998e-13
RS_417 NS_417 0 4.6727671488342185e+02
RS_418 NS_418 0 4.6727671488342185e+02
GL_417 0 NS_417 NS_418 0 1.4422859584763473e-01
GL_418 0 NS_418 NS_417 0 -1.4422859584763473e-01
GS_417_11 0 NS_417 NA_11 0 1.0694336352474016e+00
*
* Real pole n. 419
CS_419 NS_419 0 9.9999999999999998e-13
RS_419 NS_419 0 3.4413071814985372e+00
GS_419_12 0 NS_419 NA_12 0 1.0694336352474016e+00
*
* Real pole n. 420
CS_420 NS_420 0 9.9999999999999998e-13
RS_420 NS_420 0 3.0797075048869470e+01
GS_420_12 0 NS_420 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 421/422
CS_421 NS_421 0 9.9999999999999998e-13
CS_422 NS_422 0 9.9999999999999998e-13
RS_421 NS_421 0 8.9335977936087705e+00
RS_422 NS_422 0 8.9335977936087705e+00
GL_421 0 NS_421 NS_422 0 2.2441700641819512e-01
GL_422 0 NS_422 NS_421 0 -2.2441700641819512e-01
GS_421_12 0 NS_421 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 423/424
CS_423 NS_423 0 9.9999999999999998e-13
CS_424 NS_424 0 9.9999999999999998e-13
RS_423 NS_423 0 5.9158463852536897e+01
RS_424 NS_424 0 5.9158463852536897e+01
GL_423 0 NS_423 NS_424 0 2.6680991281534006e-01
GL_424 0 NS_424 NS_423 0 -2.6680991281534006e-01
GS_423_12 0 NS_423 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 425/426
CS_425 NS_425 0 9.9999999999999998e-13
CS_426 NS_426 0 9.9999999999999998e-13
RS_425 NS_425 0 9.2065834236318878e+01
RS_426 NS_426 0 9.2065834236318864e+01
GL_425 0 NS_425 NS_426 0 2.4567219632280338e-01
GL_426 0 NS_426 NS_425 0 -2.4567219632280338e-01
GS_425_12 0 NS_425 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 427/428
CS_427 NS_427 0 9.9999999999999998e-13
CS_428 NS_428 0 9.9999999999999998e-13
RS_427 NS_427 0 1.4764174191595519e+01
RS_428 NS_428 0 1.4764174191595517e+01
GL_427 0 NS_427 NS_428 0 1.4400577194218670e-02
GL_428 0 NS_428 NS_427 0 -1.4400577194218670e-02
GS_427_12 0 NS_427 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 429/430
CS_429 NS_429 0 9.9999999999999998e-13
CS_430 NS_430 0 9.9999999999999998e-13
RS_429 NS_429 0 9.7834937041354195e+01
RS_430 NS_430 0 9.7834937041354195e+01
GL_429 0 NS_429 NS_430 0 6.3371310235267833e-02
GL_430 0 NS_430 NS_429 0 -6.3371310235267833e-02
GS_429_12 0 NS_429 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 431/432
CS_431 NS_431 0 9.9999999999999998e-13
CS_432 NS_432 0 9.9999999999999998e-13
RS_431 NS_431 0 1.4785099744646029e+01
RS_432 NS_432 0 1.4785099744646031e+01
GL_431 0 NS_431 NS_432 0 1.5607347485362127e-01
GL_432 0 NS_432 NS_431 0 -1.5607347485362127e-01
GS_431_12 0 NS_431 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 433/434
CS_433 NS_433 0 9.9999999999999998e-13
CS_434 NS_434 0 9.9999999999999998e-13
RS_433 NS_433 0 1.3466736941644649e+02
RS_434 NS_434 0 1.3466736941644649e+02
GL_433 0 NS_433 NS_434 0 2.3468192685328568e-01
GL_434 0 NS_434 NS_433 0 -2.3468192685328568e-01
GS_433_12 0 NS_433 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 435/436
CS_435 NS_435 0 9.9999999999999998e-13
CS_436 NS_436 0 9.9999999999999998e-13
RS_435 NS_435 0 1.5102368550954495e+02
RS_436 NS_436 0 1.5102368550954495e+02
GL_435 0 NS_435 NS_436 0 2.2562219216120838e-01
GL_436 0 NS_436 NS_435 0 -2.2562219216120838e-01
GS_435_12 0 NS_435 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 437/438
CS_437 NS_437 0 9.9999999999999998e-13
CS_438 NS_438 0 9.9999999999999998e-13
RS_437 NS_437 0 1.6979945400908466e+02
RS_438 NS_438 0 1.6979945400908468e+02
GL_437 0 NS_437 NS_438 0 2.1538055438627146e-01
GL_438 0 NS_438 NS_437 0 -2.1538055438627146e-01
GS_437_12 0 NS_437 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 439/440
CS_439 NS_439 0 9.9999999999999998e-13
CS_440 NS_440 0 9.9999999999999998e-13
RS_439 NS_439 0 2.2834543421620666e+02
RS_440 NS_440 0 2.2834543421620666e+02
GL_439 0 NS_439 NS_440 0 2.0391309107915187e-01
GL_440 0 NS_440 NS_439 0 -2.0391309107915187e-01
GS_439_12 0 NS_439 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 441/442
CS_441 NS_441 0 9.9999999999999998e-13
CS_442 NS_442 0 9.9999999999999998e-13
RS_441 NS_441 0 3.4087022095623759e+01
RS_442 NS_442 0 3.4087022095623759e+01
GL_441 0 NS_441 NS_442 0 1.5530350392230499e-01
GL_442 0 NS_442 NS_441 0 -1.5530350392230499e-01
GS_441_12 0 NS_441 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 443/444
CS_443 NS_443 0 9.9999999999999998e-13
CS_444 NS_444 0 9.9999999999999998e-13
RS_443 NS_443 0 7.5761470378414444e+01
RS_444 NS_444 0 7.5761470378414444e+01
GL_443 0 NS_443 NS_444 0 1.6902428843873585e-01
GL_444 0 NS_444 NS_443 0 -1.6902428843873585e-01
GS_443_12 0 NS_443 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 445/446
CS_445 NS_445 0 9.9999999999999998e-13
CS_446 NS_446 0 9.9999999999999998e-13
RS_445 NS_445 0 1.1061014882057984e+02
RS_446 NS_446 0 1.1061014882057984e+02
GL_445 0 NS_445 NS_446 0 1.5628591857280719e-01
GL_446 0 NS_446 NS_445 0 -1.5628591857280719e-01
GS_445_12 0 NS_445 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 447/448
CS_447 NS_447 0 9.9999999999999998e-13
CS_448 NS_448 0 9.9999999999999998e-13
RS_447 NS_447 0 1.9636019836512071e+02
RS_448 NS_448 0 1.9636019836512071e+02
GL_447 0 NS_447 NS_448 0 1.5213319862255134e-01
GL_448 0 NS_448 NS_447 0 -1.5213319862255134e-01
GS_447_12 0 NS_447 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 449/450
CS_449 NS_449 0 9.9999999999999998e-13
CS_450 NS_450 0 9.9999999999999998e-13
RS_449 NS_449 0 4.3243187986905582e+02
RS_450 NS_450 0 4.3243187986905582e+02
GL_449 0 NS_449 NS_450 0 1.3841574306468743e-01
GL_450 0 NS_450 NS_449 0 -1.3841574306468743e-01
GS_449_12 0 NS_449 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 451/452
CS_451 NS_451 0 9.9999999999999998e-13
CS_452 NS_452 0 9.9999999999999998e-13
RS_451 NS_451 0 3.6825571251433115e+02
RS_452 NS_452 0 3.6825571251433115e+02
GL_451 0 NS_451 NS_452 0 1.3950469341450047e-01
GL_452 0 NS_452 NS_451 0 -1.3950469341450047e-01
GS_451_12 0 NS_451 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 453/454
CS_453 NS_453 0 9.9999999999999998e-13
CS_454 NS_454 0 9.9999999999999998e-13
RS_453 NS_453 0 3.0711053107765838e+02
RS_454 NS_454 0 3.0711053107765838e+02
GL_453 0 NS_453 NS_454 0 1.4553496077846845e-01
GL_454 0 NS_454 NS_453 0 -1.4553496077846845e-01
GS_453_12 0 NS_453 NA_12 0 1.0694336352474016e+00
*
* Complex pair n. 455/456
CS_455 NS_455 0 9.9999999999999998e-13
CS_456 NS_456 0 9.9999999999999998e-13
RS_455 NS_455 0 4.6727671488342185e+02
RS_456 NS_456 0 4.6727671488342185e+02
GL_455 0 NS_455 NS_456 0 1.4422859584763473e-01
GL_456 0 NS_456 NS_455 0 -1.4422859584763473e-01
GS_455_12 0 NS_455 NA_12 0 1.0694336352474016e+00
*
******************************


.ends
*******************
* End of subcircuit
*******************
