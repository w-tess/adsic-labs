**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [6 6 46] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_2_BoardVia_noStub
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 -1.8047078975622879e-02
GC_1_2 b_1 NI_1 NS_2 0 1.3361873980626082e-02
GC_1_3 b_1 NI_1 NS_3 0 4.5139176651317354e-03
GC_1_4 b_1 NI_1 NS_4 0 1.0297076947396707e-02
GC_1_5 b_1 NI_1 NS_5 0 1.6461251122929621e-02
GC_1_6 b_1 NI_1 NS_6 0 -9.2095180954144644e-03
GC_1_7 b_1 NI_1 NS_7 0 5.2857742416966428e-03
GC_1_8 b_1 NI_1 NS_8 0 5.2121539794454984e-03
GC_1_9 b_1 NI_1 NS_9 0 2.8606201150720759e-03
GC_1_10 b_1 NI_1 NS_10 0 4.6862086376231980e-03
GC_1_11 b_1 NI_1 NS_11 0 9.5130531050769563e-03
GC_1_12 b_1 NI_1 NS_12 0 1.0162429927786491e-02
GC_1_13 b_1 NI_1 NS_13 0 2.5493333539041373e-04
GC_1_14 b_1 NI_1 NS_14 0 2.0422895526801837e-04
GC_1_15 b_1 NI_1 NS_15 0 -5.5932841993935104e-05
GC_1_16 b_1 NI_1 NS_16 0 5.9054163362031938e-05
GC_1_17 b_1 NI_1 NS_17 0 1.2774975815327337e-03
GC_1_18 b_1 NI_1 NS_18 0 -3.1575387358942432e-04
GC_1_19 b_1 NI_1 NS_19 0 7.9275218213680458e-05
GC_1_20 b_1 NI_1 NS_20 0 4.3443711923828379e-05
GC_1_21 b_1 NI_1 NS_21 0 1.2177446143092376e-04
GC_1_22 b_1 NI_1 NS_22 0 -5.5606738024718727e-05
GC_1_23 b_1 NI_1 NS_23 0 -1.2512949756654050e-05
GC_1_24 b_1 NI_1 NS_24 0 -3.4953930854387469e-07
GC_1_25 b_1 NI_1 NS_25 0 -5.1232029741031630e-03
GC_1_26 b_1 NI_1 NS_26 0 6.4910551363581738e-03
GC_1_27 b_1 NI_1 NS_27 0 5.9483715614444309e-03
GC_1_28 b_1 NI_1 NS_28 0 -6.4050773905122800e-04
GC_1_29 b_1 NI_1 NS_29 0 -4.8563861193415530e-04
GC_1_30 b_1 NI_1 NS_30 0 5.1266897881240654e-04
GC_1_31 b_1 NI_1 NS_31 0 1.7377004564462460e-06
GC_1_32 b_1 NI_1 NS_32 0 4.8199204227323768e-06
GC_1_33 b_1 NI_1 NS_33 0 2.3683291538138685e-04
GC_1_34 b_1 NI_1 NS_34 0 3.2011993544221540e-05
GC_1_35 b_1 NI_1 NS_35 0 5.5081642545477103e-06
GC_1_36 b_1 NI_1 NS_36 0 1.6379441744153186e-06
GC_1_37 b_1 NI_1 NS_37 0 2.9735096195435413e-06
GC_1_38 b_1 NI_1 NS_38 0 3.1478022600746553e-06
GC_1_39 b_1 NI_1 NS_39 0 -4.0178368564975573e-04
GC_1_40 b_1 NI_1 NS_40 0 3.0192980625090712e-04
GC_1_41 b_1 NI_1 NS_41 0 -7.5805280475661559e-05
GC_1_42 b_1 NI_1 NS_42 0 -3.3816664895293360e-05
GC_1_43 b_1 NI_1 NS_43 0 -2.1225703896696590e-05
GC_1_44 b_1 NI_1 NS_44 0 1.7497587049806047e-05
GC_1_45 b_1 NI_1 NS_45 0 2.6054150235721187e-02
GC_1_46 b_1 NI_1 NS_46 0 1.6788223938157692e-02
GC_1_47 b_1 NI_1 NS_47 0 -1.9815077026460990e-02
GC_1_48 b_1 NI_1 NS_48 0 -7.4654803423593328e-03
GC_1_49 b_1 NI_1 NS_49 0 -2.6099780470199577e-02
GC_1_50 b_1 NI_1 NS_50 0 2.0041949380766848e-03
GC_1_51 b_1 NI_1 NS_51 0 3.0136121802917678e-03
GC_1_52 b_1 NI_1 NS_52 0 1.9753011331270828e-03
GC_1_53 b_1 NI_1 NS_53 0 -7.8484592257623486e-04
GC_1_54 b_1 NI_1 NS_54 0 6.1124814411728961e-04
GC_1_55 b_1 NI_1 NS_55 0 8.7608535090844472e-03
GC_1_56 b_1 NI_1 NS_56 0 -3.9534026163486821e-03
GC_1_57 b_1 NI_1 NS_57 0 -3.2892178643368952e-04
GC_1_58 b_1 NI_1 NS_58 0 8.2757902794755383e-06
GC_1_59 b_1 NI_1 NS_59 0 9.9988229121495640e-06
GC_1_60 b_1 NI_1 NS_60 0 1.5012218523085316e-05
GC_1_61 b_1 NI_1 NS_61 0 2.9955075499348981e-04
GC_1_62 b_1 NI_1 NS_62 0 -4.5263075396487234e-04
GC_1_63 b_1 NI_1 NS_63 0 -2.0269373379274258e-05
GC_1_64 b_1 NI_1 NS_64 0 -6.4687750514096430e-06
GC_1_65 b_1 NI_1 NS_65 0 -4.1229530652186405e-05
GC_1_66 b_1 NI_1 NS_66 0 5.1554757324793720e-06
GC_1_67 b_1 NI_1 NS_67 0 2.5964432440410599e-06
GC_1_68 b_1 NI_1 NS_68 0 7.9589517337639512e-07
GC_1_69 b_1 NI_1 NS_69 0 -1.1855968523987400e-03
GC_1_70 b_1 NI_1 NS_70 0 -5.7443834716666064e-03
GC_1_71 b_1 NI_1 NS_71 0 -9.8027689212128275e-05
GC_1_72 b_1 NI_1 NS_72 0 1.9907089791670585e-03
GC_1_73 b_1 NI_1 NS_73 0 5.9227408808240692e-05
GC_1_74 b_1 NI_1 NS_74 0 1.6117214921916636e-04
GC_1_75 b_1 NI_1 NS_75 0 6.3385406661192562e-07
GC_1_76 b_1 NI_1 NS_76 0 8.8002356189512373e-07
GC_1_77 b_1 NI_1 NS_77 0 4.5772227914256818e-05
GC_1_78 b_1 NI_1 NS_78 0 -8.2453266528328140e-06
GC_1_79 b_1 NI_1 NS_79 0 1.0163799348693825e-06
GC_1_80 b_1 NI_1 NS_80 0 -7.4324831272045018e-07
GC_1_81 b_1 NI_1 NS_81 0 3.5658978991974893e-06
GC_1_82 b_1 NI_1 NS_82 0 -8.3880520348053317e-07
GC_1_83 b_1 NI_1 NS_83 0 3.0577508848793290e-05
GC_1_84 b_1 NI_1 NS_84 0 9.4492715199634829e-05
GC_1_85 b_1 NI_1 NS_85 0 1.8153377291647337e-06
GC_1_86 b_1 NI_1 NS_86 0 3.5496323331631462e-05
GC_1_87 b_1 NI_1 NS_87 0 7.6865786754466219e-06
GC_1_88 b_1 NI_1 NS_88 0 4.1806570153541225e-06
GC_1_89 b_1 NI_1 NS_89 0 8.1298888220752066e-03
GC_1_90 b_1 NI_1 NS_90 0 -4.6313664333942888e-04
GC_1_91 b_1 NI_1 NS_91 0 1.1775616910082772e-02
GC_1_92 b_1 NI_1 NS_92 0 3.4756009174440367e-03
GC_1_93 b_1 NI_1 NS_93 0 -9.1264956974332137e-03
GC_1_94 b_1 NI_1 NS_94 0 -8.4944380370542884e-03
GC_1_95 b_1 NI_1 NS_95 0 1.1666689942321673e-02
GC_1_96 b_1 NI_1 NS_96 0 7.1468101097935275e-03
GC_1_97 b_1 NI_1 NS_97 0 -2.9079236264730186e-03
GC_1_98 b_1 NI_1 NS_98 0 -1.1074628460343025e-03
GC_1_99 b_1 NI_1 NS_99 0 2.7737482651150102e-03
GC_1_100 b_1 NI_1 NS_100 0 2.8643816821392054e-03
GC_1_101 b_1 NI_1 NS_101 0 5.1414858487714755e-04
GC_1_102 b_1 NI_1 NS_102 0 4.4167817349773591e-04
GC_1_103 b_1 NI_1 NS_103 0 5.6985398085413060e-05
GC_1_104 b_1 NI_1 NS_104 0 1.9751981092293864e-04
GC_1_105 b_1 NI_1 NS_105 0 1.3150881529618360e-03
GC_1_106 b_1 NI_1 NS_106 0 3.6828708635683506e-04
GC_1_107 b_1 NI_1 NS_107 0 1.5243466980848852e-04
GC_1_108 b_1 NI_1 NS_108 0 1.4876395456431965e-04
GC_1_109 b_1 NI_1 NS_109 0 2.6549024590819112e-04
GC_1_110 b_1 NI_1 NS_110 0 4.3527186433841819e-05
GC_1_111 b_1 NI_1 NS_111 0 -1.0262837575083311e-05
GC_1_112 b_1 NI_1 NS_112 0 3.3651479283446454e-06
GC_1_113 b_1 NI_1 NS_113 0 -1.9801857301250596e-02
GC_1_114 b_1 NI_1 NS_114 0 7.5551435785673488e-03
GC_1_115 b_1 NI_1 NS_115 0 1.4228094632457770e-02
GC_1_116 b_1 NI_1 NS_116 0 1.1891842589361085e-03
GC_1_117 b_1 NI_1 NS_117 0 -4.2618652470487227e-04
GC_1_118 b_1 NI_1 NS_118 0 7.0823364160501036e-06
GC_1_119 b_1 NI_1 NS_119 0 1.6111007194803199e-06
GC_1_120 b_1 NI_1 NS_120 0 3.5599396390078671e-06
GC_1_121 b_1 NI_1 NS_121 0 2.1165662609029192e-04
GC_1_122 b_1 NI_1 NS_122 0 -1.8258783416698386e-05
GC_1_123 b_1 NI_1 NS_123 0 5.1141436212614634e-06
GC_1_124 b_1 NI_1 NS_124 0 9.6168016077313257e-07
GC_1_125 b_1 NI_1 NS_125 0 3.1338806345800870e-07
GC_1_126 b_1 NI_1 NS_126 0 7.9388977764005474e-07
GC_1_127 b_1 NI_1 NS_127 0 -2.8029008656075698e-04
GC_1_128 b_1 NI_1 NS_128 0 2.8861647396669874e-04
GC_1_129 b_1 NI_1 NS_129 0 -3.5661394941241958e-05
GC_1_130 b_1 NI_1 NS_130 0 -5.7109012747122068e-05
GC_1_131 b_1 NI_1 NS_131 0 -1.7863884658282121e-05
GC_1_132 b_1 NI_1 NS_132 0 1.0868955973749419e-05
GC_1_133 b_1 NI_1 NS_133 0 6.1783341262023617e-03
GC_1_134 b_1 NI_1 NS_134 0 -3.7221244443601308e-04
GC_1_135 b_1 NI_1 NS_135 0 -2.0234199944319631e-02
GC_1_136 b_1 NI_1 NS_136 0 -3.0973193626442417e-03
GC_1_137 b_1 NI_1 NS_137 0 1.0273186404537832e-02
GC_1_138 b_1 NI_1 NS_138 0 -3.0432489324587995e-03
GC_1_139 b_1 NI_1 NS_139 0 5.8008064102922858e-03
GC_1_140 b_1 NI_1 NS_140 0 1.0544994379758621e-03
GC_1_141 b_1 NI_1 NS_141 0 1.8472440092420148e-03
GC_1_142 b_1 NI_1 NS_142 0 -5.2924024160756289e-04
GC_1_143 b_1 NI_1 NS_143 0 -7.2836452790861885e-04
GC_1_144 b_1 NI_1 NS_144 0 -8.7666286246263977e-03
GC_1_145 b_1 NI_1 NS_145 0 -2.7303355822281021e-04
GC_1_146 b_1 NI_1 NS_146 0 3.8620741870170757e-05
GC_1_147 b_1 NI_1 NS_147 0 1.7685662290304582e-04
GC_1_148 b_1 NI_1 NS_148 0 6.2209955780299036e-05
GC_1_149 b_1 NI_1 NS_149 0 5.4327097672122538e-04
GC_1_150 b_1 NI_1 NS_150 0 4.8081377505014247e-04
GC_1_151 b_1 NI_1 NS_151 0 3.4810666064125838e-05
GC_1_152 b_1 NI_1 NS_152 0 3.3290197896397506e-05
GC_1_153 b_1 NI_1 NS_153 0 6.9368235382700775e-05
GC_1_154 b_1 NI_1 NS_154 0 1.1406950112113439e-05
GC_1_155 b_1 NI_1 NS_155 0 5.3522247266642766e-06
GC_1_156 b_1 NI_1 NS_156 0 -1.9451375007430333e-06
GC_1_157 b_1 NI_1 NS_157 0 -6.4795852496178233e-03
GC_1_158 b_1 NI_1 NS_158 0 8.1058085975704280e-03
GC_1_159 b_1 NI_1 NS_159 0 4.7484983140375003e-03
GC_1_160 b_1 NI_1 NS_160 0 -3.1909267764600019e-03
GC_1_161 b_1 NI_1 NS_161 0 -1.9213544848574831e-04
GC_1_162 b_1 NI_1 NS_162 0 1.8309860619107721e-04
GC_1_163 b_1 NI_1 NS_163 0 -5.3295997558524851e-07
GC_1_164 b_1 NI_1 NS_164 0 2.6108714931024329e-07
GC_1_165 b_1 NI_1 NS_165 0 8.9411675081290340e-06
GC_1_166 b_1 NI_1 NS_166 0 4.4378722599442055e-05
GC_1_167 b_1 NI_1 NS_167 0 1.0538695980854309e-07
GC_1_168 b_1 NI_1 NS_168 0 8.1440759073888631e-07
GC_1_169 b_1 NI_1 NS_169 0 1.6344353781495764e-07
GC_1_170 b_1 NI_1 NS_170 0 1.3798537923800453e-06
GC_1_171 b_1 NI_1 NS_171 0 -5.6397528022635824e-05
GC_1_172 b_1 NI_1 NS_172 0 -1.6206890529595931e-04
GC_1_173 b_1 NI_1 NS_173 0 -5.7041757645843857e-07
GC_1_174 b_1 NI_1 NS_174 0 -1.1831905612830878e-05
GC_1_175 b_1 NI_1 NS_175 0 -1.7424126407219506e-07
GC_1_176 b_1 NI_1 NS_176 0 -6.0528681451970242e-06
GC_1_177 b_1 NI_1 NS_177 0 1.4888401712570045e-02
GC_1_178 b_1 NI_1 NS_178 0 -9.3518480534758365e-06
GC_1_179 b_1 NI_1 NS_179 0 1.2024151653626705e-02
GC_1_180 b_1 NI_1 NS_180 0 -5.2254723615882516e-03
GC_1_181 b_1 NI_1 NS_181 0 -2.3071146560527970e-03
GC_1_182 b_1 NI_1 NS_182 0 5.8586359722771052e-03
GC_1_183 b_1 NI_1 NS_183 0 1.2364954931264561e-02
GC_1_184 b_1 NI_1 NS_184 0 9.2062676968266977e-03
GC_1_185 b_1 NI_1 NS_185 0 -2.2188545995756293e-03
GC_1_186 b_1 NI_1 NS_186 0 -3.0825900370840108e-03
GC_1_187 b_1 NI_1 NS_187 0 -1.0102730895459150e-02
GC_1_188 b_1 NI_1 NS_188 0 9.6134683530376529e-03
GC_1_189 b_1 NI_1 NS_189 0 5.4911431511251525e-04
GC_1_190 b_1 NI_1 NS_190 0 4.2797708634814441e-04
GC_1_191 b_1 NI_1 NS_191 0 5.5714477042035982e-05
GC_1_192 b_1 NI_1 NS_192 0 2.1799559001127664e-04
GC_1_193 b_1 NI_1 NS_193 0 1.3139424947679480e-03
GC_1_194 b_1 NI_1 NS_194 0 2.3427081311820565e-04
GC_1_195 b_1 NI_1 NS_195 0 1.5519461050893905e-04
GC_1_196 b_1 NI_1 NS_196 0 1.4245051926242515e-04
GC_1_197 b_1 NI_1 NS_197 0 2.3535465258341613e-04
GC_1_198 b_1 NI_1 NS_198 0 5.2771923484891158e-05
GC_1_199 b_1 NI_1 NS_199 0 -9.1466667977504430e-06
GC_1_200 b_1 NI_1 NS_200 0 3.9142335685442605e-06
GC_1_201 b_1 NI_1 NS_201 0 -2.4379490423038250e-02
GC_1_202 b_1 NI_1 NS_202 0 -9.8093355717727504e-04
GC_1_203 b_1 NI_1 NS_203 0 1.5256180092878166e-02
GC_1_204 b_1 NI_1 NS_204 0 3.8108865834751409e-03
GC_1_205 b_1 NI_1 NS_205 0 -3.4039717499606591e-04
GC_1_206 b_1 NI_1 NS_206 0 -4.8567332572583600e-04
GC_1_207 b_1 NI_1 NS_207 0 9.1459998020402380e-07
GC_1_208 b_1 NI_1 NS_208 0 4.5967216745145888e-07
GC_1_209 b_1 NI_1 NS_209 0 9.9142384636878480e-05
GC_1_210 b_1 NI_1 NS_210 0 -5.3583112263144498e-05
GC_1_211 b_1 NI_1 NS_211 0 2.1456157635949741e-06
GC_1_212 b_1 NI_1 NS_212 0 3.0865102073394589e-07
GC_1_213 b_1 NI_1 NS_213 0 -1.9245036014797487e-06
GC_1_214 b_1 NI_1 NS_214 0 -1.1735224944871366e-06
GC_1_215 b_1 NI_1 NS_215 0 -6.5682388735319270e-05
GC_1_216 b_1 NI_1 NS_216 0 2.1932692681570070e-04
GC_1_217 b_1 NI_1 NS_217 0 2.0903108903736811e-05
GC_1_218 b_1 NI_1 NS_218 0 -7.0297658116458324e-05
GC_1_219 b_1 NI_1 NS_219 0 -1.1994220959436528e-05
GC_1_220 b_1 NI_1 NS_220 0 -1.4131663487940362e-06
GC_1_221 b_1 NI_1 NS_221 0 1.4112468708626265e-02
GC_1_222 b_1 NI_1 NS_222 0 -6.0820585627260827e-04
GC_1_223 b_1 NI_1 NS_223 0 -1.5409865371543579e-02
GC_1_224 b_1 NI_1 NS_224 0 6.3372079764299006e-03
GC_1_225 b_1 NI_1 NS_225 0 2.3440157145016927e-03
GC_1_226 b_1 NI_1 NS_226 0 -1.2292674427882086e-02
GC_1_227 b_1 NI_1 NS_227 0 8.6622331958593514e-03
GC_1_228 b_1 NI_1 NS_228 0 9.3590176400180707e-04
GC_1_229 b_1 NI_1 NS_229 0 -4.2273216718384499e-04
GC_1_230 b_1 NI_1 NS_230 0 -6.2490282474047382e-04
GC_1_231 b_1 NI_1 NS_231 0 -7.4366755644213658e-03
GC_1_232 b_1 NI_1 NS_232 0 -2.5616625251912270e-03
GC_1_233 b_1 NI_1 NS_233 0 -2.8290821983849632e-04
GC_1_234 b_1 NI_1 NS_234 0 9.9873141396215521e-05
GC_1_235 b_1 NI_1 NS_235 0 1.4028345289088351e-04
GC_1_236 b_1 NI_1 NS_236 0 3.7184731672339288e-05
GC_1_237 b_1 NI_1 NS_237 0 6.0003137430693929e-04
GC_1_238 b_1 NI_1 NS_238 0 1.3116124746293231e-04
GC_1_239 b_1 NI_1 NS_239 0 2.6151008574512524e-05
GC_1_240 b_1 NI_1 NS_240 0 1.5509521873307654e-05
GC_1_241 b_1 NI_1 NS_241 0 5.2609416930533179e-05
GC_1_242 b_1 NI_1 NS_242 0 -1.6342984312418218e-05
GC_1_243 b_1 NI_1 NS_243 0 7.1935138306252046e-06
GC_1_244 b_1 NI_1 NS_244 0 -5.0563598437058948e-08
GC_1_245 b_1 NI_1 NS_245 0 -3.0349579133553446e-04
GC_1_246 b_1 NI_1 NS_246 0 3.1321499703077177e-03
GC_1_247 b_1 NI_1 NS_247 0 1.9318343152081399e-03
GC_1_248 b_1 NI_1 NS_248 0 -1.7750716646077051e-03
GC_1_249 b_1 NI_1 NS_249 0 1.7999948139396895e-05
GC_1_250 b_1 NI_1 NS_250 0 -2.6283026770074434e-05
GC_1_251 b_1 NI_1 NS_251 0 -1.5737649874605132e-07
GC_1_252 b_1 NI_1 NS_252 0 1.4176124851230246e-08
GC_1_253 b_1 NI_1 NS_253 0 5.8309901269895959e-06
GC_1_254 b_1 NI_1 NS_254 0 -1.3992874587997102e-05
GC_1_255 b_1 NI_1 NS_255 0 9.3550153846168259e-08
GC_1_256 b_1 NI_1 NS_256 0 -6.2686481096018683e-07
GC_1_257 b_1 NI_1 NS_257 0 3.1536238724812709e-06
GC_1_258 b_1 NI_1 NS_258 0 2.3639585707507269e-07
GC_1_259 b_1 NI_1 NS_259 0 -2.5270305902353794e-06
GC_1_260 b_1 NI_1 NS_260 0 2.8776869288048998e-05
GC_1_261 b_1 NI_1 NS_261 0 1.3870237329924348e-05
GC_1_262 b_1 NI_1 NS_262 0 1.4507190030789509e-05
GC_1_263 b_1 NI_1 NS_263 0 6.2453973555449024e-06
GC_1_264 b_1 NI_1 NS_264 0 -1.5536764595768147e-06
GC_1_265 b_1 NI_1 NS_265 0 8.0678348141457641e-03
GC_1_266 b_1 NI_1 NS_266 0 2.4279265951733791e-04
GC_1_267 b_1 NI_1 NS_267 0 7.0724015355786941e-03
GC_1_268 b_1 NI_1 NS_268 0 -7.0940926046937879e-03
GC_1_269 b_1 NI_1 NS_269 0 3.3452930912154588e-03
GC_1_270 b_1 NI_1 NS_270 0 7.8189965493129648e-03
GC_1_271 b_1 NI_1 NS_271 0 9.6302829097826594e-03
GC_1_272 b_1 NI_1 NS_272 0 7.7632217464532671e-03
GC_1_273 b_1 NI_1 NS_273 0 2.1695161318018593e-05
GC_1_274 b_1 NI_1 NS_274 0 -3.7467283856288552e-03
GC_1_275 b_1 NI_1 NS_275 0 -1.3029598792569605e-02
GC_1_276 b_1 NI_1 NS_276 0 1.1815842226091312e-02
GC_1_277 b_1 NI_1 NS_277 0 4.2549892168000208e-04
GC_1_278 b_1 NI_1 NS_278 0 2.9282716494632435e-04
GC_1_279 b_1 NI_1 NS_279 0 3.6567343485997414e-05
GC_1_280 b_1 NI_1 NS_280 0 2.2547725912692112e-04
GC_1_281 b_1 NI_1 NS_281 0 5.2629767312833791e-04
GC_1_282 b_1 NI_1 NS_282 0 -2.7813714694770235e-04
GC_1_283 b_1 NI_1 NS_283 0 9.5387529800183244e-05
GC_1_284 b_1 NI_1 NS_284 0 1.1274327254584181e-04
GC_1_285 b_1 NI_1 NS_285 0 4.5339081751403269e-05
GC_1_286 b_1 NI_1 NS_286 0 5.4219000620817888e-05
GC_1_287 b_1 NI_1 NS_287 0 -6.6504745767958741e-06
GC_1_288 b_1 NI_1 NS_288 0 2.6857297221450307e-06
GC_1_289 b_1 NI_1 NS_289 0 -1.8209602962116735e-02
GC_1_290 b_1 NI_1 NS_290 0 -7.7990122981907804e-03
GC_1_291 b_1 NI_1 NS_291 0 9.6141322539995602e-03
GC_1_292 b_1 NI_1 NS_292 0 5.1853209234903296e-03
GC_1_293 b_1 NI_1 NS_293 0 -1.6326950250393851e-04
GC_1_294 b_1 NI_1 NS_294 0 -4.4113601250572910e-04
GC_1_295 b_1 NI_1 NS_295 0 7.8930443643209364e-07
GC_1_296 b_1 NI_1 NS_296 0 2.8147367235529219e-08
GC_1_297 b_1 NI_1 NS_297 0 4.8560994068505668e-05
GC_1_298 b_1 NI_1 NS_298 0 -5.4730653968521439e-05
GC_1_299 b_1 NI_1 NS_299 0 1.1114820923313135e-06
GC_1_300 b_1 NI_1 NS_300 0 -1.3801920749458200e-07
GC_1_301 b_1 NI_1 NS_301 0 -8.9165880659614363e-07
GC_1_302 b_1 NI_1 NS_302 0 -2.6989598376219689e-06
GC_1_303 b_1 NI_1 NS_303 0 6.8568315591389513e-05
GC_1_304 b_1 NI_1 NS_304 0 2.0889738559935357e-04
GC_1_305 b_1 NI_1 NS_305 0 1.4083727125783209e-05
GC_1_306 b_1 NI_1 NS_306 0 -2.8696275950965869e-05
GC_1_307 b_1 NI_1 NS_307 0 -3.8665155973613518e-06
GC_1_308 b_1 NI_1 NS_308 0 -1.4059424596684468e-06
GC_1_309 b_1 NI_1 NS_309 0 2.2701383137628643e-02
GC_1_310 b_1 NI_1 NS_310 0 -5.3164488024146821e-04
GC_1_311 b_1 NI_1 NS_311 0 -6.5503786045686520e-03
GC_1_312 b_1 NI_1 NS_312 0 8.2362773686277067e-03
GC_1_313 b_1 NI_1 NS_313 0 -3.6090198409885889e-03
GC_1_314 b_1 NI_1 NS_314 0 -8.8590221970589085e-03
GC_1_315 b_1 NI_1 NS_315 0 6.1402281782433126e-03
GC_1_316 b_1 NI_1 NS_316 0 4.8129312488777920e-04
GC_1_317 b_1 NI_1 NS_317 0 -1.6902783599214053e-03
GC_1_318 b_1 NI_1 NS_318 0 4.3909960252311818e-04
GC_1_319 b_1 NI_1 NS_319 0 -8.2254729575620272e-03
GC_1_320 b_1 NI_1 NS_320 0 2.8484432460413401e-03
GC_1_321 b_1 NI_1 NS_321 0 -1.6753675302598884e-04
GC_1_322 b_1 NI_1 NS_322 0 1.1463757082194408e-04
GC_1_323 b_1 NI_1 NS_323 0 1.0497005236795980e-04
GC_1_324 b_1 NI_1 NS_324 0 7.3248079190093502e-05
GC_1_325 b_1 NI_1 NS_325 0 4.3404098276911436e-05
GC_1_326 b_1 NI_1 NS_326 0 5.1326448046175427e-05
GC_1_327 b_1 NI_1 NS_327 0 -1.3610507749467718e-05
GC_1_328 b_1 NI_1 NS_328 0 2.9465331778450115e-05
GC_1_329 b_1 NI_1 NS_329 0 -7.8793111364567717e-06
GC_1_330 b_1 NI_1 NS_330 0 4.3639231679860992e-05
GC_1_331 b_1 NI_1 NS_331 0 3.3150395651007460e-06
GC_1_332 b_1 NI_1 NS_332 0 2.7916137090825528e-06
GC_1_333 b_1 NI_1 NS_333 0 -2.6241609612349980e-04
GC_1_334 b_1 NI_1 NS_334 0 -3.6640709711493261e-03
GC_1_335 b_1 NI_1 NS_335 0 1.0167936237335559e-03
GC_1_336 b_1 NI_1 NS_336 0 1.5016845663790373e-03
GC_1_337 b_1 NI_1 NS_337 0 2.3407575291024233e-04
GC_1_338 b_1 NI_1 NS_338 0 -3.3545074027293935e-04
GC_1_339 b_1 NI_1 NS_339 0 1.2063665016216471e-06
GC_1_340 b_1 NI_1 NS_340 0 -1.5445557228171482e-06
GC_1_341 b_1 NI_1 NS_341 0 -3.7386760436604566e-05
GC_1_342 b_1 NI_1 NS_342 0 -8.1394976865457761e-05
GC_1_343 b_1 NI_1 NS_343 0 -5.8536822359219638e-07
GC_1_344 b_1 NI_1 NS_344 0 -2.1526513364026869e-06
GC_1_345 b_1 NI_1 NS_345 0 2.0405916682026597e-06
GC_1_346 b_1 NI_1 NS_346 0 -2.6188172796139417e-06
GC_1_347 b_1 NI_1 NS_347 0 1.4986989963705757e-04
GC_1_348 b_1 NI_1 NS_348 0 9.1312796747941829e-05
GC_1_349 b_1 NI_1 NS_349 0 4.3196311352403608e-05
GC_1_350 b_1 NI_1 NS_350 0 4.3611220708109232e-05
GC_1_351 b_1 NI_1 NS_351 0 1.5167024618325218e-05
GC_1_352 b_1 NI_1 NS_352 0 -9.5060022847269482e-07
GC_1_353 b_1 NI_1 NS_353 0 -1.1394110043614361e-02
GC_1_354 b_1 NI_1 NS_354 0 5.3879744221281325e-05
GC_1_355 b_1 NI_1 NS_355 0 -9.8723080462374910e-04
GC_1_356 b_1 NI_1 NS_356 0 -6.7885736986834509e-04
GC_1_357 b_1 NI_1 NS_357 0 2.7015328322856986e-04
GC_1_358 b_1 NI_1 NS_358 0 -1.8137468306988265e-03
GC_1_359 b_1 NI_1 NS_359 0 9.8065716253669896e-04
GC_1_360 b_1 NI_1 NS_360 0 -2.1464622949615478e-03
GC_1_361 b_1 NI_1 NS_361 0 3.6936230799238602e-04
GC_1_362 b_1 NI_1 NS_362 0 1.3125386895614379e-03
GC_1_363 b_1 NI_1 NS_363 0 3.9409123339799630e-04
GC_1_364 b_1 NI_1 NS_364 0 -2.7742375994508836e-04
GC_1_365 b_1 NI_1 NS_365 0 3.4404789774480584e-04
GC_1_366 b_1 NI_1 NS_366 0 -2.7109771613113669e-04
GC_1_367 b_1 NI_1 NS_367 0 2.9707605304676187e-04
GC_1_368 b_1 NI_1 NS_368 0 6.0787934286053952e-04
GC_1_369 b_1 NI_1 NS_369 0 -1.9167768098630783e-03
GC_1_370 b_1 NI_1 NS_370 0 -1.5694669517797824e-03
GC_1_371 b_1 NI_1 NS_371 0 1.4566888759792151e-04
GC_1_372 b_1 NI_1 NS_372 0 9.4418302102695863e-05
GC_1_373 b_1 NI_1 NS_373 0 -7.5079176415194615e-04
GC_1_374 b_1 NI_1 NS_374 0 -2.6223496032023137e-06
GC_1_375 b_1 NI_1 NS_375 0 -1.7724531171575323e-06
GC_1_376 b_1 NI_1 NS_376 0 -4.1820800005490387e-06
GC_1_377 b_1 NI_1 NS_377 0 1.1962236119654333e-02
GC_1_378 b_1 NI_1 NS_378 0 7.5139379540347462e-03
GC_1_379 b_1 NI_1 NS_379 0 -5.7663301145365938e-03
GC_1_380 b_1 NI_1 NS_380 0 -8.4439103321084178e-03
GC_1_381 b_1 NI_1 NS_381 0 5.0316366105401133e-05
GC_1_382 b_1 NI_1 NS_382 0 2.4328749992233735e-04
GC_1_383 b_1 NI_1 NS_383 0 4.7883113127596043e-08
GC_1_384 b_1 NI_1 NS_384 0 -1.9304201919006067e-07
GC_1_385 b_1 NI_1 NS_385 0 -1.6233474382980237e-05
GC_1_386 b_1 NI_1 NS_386 0 -7.3436249902549452e-05
GC_1_387 b_1 NI_1 NS_387 0 -3.9354883773914403e-09
GC_1_388 b_1 NI_1 NS_388 0 1.2088391620714307e-07
GC_1_389 b_1 NI_1 NS_389 0 -6.8269680056045362e-07
GC_1_390 b_1 NI_1 NS_390 0 -3.5484685237805144e-06
GC_1_391 b_1 NI_1 NS_391 0 2.3502666210701279e-04
GC_1_392 b_1 NI_1 NS_392 0 4.0007149268351529e-04
GC_1_393 b_1 NI_1 NS_393 0 -1.4727562969123859e-04
GC_1_394 b_1 NI_1 NS_394 0 8.1879697462817352e-05
GC_1_395 b_1 NI_1 NS_395 0 -1.1231031129461442e-05
GC_1_396 b_1 NI_1 NS_396 0 -7.4139974408313973e-06
GC_1_397 b_1 NI_1 NS_397 0 -3.1343479687062589e-03
GC_1_398 b_1 NI_1 NS_398 0 4.3166440025267355e-05
GC_1_399 b_1 NI_1 NS_399 0 -1.5455853079215230e-05
GC_1_400 b_1 NI_1 NS_400 0 3.6118218364002911e-04
GC_1_401 b_1 NI_1 NS_401 0 -1.0071123414497713e-03
GC_1_402 b_1 NI_1 NS_402 0 -4.2339505591776035e-04
GC_1_403 b_1 NI_1 NS_403 0 -2.5534355234792277e-04
GC_1_404 b_1 NI_1 NS_404 0 -1.4776842959832056e-03
GC_1_405 b_1 NI_1 NS_405 0 2.8524762423597349e-04
GC_1_406 b_1 NI_1 NS_406 0 -5.0422578116772708e-05
GC_1_407 b_1 NI_1 NS_407 0 1.4139041255064962e-03
GC_1_408 b_1 NI_1 NS_408 0 -1.2322107141048667e-03
GC_1_409 b_1 NI_1 NS_409 0 -4.2027475770706194e-06
GC_1_410 b_1 NI_1 NS_410 0 1.8839119023427860e-04
GC_1_411 b_1 NI_1 NS_411 0 2.1091379052460286e-04
GC_1_412 b_1 NI_1 NS_412 0 -7.3898888176833312e-05
GC_1_413 b_1 NI_1 NS_413 0 -2.0294948991884178e-04
GC_1_414 b_1 NI_1 NS_414 0 6.1533548752831148e-05
GC_1_415 b_1 NI_1 NS_415 0 -8.6801400473590279e-06
GC_1_416 b_1 NI_1 NS_416 0 -1.1110998475024373e-05
GC_1_417 b_1 NI_1 NS_417 0 -2.9359761558843366e-05
GC_1_418 b_1 NI_1 NS_418 0 -5.7334880719555747e-05
GC_1_419 b_1 NI_1 NS_419 0 3.5413081315423038e-06
GC_1_420 b_1 NI_1 NS_420 0 3.0127554939014840e-06
GC_1_421 b_1 NI_1 NS_421 0 2.4421199316424971e-03
GC_1_422 b_1 NI_1 NS_422 0 3.7498088124294235e-03
GC_1_423 b_1 NI_1 NS_423 0 -1.4394589167904400e-03
GC_1_424 b_1 NI_1 NS_424 0 -2.8128705914642000e-03
GC_1_425 b_1 NI_1 NS_425 0 -1.4192475295535299e-04
GC_1_426 b_1 NI_1 NS_426 0 2.9433315895404518e-05
GC_1_427 b_1 NI_1 NS_427 0 -6.2237066143647369e-07
GC_1_428 b_1 NI_1 NS_428 0 1.3836169282128862e-07
GC_1_429 b_1 NI_1 NS_429 0 -1.6028860889443415e-05
GC_1_430 b_1 NI_1 NS_430 0 3.0736977570038202e-05
GC_1_431 b_1 NI_1 NS_431 0 -6.8950972062654289e-07
GC_1_432 b_1 NI_1 NS_432 0 7.1768388345691796e-07
GC_1_433 b_1 NI_1 NS_433 0 1.3589709023695545e-06
GC_1_434 b_1 NI_1 NS_434 0 1.0565294902679273e-06
GC_1_435 b_1 NI_1 NS_435 0 -6.0861550190567712e-05
GC_1_436 b_1 NI_1 NS_436 0 -9.6861852872016398e-05
GC_1_437 b_1 NI_1 NS_437 0 -3.3346111761257571e-07
GC_1_438 b_1 NI_1 NS_438 0 -4.3028551479207985e-05
GC_1_439 b_1 NI_1 NS_439 0 -8.2481922745260886e-06
GC_1_440 b_1 NI_1 NS_440 0 -3.2058185792641375e-06
GC_1_441 b_1 NI_1 NS_441 0 -5.2728379851390951e-03
GC_1_442 b_1 NI_1 NS_442 0 6.6652010760696951e-05
GC_1_443 b_1 NI_1 NS_443 0 -1.8650511765668830e-04
GC_1_444 b_1 NI_1 NS_444 0 -1.6783837526660901e-03
GC_1_445 b_1 NI_1 NS_445 0 1.6669619891636919e-03
GC_1_446 b_1 NI_1 NS_446 0 -3.8660493333036414e-04
GC_1_447 b_1 NI_1 NS_447 0 2.7653820693808551e-03
GC_1_448 b_1 NI_1 NS_448 0 -2.5015957562632570e-04
GC_1_449 b_1 NI_1 NS_449 0 -1.5644520406418426e-05
GC_1_450 b_1 NI_1 NS_450 0 -3.9238276287391490e-04
GC_1_451 b_1 NI_1 NS_451 0 -1.3578920610215826e-03
GC_1_452 b_1 NI_1 NS_452 0 3.8126783621767069e-03
GC_1_453 b_1 NI_1 NS_453 0 3.2378883776581515e-04
GC_1_454 b_1 NI_1 NS_454 0 -1.2353992539101901e-04
GC_1_455 b_1 NI_1 NS_455 0 2.0787701516574393e-04
GC_1_456 b_1 NI_1 NS_456 0 4.4667844758288378e-04
GC_1_457 b_1 NI_1 NS_457 0 -1.2761648388074386e-03
GC_1_458 b_1 NI_1 NS_458 0 -9.8061163894445761e-04
GC_1_459 b_1 NI_1 NS_459 0 1.1216839679871414e-04
GC_1_460 b_1 NI_1 NS_460 0 9.3592020019612698e-05
GC_1_461 b_1 NI_1 NS_461 0 -4.7341479107555328e-04
GC_1_462 b_1 NI_1 NS_462 0 2.2669963689706983e-05
GC_1_463 b_1 NI_1 NS_463 0 -5.5281583023757830e-07
GC_1_464 b_1 NI_1 NS_464 0 -1.7254423011113106e-06
GC_1_465 b_1 NI_1 NS_465 0 2.1479258693215468e-03
GC_1_466 b_1 NI_1 NS_466 0 2.2662692730022276e-03
GC_1_467 b_1 NI_1 NS_467 0 -1.3144167372655499e-03
GC_1_468 b_1 NI_1 NS_468 0 -3.3437514675795947e-03
GC_1_469 b_1 NI_1 NS_469 0 1.6784150063476518e-04
GC_1_470 b_1 NI_1 NS_470 0 -1.5986954132866861e-05
GC_1_471 b_1 NI_1 NS_471 0 2.4682982794833708e-07
GC_1_472 b_1 NI_1 NS_472 0 -6.2979471668028603e-07
GC_1_473 b_1 NI_1 NS_473 0 -1.4337043230964107e-05
GC_1_474 b_1 NI_1 NS_474 0 -7.8788469384490469e-05
GC_1_475 b_1 NI_1 NS_475 0 -2.3683908205165199e-07
GC_1_476 b_1 NI_1 NS_476 0 -2.8911465589641870e-07
GC_1_477 b_1 NI_1 NS_477 0 1.7114269742106722e-07
GC_1_478 b_1 NI_1 NS_478 0 -3.3079790040188181e-06
GC_1_479 b_1 NI_1 NS_479 0 1.9489788625287637e-04
GC_1_480 b_1 NI_1 NS_480 0 3.1959820887115874e-04
GC_1_481 b_1 NI_1 NS_481 0 -8.8378534469255054e-05
GC_1_482 b_1 NI_1 NS_482 0 5.7728659906366809e-05
GC_1_483 b_1 NI_1 NS_483 0 -6.2930208988201608e-06
GC_1_484 b_1 NI_1 NS_484 0 -3.8929526763718285e-06
GC_1_485 b_1 NI_1 NS_485 0 4.8531323672040732e-03
GC_1_486 b_1 NI_1 NS_486 0 -4.3649876182272713e-05
GC_1_487 b_1 NI_1 NS_487 0 -6.6864802960614627e-05
GC_1_488 b_1 NI_1 NS_488 0 1.5061862253044544e-03
GC_1_489 b_1 NI_1 NS_489 0 -1.7559778821092454e-03
GC_1_490 b_1 NI_1 NS_490 0 -7.3998463627203046e-04
GC_1_491 b_1 NI_1 NS_491 0 8.2701923893373610e-04
GC_1_492 b_1 NI_1 NS_492 0 -9.5862125467570771e-04
GC_1_493 b_1 NI_1 NS_493 0 2.8332973984580629e-05
GC_1_494 b_1 NI_1 NS_494 0 6.3430913103488715e-05
GC_1_495 b_1 NI_1 NS_495 0 -7.5167401952528709e-05
GC_1_496 b_1 NI_1 NS_496 0 1.2237696843845757e-03
GC_1_497 b_1 NI_1 NS_497 0 3.1295802906703283e-06
GC_1_498 b_1 NI_1 NS_498 0 1.3610040821242987e-04
GC_1_499 b_1 NI_1 NS_499 0 1.8544849033468971e-04
GC_1_500 b_1 NI_1 NS_500 0 -1.1512465199303198e-05
GC_1_501 b_1 NI_1 NS_501 0 -2.2096326155138617e-04
GC_1_502 b_1 NI_1 NS_502 0 2.0637401549837415e-04
GC_1_503 b_1 NI_1 NS_503 0 -4.5355204772623325e-06
GC_1_504 b_1 NI_1 NS_504 0 7.2572664302174422e-06
GC_1_505 b_1 NI_1 NS_505 0 2.1469900450855620e-05
GC_1_506 b_1 NI_1 NS_506 0 -6.1794067795436315e-06
GC_1_507 b_1 NI_1 NS_507 0 4.1879283530566809e-06
GC_1_508 b_1 NI_1 NS_508 0 1.3813530524267100e-06
GC_1_509 b_1 NI_1 NS_509 0 -1.7205037505914646e-03
GC_1_510 b_1 NI_1 NS_510 0 1.4659569926866577e-03
GC_1_511 b_1 NI_1 NS_511 0 8.3740845337352458e-04
GC_1_512 b_1 NI_1 NS_512 0 -1.2555801941269420e-03
GC_1_513 b_1 NI_1 NS_513 0 -1.7267001986613162e-04
GC_1_514 b_1 NI_1 NS_514 0 -2.7959000143023465e-04
GC_1_515 b_1 NI_1 NS_515 0 -1.2052302118934511e-06
GC_1_516 b_1 NI_1 NS_516 0 -1.0332950312593623e-06
GC_1_517 b_1 NI_1 NS_517 0 -7.1020870973064227e-05
GC_1_518 b_1 NI_1 NS_518 0 1.4818226572466409e-05
GC_1_519 b_1 NI_1 NS_519 0 -1.8516952569772968e-06
GC_1_520 b_1 NI_1 NS_520 0 4.7519720394401016e-07
GC_1_521 b_1 NI_1 NS_521 0 -4.6311545253186130e-07
GC_1_522 b_1 NI_1 NS_522 0 -2.0724548996688425e-07
GC_1_523 b_1 NI_1 NS_523 0 4.7433695819711404e-05
GC_1_524 b_1 NI_1 NS_524 0 -1.2704949864192241e-04
GC_1_525 b_1 NI_1 NS_525 0 3.5458474176558653e-05
GC_1_526 b_1 NI_1 NS_526 0 -3.7224988754102263e-05
GC_1_527 b_1 NI_1 NS_527 0 9.7157724399002540e-08
GC_1_528 b_1 NI_1 NS_528 0 -7.8350613330076529e-06
GD_1_1 b_1 NI_1 NA_1 0 -1.6994685476604068e-01
GD_1_2 b_1 NI_1 NA_2 0 -7.2737643139208254e-03
GD_1_3 b_1 NI_1 NA_3 0 -2.4065254918707452e-02
GD_1_4 b_1 NI_1 NA_4 0 -2.5623308108879725e-03
GD_1_5 b_1 NI_1 NA_5 0 -2.2869906298704432e-02
GD_1_6 b_1 NI_1 NA_6 0 -3.5671852665028476e-03
GD_1_7 b_1 NI_1 NA_7 0 -9.0786133963413895e-03
GD_1_8 b_1 NI_1 NA_8 0 -9.8904579298554098e-03
GD_1_9 b_1 NI_1 NA_9 0 5.9829461828021426e-03
GD_1_10 b_1 NI_1 NA_10 0 1.9716467045851073e-03
GD_1_11 b_1 NI_1 NA_11 0 2.8504604616393773e-03
GD_1_12 b_1 NI_1 NA_12 0 -3.1612752692549476e-03
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 2.6054150235727477e-02
GC_2_2 b_2 NI_2 NS_2 0 1.6788223938156870e-02
GC_2_3 b_2 NI_2 NS_3 0 -1.9815077026463832e-02
GC_2_4 b_2 NI_2 NS_4 0 -7.4654803423542023e-03
GC_2_5 b_2 NI_2 NS_5 0 -2.6099780470205947e-02
GC_2_6 b_2 NI_2 NS_6 0 2.0041949380722301e-03
GC_2_7 b_2 NI_2 NS_7 0 3.0136121802909182e-03
GC_2_8 b_2 NI_2 NS_8 0 1.9753011331232408e-03
GC_2_9 b_2 NI_2 NS_9 0 -7.8484592257605618e-04
GC_2_10 b_2 NI_2 NS_10 0 6.1124814411662239e-04
GC_2_11 b_2 NI_2 NS_11 0 8.7608535090856823e-03
GC_2_12 b_2 NI_2 NS_12 0 -3.9534026163520605e-03
GC_2_13 b_2 NI_2 NS_13 0 -3.2892178643374753e-04
GC_2_14 b_2 NI_2 NS_14 0 8.2757902795996930e-06
GC_2_15 b_2 NI_2 NS_15 0 9.9988229120235289e-06
GC_2_16 b_2 NI_2 NS_16 0 1.5012218523080896e-05
GC_2_17 b_2 NI_2 NS_17 0 2.9955075499360376e-04
GC_2_18 b_2 NI_2 NS_18 0 -4.5263075396561610e-04
GC_2_19 b_2 NI_2 NS_19 0 -2.0269373379336369e-05
GC_2_20 b_2 NI_2 NS_20 0 -6.4687750515035764e-06
GC_2_21 b_2 NI_2 NS_21 0 -4.1229530652352546e-05
GC_2_22 b_2 NI_2 NS_22 0 5.1554757321768398e-06
GC_2_23 b_2 NI_2 NS_23 0 2.5964432440468947e-06
GC_2_24 b_2 NI_2 NS_24 0 7.9589517332092822e-07
GC_2_25 b_2 NI_2 NS_25 0 -1.1855968523976405e-03
GC_2_26 b_2 NI_2 NS_26 0 -5.7443834716576396e-03
GC_2_27 b_2 NI_2 NS_27 0 -9.8027689211408216e-05
GC_2_28 b_2 NI_2 NS_28 0 1.9907089791606253e-03
GC_2_29 b_2 NI_2 NS_29 0 5.9227408808219963e-05
GC_2_30 b_2 NI_2 NS_30 0 1.6117214921890916e-04
GC_2_31 b_2 NI_2 NS_31 0 6.3385406661234924e-07
GC_2_32 b_2 NI_2 NS_32 0 8.8002356189340743e-07
GC_2_33 b_2 NI_2 NS_33 0 4.5772227914172047e-05
GC_2_34 b_2 NI_2 NS_34 0 -8.2453266528496242e-06
GC_2_35 b_2 NI_2 NS_35 0 1.0163799348665306e-06
GC_2_36 b_2 NI_2 NS_36 0 -7.4324831272093161e-07
GC_2_37 b_2 NI_2 NS_37 0 3.5658978991896860e-06
GC_2_38 b_2 NI_2 NS_38 0 -8.3880520348095023e-07
GC_2_39 b_2 NI_2 NS_39 0 3.0577508848858627e-05
GC_2_40 b_2 NI_2 NS_40 0 9.4492715199276297e-05
GC_2_41 b_2 NI_2 NS_41 0 1.8153377292163678e-06
GC_2_42 b_2 NI_2 NS_42 0 3.5496323331577448e-05
GC_2_43 b_2 NI_2 NS_43 0 7.6865786754472216e-06
GC_2_44 b_2 NI_2 NS_44 0 4.1806570153343799e-06
GC_2_45 b_2 NI_2 NS_45 0 -1.4008600562148757e-01
GC_2_46 b_2 NI_2 NS_46 0 1.7632963558765258e-02
GC_2_47 b_2 NI_2 NS_47 0 9.5238590064089263e-03
GC_2_48 b_2 NI_2 NS_48 0 1.3521040754311981e-02
GC_2_49 b_2 NI_2 NS_49 0 1.5594276588744816e-02
GC_2_50 b_2 NI_2 NS_50 0 -1.4204990532941886e-02
GC_2_51 b_2 NI_2 NS_51 0 1.6226179525247999e-03
GC_2_52 b_2 NI_2 NS_52 0 1.6812665210287068e-03
GC_2_53 b_2 NI_2 NS_53 0 -4.5405977652696733e-04
GC_2_54 b_2 NI_2 NS_54 0 5.7416874755289395e-04
GC_2_55 b_2 NI_2 NS_55 0 7.1074520791293760e-03
GC_2_56 b_2 NI_2 NS_56 0 1.2093229400524127e-03
GC_2_57 b_2 NI_2 NS_57 0 -2.3732099396169629e-05
GC_2_58 b_2 NI_2 NS_58 0 -1.7290906670258170e-04
GC_2_59 b_2 NI_2 NS_59 0 9.4200963375240309e-06
GC_2_60 b_2 NI_2 NS_60 0 -7.5367264384286340e-05
GC_2_61 b_2 NI_2 NS_61 0 2.3555669437313784e-04
GC_2_62 b_2 NI_2 NS_62 0 -5.0865227051055740e-05
GC_2_63 b_2 NI_2 NS_63 0 3.1024641195773919e-05
GC_2_64 b_2 NI_2 NS_64 0 -7.1134141076144529e-06
GC_2_65 b_2 NI_2 NS_65 0 4.4845845872393459e-05
GC_2_66 b_2 NI_2 NS_66 0 -1.9537249679662680e-05
GC_2_67 b_2 NI_2 NS_67 0 -9.9724409092317106e-07
GC_2_68 b_2 NI_2 NS_68 0 -2.1164557001458051e-06
GC_2_69 b_2 NI_2 NS_69 0 -1.8311962418613157e-03
GC_2_70 b_2 NI_2 NS_70 0 7.0353046360815087e-03
GC_2_71 b_2 NI_2 NS_71 0 1.2721201459331632e-03
GC_2_72 b_2 NI_2 NS_72 0 -3.2019270036965919e-03
GC_2_73 b_2 NI_2 NS_73 0 -1.3876171904109511e-04
GC_2_74 b_2 NI_2 NS_74 0 -3.2605284818174892e-04
GC_2_75 b_2 NI_2 NS_75 0 4.5469557344470563e-07
GC_2_76 b_2 NI_2 NS_76 0 -2.5017681815488596e-06
GC_2_77 b_2 NI_2 NS_77 0 -1.6268174391672360e-04
GC_2_78 b_2 NI_2 NS_78 0 5.4454545646035412e-05
GC_2_79 b_2 NI_2 NS_79 0 -5.8520043135856766e-06
GC_2_80 b_2 NI_2 NS_80 0 -3.0719991152577681e-06
GC_2_81 b_2 NI_2 NS_81 0 -8.4923725691935963e-06
GC_2_82 b_2 NI_2 NS_82 0 -1.2554464125919406e-05
GC_2_83 b_2 NI_2 NS_83 0 -1.2036466225581497e-04
GC_2_84 b_2 NI_2 NS_84 0 -1.2869312766000541e-04
GC_2_85 b_2 NI_2 NS_85 0 -5.9709835854079256e-05
GC_2_86 b_2 NI_2 NS_86 0 -8.6732261270408976e-05
GC_2_87 b_2 NI_2 NS_87 0 -2.7299448823644768e-05
GC_2_88 b_2 NI_2 NS_88 0 -2.6571473946958882e-05
GC_2_89 b_2 NI_2 NS_89 0 4.1353853743958538e-03
GC_2_90 b_2 NI_2 NS_90 0 -3.8950436030148693e-04
GC_2_91 b_2 NI_2 NS_91 0 -2.0786969519512602e-02
GC_2_92 b_2 NI_2 NS_92 0 -3.3764631098210335e-03
GC_2_93 b_2 NI_2 NS_93 0 1.0882611112276171e-02
GC_2_94 b_2 NI_2 NS_94 0 -3.7983016640820762e-03
GC_2_95 b_2 NI_2 NS_95 0 6.3210213390043337e-03
GC_2_96 b_2 NI_2 NS_96 0 1.0575600338919987e-03
GC_2_97 b_2 NI_2 NS_97 0 1.7290934516663930e-03
GC_2_98 b_2 NI_2 NS_98 0 1.1711422664196080e-04
GC_2_99 b_2 NI_2 NS_99 0 -8.1541195205128898e-04
GC_2_100 b_2 NI_2 NS_100 0 -8.9796307251469153e-03
GC_2_101 b_2 NI_2 NS_101 0 -2.5676279977737460e-04
GC_2_102 b_2 NI_2 NS_102 0 5.5670860307613811e-05
GC_2_103 b_2 NI_2 NS_103 0 1.8232763210359546e-04
GC_2_104 b_2 NI_2 NS_104 0 4.8224998791132962e-05
GC_2_105 b_2 NI_2 NS_105 0 5.2801459320035672e-04
GC_2_106 b_2 NI_2 NS_106 0 4.1049378120135805e-04
GC_2_107 b_2 NI_2 NS_107 0 3.6402264054781473e-05
GC_2_108 b_2 NI_2 NS_108 0 2.2720379219466765e-05
GC_2_109 b_2 NI_2 NS_109 0 7.2644729265672282e-05
GC_2_110 b_2 NI_2 NS_110 0 -2.6561525809493270e-06
GC_2_111 b_2 NI_2 NS_111 0 7.1455434930228357e-06
GC_2_112 b_2 NI_2 NS_112 0 -2.6258464294494502e-06
GC_2_113 b_2 NI_2 NS_113 0 -4.2482848656284376e-03
GC_2_114 b_2 NI_2 NS_114 0 8.4802273171719171e-03
GC_2_115 b_2 NI_2 NS_115 0 3.6436292071362728e-03
GC_2_116 b_2 NI_2 NS_116 0 -3.6565506073502506e-03
GC_2_117 b_2 NI_2 NS_117 0 -1.7806454419374429e-04
GC_2_118 b_2 NI_2 NS_118 0 1.9560305428955595e-04
GC_2_119 b_2 NI_2 NS_119 0 -5.5118032007160593e-07
GC_2_120 b_2 NI_2 NS_120 0 8.4487321428819754e-07
GC_2_121 b_2 NI_2 NS_121 0 2.3642872544096086e-05
GC_2_122 b_2 NI_2 NS_122 0 5.7969512907821284e-05
GC_2_123 b_2 NI_2 NS_123 0 -3.6087148457955340e-07
GC_2_124 b_2 NI_2 NS_124 0 8.1753374210639751e-07
GC_2_125 b_2 NI_2 NS_125 0 -1.9425296765362901e-06
GC_2_126 b_2 NI_2 NS_126 0 -3.7933020889190574e-07
GC_2_127 b_2 NI_2 NS_127 0 -4.3560450224517711e-05
GC_2_128 b_2 NI_2 NS_128 0 -1.2838865325235263e-04
GC_2_129 b_2 NI_2 NS_129 0 -7.7535494917229482e-06
GC_2_130 b_2 NI_2 NS_130 0 -2.5629333688863314e-06
GC_2_131 b_2 NI_2 NS_131 0 -3.9876177363431412e-06
GC_2_132 b_2 NI_2 NS_132 0 -5.5167005632415455e-06
GC_2_133 b_2 NI_2 NS_133 0 -4.6974782808973103e-03
GC_2_134 b_2 NI_2 NS_134 0 -1.0219314154773429e-03
GC_2_135 b_2 NI_2 NS_135 0 1.4143515812236256e-02
GC_2_136 b_2 NI_2 NS_136 0 3.3541475722943365e-03
GC_2_137 b_2 NI_2 NS_137 0 -1.6532589860792958e-02
GC_2_138 b_2 NI_2 NS_138 0 -2.9391657335722608e-03
GC_2_139 b_2 NI_2 NS_139 0 5.2421008818699169e-03
GC_2_140 b_2 NI_2 NS_140 0 -8.9796558994643483e-04
GC_2_141 b_2 NI_2 NS_141 0 -8.8370735472231355e-04
GC_2_142 b_2 NI_2 NS_142 0 5.2597544400250537e-04
GC_2_143 b_2 NI_2 NS_143 0 1.0495816932228664e-03
GC_2_144 b_2 NI_2 NS_144 0 -3.0938269122115455e-03
GC_2_145 b_2 NI_2 NS_145 0 1.1507895503849462e-04
GC_2_146 b_2 NI_2 NS_146 0 -1.2392893254721286e-04
GC_2_147 b_2 NI_2 NS_147 0 2.3712826130611588e-05
GC_2_148 b_2 NI_2 NS_148 0 -3.5725294380228548e-05
GC_2_149 b_2 NI_2 NS_149 0 1.2015434770222746e-04
GC_2_150 b_2 NI_2 NS_150 0 -2.4359365421153066e-05
GC_2_151 b_2 NI_2 NS_151 0 1.4668317054393360e-05
GC_2_152 b_2 NI_2 NS_152 0 -6.0990489158751799e-06
GC_2_153 b_2 NI_2 NS_153 0 8.0170528191388210e-06
GC_2_154 b_2 NI_2 NS_154 0 -1.9004397230468540e-05
GC_2_155 b_2 NI_2 NS_155 0 -2.5995820307242423e-06
GC_2_156 b_2 NI_2 NS_156 0 -7.0854473254627540e-07
GC_2_157 b_2 NI_2 NS_157 0 4.5887345056387866e-03
GC_2_158 b_2 NI_2 NS_158 0 7.1101836417868450e-03
GC_2_159 b_2 NI_2 NS_159 0 -1.4957572226613871e-03
GC_2_160 b_2 NI_2 NS_160 0 -3.4097038649950617e-03
GC_2_161 b_2 NI_2 NS_161 0 -2.1124898861478916e-04
GC_2_162 b_2 NI_2 NS_162 0 -7.0861499213160500e-05
GC_2_163 b_2 NI_2 NS_163 0 -4.4002827903572034e-07
GC_2_164 b_2 NI_2 NS_164 0 4.6990824273163056e-07
GC_2_165 b_2 NI_2 NS_165 0 -6.5632200379994211e-05
GC_2_166 b_2 NI_2 NS_166 0 1.0730972501743362e-04
GC_2_167 b_2 NI_2 NS_167 0 -3.6452483014592744e-06
GC_2_168 b_2 NI_2 NS_168 0 -2.4918352824915344e-06
GC_2_169 b_2 NI_2 NS_169 0 -5.8478048547249071e-06
GC_2_170 b_2 NI_2 NS_170 0 -1.2234873010122079e-05
GC_2_171 b_2 NI_2 NS_171 0 -2.5290690076036214e-04
GC_2_172 b_2 NI_2 NS_172 0 7.1593872813075182e-05
GC_2_173 b_2 NI_2 NS_173 0 -1.2524514827127114e-04
GC_2_174 b_2 NI_2 NS_174 0 -5.0326143957820503e-05
GC_2_175 b_2 NI_2 NS_175 0 -3.0547799761846020e-05
GC_2_176 b_2 NI_2 NS_176 0 -7.1780745155126437e-06
GC_2_177 b_2 NI_2 NS_177 0 1.3168575740225659e-02
GC_2_178 b_2 NI_2 NS_178 0 -5.8033216824201865e-04
GC_2_179 b_2 NI_2 NS_179 0 -1.5406741695627441e-02
GC_2_180 b_2 NI_2 NS_180 0 6.1074988667727762e-03
GC_2_181 b_2 NI_2 NS_181 0 2.5861106581127201e-03
GC_2_182 b_2 NI_2 NS_182 0 -1.2319324840468366e-02
GC_2_183 b_2 NI_2 NS_183 0 8.7210186906419955e-03
GC_2_184 b_2 NI_2 NS_184 0 9.0037929058801359e-04
GC_2_185 b_2 NI_2 NS_185 0 -4.9795602169663616e-04
GC_2_186 b_2 NI_2 NS_186 0 -5.2255038624370888e-04
GC_2_187 b_2 NI_2 NS_187 0 -7.2163140669973362e-03
GC_2_188 b_2 NI_2 NS_188 0 -2.7242077050782972e-03
GC_2_189 b_2 NI_2 NS_189 0 -2.6607579565196294e-04
GC_2_190 b_2 NI_2 NS_190 0 9.1619082533729544e-05
GC_2_191 b_2 NI_2 NS_191 0 1.4115681002778853e-04
GC_2_192 b_2 NI_2 NS_192 0 2.8471219323678057e-05
GC_2_193 b_2 NI_2 NS_193 0 5.8069371680731367e-04
GC_2_194 b_2 NI_2 NS_194 0 7.7827289760597663e-05
GC_2_195 b_2 NI_2 NS_195 0 1.7744593264281886e-05
GC_2_196 b_2 NI_2 NS_196 0 1.3644662326488314e-06
GC_2_197 b_2 NI_2 NS_197 0 2.7646981342870554e-05
GC_2_198 b_2 NI_2 NS_198 0 -2.9931298068269267e-05
GC_2_199 b_2 NI_2 NS_199 0 6.2612320659154224e-06
GC_2_200 b_2 NI_2 NS_200 0 -2.9297897086100169e-06
GC_2_201 b_2 NI_2 NS_201 0 9.2196759660362001e-04
GC_2_202 b_2 NI_2 NS_202 0 4.6350572839868988e-03
GC_2_203 b_2 NI_2 NS_203 0 1.2090088203997489e-03
GC_2_204 b_2 NI_2 NS_204 0 -2.7465139938093828e-03
GC_2_205 b_2 NI_2 NS_205 0 -1.2960474857272088e-05
GC_2_206 b_2 NI_2 NS_206 0 -5.3539126923588092e-05
GC_2_207 b_2 NI_2 NS_207 0 -5.1457033823789171e-09
GC_2_208 b_2 NI_2 NS_208 0 1.6912619308248874e-07
GC_2_209 b_2 NI_2 NS_209 0 -1.2102239999019448e-05
GC_2_210 b_2 NI_2 NS_210 0 5.5876271647372248e-06
GC_2_211 b_2 NI_2 NS_211 0 2.5318691454506547e-07
GC_2_212 b_2 NI_2 NS_212 0 -1.4145354745747211e-07
GC_2_213 b_2 NI_2 NS_213 0 2.9982820118965037e-06
GC_2_214 b_2 NI_2 NS_214 0 -1.3346114598449846e-07
GC_2_215 b_2 NI_2 NS_215 0 -4.1929143608957548e-05
GC_2_216 b_2 NI_2 NS_216 0 -4.6870406181454651e-05
GC_2_217 b_2 NI_2 NS_217 0 2.8638373402433284e-06
GC_2_218 b_2 NI_2 NS_218 0 -1.0549144923927072e-06
GC_2_219 b_2 NI_2 NS_219 0 1.7502705895595046e-06
GC_2_220 b_2 NI_2 NS_220 0 -4.5742259217860725e-06
GC_2_221 b_2 NI_2 NS_221 0 -1.8304325853747354e-02
GC_2_222 b_2 NI_2 NS_222 0 9.4343763878141013e-05
GC_2_223 b_2 NI_2 NS_223 0 1.0992279551523229e-02
GC_2_224 b_2 NI_2 NS_224 0 -8.8287399600673055e-03
GC_2_225 b_2 NI_2 NS_225 0 -1.4721970915936617e-03
GC_2_226 b_2 NI_2 NS_226 0 7.3804244445366991e-03
GC_2_227 b_2 NI_2 NS_227 0 6.5444475108929496e-03
GC_2_228 b_2 NI_2 NS_228 0 7.2497330726828852e-05
GC_2_229 b_2 NI_2 NS_229 0 -2.1772676130097425e-03
GC_2_230 b_2 NI_2 NS_230 0 -2.0344017971627385e-03
GC_2_231 b_2 NI_2 NS_231 0 -1.0511637422555295e-03
GC_2_232 b_2 NI_2 NS_232 0 4.1364617698708165e-03
GC_2_233 b_2 NI_2 NS_233 0 1.0826425534843308e-04
GC_2_234 b_2 NI_2 NS_234 0 -1.3510495797179348e-04
GC_2_235 b_2 NI_2 NS_235 0 -7.3274034286549747e-06
GC_2_236 b_2 NI_2 NS_236 0 -3.6813368376294036e-05
GC_2_237 b_2 NI_2 NS_237 0 5.9208532565269804e-05
GC_2_238 b_2 NI_2 NS_238 0 -2.3283379809020444e-04
GC_2_239 b_2 NI_2 NS_239 0 -3.4391599992912310e-06
GC_2_240 b_2 NI_2 NS_240 0 -1.1077300717411402e-05
GC_2_241 b_2 NI_2 NS_241 0 -3.5853797609917624e-05
GC_2_242 b_2 NI_2 NS_242 0 -1.2023799108250486e-05
GC_2_243 b_2 NI_2 NS_243 0 -6.5784171957099172e-06
GC_2_244 b_2 NI_2 NS_244 0 -1.1001697587888857e-06
GC_2_245 b_2 NI_2 NS_245 0 5.1981096425164760e-03
GC_2_246 b_2 NI_2 NS_246 0 7.5917200122475881e-03
GC_2_247 b_2 NI_2 NS_247 0 -2.5683500636750132e-03
GC_2_248 b_2 NI_2 NS_248 0 -3.5182470795134860e-03
GC_2_249 b_2 NI_2 NS_249 0 -3.5119961975428528e-04
GC_2_250 b_2 NI_2 NS_250 0 -5.9277701985067441e-05
GC_2_251 b_2 NI_2 NS_251 0 -1.0106058347138826e-08
GC_2_252 b_2 NI_2 NS_252 0 8.7607962482813507e-07
GC_2_253 b_2 NI_2 NS_253 0 -7.8295119980817512e-05
GC_2_254 b_2 NI_2 NS_254 0 1.6659559371618525e-04
GC_2_255 b_2 NI_2 NS_255 0 -4.0090664178990847e-06
GC_2_256 b_2 NI_2 NS_256 0 -3.1648973391936759e-06
GC_2_257 b_2 NI_2 NS_257 0 -7.6632663683464246e-06
GC_2_258 b_2 NI_2 NS_258 0 -2.0112510740782180e-05
GC_2_259 b_2 NI_2 NS_259 0 -3.6834113681123585e-04
GC_2_260 b_2 NI_2 NS_260 0 1.5609629405498014e-04
GC_2_261 b_2 NI_2 NS_261 0 -1.9882963591357432e-04
GC_2_262 b_2 NI_2 NS_262 0 -5.9439222031202788e-05
GC_2_263 b_2 NI_2 NS_263 0 -4.1363970428796061e-05
GC_2_264 b_2 NI_2 NS_264 0 -5.6111904906548138e-06
GC_2_265 b_2 NI_2 NS_265 0 2.2948301871707516e-02
GC_2_266 b_2 NI_2 NS_266 0 -5.3842917103643685e-04
GC_2_267 b_2 NI_2 NS_267 0 -6.7369915218252032e-03
GC_2_268 b_2 NI_2 NS_268 0 8.1863869839353936e-03
GC_2_269 b_2 NI_2 NS_269 0 -3.3877637453874742e-03
GC_2_270 b_2 NI_2 NS_270 0 -9.1189585495052312e-03
GC_2_271 b_2 NI_2 NS_271 0 6.4574413697182148e-03
GC_2_272 b_2 NI_2 NS_272 0 4.8890777964432806e-04
GC_2_273 b_2 NI_2 NS_273 0 -2.0439170955097140e-03
GC_2_274 b_2 NI_2 NS_274 0 9.0199755405290195e-04
GC_2_275 b_2 NI_2 NS_275 0 -8.2736238464650273e-03
GC_2_276 b_2 NI_2 NS_276 0 2.9338873651062179e-03
GC_2_277 b_2 NI_2 NS_277 0 -1.5612575571941683e-04
GC_2_278 b_2 NI_2 NS_278 0 1.1334855413045649e-04
GC_2_279 b_2 NI_2 NS_279 0 1.0636730255073439e-04
GC_2_280 b_2 NI_2 NS_280 0 6.6658769272031490e-05
GC_2_281 b_2 NI_2 NS_281 0 -6.2653489996279321e-06
GC_2_282 b_2 NI_2 NS_282 0 3.6242976870219356e-05
GC_2_283 b_2 NI_2 NS_283 0 -1.0501946086942847e-05
GC_2_284 b_2 NI_2 NS_284 0 2.5674300525147206e-05
GC_2_285 b_2 NI_2 NS_285 0 -3.6817673476874404e-06
GC_2_286 b_2 NI_2 NS_286 0 4.3958088448512716e-05
GC_2_287 b_2 NI_2 NS_287 0 3.8785826680613792e-06
GC_2_288 b_2 NI_2 NS_288 0 2.6611844246806781e-06
GC_2_289 b_2 NI_2 NS_289 0 1.1590208880735804e-03
GC_2_290 b_2 NI_2 NS_290 0 -3.2210073781198745e-03
GC_2_291 b_2 NI_2 NS_291 0 2.6143654296434133e-04
GC_2_292 b_2 NI_2 NS_292 0 1.2121985100609154e-03
GC_2_293 b_2 NI_2 NS_293 0 2.3177105225077397e-04
GC_2_294 b_2 NI_2 NS_294 0 -3.1244705689401694e-04
GC_2_295 b_2 NI_2 NS_295 0 1.5929202578394166e-06
GC_2_296 b_2 NI_2 NS_296 0 -1.1741403603297224e-06
GC_2_297 b_2 NI_2 NS_297 0 -3.7724423032074655e-05
GC_2_298 b_2 NI_2 NS_298 0 -7.5794675054950889e-05
GC_2_299 b_2 NI_2 NS_299 0 -9.7753472714100053e-07
GC_2_300 b_2 NI_2 NS_300 0 -2.3368512417510151e-06
GC_2_301 b_2 NI_2 NS_301 0 3.3777470672541973e-08
GC_2_302 b_2 NI_2 NS_302 0 -4.4193393432666547e-06
GC_2_303 b_2 NI_2 NS_303 0 1.4335024226076927e-04
GC_2_304 b_2 NI_2 NS_304 0 1.0012941665591916e-04
GC_2_305 b_2 NI_2 NS_305 0 3.2113032995881542e-05
GC_2_306 b_2 NI_2 NS_306 0 3.9293842067847096e-05
GC_2_307 b_2 NI_2 NS_307 0 1.0596578986689366e-05
GC_2_308 b_2 NI_2 NS_308 0 -2.3269419541312232e-06
GC_2_309 b_2 NI_2 NS_309 0 -1.3893730258818850e-02
GC_2_310 b_2 NI_2 NS_310 0 2.9026102260314038e-04
GC_2_311 b_2 NI_2 NS_311 0 4.8228597249886807e-03
GC_2_312 b_2 NI_2 NS_312 0 -9.7669134193473436e-03
GC_2_313 b_2 NI_2 NS_313 0 5.6062432698941091e-03
GC_2_314 b_2 NI_2 NS_314 0 6.9731523325504098e-03
GC_2_315 b_2 NI_2 NS_315 0 5.5234001046188669e-03
GC_2_316 b_2 NI_2 NS_316 0 7.3380258070920650e-04
GC_2_317 b_2 NI_2 NS_317 0 -1.9106744232108884e-03
GC_2_318 b_2 NI_2 NS_318 0 -1.1727547925272431e-03
GC_2_319 b_2 NI_2 NS_319 0 -8.2268498478394023e-04
GC_2_320 b_2 NI_2 NS_320 0 7.3480383871385533e-03
GC_2_321 b_2 NI_2 NS_321 0 6.9575961953820809e-05
GC_2_322 b_2 NI_2 NS_322 0 -9.5434784510327653e-05
GC_2_323 b_2 NI_2 NS_323 0 1.4706061031995664e-06
GC_2_324 b_2 NI_2 NS_324 0 -1.4718974485804501e-05
GC_2_325 b_2 NI_2 NS_325 0 -8.5476036403173112e-05
GC_2_326 b_2 NI_2 NS_326 0 -8.9163477564147448e-05
GC_2_327 b_2 NI_2 NS_327 0 1.1463293346872502e-06
GC_2_328 b_2 NI_2 NS_328 0 4.7508347406137928e-06
GC_2_329 b_2 NI_2 NS_329 0 3.0264435367647635e-06
GC_2_330 b_2 NI_2 NS_330 0 1.6333030724758821e-05
GC_2_331 b_2 NI_2 NS_331 0 -1.2945820052244734e-06
GC_2_332 b_2 NI_2 NS_332 0 3.6536968317555532e-07
GC_2_333 b_2 NI_2 NS_333 0 -1.3192198976325331e-03
GC_2_334 b_2 NI_2 NS_334 0 3.4185839203154391e-03
GC_2_335 b_2 NI_2 NS_335 0 3.4934756350963475e-04
GC_2_336 b_2 NI_2 NS_336 0 -1.0911559514151384e-03
GC_2_337 b_2 NI_2 NS_337 0 -1.5710296991539583e-04
GC_2_338 b_2 NI_2 NS_338 0 -1.2483946531991605e-04
GC_2_339 b_2 NI_2 NS_339 0 -2.9558702803376076e-07
GC_2_340 b_2 NI_2 NS_340 0 2.2030008634529505e-08
GC_2_341 b_2 NI_2 NS_341 0 -6.0982957870091750e-05
GC_2_342 b_2 NI_2 NS_342 0 6.4431260603476062e-05
GC_2_343 b_2 NI_2 NS_343 0 -3.0538690357748591e-06
GC_2_344 b_2 NI_2 NS_344 0 -1.2068345885272191e-06
GC_2_345 b_2 NI_2 NS_345 0 -5.2754100552014584e-06
GC_2_346 b_2 NI_2 NS_346 0 -1.2386946183512108e-05
GC_2_347 b_2 NI_2 NS_347 0 -1.2300988782440090e-04
GC_2_348 b_2 NI_2 NS_348 0 2.6460789109102542e-05
GC_2_349 b_2 NI_2 NS_349 0 -8.5507141967118704e-05
GC_2_350 b_2 NI_2 NS_350 0 -4.5749619149008469e-05
GC_2_351 b_2 NI_2 NS_351 0 -1.5451556390134935e-05
GC_2_352 b_2 NI_2 NS_352 0 -3.2006998600218636e-06
GC_2_353 b_2 NI_2 NS_353 0 -3.0548453918575785e-03
GC_2_354 b_2 NI_2 NS_354 0 4.2903336641686789e-05
GC_2_355 b_2 NI_2 NS_355 0 -9.6647408528049485e-06
GC_2_356 b_2 NI_2 NS_356 0 3.6005487693615895e-04
GC_2_357 b_2 NI_2 NS_357 0 -9.9797222235524659e-04
GC_2_358 b_2 NI_2 NS_358 0 -4.1025550018221378e-04
GC_2_359 b_2 NI_2 NS_359 0 -2.4854498401011581e-04
GC_2_360 b_2 NI_2 NS_360 0 -1.4564868200065591e-03
GC_2_361 b_2 NI_2 NS_361 0 3.1072139561217054e-04
GC_2_362 b_2 NI_2 NS_362 0 -4.1918890119439169e-05
GC_2_363 b_2 NI_2 NS_363 0 1.4124705031723114e-03
GC_2_364 b_2 NI_2 NS_364 0 -1.1653485419026869e-03
GC_2_365 b_2 NI_2 NS_365 0 -1.0494437660220253e-05
GC_2_366 b_2 NI_2 NS_366 0 1.8459527648338465e-04
GC_2_367 b_2 NI_2 NS_367 0 2.1211595109365235e-04
GC_2_368 b_2 NI_2 NS_368 0 -8.7597575019128350e-05
GC_2_369 b_2 NI_2 NS_369 0 -1.8971725494097431e-04
GC_2_370 b_2 NI_2 NS_370 0 1.2548583488421593e-04
GC_2_371 b_2 NI_2 NS_371 0 -1.8410270438319140e-05
GC_2_372 b_2 NI_2 NS_372 0 -1.5639364519903198e-05
GC_2_373 b_2 NI_2 NS_373 0 -4.4386195558264603e-06
GC_2_374 b_2 NI_2 NS_374 0 -5.0753899602943496e-05
GC_2_375 b_2 NI_2 NS_375 0 4.7062720113860348e-06
GC_2_376 b_2 NI_2 NS_376 0 2.4035829340799445e-06
GC_2_377 b_2 NI_2 NS_377 0 2.3765047109728030e-03
GC_2_378 b_2 NI_2 NS_378 0 3.0204123580647958e-03
GC_2_379 b_2 NI_2 NS_379 0 -1.4545168383704270e-03
GC_2_380 b_2 NI_2 NS_380 0 -2.2237740734171092e-03
GC_2_381 b_2 NI_2 NS_381 0 -1.4344081759101821e-04
GC_2_382 b_2 NI_2 NS_382 0 4.4317697326695393e-05
GC_2_383 b_2 NI_2 NS_383 0 -7.7608163436797340e-07
GC_2_384 b_2 NI_2 NS_384 0 4.6675061898144092e-07
GC_2_385 b_2 NI_2 NS_385 0 8.0425714901415033e-08
GC_2_386 b_2 NI_2 NS_386 0 2.8073070446840358e-05
GC_2_387 b_2 NI_2 NS_387 0 -9.9666977822677929e-07
GC_2_388 b_2 NI_2 NS_388 0 1.1224869086852922e-06
GC_2_389 b_2 NI_2 NS_389 0 1.7158802719719035e-06
GC_2_390 b_2 NI_2 NS_390 0 6.0925076513503129e-07
GC_2_391 b_2 NI_2 NS_391 0 -1.0052660390036319e-04
GC_2_392 b_2 NI_2 NS_392 0 -8.9327236264735851e-05
GC_2_393 b_2 NI_2 NS_393 0 -4.9561199467249501e-06
GC_2_394 b_2 NI_2 NS_394 0 -5.4431559589148851e-05
GC_2_395 b_2 NI_2 NS_395 0 -6.9059987283785738e-06
GC_2_396 b_2 NI_2 NS_396 0 1.4081668083384394e-06
GC_2_397 b_2 NI_2 NS_397 0 -7.4712241648775355e-03
GC_2_398 b_2 NI_2 NS_398 0 -3.7561783335167365e-06
GC_2_399 b_2 NI_2 NS_399 0 -7.0776931132161716e-04
GC_2_400 b_2 NI_2 NS_400 0 -3.6537222418061524e-04
GC_2_401 b_2 NI_2 NS_401 0 1.3974827401094892e-04
GC_2_402 b_2 NI_2 NS_402 0 -9.7990084198358910e-04
GC_2_403 b_2 NI_2 NS_403 0 -5.5936302972017762e-05
GC_2_404 b_2 NI_2 NS_404 0 -1.2390964501964160e-03
GC_2_405 b_2 NI_2 NS_405 0 9.5009474298937398e-04
GC_2_406 b_2 NI_2 NS_406 0 7.0719923835694599e-04
GC_2_407 b_2 NI_2 NS_407 0 1.1643597078637722e-03
GC_2_408 b_2 NI_2 NS_408 0 -8.1019452495939570e-04
GC_2_409 b_2 NI_2 NS_409 0 -6.5949394401336895e-05
GC_2_410 b_2 NI_2 NS_410 0 -7.0904955867120438e-05
GC_2_411 b_2 NI_2 NS_411 0 2.7971431652467720e-05
GC_2_412 b_2 NI_2 NS_412 0 -2.9507957953521657e-05
GC_2_413 b_2 NI_2 NS_413 0 -1.4569953788208924e-04
GC_2_414 b_2 NI_2 NS_414 0 1.9184084497495891e-04
GC_2_415 b_2 NI_2 NS_415 0 -9.9678491836806400e-06
GC_2_416 b_2 NI_2 NS_416 0 1.8883028600059826e-05
GC_2_417 b_2 NI_2 NS_417 0 -4.7106866882105551e-06
GC_2_418 b_2 NI_2 NS_418 0 6.4296425312806792e-05
GC_2_419 b_2 NI_2 NS_419 0 -7.9851578341811593e-07
GC_2_420 b_2 NI_2 NS_420 0 -2.0953949566777071e-07
GC_2_421 b_2 NI_2 NS_421 0 3.4019245258355979e-03
GC_2_422 b_2 NI_2 NS_422 0 -4.2108099289034501e-03
GC_2_423 b_2 NI_2 NS_423 0 -1.9831653689060518e-03
GC_2_424 b_2 NI_2 NS_424 0 2.3988985359626289e-03
GC_2_425 b_2 NI_2 NS_425 0 1.3333553247125515e-04
GC_2_426 b_2 NI_2 NS_426 0 7.1231993320901345e-05
GC_2_427 b_2 NI_2 NS_427 0 2.1726896164727731e-06
GC_2_428 b_2 NI_2 NS_428 0 4.9065804508798785e-07
GC_2_429 b_2 NI_2 NS_429 0 1.8764448668074476e-05
GC_2_430 b_2 NI_2 NS_430 0 -6.6746659652566919e-05
GC_2_431 b_2 NI_2 NS_431 0 3.8683657990560323e-06
GC_2_432 b_2 NI_2 NS_432 0 7.2832691611752922e-06
GC_2_433 b_2 NI_2 NS_433 0 -9.5787296962117968e-06
GC_2_434 b_2 NI_2 NS_434 0 -2.2926818877180860e-05
GC_2_435 b_2 NI_2 NS_435 0 -1.7534704644637993e-05
GC_2_436 b_2 NI_2 NS_436 0 2.5946716169120539e-04
GC_2_437 b_2 NI_2 NS_437 0 -1.8547747699624301e-04
GC_2_438 b_2 NI_2 NS_438 0 1.3937575907648981e-06
GC_2_439 b_2 NI_2 NS_439 0 4.3717681186858685e-05
GC_2_440 b_2 NI_2 NS_440 0 6.0599615467949236e-05
GC_2_441 b_2 NI_2 NS_441 0 4.7363613247105628e-03
GC_2_442 b_2 NI_2 NS_442 0 -4.3241768768392019e-05
GC_2_443 b_2 NI_2 NS_443 0 -7.5964936884036652e-05
GC_2_444 b_2 NI_2 NS_444 0 1.5091969840030509e-03
GC_2_445 b_2 NI_2 NS_445 0 -1.7719636936816159e-03
GC_2_446 b_2 NI_2 NS_446 0 -7.6151044981323849e-04
GC_2_447 b_2 NI_2 NS_447 0 8.3298023251964859e-04
GC_2_448 b_2 NI_2 NS_448 0 -9.9704595298670692e-04
GC_2_449 b_2 NI_2 NS_449 0 1.1335302015566583e-04
GC_2_450 b_2 NI_2 NS_450 0 1.4084194661344551e-04
GC_2_451 b_2 NI_2 NS_451 0 -3.9469324108687037e-05
GC_2_452 b_2 NI_2 NS_452 0 1.2378843102866502e-03
GC_2_453 b_2 NI_2 NS_453 0 2.5020193866724014e-07
GC_2_454 b_2 NI_2 NS_454 0 1.3294696394776883e-04
GC_2_455 b_2 NI_2 NS_455 0 1.8171066811793396e-04
GC_2_456 b_2 NI_2 NS_456 0 -3.1244219555554999e-05
GC_2_457 b_2 NI_2 NS_457 0 -1.9332152614710330e-04
GC_2_458 b_2 NI_2 NS_458 0 2.7287839375829089e-04
GC_2_459 b_2 NI_2 NS_459 0 -6.9931841373738263e-07
GC_2_460 b_2 NI_2 NS_460 0 7.5432030939670111e-06
GC_2_461 b_2 NI_2 NS_461 0 3.5995035306485461e-05
GC_2_462 b_2 NI_2 NS_462 0 -6.6370412536265992e-06
GC_2_463 b_2 NI_2 NS_463 0 5.4957730258634839e-06
GC_2_464 b_2 NI_2 NS_464 0 1.6960362651062392e-06
GC_2_465 b_2 NI_2 NS_465 0 -1.8441734751115501e-03
GC_2_466 b_2 NI_2 NS_466 0 7.2547656387353236e-04
GC_2_467 b_2 NI_2 NS_467 0 8.8415464303359063e-04
GC_2_468 b_2 NI_2 NS_468 0 -7.2362249586577416e-04
GC_2_469 b_2 NI_2 NS_469 0 -1.7370537981510593e-04
GC_2_470 b_2 NI_2 NS_470 0 -2.5174035245557495e-04
GC_2_471 b_2 NI_2 NS_471 0 -1.1650132152928826e-06
GC_2_472 b_2 NI_2 NS_472 0 -1.1275636457535527e-06
GC_2_473 b_2 NI_2 NS_473 0 -5.4668740162236290e-05
GC_2_474 b_2 NI_2 NS_474 0 1.6240973990150194e-05
GC_2_475 b_2 NI_2 NS_475 0 -1.0587979381144961e-06
GC_2_476 b_2 NI_2 NS_476 0 -3.2037016818829446e-08
GC_2_477 b_2 NI_2 NS_477 0 -2.8400643513660865e-06
GC_2_478 b_2 NI_2 NS_478 0 -1.8549790021026209e-06
GC_2_479 b_2 NI_2 NS_479 0 5.7932958849694231e-05
GC_2_480 b_2 NI_2 NS_480 0 -1.1120971013706280e-04
GC_2_481 b_2 NI_2 NS_481 0 2.0166841556902499e-05
GC_2_482 b_2 NI_2 NS_482 0 -3.6151431612873995e-05
GC_2_483 b_2 NI_2 NS_483 0 5.9349068284453076e-06
GC_2_484 b_2 NI_2 NS_484 0 -6.0312211614388469e-06
GC_2_485 b_2 NI_2 NS_485 0 -7.0009713482852877e-03
GC_2_486 b_2 NI_2 NS_486 0 4.8134337560931908e-05
GC_2_487 b_2 NI_2 NS_487 0 -5.2245231104693730e-04
GC_2_488 b_2 NI_2 NS_488 0 -1.7389684517120324e-03
GC_2_489 b_2 NI_2 NS_489 0 1.7859563375143724e-03
GC_2_490 b_2 NI_2 NS_490 0 -4.9223521168674956e-04
GC_2_491 b_2 NI_2 NS_491 0 1.2938659980273675e-03
GC_2_492 b_2 NI_2 NS_492 0 -9.0056138653311804e-04
GC_2_493 b_2 NI_2 NS_493 0 -2.5114284586269482e-04
GC_2_494 b_2 NI_2 NS_494 0 2.5924648839054185e-04
GC_2_495 b_2 NI_2 NS_495 0 1.7657872136180250e-03
GC_2_496 b_2 NI_2 NS_496 0 1.3062342906769797e-03
GC_2_497 b_2 NI_2 NS_497 0 -2.4702266291884128e-05
GC_2_498 b_2 NI_2 NS_498 0 -6.4663827869055834e-05
GC_2_499 b_2 NI_2 NS_499 0 2.6834901486777538e-05
GC_2_500 b_2 NI_2 NS_500 0 -2.3854992740695017e-05
GC_2_501 b_2 NI_2 NS_501 0 -8.3833893349802359e-05
GC_2_502 b_2 NI_2 NS_502 0 1.5331454557928611e-04
GC_2_503 b_2 NI_2 NS_503 0 -1.8534900347083444e-06
GC_2_504 b_2 NI_2 NS_504 0 1.0180698426887929e-05
GC_2_505 b_2 NI_2 NS_505 0 4.3862392018009432e-06
GC_2_506 b_2 NI_2 NS_506 0 3.0936550171997705e-05
GC_2_507 b_2 NI_2 NS_507 0 -6.2342257391899419e-07
GC_2_508 b_2 NI_2 NS_508 0 2.2712755022244840e-07
GC_2_509 b_2 NI_2 NS_509 0 8.0486074696440300e-04
GC_2_510 b_2 NI_2 NS_510 0 -8.8262624674594363e-05
GC_2_511 b_2 NI_2 NS_511 0 -4.4552090311688523e-04
GC_2_512 b_2 NI_2 NS_512 0 4.3729240437113552e-04
GC_2_513 b_2 NI_2 NS_513 0 1.1171733688156650e-05
GC_2_514 b_2 NI_2 NS_514 0 -2.5726433397813925e-05
GC_2_515 b_2 NI_2 NS_515 0 7.6346496527715050e-07
GC_2_516 b_2 NI_2 NS_516 0 -2.9276901755752163e-08
GC_2_517 b_2 NI_2 NS_517 0 -8.9731485202120356e-06
GC_2_518 b_2 NI_2 NS_518 0 -1.5131074961270372e-05
GC_2_519 b_2 NI_2 NS_519 0 5.3457667862960110e-07
GC_2_520 b_2 NI_2 NS_520 0 3.1692041975415030e-06
GC_2_521 b_2 NI_2 NS_521 0 -5.5403055254994188e-06
GC_2_522 b_2 NI_2 NS_522 0 -1.3507680947926551e-05
GC_2_523 b_2 NI_2 NS_523 0 -2.4375028596931138e-05
GC_2_524 b_2 NI_2 NS_524 0 8.9816869254378881e-05
GC_2_525 b_2 NI_2 NS_525 0 -9.2256127156705364e-05
GC_2_526 b_2 NI_2 NS_526 0 -1.3513340797080998e-05
GC_2_527 b_2 NI_2 NS_527 0 1.6340525871743286e-05
GC_2_528 b_2 NI_2 NS_528 0 2.5546316554706231e-05
GD_2_1 b_2 NI_2 NA_1 0 -7.2737643139165475e-03
GD_2_2 b_2 NI_2 NA_2 0 1.2974654951848591e-01
GD_2_3 b_2 NI_2 NA_3 0 -2.4079607662927200e-03
GD_2_4 b_2 NI_2 NA_4 0 -1.5147017228272035e-03
GD_2_5 b_2 NI_2 NA_5 0 -3.6721389996685603e-03
GD_2_6 b_2 NI_2 NA_6 0 1.3532982709456524e-03
GD_2_7 b_2 NI_2 NA_7 0 -1.1073250957355342e-02
GD_2_8 b_2 NI_2 NA_8 0 1.4622702056562311e-03
GD_2_9 b_2 NI_2 NA_9 0 1.9149126078376935e-03
GD_2_10 b_2 NI_2 NA_10 0 5.2730083733379621e-03
GD_2_11 b_2 NI_2 NA_11 0 -3.1761320459139184e-03
GD_2_12 b_2 NI_2 NA_12 0 2.9574426790477948e-03
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 8.1298888220935183e-03
GC_3_2 b_3 NI_3 NS_2 0 -4.6313664333959834e-04
GC_3_3 b_3 NI_3 NS_3 0 1.1775616910083705e-02
GC_3_4 b_3 NI_3 NS_4 0 3.4756009174450688e-03
GC_3_5 b_3 NI_3 NS_5 0 -9.1264956974341695e-03
GC_3_6 b_3 NI_3 NS_6 0 -8.4944380370523057e-03
GC_3_7 b_3 NI_3 NS_7 0 1.1666689942321109e-02
GC_3_8 b_3 NI_3 NS_8 0 7.1468101097944877e-03
GC_3_9 b_3 NI_3 NS_9 0 -2.9079236264750556e-03
GC_3_10 b_3 NI_3 NS_10 0 -1.1074628460339111e-03
GC_3_11 b_3 NI_3 NS_11 0 2.7737482651146420e-03
GC_3_12 b_3 NI_3 NS_12 0 2.8643816821407055e-03
GC_3_13 b_3 NI_3 NS_13 0 5.1414858487716501e-04
GC_3_14 b_3 NI_3 NS_14 0 4.4167817349768202e-04
GC_3_15 b_3 NI_3 NS_15 0 5.6985398085405308e-05
GC_3_16 b_3 NI_3 NS_16 0 1.9751981092291029e-04
GC_3_17 b_3 NI_3 NS_17 0 1.3150881529620248e-03
GC_3_18 b_3 NI_3 NS_18 0 3.6828708635688342e-04
GC_3_19 b_3 NI_3 NS_19 0 1.5243466980850202e-04
GC_3_20 b_3 NI_3 NS_20 0 1.4876395456431049e-04
GC_3_21 b_3 NI_3 NS_21 0 2.6549024590820749e-04
GC_3_22 b_3 NI_3 NS_22 0 4.3527186433795402e-05
GC_3_23 b_3 NI_3 NS_23 0 -1.0262837575082627e-05
GC_3_24 b_3 NI_3 NS_24 0 3.3651479283350079e-06
GC_3_25 b_3 NI_3 NS_25 0 -1.9801857301253077e-02
GC_3_26 b_3 NI_3 NS_26 0 7.5551435785730838e-03
GC_3_27 b_3 NI_3 NS_27 0 1.4228094632459330e-02
GC_3_28 b_3 NI_3 NS_28 0 1.1891842589333466e-03
GC_3_29 b_3 NI_3 NS_29 0 -4.2618652470525088e-04
GC_3_30 b_3 NI_3 NS_30 0 7.0823364159519282e-06
GC_3_31 b_3 NI_3 NS_31 0 1.6111007194781610e-06
GC_3_32 b_3 NI_3 NS_32 0 3.5599396390083555e-06
GC_3_33 b_3 NI_3 NS_33 0 2.1165662609025086e-04
GC_3_34 b_3 NI_3 NS_34 0 -1.8258783416623498e-05
GC_3_35 b_3 NI_3 NS_35 0 5.1141436212598160e-06
GC_3_36 b_3 NI_3 NS_36 0 9.6168016077468899e-07
GC_3_37 b_3 NI_3 NS_37 0 3.1338806345524002e-07
GC_3_38 b_3 NI_3 NS_38 0 7.9388977764251759e-07
GC_3_39 b_3 NI_3 NS_39 0 -2.8029008656081775e-04
GC_3_40 b_3 NI_3 NS_40 0 2.8861647396649003e-04
GC_3_41 b_3 NI_3 NS_41 0 -3.5661394941243219e-05
GC_3_42 b_3 NI_3 NS_42 0 -5.7109012747172965e-05
GC_3_43 b_3 NI_3 NS_43 0 -1.7863884658288473e-05
GC_3_44 b_3 NI_3 NS_44 0 1.0868955973740452e-05
GC_3_45 b_3 NI_3 NS_45 0 4.1353853743977802e-03
GC_3_46 b_3 NI_3 NS_46 0 -3.8950436030153691e-04
GC_3_47 b_3 NI_3 NS_47 0 -2.0786969519512939e-02
GC_3_48 b_3 NI_3 NS_48 0 -3.3764631098210773e-03
GC_3_49 b_3 NI_3 NS_49 0 1.0882611112276237e-02
GC_3_50 b_3 NI_3 NS_50 0 -3.7983016640827220e-03
GC_3_51 b_3 NI_3 NS_51 0 6.3210213390045428e-03
GC_3_52 b_3 NI_3 NS_52 0 1.0575600338915193e-03
GC_3_53 b_3 NI_3 NS_53 0 1.7290934516665741e-03
GC_3_54 b_3 NI_3 NS_54 0 1.1711422664489524e-04
GC_3_55 b_3 NI_3 NS_55 0 -8.1541195205052559e-04
GC_3_56 b_3 NI_3 NS_56 0 -8.9796307251480117e-03
GC_3_57 b_3 NI_3 NS_57 0 -2.5676279977738527e-04
GC_3_58 b_3 NI_3 NS_58 0 5.5670860307670095e-05
GC_3_59 b_3 NI_3 NS_59 0 1.8232763210353732e-04
GC_3_60 b_3 NI_3 NS_60 0 4.8224998791142862e-05
GC_3_61 b_3 NI_3 NS_61 0 5.2801459320032593e-04
GC_3_62 b_3 NI_3 NS_62 0 4.1049378120103485e-04
GC_3_63 b_3 NI_3 NS_63 0 3.6402264054753365e-05
GC_3_64 b_3 NI_3 NS_64 0 2.2720379219436885e-05
GC_3_65 b_3 NI_3 NS_65 0 7.2644729265617774e-05
GC_3_66 b_3 NI_3 NS_66 0 -2.6561525810010667e-06
GC_3_67 b_3 NI_3 NS_67 0 7.1455434930235845e-06
GC_3_68 b_3 NI_3 NS_68 0 -2.6258464294509045e-06
GC_3_69 b_3 NI_3 NS_69 0 -4.2482848656218214e-03
GC_3_70 b_3 NI_3 NS_70 0 8.4802273171720351e-03
GC_3_71 b_3 NI_3 NS_71 0 3.6436292071331680e-03
GC_3_72 b_3 NI_3 NS_72 0 -3.6565506073507428e-03
GC_3_73 b_3 NI_3 NS_73 0 -1.7806454419369135e-04
GC_3_74 b_3 NI_3 NS_74 0 1.9560305429019401e-04
GC_3_75 b_3 NI_3 NS_75 0 -5.5118032006927998e-07
GC_3_76 b_3 NI_3 NS_76 0 8.4487321429201342e-07
GC_3_77 b_3 NI_3 NS_77 0 2.3642872544252987e-05
GC_3_78 b_3 NI_3 NS_78 0 5.7969512907821372e-05
GC_3_79 b_3 NI_3 NS_79 0 -3.6087148457585462e-07
GC_3_80 b_3 NI_3 NS_80 0 8.1753374210547732e-07
GC_3_81 b_3 NI_3 NS_81 0 -1.9425296765333810e-06
GC_3_82 b_3 NI_3 NS_82 0 -3.7933020889209860e-07
GC_3_83 b_3 NI_3 NS_83 0 -4.3560450224626701e-05
GC_3_84 b_3 NI_3 NS_84 0 -1.2838865325217510e-04
GC_3_85 b_3 NI_3 NS_85 0 -7.7535494917729892e-06
GC_3_86 b_3 NI_3 NS_86 0 -2.5629333688322852e-06
GC_3_87 b_3 NI_3 NS_87 0 -3.9876177363401885e-06
GC_3_88 b_3 NI_3 NS_88 0 -5.5167005632254959e-06
GC_3_89 b_3 NI_3 NS_89 0 -1.3825734607730351e-02
GC_3_90 b_3 NI_3 NS_90 0 1.3949736747738624e-02
GC_3_91 b_3 NI_3 NS_91 0 1.3443994015635528e-02
GC_3_92 b_3 NI_3 NS_92 0 2.8884592788084871e-03
GC_3_93 b_3 NI_3 NS_93 0 1.8659211346886171e-02
GC_3_94 b_3 NI_3 NS_94 0 -7.8978521960721933e-04
GC_3_95 b_3 NI_3 NS_95 0 1.4666656852023240e-02
GC_3_96 b_3 NI_3 NS_96 0 1.2858489302541694e-02
GC_3_97 b_3 NI_3 NS_97 0 2.5815277743514277e-03
GC_3_98 b_3 NI_3 NS_98 0 3.0567215644103350e-03
GC_3_99 b_3 NI_3 NS_99 0 -2.1482889850685289e-03
GC_3_100 b_3 NI_3 NS_100 0 1.8557707088420441e-02
GC_3_101 b_3 NI_3 NS_101 0 6.0685528564230582e-04
GC_3_102 b_3 NI_3 NS_102 0 4.5197175718815762e-04
GC_3_103 b_3 NI_3 NS_103 0 -3.4134346922265990e-06
GC_3_104 b_3 NI_3 NS_104 0 2.3373764299310600e-04
GC_3_105 b_3 NI_3 NS_105 0 2.0955849288964495e-03
GC_3_106 b_3 NI_3 NS_106 0 -5.6072423795650559e-04
GC_3_107 b_3 NI_3 NS_107 0 1.8453483330579072e-04
GC_3_108 b_3 NI_3 NS_108 0 1.3828215306845143e-04
GC_3_109 b_3 NI_3 NS_109 0 2.2198664866622373e-04
GC_3_110 b_3 NI_3 NS_110 0 -5.7446917270155169e-05
GC_3_111 b_3 NI_3 NS_111 0 -1.9424696358270738e-05
GC_3_112 b_3 NI_3 NS_112 0 2.6716947433710981e-06
GC_3_113 b_3 NI_3 NS_113 0 -1.8170187543826172e-02
GC_3_114 b_3 NI_3 NS_114 0 1.7373059893334120e-03
GC_3_115 b_3 NI_3 NS_115 0 1.3951734051196771e-02
GC_3_116 b_3 NI_3 NS_116 0 3.1643583292137126e-03
GC_3_117 b_3 NI_3 NS_117 0 -7.6251975805356677e-04
GC_3_118 b_3 NI_3 NS_118 0 2.6970870442313171e-04
GC_3_119 b_3 NI_3 NS_119 0 2.5038210343030061e-06
GC_3_120 b_3 NI_3 NS_120 0 6.6504750708737150e-06
GC_3_121 b_3 NI_3 NS_121 0 3.5631160951483552e-04
GC_3_122 b_3 NI_3 NS_122 0 1.1522462673935510e-05
GC_3_123 b_3 NI_3 NS_123 0 8.0008168798941005e-06
GC_3_124 b_3 NI_3 NS_124 0 2.6527859483940873e-06
GC_3_125 b_3 NI_3 NS_125 0 6.4552650206920323e-06
GC_3_126 b_3 NI_3 NS_126 0 3.2976570271709442e-06
GC_3_127 b_3 NI_3 NS_127 0 -5.4277859039638743e-04
GC_3_128 b_3 NI_3 NS_128 0 6.3406073684512624e-04
GC_3_129 b_3 NI_3 NS_129 0 -1.1215077809030826e-04
GC_3_130 b_3 NI_3 NS_130 0 -8.1009608512948184e-05
GC_3_131 b_3 NI_3 NS_131 0 -3.7296206383344493e-05
GC_3_132 b_3 NI_3 NS_132 0 2.8541065043783924e-05
GC_3_133 b_3 NI_3 NS_133 0 4.7915361593402379e-02
GC_3_134 b_3 NI_3 NS_134 0 1.5971319761536287e-02
GC_3_135 b_3 NI_3 NS_135 0 -2.8757406935924212e-02
GC_3_136 b_3 NI_3 NS_136 0 1.3753326472976928e-03
GC_3_137 b_3 NI_3 NS_137 0 -2.8512400701537453e-02
GC_3_138 b_3 NI_3 NS_138 0 -9.2423545748934067e-03
GC_3_139 b_3 NI_3 NS_139 0 8.8978499327095235e-03
GC_3_140 b_3 NI_3 NS_140 0 2.8427078151400300e-03
GC_3_141 b_3 NI_3 NS_141 0 -2.3982359899307197e-03
GC_3_142 b_3 NI_3 NS_142 0 1.3191073929989287e-03
GC_3_143 b_3 NI_3 NS_143 0 2.7612534311523897e-04
GC_3_144 b_3 NI_3 NS_144 0 -3.0765627564851516e-03
GC_3_145 b_3 NI_3 NS_145 0 -4.6989798781392196e-04
GC_3_146 b_3 NI_3 NS_146 0 5.9846086908799712e-05
GC_3_147 b_3 NI_3 NS_147 0 1.1752663190361015e-04
GC_3_148 b_3 NI_3 NS_148 0 8.9982018292484017e-05
GC_3_149 b_3 NI_3 NS_149 0 4.6686419118881911e-04
GC_3_150 b_3 NI_3 NS_150 0 -2.9547342423261495e-04
GC_3_151 b_3 NI_3 NS_151 0 -3.2020721364017119e-05
GC_3_152 b_3 NI_3 NS_152 0 3.0370737140745293e-05
GC_3_153 b_3 NI_3 NS_153 0 -7.0959973586951275e-05
GC_3_154 b_3 NI_3 NS_154 0 6.5733461988627247e-05
GC_3_155 b_3 NI_3 NS_155 0 1.8652103399200443e-06
GC_3_156 b_3 NI_3 NS_156 0 3.3938819522022803e-06
GC_3_157 b_3 NI_3 NS_157 0 1.0171114916568565e-03
GC_3_158 b_3 NI_3 NS_158 0 -9.9018848429361511e-03
GC_3_159 b_3 NI_3 NS_159 0 4.0056175156228799e-05
GC_3_160 b_3 NI_3 NS_160 0 3.7603968721586483e-03
GC_3_161 b_3 NI_3 NS_161 0 4.8108134468997178e-04
GC_3_162 b_3 NI_3 NS_162 0 8.1544504918093139e-05
GC_3_163 b_3 NI_3 NS_163 0 4.1785650785543151e-06
GC_3_164 b_3 NI_3 NS_164 0 2.4976324097938082e-07
GC_3_165 b_3 NI_3 NS_165 0 6.5642130290653286e-05
GC_3_166 b_3 NI_3 NS_166 0 -1.3022910004816007e-04
GC_3_167 b_3 NI_3 NS_167 0 9.2945611738753442e-07
GC_3_168 b_3 NI_3 NS_168 0 -3.5380960473476509e-06
GC_3_169 b_3 NI_3 NS_169 0 2.6304728595304730e-06
GC_3_170 b_3 NI_3 NS_170 0 -5.9534095891791335e-06
GC_3_171 b_3 NI_3 NS_171 0 1.6244642535537008e-04
GC_3_172 b_3 NI_3 NS_172 0 2.9614850722682568e-04
GC_3_173 b_3 NI_3 NS_173 0 2.4506662464002768e-05
GC_3_174 b_3 NI_3 NS_174 0 1.2283545652848078e-04
GC_3_175 b_3 NI_3 NS_175 0 2.0681887042165700e-05
GC_3_176 b_3 NI_3 NS_176 0 9.6888730823881597e-06
GC_3_177 b_3 NI_3 NS_177 0 1.4223626652669791e-02
GC_3_178 b_3 NI_3 NS_178 0 -3.0973857615630891e-04
GC_3_179 b_3 NI_3 NS_179 0 1.5676679373708331e-02
GC_3_180 b_3 NI_3 NS_180 0 -1.5966002381456346e-03
GC_3_181 b_3 NI_3 NS_181 0 -5.5294404200655787e-03
GC_3_182 b_3 NI_3 NS_182 0 -3.2743694507689669e-03
GC_3_183 b_3 NI_3 NS_183 0 1.7870505406364982e-02
GC_3_184 b_3 NI_3 NS_184 0 1.2336324544689961e-02
GC_3_185 b_3 NI_3 NS_185 0 -2.5331500892898404e-03
GC_3_186 b_3 NI_3 NS_186 0 -4.1354013608289686e-03
GC_3_187 b_3 NI_3 NS_187 0 -5.3452539779920340e-03
GC_3_188 b_3 NI_3 NS_188 0 1.2018818856237548e-02
GC_3_189 b_3 NI_3 NS_189 0 7.1888857076216972e-04
GC_3_190 b_3 NI_3 NS_190 0 5.6256742630853896e-04
GC_3_191 b_3 NI_3 NS_191 0 9.4834554646512319e-05
GC_3_192 b_3 NI_3 NS_192 0 3.6208466296416510e-04
GC_3_193 b_3 NI_3 NS_193 0 1.4786223860527783e-03
GC_3_194 b_3 NI_3 NS_194 0 1.8745457771899454e-04
GC_3_195 b_3 NI_3 NS_195 0 2.1471686980834587e-04
GC_3_196 b_3 NI_3 NS_196 0 2.2927059446920748e-04
GC_3_197 b_3 NI_3 NS_197 0 2.9202131855305487e-04
GC_3_198 b_3 NI_3 NS_198 0 1.0185886520755504e-04
GC_3_199 b_3 NI_3 NS_199 0 -1.3096785416745952e-05
GC_3_200 b_3 NI_3 NS_200 0 7.8082902261856918e-06
GC_3_201 b_3 NI_3 NS_201 0 -3.3455247963898267e-02
GC_3_202 b_3 NI_3 NS_202 0 2.6928649732196356e-03
GC_3_203 b_3 NI_3 NS_203 0 2.1120487428676612e-02
GC_3_204 b_3 NI_3 NS_204 0 4.4461598615990802e-03
GC_3_205 b_3 NI_3 NS_205 0 -6.7251109925026804e-04
GC_3_206 b_3 NI_3 NS_206 0 -3.3691729564910269e-04
GC_3_207 b_3 NI_3 NS_207 0 1.4897808941421375e-06
GC_3_208 b_3 NI_3 NS_208 0 3.1634383184073555e-06
GC_3_209 b_3 NI_3 NS_209 0 2.1952963034635838e-04
GC_3_210 b_3 NI_3 NS_210 0 -3.6443569460324473e-05
GC_3_211 b_3 NI_3 NS_211 0 5.4073168165234857e-06
GC_3_212 b_3 NI_3 NS_212 0 1.0081925557529669e-06
GC_3_213 b_3 NI_3 NS_213 0 -1.0329908378027488e-06
GC_3_214 b_3 NI_3 NS_214 0 -6.2435838122103189e-07
GC_3_215 b_3 NI_3 NS_215 0 -1.8707043302684733e-04
GC_3_216 b_3 NI_3 NS_216 0 3.7590705331153317e-04
GC_3_217 b_3 NI_3 NS_217 0 -1.2789170263152870e-05
GC_3_218 b_3 NI_3 NS_218 0 -8.9008967628666482e-05
GC_3_219 b_3 NI_3 NS_219 0 -2.0760710127972431e-05
GC_3_220 b_3 NI_3 NS_220 0 4.9325651137484561e-06
GC_3_221 b_3 NI_3 NS_221 0 2.1741675366189695e-02
GC_3_222 b_3 NI_3 NS_222 0 -7.0767733720997618e-04
GC_3_223 b_3 NI_3 NS_223 0 -2.4103492833784480e-02
GC_3_224 b_3 NI_3 NS_224 0 2.0857034181920894e-03
GC_3_225 b_3 NI_3 NS_225 0 7.8016341299955317e-03
GC_3_226 b_3 NI_3 NS_226 0 -8.9897627851678718e-03
GC_3_227 b_3 NI_3 NS_227 0 1.0382015344121687e-02
GC_3_228 b_3 NI_3 NS_228 0 1.0956933802612930e-03
GC_3_229 b_3 NI_3 NS_229 0 -2.1120333646275075e-05
GC_3_230 b_3 NI_3 NS_230 0 1.0438424227267565e-03
GC_3_231 b_3 NI_3 NS_231 0 -5.6257911855357532e-03
GC_3_232 b_3 NI_3 NS_232 0 -6.4630736150212333e-03
GC_3_233 b_3 NI_3 NS_233 0 -3.6620978047084647e-04
GC_3_234 b_3 NI_3 NS_234 0 1.7291379601823913e-04
GC_3_235 b_3 NI_3 NS_235 0 2.1628794752751208e-04
GC_3_236 b_3 NI_3 NS_236 0 1.0406288522359852e-04
GC_3_237 b_3 NI_3 NS_237 0 5.1664554234098455e-04
GC_3_238 b_3 NI_3 NS_238 0 3.2572089182577641e-04
GC_3_239 b_3 NI_3 NS_239 0 3.0771089761707460e-05
GC_3_240 b_3 NI_3 NS_240 0 4.4270873586857578e-05
GC_3_241 b_3 NI_3 NS_241 0 7.3720422870342101e-05
GC_3_242 b_3 NI_3 NS_242 0 9.8804042275413918e-06
GC_3_243 b_3 NI_3 NS_243 0 8.8736175996251663e-06
GC_3_244 b_3 NI_3 NS_244 0 -4.4111079800970683e-07
GC_3_245 b_3 NI_3 NS_245 0 -4.0603204597325325e-03
GC_3_246 b_3 NI_3 NS_246 0 6.9355308562863765e-03
GC_3_247 b_3 NI_3 NS_247 0 4.2510532902142262e-03
GC_3_248 b_3 NI_3 NS_248 0 -3.0466215039097197e-03
GC_3_249 b_3 NI_3 NS_249 0 -9.3510920506006452e-05
GC_3_250 b_3 NI_3 NS_250 0 3.0181678768575303e-05
GC_3_251 b_3 NI_3 NS_251 0 -1.2736045548841011e-07
GC_3_252 b_3 NI_3 NS_252 0 -2.3136946864205961e-08
GC_3_253 b_3 NI_3 NS_253 0 6.4282585786969694e-06
GC_3_254 b_3 NI_3 NS_254 0 1.2877456111551223e-05
GC_3_255 b_3 NI_3 NS_255 0 -5.3253719615631635e-07
GC_3_256 b_3 NI_3 NS_256 0 -2.3353212463985216e-07
GC_3_257 b_3 NI_3 NS_257 0 -1.4391840947799488e-06
GC_3_258 b_3 NI_3 NS_258 0 -2.3459791001721972e-06
GC_3_259 b_3 NI_3 NS_259 0 1.8411541441817349e-05
GC_3_260 b_3 NI_3 NS_260 0 5.8513725805609235e-06
GC_3_261 b_3 NI_3 NS_261 0 7.0700508735435422e-06
GC_3_262 b_3 NI_3 NS_262 0 2.3792649206594840e-05
GC_3_263 b_3 NI_3 NS_263 0 1.7612973072003936e-06
GC_3_264 b_3 NI_3 NS_264 0 -4.1088855641296963e-06
GC_3_265 b_3 NI_3 NS_265 0 9.9818664266472356e-03
GC_3_266 b_3 NI_3 NS_266 0 1.5045400667278486e-04
GC_3_267 b_3 NI_3 NS_267 0 1.1789443444855486e-02
GC_3_268 b_3 NI_3 NS_268 0 -5.2505934137347544e-03
GC_3_269 b_3 NI_3 NS_269 0 -1.9371351844908013e-03
GC_3_270 b_3 NI_3 NS_270 0 4.9258926213427571e-03
GC_3_271 b_3 NI_3 NS_271 0 1.2517409746386913e-02
GC_3_272 b_3 NI_3 NS_272 0 8.9652562394798435e-03
GC_3_273 b_3 NI_3 NS_273 0 -1.9239124801317222e-03
GC_3_274 b_3 NI_3 NS_274 0 -2.4865856789162265e-03
GC_3_275 b_3 NI_3 NS_275 0 -9.7661868281680650e-03
GC_3_276 b_3 NI_3 NS_276 0 8.8928008328628960e-03
GC_3_277 b_3 NI_3 NS_277 0 5.8049079826563905e-04
GC_3_278 b_3 NI_3 NS_278 0 3.7355971365069386e-04
GC_3_279 b_3 NI_3 NS_279 0 1.2603095789338282e-04
GC_3_280 b_3 NI_3 NS_280 0 2.9540492461346249e-04
GC_3_281 b_3 NI_3 NS_281 0 9.7537432970563041e-04
GC_3_282 b_3 NI_3 NS_282 0 -9.0222303389438088e-05
GC_3_283 b_3 NI_3 NS_283 0 1.9116872871042425e-04
GC_3_284 b_3 NI_3 NS_284 0 1.5172835083544702e-04
GC_3_285 b_3 NI_3 NS_285 0 1.1166578991576264e-04
GC_3_286 b_3 NI_3 NS_286 0 1.4012369637789382e-05
GC_3_287 b_3 NI_3 NS_287 0 -5.6488213994867477e-06
GC_3_288 b_3 NI_3 NS_288 0 2.2481555752385798e-06
GC_3_289 b_3 NI_3 NS_289 0 -2.0697010641674653e-02
GC_3_290 b_3 NI_3 NS_290 0 4.1956786199619049e-04
GC_3_291 b_3 NI_3 NS_291 0 1.3340586991600638e-02
GC_3_292 b_3 NI_3 NS_292 0 2.3195750793341590e-03
GC_3_293 b_3 NI_3 NS_293 0 -3.0587828970185781e-04
GC_3_294 b_3 NI_3 NS_294 0 -4.5083622758731150e-04
GC_3_295 b_3 NI_3 NS_295 0 9.6451887130752166e-07
GC_3_296 b_3 NI_3 NS_296 0 5.6514710221454092e-07
GC_3_297 b_3 NI_3 NS_297 0 9.5799145236937422e-05
GC_3_298 b_3 NI_3 NS_298 0 -6.0553483481303252e-05
GC_3_299 b_3 NI_3 NS_299 0 1.8789972871154825e-06
GC_3_300 b_3 NI_3 NS_300 0 3.9977701151920802e-07
GC_3_301 b_3 NI_3 NS_301 0 -1.2005928945910056e-06
GC_3_302 b_3 NI_3 NS_302 0 -1.9855078906174725e-06
GC_3_303 b_3 NI_3 NS_303 0 -9.4007608697232070e-06
GC_3_304 b_3 NI_3 NS_304 0 2.6929478439757267e-04
GC_3_305 b_3 NI_3 NS_305 0 -7.9152312476896792e-06
GC_3_306 b_3 NI_3 NS_306 0 -5.6596677515233401e-05
GC_3_307 b_3 NI_3 NS_307 0 -1.3865358019719997e-05
GC_3_308 b_3 NI_3 NS_308 0 -1.0496156926827372e-06
GC_3_309 b_3 NI_3 NS_309 0 1.0514065926683335e-02
GC_3_310 b_3 NI_3 NS_310 0 -5.4058377238724051e-04
GC_3_311 b_3 NI_3 NS_311 0 -1.5154914903478879e-02
GC_3_312 b_3 NI_3 NS_312 0 5.6633492917475582e-03
GC_3_313 b_3 NI_3 NS_313 0 2.8294697761629497e-03
GC_3_314 b_3 NI_3 NS_314 0 -1.2088446004758299e-02
GC_3_315 b_3 NI_3 NS_315 0 8.3137025276588811e-03
GC_3_316 b_3 NI_3 NS_316 0 6.6309770995876601e-04
GC_3_317 b_3 NI_3 NS_317 0 -3.4484997010453744e-04
GC_3_318 b_3 NI_3 NS_318 0 -2.8598223431094559e-05
GC_3_319 b_3 NI_3 NS_319 0 -6.7348291807615935e-03
GC_3_320 b_3 NI_3 NS_320 0 -3.2229970949927663e-03
GC_3_321 b_3 NI_3 NS_321 0 -2.4894218878713723e-04
GC_3_322 b_3 NI_3 NS_322 0 1.1680764457510104e-04
GC_3_323 b_3 NI_3 NS_323 0 1.7347978838582275e-04
GC_3_324 b_3 NI_3 NS_324 0 4.1149025659726604e-05
GC_3_325 b_3 NI_3 NS_325 0 4.6942272912431750e-04
GC_3_326 b_3 NI_3 NS_326 0 1.4013402084152204e-04
GC_3_327 b_3 NI_3 NS_327 0 1.2727223475254973e-06
GC_3_328 b_3 NI_3 NS_328 0 1.1211335419864816e-05
GC_3_329 b_3 NI_3 NS_329 0 -3.7678167085417257e-07
GC_3_330 b_3 NI_3 NS_330 0 -1.4114224300075281e-05
GC_3_331 b_3 NI_3 NS_331 0 3.0806649660894553e-06
GC_3_332 b_3 NI_3 NS_332 0 -5.3051361945933962e-07
GC_3_333 b_3 NI_3 NS_333 0 2.3954362665705550e-03
GC_3_334 b_3 NI_3 NS_334 0 3.3323572354617974e-03
GC_3_335 b_3 NI_3 NS_335 0 5.1032123516019914e-04
GC_3_336 b_3 NI_3 NS_336 0 -2.1558234051126455e-03
GC_3_337 b_3 NI_3 NS_337 0 6.6241398565062049e-05
GC_3_338 b_3 NI_3 NS_338 0 5.4420217290948517e-05
GC_3_339 b_3 NI_3 NS_339 0 6.4337507987730588e-07
GC_3_340 b_3 NI_3 NS_340 0 4.1806208402951689e-07
GC_3_341 b_3 NI_3 NS_341 0 2.2552325329624595e-05
GC_3_342 b_3 NI_3 NS_342 0 -7.9382844953445705e-06
GC_3_343 b_3 NI_3 NS_343 0 2.1940902841156775e-07
GC_3_344 b_3 NI_3 NS_344 0 -1.4624724365574025e-07
GC_3_345 b_3 NI_3 NS_345 0 2.9189598158209083e-07
GC_3_346 b_3 NI_3 NS_346 0 -1.2057456190553936e-06
GC_3_347 b_3 NI_3 NS_347 0 -4.4287581135649081e-05
GC_3_348 b_3 NI_3 NS_348 0 5.0083392130126345e-05
GC_3_349 b_3 NI_3 NS_349 0 -8.6788980108762931e-06
GC_3_350 b_3 NI_3 NS_350 0 3.3894161815937742e-05
GC_3_351 b_3 NI_3 NS_351 0 3.5248380954808508e-06
GC_3_352 b_3 NI_3 NS_352 0 2.2051796556769641e-06
GC_3_353 b_3 NI_3 NS_353 0 -1.6010149182668500e-02
GC_3_354 b_3 NI_3 NS_354 0 8.4556712492892764e-05
GC_3_355 b_3 NI_3 NS_355 0 -1.0880593474425024e-03
GC_3_356 b_3 NI_3 NS_356 0 -1.3722877455202456e-03
GC_3_357 b_3 NI_3 NS_357 0 7.2095672858100794e-04
GC_3_358 b_3 NI_3 NS_358 0 -2.0089286349000228e-03
GC_3_359 b_3 NI_3 NS_359 0 1.8327073446930469e-03
GC_3_360 b_3 NI_3 NS_360 0 -2.4202876331503227e-03
GC_3_361 b_3 NI_3 NS_361 0 7.5045369873770723e-04
GC_3_362 b_3 NI_3 NS_362 0 9.8520254495161911e-04
GC_3_363 b_3 NI_3 NS_363 0 -6.7278517476796872e-04
GC_3_364 b_3 NI_3 NS_364 0 6.0838331308309124e-04
GC_3_365 b_3 NI_3 NS_365 0 4.6813767728830409e-04
GC_3_366 b_3 NI_3 NS_366 0 -3.4954146279999877e-04
GC_3_367 b_3 NI_3 NS_367 0 4.0783402292011653e-04
GC_3_368 b_3 NI_3 NS_368 0 8.7236767648586687e-04
GC_3_369 b_3 NI_3 NS_369 0 -2.7876297777501562e-03
GC_3_370 b_3 NI_3 NS_370 0 -2.2314859015542836e-03
GC_3_371 b_3 NI_3 NS_371 0 2.0925991794825481e-04
GC_3_372 b_3 NI_3 NS_372 0 1.4856713555089823e-04
GC_3_373 b_3 NI_3 NS_373 0 -1.0575707871659915e-03
GC_3_374 b_3 NI_3 NS_374 0 9.2076646970828329e-07
GC_3_375 b_3 NI_3 NS_375 0 -2.5480238822899758e-06
GC_3_376 b_3 NI_3 NS_376 0 -3.7622174150004497e-06
GC_3_377 b_3 NI_3 NS_377 0 1.5846693001629501e-02
GC_3_378 b_3 NI_3 NS_378 0 8.8977282823703447e-03
GC_3_379 b_3 NI_3 NS_379 0 -7.8134765697878139e-03
GC_3_380 b_3 NI_3 NS_380 0 -1.1117849172032195e-02
GC_3_381 b_3 NI_3 NS_381 0 -2.0510235383942845e-05
GC_3_382 b_3 NI_3 NS_382 0 5.3591418898104768e-04
GC_3_383 b_3 NI_3 NS_383 0 5.5993450234157323e-08
GC_3_384 b_3 NI_3 NS_384 0 4.5085408719189517e-08
GC_3_385 b_3 NI_3 NS_385 0 -1.2243503354682328e-05
GC_3_386 b_3 NI_3 NS_386 0 -9.8372915013640973e-05
GC_3_387 b_3 NI_3 NS_387 0 4.3589435743686852e-07
GC_3_388 b_3 NI_3 NS_388 0 6.3551889308878739e-07
GC_3_389 b_3 NI_3 NS_389 0 -1.5228888850347835e-07
GC_3_390 b_3 NI_3 NS_390 0 -4.7680094947881860e-06
GC_3_391 b_3 NI_3 NS_391 0 3.2025091371565403e-04
GC_3_392 b_3 NI_3 NS_392 0 5.9623175434196445e-04
GC_3_393 b_3 NI_3 NS_393 0 -2.2013619201618334e-04
GC_3_394 b_3 NI_3 NS_394 0 1.1583315698659160e-04
GC_3_395 b_3 NI_3 NS_395 0 -1.8662076386431280e-05
GC_3_396 b_3 NI_3 NS_396 0 -8.2192323719456198e-06
GC_3_397 b_3 NI_3 NS_397 0 -3.2927922961638700e-03
GC_3_398 b_3 NI_3 NS_398 0 2.2446999109706871e-05
GC_3_399 b_3 NI_3 NS_399 0 -2.3649087140605989e-04
GC_3_400 b_3 NI_3 NS_400 0 1.1270724318279439e-03
GC_3_401 b_3 NI_3 NS_401 0 -1.9781904552553125e-03
GC_3_402 b_3 NI_3 NS_402 0 -1.0394287052698156e-03
GC_3_403 b_3 NI_3 NS_403 0 -1.1642155414616026e-04
GC_3_404 b_3 NI_3 NS_404 0 -2.1027193702562834e-03
GC_3_405 b_3 NI_3 NS_405 0 5.4967923160493528e-04
GC_3_406 b_3 NI_3 NS_406 0 4.3256135722494671e-04
GC_3_407 b_3 NI_3 NS_407 0 1.0728716969328591e-03
GC_3_408 b_3 NI_3 NS_408 0 -1.4856778190178816e-03
GC_3_409 b_3 NI_3 NS_409 0 -2.5758262341967766e-05
GC_3_410 b_3 NI_3 NS_410 0 2.8541115645756404e-04
GC_3_411 b_3 NI_3 NS_411 0 2.8697881013268578e-04
GC_3_412 b_3 NI_3 NS_412 0 -8.1332166019807737e-05
GC_3_413 b_3 NI_3 NS_413 0 -4.2960364440455107e-04
GC_3_414 b_3 NI_3 NS_414 0 3.7185475766022679e-05
GC_3_415 b_3 NI_3 NS_415 0 -2.1485800825336442e-05
GC_3_416 b_3 NI_3 NS_416 0 -1.3805957371859979e-06
GC_3_417 b_3 NI_3 NS_417 0 -5.7868421056367109e-05
GC_3_418 b_3 NI_3 NS_418 0 -4.1755665060971059e-05
GC_3_419 b_3 NI_3 NS_419 0 4.8360285740504658e-06
GC_3_420 b_3 NI_3 NS_420 0 4.8951747508091937e-06
GC_3_421 b_3 NI_3 NS_421 0 4.7302599547250235e-03
GC_3_422 b_3 NI_3 NS_422 0 2.0426220108515896e-03
GC_3_423 b_3 NI_3 NS_423 0 -2.8695060019956146e-03
GC_3_424 b_3 NI_3 NS_424 0 -2.1824961772422798e-03
GC_3_425 b_3 NI_3 NS_425 0 -1.0021021831686385e-04
GC_3_426 b_3 NI_3 NS_426 0 1.3801248494341171e-05
GC_3_427 b_3 NI_3 NS_427 0 -6.5732898542746740e-07
GC_3_428 b_3 NI_3 NS_428 0 -3.0161191679736624e-07
GC_3_429 b_3 NI_3 NS_429 0 -1.2367332438227706e-05
GC_3_430 b_3 NI_3 NS_430 0 4.0147865683002198e-05
GC_3_431 b_3 NI_3 NS_431 0 1.0315818908457609e-06
GC_3_432 b_3 NI_3 NS_432 0 4.3900986527226275e-07
GC_3_433 b_3 NI_3 NS_433 0 -1.8678496968872799e-06
GC_3_434 b_3 NI_3 NS_434 0 -1.1860836047516723e-06
GC_3_435 b_3 NI_3 NS_435 0 -5.2268710855586364e-05
GC_3_436 b_3 NI_3 NS_436 0 -2.9095808706970414e-05
GC_3_437 b_3 NI_3 NS_437 0 -1.8127078908078359e-05
GC_3_438 b_3 NI_3 NS_438 0 -1.5549735082517286e-05
GC_3_439 b_3 NI_3 NS_439 0 4.3221708449817870e-06
GC_3_440 b_3 NI_3 NS_440 0 1.7151045971610601e-07
GC_3_441 b_3 NI_3 NS_441 0 -8.0348016256092270e-03
GC_3_442 b_3 NI_3 NS_442 0 1.0429383636467543e-04
GC_3_443 b_3 NI_3 NS_443 0 5.9391707802425829e-04
GC_3_444 b_3 NI_3 NS_444 0 -2.3916223286929855e-03
GC_3_445 b_3 NI_3 NS_445 0 1.3647430122116352e-03
GC_3_446 b_3 NI_3 NS_446 0 1.3617959295743112e-04
GC_3_447 b_3 NI_3 NS_447 0 3.5000027138475851e-03
GC_3_448 b_3 NI_3 NS_448 0 -1.1114017620298404e-04
GC_3_449 b_3 NI_3 NS_449 0 1.4459670201228170e-04
GC_3_450 b_3 NI_3 NS_450 0 1.5316438455604780e-04
GC_3_451 b_3 NI_3 NS_451 0 -2.7995810230831502e-03
GC_3_452 b_3 NI_3 NS_452 0 3.3982189247359755e-03
GC_3_453 b_3 NI_3 NS_453 0 4.2530722700843379e-04
GC_3_454 b_3 NI_3 NS_454 0 -1.6037878302582552e-04
GC_3_455 b_3 NI_3 NS_455 0 2.9696162102112368e-04
GC_3_456 b_3 NI_3 NS_456 0 6.1054349855272619e-04
GC_3_457 b_3 NI_3 NS_457 0 -1.7227385516026253e-03
GC_3_458 b_3 NI_3 NS_458 0 -1.3974823703959082e-03
GC_3_459 b_3 NI_3 NS_459 0 1.6234919172520480e-04
GC_3_460 b_3 NI_3 NS_460 0 1.2334858519874283e-04
GC_3_461 b_3 NI_3 NS_461 0 -6.9908029337138321e-04
GC_3_462 b_3 NI_3 NS_462 0 1.9751111344512685e-05
GC_3_463 b_3 NI_3 NS_463 0 -5.8763602407442118e-07
GC_3_464 b_3 NI_3 NS_464 0 -6.5881360554105371e-08
GC_3_465 b_3 NI_3 NS_465 0 6.4245482704139009e-03
GC_3_466 b_3 NI_3 NS_466 0 4.2081817224467917e-03
GC_3_467 b_3 NI_3 NS_467 0 -3.2245895015618415e-03
GC_3_468 b_3 NI_3 NS_468 0 -6.0058478263659400e-03
GC_3_469 b_3 NI_3 NS_469 0 4.7623577950774595e-05
GC_3_470 b_3 NI_3 NS_470 0 1.9860905205659461e-04
GC_3_471 b_3 NI_3 NS_471 0 3.7434772286744391e-07
GC_3_472 b_3 NI_3 NS_472 0 -3.9527667857787822e-07
GC_3_473 b_3 NI_3 NS_473 0 -3.4600673598509526e-06
GC_3_474 b_3 NI_3 NS_474 0 -9.3206189895150211e-05
GC_3_475 b_3 NI_3 NS_475 0 1.5136865835435192e-08
GC_3_476 b_3 NI_3 NS_476 0 -2.5600280302233607e-07
GC_3_477 b_3 NI_3 NS_477 0 -1.1334647212819928e-06
GC_3_478 b_3 NI_3 NS_478 0 -3.8905051214204694e-06
GC_3_479 b_3 NI_3 NS_479 0 2.2688940327503983e-04
GC_3_480 b_3 NI_3 NS_480 0 4.1172440467019425e-04
GC_3_481 b_3 NI_3 NS_481 0 -1.3790953426108768e-04
GC_3_482 b_3 NI_3 NS_482 0 7.5855376296043016e-05
GC_3_483 b_3 NI_3 NS_483 0 -1.2034996968776552e-05
GC_3_484 b_3 NI_3 NS_484 0 -5.7495618201676371e-06
GC_3_485 b_3 NI_3 NS_485 0 1.8353629104700040e-03
GC_3_486 b_3 NI_3 NS_486 0 -8.1496573541571882e-05
GC_3_487 b_3 NI_3 NS_487 0 -1.4246904317904547e-03
GC_3_488 b_3 NI_3 NS_488 0 2.3503729805299657e-03
GC_3_489 b_3 NI_3 NS_489 0 -2.0309473490100470e-03
GC_3_490 b_3 NI_3 NS_490 0 -2.5779773943458055e-03
GC_3_491 b_3 NI_3 NS_491 0 1.3478924619197427e-03
GC_3_492 b_3 NI_3 NS_492 0 -1.4137399015678493e-03
GC_3_493 b_3 NI_3 NS_493 0 -1.6671024045145310e-05
GC_3_494 b_3 NI_3 NS_494 0 3.0109292261389575e-04
GC_3_495 b_3 NI_3 NS_495 0 -8.3429487393368244e-04
GC_3_496 b_3 NI_3 NS_496 0 -1.6100691876835021e-04
GC_3_497 b_3 NI_3 NS_497 0 -5.0045096989815016e-05
GC_3_498 b_3 NI_3 NS_498 0 1.9961663943035302e-04
GC_3_499 b_3 NI_3 NS_499 0 2.2201615080162941e-04
GC_3_500 b_3 NI_3 NS_500 0 -3.2028405179766663e-05
GC_3_501 b_3 NI_3 NS_501 0 -2.5660035049352960e-04
GC_3_502 b_3 NI_3 NS_502 0 3.4517837272104223e-05
GC_3_503 b_3 NI_3 NS_503 0 -2.6981829216080875e-05
GC_3_504 b_3 NI_3 NS_504 0 -4.7971095406651899e-06
GC_3_505 b_3 NI_3 NS_505 0 -2.0765423613329695e-05
GC_3_506 b_3 NI_3 NS_506 0 -1.8735738993391274e-05
GC_3_507 b_3 NI_3 NS_507 0 2.9422995686381803e-06
GC_3_508 b_3 NI_3 NS_508 0 1.6729852798682420e-06
GC_3_509 b_3 NI_3 NS_509 0 2.6680134013143367e-03
GC_3_510 b_3 NI_3 NS_510 0 1.0553606427033224e-03
GC_3_511 b_3 NI_3 NS_511 0 -1.3904690700025379e-03
GC_3_512 b_3 NI_3 NS_512 0 -1.4499572984550341e-03
GC_3_513 b_3 NI_3 NS_513 0 -3.5086163313818228e-05
GC_3_514 b_3 NI_3 NS_514 0 -5.9577560389251098e-05
GC_3_515 b_3 NI_3 NS_515 0 -4.1939740353587795e-07
GC_3_516 b_3 NI_3 NS_516 0 -4.0902891029164559e-07
GC_3_517 b_3 NI_3 NS_517 0 -1.1418185354749896e-05
GC_3_518 b_3 NI_3 NS_518 0 1.0428347168362962e-05
GC_3_519 b_3 NI_3 NS_519 0 -2.6985344143655277e-07
GC_3_520 b_3 NI_3 NS_520 0 4.0623754427013945e-07
GC_3_521 b_3 NI_3 NS_521 0 -9.5997446118416732e-07
GC_3_522 b_3 NI_3 NS_522 0 -1.2878619097707974e-06
GC_3_523 b_3 NI_3 NS_523 0 -1.8954257541954429e-05
GC_3_524 b_3 NI_3 NS_524 0 -3.4595309187475390e-05
GC_3_525 b_3 NI_3 NS_525 0 1.1022922227450960e-05
GC_3_526 b_3 NI_3 NS_526 0 -9.1976516587123689e-06
GC_3_527 b_3 NI_3 NS_527 0 5.5940253281885001e-06
GC_3_528 b_3 NI_3 NS_528 0 -8.7726319169230972e-07
GD_3_1 b_3 NI_3 NA_1 0 -2.4065254918726079e-02
GD_3_2 b_3 NI_3 NA_2 0 -2.4079607663055596e-03
GD_3_3 b_3 NI_3 NA_3 0 -1.8278252519559415e-01
GD_3_4 b_3 NI_3 NA_4 0 -1.7485402243864127e-02
GD_3_5 b_3 NI_3 NA_5 0 -3.0752557099565085e-02
GD_3_6 b_3 NI_3 NA_6 0 -1.3246278655179388e-02
GD_3_7 b_3 NI_3 NA_7 0 -2.0609250360912140e-02
GD_3_8 b_3 NI_3 NA_8 0 -2.8358596812269074e-03
GD_3_9 b_3 NI_3 NA_9 0 9.8570499901989312e-03
GD_3_10 b_3 NI_3 NA_10 0 2.6616533358836208e-03
GD_3_11 b_3 NI_3 NA_11 0 3.4474710667440731e-03
GD_3_12 b_3 NI_3 NA_12 0 2.3832794159979101e-04
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 6.1783341262029723e-03
GC_4_2 b_4 NI_4 NS_2 0 -3.7221244443596261e-04
GC_4_3 b_4 NI_4 NS_3 0 -2.0234199944319471e-02
GC_4_4 b_4 NI_4 NS_4 0 -3.0973193626438939e-03
GC_4_5 b_4 NI_4 NS_5 0 1.0273186404537362e-02
GC_4_6 b_4 NI_4 NS_6 0 -3.0432489324587540e-03
GC_4_7 b_4 NI_4 NS_7 0 5.8008064102920464e-03
GC_4_8 b_4 NI_4 NS_8 0 1.0544994379757121e-03
GC_4_9 b_4 NI_4 NS_9 0 1.8472440092425694e-03
GC_4_10 b_4 NI_4 NS_10 0 -5.2924024160640442e-04
GC_4_11 b_4 NI_4 NS_11 0 -7.2836452790909698e-04
GC_4_12 b_4 NI_4 NS_12 0 -8.7666286246266302e-03
GC_4_13 b_4 NI_4 NS_13 0 -2.7303355822279275e-04
GC_4_14 b_4 NI_4 NS_14 0 3.8620741870171360e-05
GC_4_15 b_4 NI_4 NS_15 0 1.7685662290313465e-04
GC_4_16 b_4 NI_4 NS_16 0 6.2209955780342634e-05
GC_4_17 b_4 NI_4 NS_17 0 5.4327097672080557e-04
GC_4_18 b_4 NI_4 NS_18 0 4.8081377505043829e-04
GC_4_19 b_4 NI_4 NS_19 0 3.4810666064097418e-05
GC_4_20 b_4 NI_4 NS_20 0 3.3290197896480915e-05
GC_4_21 b_4 NI_4 NS_21 0 6.9368235382617210e-05
GC_4_22 b_4 NI_4 NS_22 0 1.1406950112367583e-05
GC_4_23 b_4 NI_4 NS_23 0 5.3522247266539885e-06
GC_4_24 b_4 NI_4 NS_24 0 -1.9451375006848099e-06
GC_4_25 b_4 NI_4 NS_25 0 -6.4795852496093657e-03
GC_4_26 b_4 NI_4 NS_26 0 8.1058085975647051e-03
GC_4_27 b_4 NI_4 NS_27 0 4.7484983140312917e-03
GC_4_28 b_4 NI_4 NS_28 0 -3.1909267764570039e-03
GC_4_29 b_4 NI_4 NS_29 0 -1.9213544848577357e-04
GC_4_30 b_4 NI_4 NS_30 0 1.8309860619135753e-04
GC_4_31 b_4 NI_4 NS_31 0 -5.3295997558411010e-07
GC_4_32 b_4 NI_4 NS_32 0 2.6108714931117942e-07
GC_4_33 b_4 NI_4 NS_33 0 8.9411675081872319e-06
GC_4_34 b_4 NI_4 NS_34 0 4.4378722599479839e-05
GC_4_35 b_4 NI_4 NS_35 0 1.0538695980969583e-07
GC_4_36 b_4 NI_4 NS_36 0 8.1440759073995813e-07
GC_4_37 b_4 NI_4 NS_37 0 1.6344353782001432e-07
GC_4_38 b_4 NI_4 NS_38 0 1.3798537923857795e-06
GC_4_39 b_4 NI_4 NS_39 0 -5.6397528022989057e-05
GC_4_40 b_4 NI_4 NS_40 0 -1.6206890529575724e-04
GC_4_41 b_4 NI_4 NS_41 0 -5.7041757654037006e-07
GC_4_42 b_4 NI_4 NS_42 0 -1.1831905612843739e-05
GC_4_43 b_4 NI_4 NS_43 0 -1.7424126409177897e-07
GC_4_44 b_4 NI_4 NS_44 0 -6.0528681451814752e-06
GC_4_45 b_4 NI_4 NS_45 0 -4.6974782809280132e-03
GC_4_46 b_4 NI_4 NS_46 0 -1.0219314154766006e-03
GC_4_47 b_4 NI_4 NS_47 0 1.4143515812236260e-02
GC_4_48 b_4 NI_4 NS_48 0 3.3541475722908389e-03
GC_4_49 b_4 NI_4 NS_49 0 -1.6532589860789499e-02
GC_4_50 b_4 NI_4 NS_50 0 -2.9391657335733927e-03
GC_4_51 b_4 NI_4 NS_51 0 5.2421008818710133e-03
GC_4_52 b_4 NI_4 NS_52 0 -8.9796558994732702e-04
GC_4_53 b_4 NI_4 NS_53 0 -8.8370735471972328e-04
GC_4_54 b_4 NI_4 NS_54 0 5.2597544400287757e-04
GC_4_55 b_4 NI_4 NS_55 0 1.0495816932239628e-03
GC_4_56 b_4 NI_4 NS_56 0 -3.0938269122137425e-03
GC_4_57 b_4 NI_4 NS_57 0 1.1507895503848395e-04
GC_4_58 b_4 NI_4 NS_58 0 -1.2392893254714273e-04
GC_4_59 b_4 NI_4 NS_59 0 2.3712826130554969e-05
GC_4_60 b_4 NI_4 NS_60 0 -3.5725294380198096e-05
GC_4_61 b_4 NI_4 NS_61 0 1.2015434770202043e-04
GC_4_62 b_4 NI_4 NS_62 0 -2.4359365421515470e-05
GC_4_63 b_4 NI_4 NS_63 0 1.4668317054347507e-05
GC_4_64 b_4 NI_4 NS_64 0 -6.0990489158875720e-06
GC_4_65 b_4 NI_4 NS_65 0 8.0170528190423660e-06
GC_4_66 b_4 NI_4 NS_66 0 -1.9004397230473473e-05
GC_4_67 b_4 NI_4 NS_67 0 -2.5995820307280302e-06
GC_4_68 b_4 NI_4 NS_68 0 -7.0854473254512714e-07
GC_4_69 b_4 NI_4 NS_69 0 4.5887345056465668e-03
GC_4_70 b_4 NI_4 NS_70 0 7.1101836417827970e-03
GC_4_71 b_4 NI_4 NS_71 0 -1.4957572226655337e-03
GC_4_72 b_4 NI_4 NS_72 0 -3.4097038649938162e-03
GC_4_73 b_4 NI_4 NS_73 0 -2.1124898861449068e-04
GC_4_74 b_4 NI_4 NS_74 0 -7.0861499212812105e-05
GC_4_75 b_4 NI_4 NS_75 0 -4.4002827903363854e-07
GC_4_76 b_4 NI_4 NS_76 0 4.6990824273337577e-07
GC_4_77 b_4 NI_4 NS_77 0 -6.5632200379890507e-05
GC_4_78 b_4 NI_4 NS_78 0 1.0730972501738933e-04
GC_4_79 b_4 NI_4 NS_79 0 -3.6452483014564038e-06
GC_4_80 b_4 NI_4 NS_80 0 -2.4918352824924615e-06
GC_4_81 b_4 NI_4 NS_81 0 -5.8478048547213910e-06
GC_4_82 b_4 NI_4 NS_82 0 -1.2234873010122276e-05
GC_4_83 b_4 NI_4 NS_83 0 -2.5290690076043668e-04
GC_4_84 b_4 NI_4 NS_84 0 7.1593872813307933e-05
GC_4_85 b_4 NI_4 NS_85 0 -1.2524514827130293e-04
GC_4_86 b_4 NI_4 NS_86 0 -5.0326143957762851e-05
GC_4_87 b_4 NI_4 NS_87 0 -3.0547799761842503e-05
GC_4_88 b_4 NI_4 NS_88 0 -7.1780745154985500e-06
GC_4_89 b_4 NI_4 NS_89 0 4.7915361593392665e-02
GC_4_90 b_4 NI_4 NS_90 0 1.5971319761536505e-02
GC_4_91 b_4 NI_4 NS_91 0 -2.8757406935924198e-02
GC_4_92 b_4 NI_4 NS_92 0 1.3753326472961973e-03
GC_4_93 b_4 NI_4 NS_93 0 -2.8512400701535802e-02
GC_4_94 b_4 NI_4 NS_94 0 -9.2423545748938126e-03
GC_4_95 b_4 NI_4 NS_95 0 8.8978499327101428e-03
GC_4_96 b_4 NI_4 NS_96 0 2.8427078151398301e-03
GC_4_97 b_4 NI_4 NS_97 0 -2.3982359899299460e-03
GC_4_98 b_4 NI_4 NS_98 0 1.3191073929996870e-03
GC_4_99 b_4 NI_4 NS_99 0 2.7612534311584200e-04
GC_4_100 b_4 NI_4 NS_100 0 -3.0765627564858572e-03
GC_4_101 b_4 NI_4 NS_101 0 -4.6989798781391551e-04
GC_4_102 b_4 NI_4 NS_102 0 5.9846086908823409e-05
GC_4_103 b_4 NI_4 NS_103 0 1.1752663190356849e-04
GC_4_104 b_4 NI_4 NS_104 0 8.9982018292506378e-05
GC_4_105 b_4 NI_4 NS_105 0 4.6686419118877086e-04
GC_4_106 b_4 NI_4 NS_106 0 -2.9547342423287879e-04
GC_4_107 b_4 NI_4 NS_107 0 -3.2020721364036669e-05
GC_4_108 b_4 NI_4 NS_108 0 3.0370737140724568e-05
GC_4_109 b_4 NI_4 NS_109 0 -7.0959973587001406e-05
GC_4_110 b_4 NI_4 NS_110 0 6.5733461988587958e-05
GC_4_111 b_4 NI_4 NS_111 0 1.8652103399172036e-06
GC_4_112 b_4 NI_4 NS_112 0 3.3938819521982248e-06
GC_4_113 b_4 NI_4 NS_113 0 1.0171114916605359e-03
GC_4_114 b_4 NI_4 NS_114 0 -9.9018848429358684e-03
GC_4_115 b_4 NI_4 NS_115 0 4.0056175154542255e-05
GC_4_116 b_4 NI_4 NS_116 0 3.7603968721580056e-03
GC_4_117 b_4 NI_4 NS_117 0 4.8108134469001325e-04
GC_4_118 b_4 NI_4 NS_118 0 8.1544504918310020e-05
GC_4_119 b_4 NI_4 NS_119 0 4.1785650785547844e-06
GC_4_120 b_4 NI_4 NS_120 0 2.4976324098048355e-07
GC_4_121 b_4 NI_4 NS_121 0 6.5642130290714028e-05
GC_4_122 b_4 NI_4 NS_122 0 -1.3022910004815538e-04
GC_4_123 b_4 NI_4 NS_123 0 9.2945611738956041e-07
GC_4_124 b_4 NI_4 NS_124 0 -3.5380960473484255e-06
GC_4_125 b_4 NI_4 NS_125 0 2.6304728595304260e-06
GC_4_126 b_4 NI_4 NS_126 0 -5.9534095891798136e-06
GC_4_127 b_4 NI_4 NS_127 0 1.6244642535533831e-04
GC_4_128 b_4 NI_4 NS_128 0 2.9614850722689355e-04
GC_4_129 b_4 NI_4 NS_129 0 2.4506662463982954e-05
GC_4_130 b_4 NI_4 NS_130 0 1.2283545652850428e-04
GC_4_131 b_4 NI_4 NS_131 0 2.0681887042166642e-05
GC_4_132 b_4 NI_4 NS_132 0 9.6888730823957779e-06
GC_4_133 b_4 NI_4 NS_133 0 -1.3920303386949562e-01
GC_4_134 b_4 NI_4 NS_134 0 1.7536159600762654e-02
GC_4_135 b_4 NI_4 NS_135 0 1.6547474721776621e-02
GC_4_136 b_4 NI_4 NS_136 0 5.2069216487723394e-03
GC_4_137 b_4 NI_4 NS_137 0 1.7153371397962826e-02
GC_4_138 b_4 NI_4 NS_138 0 -3.0586379387722200e-03
GC_4_139 b_4 NI_4 NS_139 0 4.8263583274810173e-03
GC_4_140 b_4 NI_4 NS_140 0 3.0318501898803020e-03
GC_4_141 b_4 NI_4 NS_141 0 -1.6834751390653042e-03
GC_4_142 b_4 NI_4 NS_142 0 -3.4545582649013110e-04
GC_4_143 b_4 NI_4 NS_143 0 2.8116069952871356e-03
GC_4_144 b_4 NI_4 NS_144 0 8.6550217557674006e-03
GC_4_145 b_4 NI_4 NS_145 0 1.2202808854114844e-04
GC_4_146 b_4 NI_4 NS_146 0 -3.3639326975896938e-04
GC_4_147 b_4 NI_4 NS_147 0 1.0878385190993068e-04
GC_4_148 b_4 NI_4 NS_148 0 -7.8652998236720679e-05
GC_4_149 b_4 NI_4 NS_149 0 1.9906503458430659e-04
GC_4_150 b_4 NI_4 NS_150 0 3.7445505666876142e-04
GC_4_151 b_4 NI_4 NS_151 0 6.6044112628740637e-05
GC_4_152 b_4 NI_4 NS_152 0 4.1799437572950229e-05
GC_4_153 b_4 NI_4 NS_153 0 1.4563418853401301e-04
GC_4_154 b_4 NI_4 NS_154 0 6.2844236386684570e-05
GC_4_155 b_4 NI_4 NS_155 0 7.4982829797475210e-06
GC_4_156 b_4 NI_4 NS_156 0 5.6070388432665010e-07
GC_4_157 b_4 NI_4 NS_157 0 -1.4002130988554551e-02
GC_4_158 b_4 NI_4 NS_158 0 2.7444923088956971e-03
GC_4_159 b_4 NI_4 NS_159 0 7.1392474814801141e-03
GC_4_160 b_4 NI_4 NS_160 0 -1.3419449388691801e-04
GC_4_161 b_4 NI_4 NS_161 0 1.6756396193948702e-04
GC_4_162 b_4 NI_4 NS_162 0 -7.5317381189753552e-04
GC_4_163 b_4 NI_4 NS_163 0 2.5402336760412954e-06
GC_4_164 b_4 NI_4 NS_164 0 -6.2513522732751942e-06
GC_4_165 b_4 NI_4 NS_165 0 -2.4008680968760359e-04
GC_4_166 b_4 NI_4 NS_166 0 -6.0285765774914559e-05
GC_4_167 b_4 NI_4 NS_167 0 -1.0174039044215600e-05
GC_4_168 b_4 NI_4 NS_168 0 -5.7934391422878525e-06
GC_4_169 b_4 NI_4 NS_169 0 -1.6403908828667873e-05
GC_4_170 b_4 NI_4 NS_170 0 -1.8008969676051627e-05
GC_4_171 b_4 NI_4 NS_171 0 2.9449499563651292e-04
GC_4_172 b_4 NI_4 NS_172 0 -2.2165914504604101e-04
GC_4_173 b_4 NI_4 NS_173 0 3.2259452728199260e-05
GC_4_174 b_4 NI_4 NS_174 0 -6.2443789527045059e-05
GC_4_175 b_4 NI_4 NS_175 0 -5.2199770842255313e-06
GC_4_176 b_4 NI_4 NS_176 0 -3.6033555226604241e-05
GC_4_177 b_4 NI_4 NS_177 0 2.3731797583398412e-02
GC_4_178 b_4 NI_4 NS_178 0 -6.8737816589678729e-04
GC_4_179 b_4 NI_4 NS_179 0 -2.3312772142038026e-02
GC_4_180 b_4 NI_4 NS_180 0 2.3683052860111646e-03
GC_4_181 b_4 NI_4 NS_181 0 6.9937006472242163e-03
GC_4_182 b_4 NI_4 NS_182 0 -7.8656554449943773e-03
GC_4_183 b_4 NI_4 NS_183 0 9.4988523529740774e-03
GC_4_184 b_4 NI_4 NS_184 0 1.1614966947256153e-03
GC_4_185 b_4 NI_4 NS_185 0 4.9102612108336608e-04
GC_4_186 b_4 NI_4 NS_186 0 -2.0256388299625728e-04
GC_4_187 b_4 NI_4 NS_187 0 -5.5465540601658692e-03
GC_4_188 b_4 NI_4 NS_188 0 -6.2304125614246701e-03
GC_4_189 b_4 NI_4 NS_189 0 -3.6182960680650655e-04
GC_4_190 b_4 NI_4 NS_190 0 1.2215214311369336e-04
GC_4_191 b_4 NI_4 NS_191 0 2.2689121808554057e-04
GC_4_192 b_4 NI_4 NS_192 0 1.1752221737145743e-04
GC_4_193 b_4 NI_4 NS_193 0 4.8381932649895095e-04
GC_4_194 b_4 NI_4 NS_194 0 4.4802084589286599e-04
GC_4_195 b_4 NI_4 NS_195 0 2.1910150579894648e-05
GC_4_196 b_4 NI_4 NS_196 0 5.0194384300517774e-05
GC_4_197 b_4 NI_4 NS_197 0 5.0621512277067739e-05
GC_4_198 b_4 NI_4 NS_198 0 3.8357660167284085e-05
GC_4_199 b_4 NI_4 NS_199 0 6.6445647171846630e-06
GC_4_200 b_4 NI_4 NS_200 0 -9.1141460657075972e-07
GC_4_201 b_4 NI_4 NS_201 0 -6.9426537039496963e-03
GC_4_202 b_4 NI_4 NS_202 0 6.8792585183355187e-03
GC_4_203 b_4 NI_4 NS_203 0 5.3326640337012666e-03
GC_4_204 b_4 NI_4 NS_204 0 -2.8012514994296624e-03
GC_4_205 b_4 NI_4 NS_205 0 -1.4489818698107602e-04
GC_4_206 b_4 NI_4 NS_206 0 -1.1619450505354011e-04
GC_4_207 b_4 NI_4 NS_207 0 -6.9631312121455955e-07
GC_4_208 b_4 NI_4 NS_208 0 -7.0569651269516791e-07
GC_4_209 b_4 NI_4 NS_209 0 -4.4808564670496941e-05
GC_4_210 b_4 NI_4 NS_210 0 1.3313462032052399e-05
GC_4_211 b_4 NI_4 NS_211 0 -5.6874425470323700e-07
GC_4_212 b_4 NI_4 NS_212 0 -4.7174075894096939e-07
GC_4_213 b_4 NI_4 NS_213 0 1.4841532144196451e-06
GC_4_214 b_4 NI_4 NS_214 0 -5.5173332224178546e-07
GC_4_215 b_4 NI_4 NS_215 0 -5.1394537498217223e-06
GC_4_216 b_4 NI_4 NS_216 0 -1.4136568661154218e-04
GC_4_217 b_4 NI_4 NS_217 0 1.7516337384489605e-05
GC_4_218 b_4 NI_4 NS_218 0 -4.7466701182914065e-06
GC_4_219 b_4 NI_4 NS_219 0 3.7683475675864236e-06
GC_4_220 b_4 NI_4 NS_220 0 -9.7165309732813391e-06
GC_4_221 b_4 NI_4 NS_221 0 -1.9416588524813930e-02
GC_4_222 b_4 NI_4 NS_222 0 -7.4615686067082757e-04
GC_4_223 b_4 NI_4 NS_223 0 1.6105158561742553e-02
GC_4_224 b_4 NI_4 NS_224 0 -3.7351583856860488e-03
GC_4_225 b_4 NI_4 NS_225 0 -1.1137222575644682e-02
GC_4_226 b_4 NI_4 NS_226 0 3.9185227344128143e-04
GC_4_227 b_4 NI_4 NS_227 0 9.2206345693903284e-03
GC_4_228 b_4 NI_4 NS_228 0 -6.8232812035304996e-04
GC_4_229 b_4 NI_4 NS_229 0 -2.0524747598409730e-03
GC_4_230 b_4 NI_4 NS_230 0 5.4581271167265147e-05
GC_4_231 b_4 NI_4 NS_231 0 1.6080614885647505e-03
GC_4_232 b_4 NI_4 NS_232 0 1.3979481233098575e-03
GC_4_233 b_4 NI_4 NS_233 0 1.4224350608191733e-04
GC_4_234 b_4 NI_4 NS_234 0 -1.5902372605878219e-04
GC_4_235 b_4 NI_4 NS_235 0 1.9868385411405966e-06
GC_4_236 b_4 NI_4 NS_236 0 -2.8882779192626527e-05
GC_4_237 b_4 NI_4 NS_237 0 1.0048275540900642e-05
GC_4_238 b_4 NI_4 NS_238 0 -1.9636976086269926e-04
GC_4_239 b_4 NI_4 NS_239 0 1.5656797142910445e-06
GC_4_240 b_4 NI_4 NS_240 0 -7.4218636671011277e-06
GC_4_241 b_4 NI_4 NS_241 0 -2.0270584794920965e-05
GC_4_242 b_4 NI_4 NS_242 0 -1.2449759347751652e-05
GC_4_243 b_4 NI_4 NS_243 0 -5.0121853052881416e-06
GC_4_244 b_4 NI_4 NS_244 0 -5.9828597427323917e-07
GC_4_245 b_4 NI_4 NS_245 0 6.5906380909841779e-03
GC_4_246 b_4 NI_4 NS_246 0 9.3893546746943168e-03
GC_4_247 b_4 NI_4 NS_247 0 -2.6109538946938785e-03
GC_4_248 b_4 NI_4 NS_248 0 -4.2191037536819433e-03
GC_4_249 b_4 NI_4 NS_249 0 -3.7390052448452009e-04
GC_4_250 b_4 NI_4 NS_250 0 6.5001597106449500e-05
GC_4_251 b_4 NI_4 NS_251 0 -8.1958710179318766e-07
GC_4_252 b_4 NI_4 NS_252 0 1.8565788423577497e-06
GC_4_253 b_4 NI_4 NS_253 0 -3.5962724070221247e-05
GC_4_254 b_4 NI_4 NS_254 0 1.8810658404861530e-04
GC_4_255 b_4 NI_4 NS_255 0 -4.9033932065428580e-06
GC_4_256 b_4 NI_4 NS_256 0 -2.9326992908922311e-06
GC_4_257 b_4 NI_4 NS_257 0 -9.3865262007795329e-06
GC_4_258 b_4 NI_4 NS_258 0 -2.0049992673941715e-05
GC_4_259 b_4 NI_4 NS_259 0 -3.9349276260887162e-04
GC_4_260 b_4 NI_4 NS_260 0 1.9876592317713399e-04
GC_4_261 b_4 NI_4 NS_261 0 -2.2250355242589852e-04
GC_4_262 b_4 NI_4 NS_262 0 -4.3800112377538442e-05
GC_4_263 b_4 NI_4 NS_263 0 -4.0917490127276284e-05
GC_4_264 b_4 NI_4 NS_264 0 2.1432972345356279e-06
GC_4_265 b_4 NI_4 NS_265 0 1.0839454610260396e-02
GC_4_266 b_4 NI_4 NS_266 0 -5.3461293774426967e-04
GC_4_267 b_4 NI_4 NS_267 0 -1.5028118722613899e-02
GC_4_268 b_4 NI_4 NS_268 0 5.6909028619659728e-03
GC_4_269 b_4 NI_4 NS_269 0 2.7206587581673539e-03
GC_4_270 b_4 NI_4 NS_270 0 -1.1950861421299913e-02
GC_4_271 b_4 NI_4 NS_271 0 8.2375395800577175e-03
GC_4_272 b_4 NI_4 NS_272 0 6.6318010624181220e-04
GC_4_273 b_4 NI_4 NS_273 0 -3.8060551260101345e-04
GC_4_274 b_4 NI_4 NS_274 0 -2.9349273032690308e-04
GC_4_275 b_4 NI_4 NS_275 0 -6.5977941874391577e-03
GC_4_276 b_4 NI_4 NS_276 0 -3.1244351094457524e-03
GC_4_277 b_4 NI_4 NS_277 0 -2.5715150274552111e-04
GC_4_278 b_4 NI_4 NS_278 0 9.7651956192471343e-05
GC_4_279 b_4 NI_4 NS_279 0 1.6653327221127052e-04
GC_4_280 b_4 NI_4 NS_280 0 4.3650736593703421e-05
GC_4_281 b_4 NI_4 NS_281 0 4.6034031160139394e-04
GC_4_282 b_4 NI_4 NS_282 0 1.4668897178766733e-04
GC_4_283 b_4 NI_4 NS_283 0 7.0401105503321327e-06
GC_4_284 b_4 NI_4 NS_284 0 1.2265873582733690e-05
GC_4_285 b_4 NI_4 NS_285 0 2.7506507008594179e-06
GC_4_286 b_4 NI_4 NS_286 0 -9.0069109490700809e-06
GC_4_287 b_4 NI_4 NS_287 0 2.6628682629336601e-06
GC_4_288 b_4 NI_4 NS_288 0 -7.2013677696733491e-07
GC_4_289 b_4 NI_4 NS_289 0 2.0783219740454872e-03
GC_4_290 b_4 NI_4 NS_290 0 3.8165485799007432e-03
GC_4_291 b_4 NI_4 NS_291 0 5.8530761632480768e-04
GC_4_292 b_4 NI_4 NS_292 0 -2.3275328653761139e-03
GC_4_293 b_4 NI_4 NS_293 0 2.3189892290291030e-05
GC_4_294 b_4 NI_4 NS_294 0 -7.8370425883142903e-06
GC_4_295 b_4 NI_4 NS_295 0 8.2022390712449246e-07
GC_4_296 b_4 NI_4 NS_296 0 3.7928308725363911e-07
GC_4_297 b_4 NI_4 NS_297 0 1.2016034993356524e-06
GC_4_298 b_4 NI_4 NS_298 0 -7.0171390258793673e-06
GC_4_299 b_4 NI_4 NS_299 0 -4.3696738136953422e-08
GC_4_300 b_4 NI_4 NS_300 0 -2.0550641233919350e-07
GC_4_301 b_4 NI_4 NS_301 0 -1.2705087366217487e-07
GC_4_302 b_4 NI_4 NS_302 0 -1.2096128330736259e-06
GC_4_303 b_4 NI_4 NS_303 0 -6.3494731446231761e-05
GC_4_304 b_4 NI_4 NS_304 0 1.9663962922331154e-05
GC_4_305 b_4 NI_4 NS_305 0 -1.4824933676542419e-05
GC_4_306 b_4 NI_4 NS_306 0 1.9191652089817378e-05
GC_4_307 b_4 NI_4 NS_307 0 -1.1583797215160577e-07
GC_4_308 b_4 NI_4 NS_308 0 3.8801410407635293e-07
GC_4_309 b_4 NI_4 NS_309 0 -1.4671280403440276e-02
GC_4_310 b_4 NI_4 NS_310 0 -3.9612008525046709e-05
GC_4_311 b_4 NI_4 NS_311 0 1.0735646632766140e-02
GC_4_312 b_4 NI_4 NS_312 0 -8.0555438698393707e-03
GC_4_313 b_4 NI_4 NS_313 0 -2.2205184117429001e-03
GC_4_314 b_4 NI_4 NS_314 0 7.4174858857322702e-03
GC_4_315 b_4 NI_4 NS_315 0 5.8634918567739332e-03
GC_4_316 b_4 NI_4 NS_316 0 3.2191624986009937e-05
GC_4_317 b_4 NI_4 NS_317 0 -1.0338921838662786e-03
GC_4_318 b_4 NI_4 NS_318 0 -4.5070260360612390e-06
GC_4_319 b_4 NI_4 NS_319 0 -1.3392216981334445e-03
GC_4_320 b_4 NI_4 NS_320 0 3.8124200847934331e-03
GC_4_321 b_4 NI_4 NS_321 0 1.1933038061480611e-04
GC_4_322 b_4 NI_4 NS_322 0 -1.4633060599072113e-04
GC_4_323 b_4 NI_4 NS_323 0 2.3851015762184980e-05
GC_4_324 b_4 NI_4 NS_324 0 -3.7598973388039749e-05
GC_4_325 b_4 NI_4 NS_325 0 6.4637648404689449e-05
GC_4_326 b_4 NI_4 NS_326 0 -6.4426350145257443e-05
GC_4_327 b_4 NI_4 NS_327 0 6.6625356829774453e-06
GC_4_328 b_4 NI_4 NS_328 0 -8.2070104991864210e-07
GC_4_329 b_4 NI_4 NS_329 0 4.4391318305286392e-06
GC_4_330 b_4 NI_4 NS_330 0 1.7479473788119744e-06
GC_4_331 b_4 NI_4 NS_331 0 -1.2042987845861928e-06
GC_4_332 b_4 NI_4 NS_332 0 2.0397137255373817e-07
GC_4_333 b_4 NI_4 NS_333 0 1.4559893821823591e-03
GC_4_334 b_4 NI_4 NS_334 0 3.7260726853085117e-03
GC_4_335 b_4 NI_4 NS_335 0 -5.2046170624824939e-04
GC_4_336 b_4 NI_4 NS_336 0 -1.6075189593970473e-03
GC_4_337 b_4 NI_4 NS_337 0 -2.2441269655422628e-04
GC_4_338 b_4 NI_4 NS_338 0 -5.5430691673994667e-05
GC_4_339 b_4 NI_4 NS_339 0 -1.4782810094042430e-07
GC_4_340 b_4 NI_4 NS_340 0 5.4686732273381296e-07
GC_4_341 b_4 NI_4 NS_341 0 -3.2622666533570437e-05
GC_4_342 b_4 NI_4 NS_342 0 8.0490468727831515e-05
GC_4_343 b_4 NI_4 NS_343 0 -3.0471003588226586e-06
GC_4_344 b_4 NI_4 NS_344 0 1.9903398821038182e-07
GC_4_345 b_4 NI_4 NS_345 0 -6.1210686508483214e-06
GC_4_346 b_4 NI_4 NS_346 0 -1.2557782516334140e-05
GC_4_347 b_4 NI_4 NS_347 0 -1.4722852605903800e-04
GC_4_348 b_4 NI_4 NS_348 0 7.5941640691606238e-05
GC_4_349 b_4 NI_4 NS_349 0 -1.0485339413303402e-04
GC_4_350 b_4 NI_4 NS_350 0 -2.9691151766658134e-05
GC_4_351 b_4 NI_4 NS_351 0 -1.4870896669027445e-05
GC_4_352 b_4 NI_4 NS_352 0 2.6716918566058923e-06
GC_4_353 b_4 NI_4 NS_353 0 -2.7665593770409792e-03
GC_4_354 b_4 NI_4 NS_354 0 2.3848676764825210e-05
GC_4_355 b_4 NI_4 NS_355 0 -1.8665108248698398e-04
GC_4_356 b_4 NI_4 NS_356 0 1.0958629566776500e-03
GC_4_357 b_4 NI_4 NS_357 0 -1.9192392406507817e-03
GC_4_358 b_4 NI_4 NS_358 0 -9.4797577629977977e-04
GC_4_359 b_4 NI_4 NS_359 0 -1.1950401653712082e-04
GC_4_360 b_4 NI_4 NS_360 0 -2.0095925560261524e-03
GC_4_361 b_4 NI_4 NS_361 0 4.0981862017100271e-04
GC_4_362 b_4 NI_4 NS_362 0 4.1401935073133732e-04
GC_4_363 b_4 NI_4 NS_363 0 1.1378844060146943e-03
GC_4_364 b_4 NI_4 NS_364 0 -1.4196426355699448e-03
GC_4_365 b_4 NI_4 NS_365 0 -4.2762759547660602e-05
GC_4_366 b_4 NI_4 NS_366 0 2.8376264063790656e-04
GC_4_367 b_4 NI_4 NS_367 0 2.8615083716652289e-04
GC_4_368 b_4 NI_4 NS_368 0 -5.5018807482906848e-05
GC_4_369 b_4 NI_4 NS_369 0 -4.1482032653985276e-04
GC_4_370 b_4 NI_4 NS_370 0 -8.4882455951384262e-06
GC_4_371 b_4 NI_4 NS_371 0 -3.0721451216125918e-05
GC_4_372 b_4 NI_4 NS_372 0 -5.5385538692438541e-06
GC_4_373 b_4 NI_4 NS_373 0 -4.5921017934874136e-05
GC_4_374 b_4 NI_4 NS_374 0 -3.8872736723838785e-05
GC_4_375 b_4 NI_4 NS_375 0 3.7805612151618814e-06
GC_4_376 b_4 NI_4 NS_376 0 2.6211297484510189e-06
GC_4_377 b_4 NI_4 NS_377 0 4.1537484152277329e-03
GC_4_378 b_4 NI_4 NS_378 0 2.5532816055456532e-03
GC_4_379 b_4 NI_4 NS_379 0 -2.4389329149135694e-03
GC_4_380 b_4 NI_4 NS_380 0 -2.4427823384908114e-03
GC_4_381 b_4 NI_4 NS_381 0 -7.8708910054863803e-05
GC_4_382 b_4 NI_4 NS_382 0 3.4115984232228678e-05
GC_4_383 b_4 NI_4 NS_383 0 -3.5747683842790258e-07
GC_4_384 b_4 NI_4 NS_384 0 4.2833342486027282e-07
GC_4_385 b_4 NI_4 NS_385 0 1.4781630109286049e-06
GC_4_386 b_4 NI_4 NS_386 0 1.8509713307829363e-05
GC_4_387 b_4 NI_4 NS_387 0 -1.0610956312302958e-06
GC_4_388 b_4 NI_4 NS_388 0 5.6424242368555149e-07
GC_4_389 b_4 NI_4 NS_389 0 2.4592730295414182e-06
GC_4_390 b_4 NI_4 NS_390 0 -5.5099077374957406e-07
GC_4_391 b_4 NI_4 NS_391 0 -7.7184383044966038e-05
GC_4_392 b_4 NI_4 NS_392 0 -4.2278010238347345e-05
GC_4_393 b_4 NI_4 NS_393 0 6.1210227458160148e-06
GC_4_394 b_4 NI_4 NS_394 0 -4.0132187195273423e-05
GC_4_395 b_4 NI_4 NS_395 0 -2.5192484268093125e-06
GC_4_396 b_4 NI_4 NS_396 0 3.9560717926345516e-06
GC_4_397 b_4 NI_4 NS_397 0 -8.5331280581767976e-03
GC_4_398 b_4 NI_4 NS_398 0 -1.0516661592721685e-05
GC_4_399 b_4 NI_4 NS_399 0 -7.3311588018831644e-04
GC_4_400 b_4 NI_4 NS_400 0 -9.8325201273698898e-04
GC_4_401 b_4 NI_4 NS_401 0 7.0731758696445919e-04
GC_4_402 b_4 NI_4 NS_402 0 -7.7756952199149949e-04
GC_4_403 b_4 NI_4 NS_403 0 2.9114187515443397e-04
GC_4_404 b_4 NI_4 NS_404 0 -1.3867303364479473e-03
GC_4_405 b_4 NI_4 NS_405 0 7.7151127018122061e-04
GC_4_406 b_4 NI_4 NS_406 0 5.1468907704995922e-04
GC_4_407 b_4 NI_4 NS_407 0 1.5440900687517475e-03
GC_4_408 b_4 NI_4 NS_408 0 -8.0100793033536458e-05
GC_4_409 b_4 NI_4 NS_409 0 -9.5371414495039534e-05
GC_4_410 b_4 NI_4 NS_410 0 -1.0126519495775053e-04
GC_4_411 b_4 NI_4 NS_411 0 4.9773257698547085e-05
GC_4_412 b_4 NI_4 NS_412 0 -3.2382803585580513e-05
GC_4_413 b_4 NI_4 NS_413 0 -2.3576028298914474e-04
GC_4_414 b_4 NI_4 NS_414 0 2.5376975570766001e-04
GC_4_415 b_4 NI_4 NS_415 0 -1.5147555002123626e-05
GC_4_416 b_4 NI_4 NS_416 0 2.0079655066202029e-05
GC_4_417 b_4 NI_4 NS_417 0 -1.0025987308452900e-05
GC_4_418 b_4 NI_4 NS_418 0 6.4482059525600185e-05
GC_4_419 b_4 NI_4 NS_419 0 -1.0112959989639134e-06
GC_4_420 b_4 NI_4 NS_420 0 8.2034676378534758e-07
GC_4_421 b_4 NI_4 NS_421 0 3.1247846538010890e-03
GC_4_422 b_4 NI_4 NS_422 0 -3.6680387661261137e-03
GC_4_423 b_4 NI_4 NS_423 0 -1.9512084999396462e-03
GC_4_424 b_4 NI_4 NS_424 0 2.0885538930697873e-03
GC_4_425 b_4 NI_4 NS_425 0 1.3427825866398830e-04
GC_4_426 b_4 NI_4 NS_426 0 4.2675392347385782e-05
GC_4_427 b_4 NI_4 NS_427 0 2.6833776912091325e-06
GC_4_428 b_4 NI_4 NS_428 0 -6.4199301991460374e-08
GC_4_429 b_4 NI_4 NS_429 0 4.3939776092155980e-06
GC_4_430 b_4 NI_4 NS_430 0 -6.9435384285643198e-05
GC_4_431 b_4 NI_4 NS_431 0 2.0288190571396079e-06
GC_4_432 b_4 NI_4 NS_432 0 7.7012501325876480e-06
GC_4_433 b_4 NI_4 NS_433 0 -1.2189802455312925e-05
GC_4_434 b_4 NI_4 NS_434 0 -2.3754595997814255e-05
GC_4_435 b_4 NI_4 NS_435 0 -1.7232529037283719e-06
GC_4_436 b_4 NI_4 NS_436 0 2.4439492784716774e-04
GC_4_437 b_4 NI_4 NS_437 0 -1.9289596321363648e-04
GC_4_438 b_4 NI_4 NS_438 0 1.1336651881727515e-05
GC_4_439 b_4 NI_4 NS_439 0 4.5914347452882046e-05
GC_4_440 b_4 NI_4 NS_440 0 5.6879649750137065e-05
GC_4_441 b_4 NI_4 NS_441 0 1.4921896653354481e-03
GC_4_442 b_4 NI_4 NS_442 0 -7.3701568479641133e-05
GC_4_443 b_4 NI_4 NS_443 0 -1.3799814826982574e-03
GC_4_444 b_4 NI_4 NS_444 0 2.3205548654006490e-03
GC_4_445 b_4 NI_4 NS_445 0 -2.0577647646854253e-03
GC_4_446 b_4 NI_4 NS_446 0 -2.5299259057886890e-03
GC_4_447 b_4 NI_4 NS_447 0 1.2822182235883157e-03
GC_4_448 b_4 NI_4 NS_448 0 -1.4481010212282360e-03
GC_4_449 b_4 NI_4 NS_449 0 7.2089642200827016e-05
GC_4_450 b_4 NI_4 NS_450 0 2.5265585995108621e-04
GC_4_451 b_4 NI_4 NS_451 0 -7.4074317217844834e-04
GC_4_452 b_4 NI_4 NS_452 0 -2.2708897649557103e-04
GC_4_453 b_4 NI_4 NS_453 0 -6.2349947589700414e-05
GC_4_454 b_4 NI_4 NS_454 0 1.9775896212615381e-04
GC_4_455 b_4 NI_4 NS_455 0 2.1171199336411257e-04
GC_4_456 b_4 NI_4 NS_456 0 -2.2826327195565751e-05
GC_4_457 b_4 NI_4 NS_457 0 -2.4338650775552554e-04
GC_4_458 b_4 NI_4 NS_458 0 2.3359700509903906e-05
GC_4_459 b_4 NI_4 NS_459 0 -2.2076438628925180e-05
GC_4_460 b_4 NI_4 NS_460 0 -9.7713130260413373e-07
GC_4_461 b_4 NI_4 NS_461 0 -2.6245403640477522e-05
GC_4_462 b_4 NI_4 NS_462 0 -2.0576384791722602e-05
GC_4_463 b_4 NI_4 NS_463 0 2.7482735030447768e-06
GC_4_464 b_4 NI_4 NS_464 0 1.5709595852618714e-06
GC_4_465 b_4 NI_4 NS_465 0 2.4459695952422367e-03
GC_4_466 b_4 NI_4 NS_466 0 9.3397809426008403e-04
GC_4_467 b_4 NI_4 NS_467 0 -1.2354338004379475e-03
GC_4_468 b_4 NI_4 NS_468 0 -1.3629753273072345e-03
GC_4_469 b_4 NI_4 NS_469 0 -4.6651084354816133e-05
GC_4_470 b_4 NI_4 NS_470 0 -4.6352399645721999e-05
GC_4_471 b_4 NI_4 NS_471 0 -4.4755862498990862e-07
GC_4_472 b_4 NI_4 NS_472 0 -3.9746316546544546e-07
GC_4_473 b_4 NI_4 NS_473 0 -2.9955710982370004e-06
GC_4_474 b_4 NI_4 NS_474 0 -1.0244671923138588e-06
GC_4_475 b_4 NI_4 NS_475 0 -4.4739827057647577e-08
GC_4_476 b_4 NI_4 NS_476 0 1.4190673748532317e-07
GC_4_477 b_4 NI_4 NS_477 0 -1.2784652833571045e-06
GC_4_478 b_4 NI_4 NS_478 0 -1.8597080253317637e-06
GC_4_479 b_4 NI_4 NS_479 0 -7.4426597111902309e-06
GC_4_480 b_4 NI_4 NS_480 0 -2.4977904503349706e-05
GC_4_481 b_4 NI_4 NS_481 0 3.7800083238733456e-06
GC_4_482 b_4 NI_4 NS_482 0 -1.3306520796267857e-05
GC_4_483 b_4 NI_4 NS_483 0 7.0591667677483760e-06
GC_4_484 b_4 NI_4 NS_484 0 7.2630885012123906e-07
GC_4_485 b_4 NI_4 NS_485 0 -7.7201038696780820e-03
GC_4_486 b_4 NI_4 NS_486 0 4.6036720890797981e-05
GC_4_487 b_4 NI_4 NS_487 0 3.5600840642812379e-04
GC_4_488 b_4 NI_4 NS_488 0 -2.5848364737931680e-03
GC_4_489 b_4 NI_4 NS_489 0 1.6943161427047184e-03
GC_4_490 b_4 NI_4 NS_490 0 7.6434861516943198e-04
GC_4_491 b_4 NI_4 NS_491 0 1.4074003772133810e-03
GC_4_492 b_4 NI_4 NS_492 0 -8.6544116223041540e-04
GC_4_493 b_4 NI_4 NS_493 0 -9.6882068984245777e-05
GC_4_494 b_4 NI_4 NS_494 0 1.2011801859447194e-04
GC_4_495 b_4 NI_4 NS_495 0 1.1859183568404849e-03
GC_4_496 b_4 NI_4 NS_496 0 1.5431610557081830e-03
GC_4_497 b_4 NI_4 NS_497 0 -4.1974202777350739e-05
GC_4_498 b_4 NI_4 NS_498 0 -9.4653538199357574e-05
GC_4_499 b_4 NI_4 NS_499 0 3.5520558136243967e-05
GC_4_500 b_4 NI_4 NS_500 0 -3.7570138263622239e-05
GC_4_501 b_4 NI_4 NS_501 0 -9.8097146162925627e-05
GC_4_502 b_4 NI_4 NS_502 0 1.3440293197902183e-04
GC_4_503 b_4 NI_4 NS_503 0 -6.8715956153658541e-06
GC_4_504 b_4 NI_4 NS_504 0 7.5586943958995620e-06
GC_4_505 b_4 NI_4 NS_505 0 -4.8165201091137391e-06
GC_4_506 b_4 NI_4 NS_506 0 2.9354694888458654e-05
GC_4_507 b_4 NI_4 NS_507 0 -6.8688023788085871e-07
GC_4_508 b_4 NI_4 NS_508 0 8.7973206880575776e-07
GC_4_509 b_4 NI_4 NS_509 0 1.4015214406351770e-03
GC_4_510 b_4 NI_4 NS_510 0 -1.1639793122911642e-04
GC_4_511 b_4 NI_4 NS_511 0 -8.8610296437829656e-04
GC_4_512 b_4 NI_4 NS_512 0 2.7449358098695565e-04
GC_4_513 b_4 NI_4 NS_513 0 -5.3103544993882153e-05
GC_4_514 b_4 NI_4 NS_514 0 -2.1662731189988687e-05
GC_4_515 b_4 NI_4 NS_515 0 9.2333175601571110e-07
GC_4_516 b_4 NI_4 NS_516 0 -1.5294455979151858e-07
GC_4_517 b_4 NI_4 NS_517 0 -1.6339952787396022e-05
GC_4_518 b_4 NI_4 NS_518 0 -1.7237379828855198e-07
GC_4_519 b_4 NI_4 NS_519 0 -1.4771839486870639e-08
GC_4_520 b_4 NI_4 NS_520 0 4.6930604172613299e-06
GC_4_521 b_4 NI_4 NS_521 0 -6.8323688717622918e-06
GC_4_522 b_4 NI_4 NS_522 0 -1.3826781834092318e-05
GC_4_523 b_4 NI_4 NS_523 0 -3.6423461675170512e-05
GC_4_524 b_4 NI_4 NS_524 0 9.3394881876908461e-05
GC_4_525 b_4 NI_4 NS_525 0 -1.0377461268377010e-04
GC_4_526 b_4 NI_4 NS_526 0 -5.4861100466026217e-06
GC_4_527 b_4 NI_4 NS_527 0 1.7053330716744281e-05
GC_4_528 b_4 NI_4 NS_528 0 2.5300965507758096e-05
GD_4_1 b_4 NI_4 NA_1 0 -2.5623308108916982e-03
GD_4_2 b_4 NI_4 NA_2 0 -1.5147017228053098e-03
GD_4_3 b_4 NI_4 NA_3 0 -1.7485402243861560e-02
GD_4_4 b_4 NI_4 NA_4 0 1.3027808524336942e-01
GD_4_5 b_4 NI_4 NA_5 0 -1.2057227942234518e-02
GD_4_6 b_4 NI_4 NA_6 0 8.8946856249420044e-04
GD_4_7 b_4 NI_4 NA_7 0 -2.6662571492012538e-03
GD_4_8 b_4 NI_4 NA_8 0 8.7422291377659965e-04
GD_4_9 b_4 NI_4 NA_9 0 2.1561735887638050e-03
GD_4_10 b_4 NI_4 NA_10 0 5.7861508507420492e-03
GD_4_11 b_4 NI_4 NA_11 0 5.7763564578198047e-04
GD_4_12 b_4 NI_4 NA_12 0 3.1074003222985617e-03
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 1.4888401712574677e-02
GC_5_2 b_5 NI_5 NS_2 0 -9.3518480534754689e-06
GC_5_3 b_5 NI_5 NS_3 0 1.2024151653626969e-02
GC_5_4 b_5 NI_5 NS_4 0 -5.2254723615874970e-03
GC_5_5 b_5 NI_5 NS_5 0 -2.3071146560534749e-03
GC_5_6 b_5 NI_5 NS_6 0 5.8586359722770905e-03
GC_5_7 b_5 NI_5 NS_7 0 1.2364954931264653e-02
GC_5_8 b_5 NI_5 NS_8 0 9.2062676968267913e-03
GC_5_9 b_5 NI_5 NS_9 0 -2.2188545995761510e-03
GC_5_10 b_5 NI_5 NS_10 0 -3.0825900370844293e-03
GC_5_11 b_5 NI_5 NS_11 0 -1.0102730895459098e-02
GC_5_12 b_5 NI_5 NS_12 0 9.6134683530379478e-03
GC_5_13 b_5 NI_5 NS_13 0 5.4911431511253954e-04
GC_5_14 b_5 NI_5 NS_14 0 4.2797708634814241e-04
GC_5_15 b_5 NI_5 NS_15 0 5.5714477042071903e-05
GC_5_16 b_5 NI_5 NS_16 0 2.1799559001127190e-04
GC_5_17 b_5 NI_5 NS_17 0 1.3139424947679968e-03
GC_5_18 b_5 NI_5 NS_18 0 2.3427081311815391e-04
GC_5_19 b_5 NI_5 NS_19 0 1.5519461050894200e-04
GC_5_20 b_5 NI_5 NS_20 0 1.4245051926240463e-04
GC_5_21 b_5 NI_5 NS_21 0 2.3535465258338402e-04
GC_5_22 b_5 NI_5 NS_22 0 5.2771923484806170e-05
GC_5_23 b_5 NI_5 NS_23 0 -9.1466667977531992e-06
GC_5_24 b_5 NI_5 NS_24 0 3.9142335685262442e-06
GC_5_25 b_5 NI_5 NS_25 0 -2.4379490423040096e-02
GC_5_26 b_5 NI_5 NS_26 0 -9.8093355717295645e-04
GC_5_27 b_5 NI_5 NS_27 0 1.5256180092879542e-02
GC_5_28 b_5 NI_5 NS_28 0 3.8108865834726906e-03
GC_5_29 b_5 NI_5 NS_29 0 -3.4039717499623196e-04
GC_5_30 b_5 NI_5 NS_30 0 -4.8567332572604683e-04
GC_5_31 b_5 NI_5 NS_31 0 9.1459998020267913e-07
GC_5_32 b_5 NI_5 NS_32 0 4.5967216745026346e-07
GC_5_33 b_5 NI_5 NS_33 0 9.9142384636810609e-05
GC_5_34 b_5 NI_5 NS_34 0 -5.3583112263115069e-05
GC_5_35 b_5 NI_5 NS_35 0 2.1456157635928747e-06
GC_5_36 b_5 NI_5 NS_36 0 3.0865102073509870e-07
GC_5_37 b_5 NI_5 NS_37 0 -1.9245036014831232e-06
GC_5_38 b_5 NI_5 NS_38 0 -1.1735224944863787e-06
GC_5_39 b_5 NI_5 NS_39 0 -6.5682388735307777e-05
GC_5_40 b_5 NI_5 NS_40 0 2.1932692681551617e-04
GC_5_41 b_5 NI_5 NS_41 0 2.0903108903751031e-05
GC_5_42 b_5 NI_5 NS_42 0 -7.0297658116498751e-05
GC_5_43 b_5 NI_5 NS_43 0 -1.1994220959439512e-05
GC_5_44 b_5 NI_5 NS_44 0 -1.4131663488031825e-06
GC_5_45 b_5 NI_5 NS_45 0 1.3168575740214416e-02
GC_5_46 b_5 NI_5 NS_46 0 -5.8033216824185385e-04
GC_5_47 b_5 NI_5 NS_47 0 -1.5406741695628126e-02
GC_5_48 b_5 NI_5 NS_48 0 6.1074988667710450e-03
GC_5_49 b_5 NI_5 NS_49 0 2.5861106581148191e-03
GC_5_50 b_5 NI_5 NS_50 0 -1.2319324840469657e-02
GC_5_51 b_5 NI_5 NS_51 0 8.7210186906431092e-03
GC_5_52 b_5 NI_5 NS_52 0 9.0037929058741305e-04
GC_5_53 b_5 NI_5 NS_53 0 -4.9795602169660168e-04
GC_5_54 b_5 NI_5 NS_54 0 -5.2255038624303993e-04
GC_5_55 b_5 NI_5 NS_55 0 -7.2163140669954575e-03
GC_5_56 b_5 NI_5 NS_56 0 -2.7242077050791706e-03
GC_5_57 b_5 NI_5 NS_57 0 -2.6607579565203227e-04
GC_5_58 b_5 NI_5 NS_58 0 9.1619082533784431e-05
GC_5_59 b_5 NI_5 NS_59 0 1.4115681002774819e-04
GC_5_60 b_5 NI_5 NS_60 0 2.8471219323628858e-05
GC_5_61 b_5 NI_5 NS_61 0 5.8069371680756260e-04
GC_5_62 b_5 NI_5 NS_62 0 7.7827289760374371e-05
GC_5_63 b_5 NI_5 NS_63 0 1.7744593264287836e-05
GC_5_64 b_5 NI_5 NS_64 0 1.3644662326178211e-06
GC_5_65 b_5 NI_5 NS_65 0 2.7646981342877195e-05
GC_5_66 b_5 NI_5 NS_66 0 -2.9931298068326611e-05
GC_5_67 b_5 NI_5 NS_67 0 6.2612320659185344e-06
GC_5_68 b_5 NI_5 NS_68 0 -2.9297897086094896e-06
GC_5_69 b_5 NI_5 NS_69 0 9.2196759660724981e-04
GC_5_70 b_5 NI_5 NS_70 0 4.6350572839900994e-03
GC_5_71 b_5 NI_5 NS_71 0 1.2090088203982870e-03
GC_5_72 b_5 NI_5 NS_72 0 -2.7465139938112333e-03
GC_5_73 b_5 NI_5 NS_73 0 -1.2960474857446253e-05
GC_5_74 b_5 NI_5 NS_74 0 -5.3539126923437902e-05
GC_5_75 b_5 NI_5 NS_75 0 -5.1457033835131786e-09
GC_5_76 b_5 NI_5 NS_76 0 1.6912619308356918e-07
GC_5_77 b_5 NI_5 NS_77 0 -1.2102239998992327e-05
GC_5_78 b_5 NI_5 NS_78 0 5.5876271647961732e-06
GC_5_79 b_5 NI_5 NS_79 0 2.5318691454580117e-07
GC_5_80 b_5 NI_5 NS_80 0 -1.4145354745589652e-07
GC_5_81 b_5 NI_5 NS_81 0 2.9982820118976946e-06
GC_5_82 b_5 NI_5 NS_82 0 -1.3346114598210794e-07
GC_5_83 b_5 NI_5 NS_83 0 -4.1929143609115300e-05
GC_5_84 b_5 NI_5 NS_84 0 -4.6870406181453323e-05
GC_5_85 b_5 NI_5 NS_85 0 2.8638373402039862e-06
GC_5_86 b_5 NI_5 NS_86 0 -1.0549144924066329e-06
GC_5_87 b_5 NI_5 NS_87 0 1.7502705895507350e-06
GC_5_88 b_5 NI_5 NS_88 0 -4.5742259217823701e-06
GC_5_89 b_5 NI_5 NS_89 0 1.4223626652689683e-02
GC_5_90 b_5 NI_5 NS_90 0 -3.0973857615682385e-04
GC_5_91 b_5 NI_5 NS_91 0 1.5676679373708282e-02
GC_5_92 b_5 NI_5 NS_92 0 -1.5966002381428369e-03
GC_5_93 b_5 NI_5 NS_93 0 -5.5294404200685468e-03
GC_5_94 b_5 NI_5 NS_94 0 -3.2743694507681356e-03
GC_5_95 b_5 NI_5 NS_95 0 1.7870505406363719e-02
GC_5_96 b_5 NI_5 NS_96 0 1.2336324544690533e-02
GC_5_97 b_5 NI_5 NS_97 0 -2.5331500892905720e-03
GC_5_98 b_5 NI_5 NS_98 0 -4.1354013608286069e-03
GC_5_99 b_5 NI_5 NS_99 0 -5.3452539779942267e-03
GC_5_100 b_5 NI_5 NS_100 0 1.2018818856238282e-02
GC_5_101 b_5 NI_5 NS_101 0 7.1888857076226806e-04
GC_5_102 b_5 NI_5 NS_102 0 5.6256742630847391e-04
GC_5_103 b_5 NI_5 NS_103 0 9.4834554646488914e-05
GC_5_104 b_5 NI_5 NS_104 0 3.6208466296423135e-04
GC_5_105 b_5 NI_5 NS_105 0 1.4786223860525172e-03
GC_5_106 b_5 NI_5 NS_106 0 1.8745457771889059e-04
GC_5_107 b_5 NI_5 NS_107 0 2.1471686980832866e-04
GC_5_108 b_5 NI_5 NS_108 0 2.2927059446919496e-04
GC_5_109 b_5 NI_5 NS_109 0 2.9202131855307303e-04
GC_5_110 b_5 NI_5 NS_110 0 1.0185886520753988e-04
GC_5_111 b_5 NI_5 NS_111 0 -1.3096785416743770e-05
GC_5_112 b_5 NI_5 NS_112 0 7.8082902261855851e-06
GC_5_113 b_5 NI_5 NS_113 0 -3.3455247963899842e-02
GC_5_114 b_5 NI_5 NS_114 0 2.6928649732189149e-03
GC_5_115 b_5 NI_5 NS_115 0 2.1120487428677236e-02
GC_5_116 b_5 NI_5 NS_116 0 4.4461598615994583e-03
GC_5_117 b_5 NI_5 NS_117 0 -6.7251109925018997e-04
GC_5_118 b_5 NI_5 NS_118 0 -3.3691729564912140e-04
GC_5_119 b_5 NI_5 NS_119 0 1.4897808941446102e-06
GC_5_120 b_5 NI_5 NS_120 0 3.1634383184063627e-06
GC_5_121 b_5 NI_5 NS_121 0 2.1952963034634006e-04
GC_5_122 b_5 NI_5 NS_122 0 -3.6443569460360740e-05
GC_5_123 b_5 NI_5 NS_123 0 5.4073168165224134e-06
GC_5_124 b_5 NI_5 NS_124 0 1.0081925557522484e-06
GC_5_125 b_5 NI_5 NS_125 0 -1.0329908378039173e-06
GC_5_126 b_5 NI_5 NS_126 0 -6.2435838122072759e-07
GC_5_127 b_5 NI_5 NS_127 0 -1.8707043302679038e-04
GC_5_128 b_5 NI_5 NS_128 0 3.7590705331149419e-04
GC_5_129 b_5 NI_5 NS_129 0 -1.2789170263135766e-05
GC_5_130 b_5 NI_5 NS_130 0 -8.9008967628663013e-05
GC_5_131 b_5 NI_5 NS_131 0 -2.0760710127965729e-05
GC_5_132 b_5 NI_5 NS_132 0 4.9325651137451958e-06
GC_5_133 b_5 NI_5 NS_133 0 2.3731797583464789e-02
GC_5_134 b_5 NI_5 NS_134 0 -6.8737816589820489e-04
GC_5_135 b_5 NI_5 NS_135 0 -2.3312772142037089e-02
GC_5_136 b_5 NI_5 NS_136 0 2.3683052860188989e-03
GC_5_137 b_5 NI_5 NS_137 0 6.9937006472160172e-03
GC_5_138 b_5 NI_5 NS_138 0 -7.8656554449908767e-03
GC_5_139 b_5 NI_5 NS_139 0 9.4988523529708439e-03
GC_5_140 b_5 NI_5 NS_140 0 1.1614966947277676e-03
GC_5_141 b_5 NI_5 NS_141 0 4.9102612107924850e-04
GC_5_142 b_5 NI_5 NS_142 0 -2.0256388299569623e-04
GC_5_143 b_5 NI_5 NS_143 0 -5.5465540601703318e-03
GC_5_144 b_5 NI_5 NS_144 0 -6.2304125614212136e-03
GC_5_145 b_5 NI_5 NS_145 0 -3.6182960680632430e-04
GC_5_146 b_5 NI_5 NS_146 0 1.2215214311354626e-04
GC_5_147 b_5 NI_5 NS_147 0 2.2689121808559866e-04
GC_5_148 b_5 NI_5 NS_148 0 1.1752221737158104e-04
GC_5_149 b_5 NI_5 NS_149 0 4.8381932649853933e-04
GC_5_150 b_5 NI_5 NS_150 0 4.4802084589302867e-04
GC_5_151 b_5 NI_5 NS_151 0 2.1910150579846578e-05
GC_5_152 b_5 NI_5 NS_152 0 5.0194384300520010e-05
GC_5_153 b_5 NI_5 NS_153 0 5.0621512276930682e-05
GC_5_154 b_5 NI_5 NS_154 0 3.8357660167188370e-05
GC_5_155 b_5 NI_5 NS_155 0 6.6445647171609393e-06
GC_5_156 b_5 NI_5 NS_156 0 -9.1141460660290441e-07
GC_5_157 b_5 NI_5 NS_157 0 -6.9426537039580351e-03
GC_5_158 b_5 NI_5 NS_158 0 6.8792585183445939e-03
GC_5_159 b_5 NI_5 NS_159 0 5.3326640337055583e-03
GC_5_160 b_5 NI_5 NS_160 0 -2.8012514994348544e-03
GC_5_161 b_5 NI_5 NS_161 0 -1.4489818698143174e-04
GC_5_162 b_5 NI_5 NS_162 0 -1.1619450505402069e-04
GC_5_163 b_5 NI_5 NS_163 0 -6.9631312121556148e-07
GC_5_164 b_5 NI_5 NS_164 0 -7.0569651269883619e-07
GC_5_165 b_5 NI_5 NS_165 0 -4.4808564670670243e-05
GC_5_166 b_5 NI_5 NS_166 0 1.3313462032084276e-05
GC_5_167 b_5 NI_5 NS_167 0 -5.6874425470715432e-07
GC_5_168 b_5 NI_5 NS_168 0 -4.7174075893895154e-07
GC_5_169 b_5 NI_5 NS_169 0 1.4841532144087237e-06
GC_5_170 b_5 NI_5 NS_170 0 -5.5173332224228256e-07
GC_5_171 b_5 NI_5 NS_171 0 -5.1394537496665890e-06
GC_5_172 b_5 NI_5 NS_172 0 -1.4136568661208556e-04
GC_5_173 b_5 NI_5 NS_173 0 1.7516337384570988e-05
GC_5_174 b_5 NI_5 NS_174 0 -4.7466701183845826e-06
GC_5_175 b_5 NI_5 NS_175 0 3.7683475675861225e-06
GC_5_176 b_5 NI_5 NS_176 0 -9.7165309733130402e-06
GC_5_177 b_5 NI_5 NS_177 0 -1.0880179654136939e-02
GC_5_178 b_5 NI_5 NS_178 0 1.3580154587373534e-02
GC_5_179 b_5 NI_5 NS_179 0 1.2747777248338671e-02
GC_5_180 b_5 NI_5 NS_180 0 2.7463409626272439e-03
GC_5_181 b_5 NI_5 NS_181 0 1.8113032263587722e-02
GC_5_182 b_5 NI_5 NS_182 0 -3.4358758593928539e-04
GC_5_183 b_5 NI_5 NS_183 0 1.4295838267246681e-02
GC_5_184 b_5 NI_5 NS_184 0 1.1814767056003813e-02
GC_5_185 b_5 NI_5 NS_185 0 2.4711061988890001e-03
GC_5_186 b_5 NI_5 NS_186 0 2.9826159184973633e-03
GC_5_187 b_5 NI_5 NS_187 0 -1.7464923585892511e-03
GC_5_188 b_5 NI_5 NS_188 0 1.9013021957185443e-02
GC_5_189 b_5 NI_5 NS_189 0 6.7285423641640345e-04
GC_5_190 b_5 NI_5 NS_190 0 4.2824758733213148e-04
GC_5_191 b_5 NI_5 NS_191 0 2.7753530697632202e-05
GC_5_192 b_5 NI_5 NS_192 0 3.3278239306725968e-04
GC_5_193 b_5 NI_5 NS_193 0 1.7947123443067092e-03
GC_5_194 b_5 NI_5 NS_194 0 -5.4422633364382283e-04
GC_5_195 b_5 NI_5 NS_195 0 1.8352781875680363e-04
GC_5_196 b_5 NI_5 NS_196 0 1.6760157809759423e-04
GC_5_197 b_5 NI_5 NS_197 0 1.4472489321885404e-04
GC_5_198 b_5 NI_5 NS_198 0 1.7785890342945661e-05
GC_5_199 b_5 NI_5 NS_199 0 -2.0121415438617585e-05
GC_5_200 b_5 NI_5 NS_200 0 6.1134130507823420e-06
GC_5_201 b_5 NI_5 NS_201 0 -1.8591319726062382e-02
GC_5_202 b_5 NI_5 NS_202 0 1.8863525282902232e-03
GC_5_203 b_5 NI_5 NS_203 0 1.4009035267740574e-02
GC_5_204 b_5 NI_5 NS_204 0 2.7045327481041168e-03
GC_5_205 b_5 NI_5 NS_205 0 -6.8394798957541311e-04
GC_5_206 b_5 NI_5 NS_206 0 1.4657695860589411e-04
GC_5_207 b_5 NI_5 NS_207 0 2.6301191894411378e-06
GC_5_208 b_5 NI_5 NS_208 0 5.9359233725478811e-06
GC_5_209 b_5 NI_5 NS_209 0 3.2973425316314207e-04
GC_5_210 b_5 NI_5 NS_210 0 -1.5192380963136210e-05
GC_5_211 b_5 NI_5 NS_211 0 7.2232170478647811e-06
GC_5_212 b_5 NI_5 NS_212 0 2.0843205540915074e-06
GC_5_213 b_5 NI_5 NS_213 0 4.9824310881155480e-06
GC_5_214 b_5 NI_5 NS_214 0 2.5733825275527848e-06
GC_5_215 b_5 NI_5 NS_215 0 -4.5089820396847387e-04
GC_5_216 b_5 NI_5 NS_216 0 6.2702607803068904e-04
GC_5_217 b_5 NI_5 NS_217 0 -9.1305403650220109e-05
GC_5_218 b_5 NI_5 NS_218 0 -6.1418462292856991e-05
GC_5_219 b_5 NI_5 NS_219 0 -3.2474635023102361e-05
GC_5_220 b_5 NI_5 NS_220 0 2.1571867245994379e-05
GC_5_221 b_5 NI_5 NS_221 0 4.7547290818100774e-02
GC_5_222 b_5 NI_5 NS_222 0 1.6148575703483919e-02
GC_5_223 b_5 NI_5 NS_223 0 -2.8784676938770088e-02
GC_5_224 b_5 NI_5 NS_224 0 1.3904415597772188e-03
GC_5_225 b_5 NI_5 NS_225 0 -2.8618554001337882e-02
GC_5_226 b_5 NI_5 NS_226 0 -9.2802340156129971e-03
GC_5_227 b_5 NI_5 NS_227 0 9.6204946360265893e-03
GC_5_228 b_5 NI_5 NS_228 0 2.5770766881007341e-03
GC_5_229 b_5 NI_5 NS_229 0 -2.6261267865950403e-03
GC_5_230 b_5 NI_5 NS_230 0 9.3809662928540780e-05
GC_5_231 b_5 NI_5 NS_231 0 1.3380579702185627e-03
GC_5_232 b_5 NI_5 NS_232 0 -2.9466270797792169e-03
GC_5_233 b_5 NI_5 NS_233 0 -5.0555633589759706e-04
GC_5_234 b_5 NI_5 NS_234 0 1.1060588345052210e-04
GC_5_235 b_5 NI_5 NS_235 0 1.3619834283357224e-04
GC_5_236 b_5 NI_5 NS_236 0 4.0475384268751084e-05
GC_5_237 b_5 NI_5 NS_237 0 6.9117352146411614e-04
GC_5_238 b_5 NI_5 NS_238 0 -3.7665960616920706e-04
GC_5_239 b_5 NI_5 NS_239 0 -3.3764247233581772e-06
GC_5_240 b_5 NI_5 NS_240 0 1.0564266413811194e-05
GC_5_241 b_5 NI_5 NS_241 0 -9.0504273427051643e-06
GC_5_242 b_5 NI_5 NS_242 0 -1.2975905285806852e-05
GC_5_243 b_5 NI_5 NS_243 0 7.7709107487676668e-06
GC_5_244 b_5 NI_5 NS_244 0 8.7534026358240403e-07
GC_5_245 b_5 NI_5 NS_245 0 -1.5794618792187799e-03
GC_5_246 b_5 NI_5 NS_246 0 -3.8550470293181416e-03
GC_5_247 b_5 NI_5 NS_247 0 1.4547170328684373e-03
GC_5_248 b_5 NI_5 NS_248 0 5.2850931172475336e-04
GC_5_249 b_5 NI_5 NS_249 0 1.1220256898866285e-04
GC_5_250 b_5 NI_5 NS_250 0 -5.3923010191859420e-05
GC_5_251 b_5 NI_5 NS_251 0 1.3133507411609197e-06
GC_5_252 b_5 NI_5 NS_252 0 1.1915904730938004e-07
GC_5_253 b_5 NI_5 NS_253 0 -8.9935687520356617e-06
GC_5_254 b_5 NI_5 NS_254 0 -5.5497877731438435e-05
GC_5_255 b_5 NI_5 NS_255 0 6.9625767762929805e-07
GC_5_256 b_5 NI_5 NS_256 0 -1.8260244037075153e-06
GC_5_257 b_5 NI_5 NS_257 0 6.6504835290214502e-06
GC_5_258 b_5 NI_5 NS_258 0 -2.9212251284478955e-06
GC_5_259 b_5 NI_5 NS_259 0 5.4536072809828310e-05
GC_5_260 b_5 NI_5 NS_260 0 1.3167163820865599e-04
GC_5_261 b_5 NI_5 NS_261 0 1.9319945599628082e-05
GC_5_262 b_5 NI_5 NS_262 0 2.7113163285924467e-05
GC_5_263 b_5 NI_5 NS_263 0 1.0086511961617392e-05
GC_5_264 b_5 NI_5 NS_264 0 -1.5525391085485546e-06
GC_5_265 b_5 NI_5 NS_265 0 5.6120539298638262e-03
GC_5_266 b_5 NI_5 NS_266 0 -5.1913700960193895e-04
GC_5_267 b_5 NI_5 NS_267 0 1.1152832382888320e-02
GC_5_268 b_5 NI_5 NS_268 0 3.3286876797490837e-03
GC_5_269 b_5 NI_5 NS_269 0 -8.8802452741710593e-03
GC_5_270 b_5 NI_5 NS_270 0 -8.9204509768656525e-03
GC_5_271 b_5 NI_5 NS_271 0 1.1593344810250782e-02
GC_5_272 b_5 NI_5 NS_272 0 6.5240857665460937e-03
GC_5_273 b_5 NI_5 NS_273 0 -2.6330008472453840e-03
GC_5_274 b_5 NI_5 NS_274 0 -1.1657371882252392e-03
GC_5_275 b_5 NI_5 NS_275 0 2.8837397276935714e-03
GC_5_276 b_5 NI_5 NS_276 0 2.9234219270483884e-03
GC_5_277 b_5 NI_5 NS_277 0 5.7649672114961324e-04
GC_5_278 b_5 NI_5 NS_278 0 3.7833629962891343e-04
GC_5_279 b_5 NI_5 NS_279 0 1.2742624069944652e-04
GC_5_280 b_5 NI_5 NS_280 0 3.4203965796307311e-04
GC_5_281 b_5 NI_5 NS_281 0 7.7293193933663130e-04
GC_5_282 b_5 NI_5 NS_282 0 -6.4517690610389655e-05
GC_5_283 b_5 NI_5 NS_283 0 1.8599392982159943e-04
GC_5_284 b_5 NI_5 NS_284 0 1.6984865408427730e-04
GC_5_285 b_5 NI_5 NS_285 0 8.7402876868516898e-05
GC_5_286 b_5 NI_5 NS_286 0 3.6761398473695930e-05
GC_5_287 b_5 NI_5 NS_287 0 -8.5234104693584552e-06
GC_5_288 b_5 NI_5 NS_288 0 1.9060167792756390e-06
GC_5_289 b_5 NI_5 NS_289 0 -1.7137304426203596e-02
GC_5_290 b_5 NI_5 NS_290 0 9.6737302919309796e-03
GC_5_291 b_5 NI_5 NS_291 0 1.2689828848668511e-02
GC_5_292 b_5 NI_5 NS_292 0 -1.1129100038079047e-03
GC_5_293 b_5 NI_5 NS_293 0 -4.3328715421870776e-04
GC_5_294 b_5 NI_5 NS_294 0 -2.1162014479221880e-05
GC_5_295 b_5 NI_5 NS_295 0 1.2982407320329742e-06
GC_5_296 b_5 NI_5 NS_296 0 2.8962947404319530e-06
GC_5_297 b_5 NI_5 NS_297 0 1.8336278332947950e-04
GC_5_298 b_5 NI_5 NS_298 0 -2.1362352079785455e-05
GC_5_299 b_5 NI_5 NS_299 0 4.3755483143861848e-06
GC_5_300 b_5 NI_5 NS_300 0 1.0716257489351799e-06
GC_5_301 b_5 NI_5 NS_301 0 -4.9215837127030853e-09
GC_5_302 b_5 NI_5 NS_302 0 -8.4765074293709927e-08
GC_5_303 b_5 NI_5 NS_303 0 -1.8712977959623792e-04
GC_5_304 b_5 NI_5 NS_304 0 3.0580470557332412e-04
GC_5_305 b_5 NI_5 NS_305 0 -5.6725967090318061e-05
GC_5_306 b_5 NI_5 NS_306 0 -4.3286565094221368e-05
GC_5_307 b_5 NI_5 NS_307 0 -1.9141010544136533e-05
GC_5_308 b_5 NI_5 NS_308 0 5.9946355818492034e-06
GC_5_309 b_5 NI_5 NS_309 0 5.3117525550891919e-03
GC_5_310 b_5 NI_5 NS_310 0 -3.4365694724857273e-04
GC_5_311 b_5 NI_5 NS_311 0 -1.9971882412578891e-02
GC_5_312 b_5 NI_5 NS_312 0 -3.0245411875664901e-03
GC_5_313 b_5 NI_5 NS_313 0 9.7982095617133776e-03
GC_5_314 b_5 NI_5 NS_314 0 -2.9828054633968628e-03
GC_5_315 b_5 NI_5 NS_315 0 5.6535050806052149e-03
GC_5_316 b_5 NI_5 NS_316 0 5.5762876877636907e-04
GC_5_317 b_5 NI_5 NS_317 0 2.2363204799443750e-03
GC_5_318 b_5 NI_5 NS_318 0 -3.9035827238457501e-04
GC_5_319 b_5 NI_5 NS_319 0 -2.0827490630965018e-04
GC_5_320 b_5 NI_5 NS_320 0 -8.9815090995554406e-03
GC_5_321 b_5 NI_5 NS_321 0 -2.5813605053039927e-04
GC_5_322 b_5 NI_5 NS_322 0 1.0030187056167708e-04
GC_5_323 b_5 NI_5 NS_323 0 2.2578959543764348e-04
GC_5_324 b_5 NI_5 NS_324 0 5.2177047703626570e-05
GC_5_325 b_5 NI_5 NS_325 0 4.3582627497245615e-04
GC_5_326 b_5 NI_5 NS_326 0 4.4577164807046928e-04
GC_5_327 b_5 NI_5 NS_327 0 2.2967443813777994e-05
GC_5_328 b_5 NI_5 NS_328 0 2.7912270853017545e-05
GC_5_329 b_5 NI_5 NS_329 0 5.6546243808870781e-05
GC_5_330 b_5 NI_5 NS_330 0 -6.4920680256422479e-06
GC_5_331 b_5 NI_5 NS_331 0 6.2764557963505549e-06
GC_5_332 b_5 NI_5 NS_332 0 -1.7734222969901383e-06
GC_5_333 b_5 NI_5 NS_333 0 -5.8493308428206880e-03
GC_5_334 b_5 NI_5 NS_334 0 8.9112016487685863e-03
GC_5_335 b_5 NI_5 NS_335 0 4.2883855088104456e-03
GC_5_336 b_5 NI_5 NS_336 0 -3.9254650144841053e-03
GC_5_337 b_5 NI_5 NS_337 0 -2.2543551512417683e-04
GC_5_338 b_5 NI_5 NS_338 0 1.6173885610339215e-04
GC_5_339 b_5 NI_5 NS_339 0 -8.9621890538372060e-07
GC_5_340 b_5 NI_5 NS_340 0 4.5080165507996325e-07
GC_5_341 b_5 NI_5 NS_341 0 -7.1820357026994300e-06
GC_5_342 b_5 NI_5 NS_342 0 5.0950835896534423e-05
GC_5_343 b_5 NI_5 NS_343 0 -1.6752471426881163e-07
GC_5_344 b_5 NI_5 NS_344 0 6.1315702703244971e-07
GC_5_345 b_5 NI_5 NS_345 0 8.9882225358147035e-07
GC_5_346 b_5 NI_5 NS_346 0 8.3013983883210874e-07
GC_5_347 b_5 NI_5 NS_347 0 -7.4655509108790996e-05
GC_5_348 b_5 NI_5 NS_348 0 -1.7674251278419740e-04
GC_5_349 b_5 NI_5 NS_349 0 -2.8288028214384025e-06
GC_5_350 b_5 NI_5 NS_350 0 -2.9368078386411271e-05
GC_5_351 b_5 NI_5 NS_351 0 -2.6804632783804232e-06
GC_5_352 b_5 NI_5 NS_352 0 -7.6383025819216025e-06
GC_5_353 b_5 NI_5 NS_353 0 -1.6158609900310664e-02
GC_5_354 b_5 NI_5 NS_354 0 9.1107310938880960e-05
GC_5_355 b_5 NI_5 NS_355 0 -4.3254019157889400e-04
GC_5_356 b_5 NI_5 NS_356 0 -1.8778414691806881e-03
GC_5_357 b_5 NI_5 NS_357 0 8.0261132069984749e-04
GC_5_358 b_5 NI_5 NS_358 0 -1.0036537689308688e-03
GC_5_359 b_5 NI_5 NS_359 0 2.0572436509997505e-03
GC_5_360 b_5 NI_5 NS_360 0 -1.5296001819546494e-03
GC_5_361 b_5 NI_5 NS_361 0 1.4875913351313262e-03
GC_5_362 b_5 NI_5 NS_362 0 5.0912717544941374e-04
GC_5_363 b_5 NI_5 NS_363 0 -2.8274675581329016e-03
GC_5_364 b_5 NI_5 NS_364 0 9.4844968661075108e-04
GC_5_365 b_5 NI_5 NS_365 0 4.8312754789078707e-04
GC_5_366 b_5 NI_5 NS_366 0 -3.3369915002472237e-04
GC_5_367 b_5 NI_5 NS_367 0 3.9123081488919324e-04
GC_5_368 b_5 NI_5 NS_368 0 8.9631101666165004e-04
GC_5_369 b_5 NI_5 NS_369 0 -2.8039633253659391e-03
GC_5_370 b_5 NI_5 NS_370 0 -2.3539979806315842e-03
GC_5_371 b_5 NI_5 NS_371 0 2.0109589934053833e-04
GC_5_372 b_5 NI_5 NS_372 0 1.4905611231955964e-04
GC_5_373 b_5 NI_5 NS_373 0 -1.0499536289492752e-03
GC_5_374 b_5 NI_5 NS_374 0 2.7558435783084639e-05
GC_5_375 b_5 NI_5 NS_375 0 -5.6646409242034266e-06
GC_5_376 b_5 NI_5 NS_376 0 -1.1322788231030885e-06
GC_5_377 b_5 NI_5 NS_377 0 1.5717068484343861e-02
GC_5_378 b_5 NI_5 NS_378 0 6.6254528864057990e-03
GC_5_379 b_5 NI_5 NS_379 0 -7.9304325621462717e-03
GC_5_380 b_5 NI_5 NS_380 0 -1.0255598463578866e-02
GC_5_381 b_5 NI_5 NS_381 0 -1.0155421041068711e-04
GC_5_382 b_5 NI_5 NS_382 0 5.9377354495698982e-04
GC_5_383 b_5 NI_5 NS_383 0 3.2944058727498684e-07
GC_5_384 b_5 NI_5 NS_384 0 2.3782145447755469e-07
GC_5_385 b_5 NI_5 NS_385 0 4.5743571821127855e-06
GC_5_386 b_5 NI_5 NS_386 0 -1.0484008446771693e-04
GC_5_387 b_5 NI_5 NS_387 0 3.4052897278504705e-07
GC_5_388 b_5 NI_5 NS_388 0 2.3972188554717713e-07
GC_5_389 b_5 NI_5 NS_389 0 -1.4652513307622286e-07
GC_5_390 b_5 NI_5 NS_390 0 -4.4748074803805727e-06
GC_5_391 b_5 NI_5 NS_391 0 3.0142477753232510e-04
GC_5_392 b_5 NI_5 NS_392 0 6.2621930701080482e-04
GC_5_393 b_5 NI_5 NS_393 0 -2.1232441495842505e-04
GC_5_394 b_5 NI_5 NS_394 0 1.0183783725932148e-04
GC_5_395 b_5 NI_5 NS_395 0 -1.9757008162512120e-05
GC_5_396 b_5 NI_5 NS_396 0 -9.2648038572561518e-06
GC_5_397 b_5 NI_5 NS_397 0 4.0771973492119679e-05
GC_5_398 b_5 NI_5 NS_398 0 -5.3422053168745934e-05
GC_5_399 b_5 NI_5 NS_399 0 -7.0358329661485966e-04
GC_5_400 b_5 NI_5 NS_400 0 2.0787877769915383e-03
GC_5_401 b_5 NI_5 NS_401 0 -2.5979038424229521e-03
GC_5_402 b_5 NI_5 NS_402 0 -1.6917059050189742e-03
GC_5_403 b_5 NI_5 NS_403 0 2.4394388692914554e-04
GC_5_404 b_5 NI_5 NS_404 0 -1.8902433044405760e-03
GC_5_405 b_5 NI_5 NS_405 0 1.7570369836857675e-06
GC_5_406 b_5 NI_5 NS_406 0 6.5621977445851651e-04
GC_5_407 b_5 NI_5 NS_407 0 -7.5300677769659665e-05
GC_5_408 b_5 NI_5 NS_408 0 -1.4134034929754050e-03
GC_5_409 b_5 NI_5 NS_409 0 -5.8893405805835468e-05
GC_5_410 b_5 NI_5 NS_410 0 3.1286283695248091e-04
GC_5_411 b_5 NI_5 NS_411 0 2.7373746834261439e-04
GC_5_412 b_5 NI_5 NS_412 0 -7.2621914665411223e-05
GC_5_413 b_5 NI_5 NS_413 0 -4.7303299005451441e-04
GC_5_414 b_5 NI_5 NS_414 0 -8.6860354969608549e-05
GC_5_415 b_5 NI_5 NS_415 0 -3.6753425372914035e-05
GC_5_416 b_5 NI_5 NS_416 0 -6.1355427865210463e-06
GC_5_417 b_5 NI_5 NS_417 0 -8.7028929771070906e-05
GC_5_418 b_5 NI_5 NS_418 0 -4.5614640458506617e-05
GC_5_419 b_5 NI_5 NS_419 0 4.9433072544480025e-06
GC_5_420 b_5 NI_5 NS_420 0 5.7013348990148853e-06
GC_5_421 b_5 NI_5 NS_421 0 6.0732001898286614e-03
GC_5_422 b_5 NI_5 NS_422 0 1.7476508141283384e-03
GC_5_423 b_5 NI_5 NS_423 0 -3.6093772074839992e-03
GC_5_424 b_5 NI_5 NS_424 0 -2.1348596486408127e-03
GC_5_425 b_5 NI_5 NS_425 0 3.1621814982850677e-05
GC_5_426 b_5 NI_5 NS_426 0 5.8924596118656960e-05
GC_5_427 b_5 NI_5 NS_427 0 -1.3506942149855566e-08
GC_5_428 b_5 NI_5 NS_428 0 4.8192706716479834e-07
GC_5_429 b_5 NI_5 NS_429 0 1.4552337178186976e-05
GC_5_430 b_5 NI_5 NS_430 0 -1.0268437044575696e-05
GC_5_431 b_5 NI_5 NS_431 0 -9.9978850373837202e-07
GC_5_432 b_5 NI_5 NS_432 0 5.8136052987070945e-07
GC_5_433 b_5 NI_5 NS_433 0 4.2496792251387462e-06
GC_5_434 b_5 NI_5 NS_434 0 -2.6335934197491776e-07
GC_5_435 b_5 NI_5 NS_435 0 -9.9741770373476334e-05
GC_5_436 b_5 NI_5 NS_436 0 -1.5869860359630127e-05
GC_5_437 b_5 NI_5 NS_437 0 -1.0699217883589780e-05
GC_5_438 b_5 NI_5 NS_438 0 -4.5737371146903026e-05
GC_5_439 b_5 NI_5 NS_439 0 -7.2236696280725936e-06
GC_5_440 b_5 NI_5 NS_440 0 5.3444761754046504e-06
GC_5_441 b_5 NI_5 NS_441 0 -7.5740530056836912e-03
GC_5_442 b_5 NI_5 NS_442 0 4.6628792659404756e-05
GC_5_443 b_5 NI_5 NS_443 0 1.9120424654356810e-03
GC_5_444 b_5 NI_5 NS_444 0 -1.5857972592648148e-03
GC_5_445 b_5 NI_5 NS_445 0 -1.1333027495970031e-03
GC_5_446 b_5 NI_5 NS_446 0 6.7014673491480484e-04
GC_5_447 b_5 NI_5 NS_447 0 2.4906704766540794e-03
GC_5_448 b_5 NI_5 NS_448 0 -6.4707425706389589e-05
GC_5_449 b_5 NI_5 NS_449 0 2.1093494273953650e-04
GC_5_450 b_5 NI_5 NS_450 0 8.1204703072574322e-04
GC_5_451 b_5 NI_5 NS_451 0 -3.3539868012653871e-03
GC_5_452 b_5 NI_5 NS_452 0 1.2068615863944978e-04
GC_5_453 b_5 NI_5 NS_453 0 4.2555997092495810e-04
GC_5_454 b_5 NI_5 NS_454 0 -1.7587611308956917e-04
GC_5_455 b_5 NI_5 NS_455 0 2.9436829290263350e-04
GC_5_456 b_5 NI_5 NS_456 0 6.1362507272142753e-04
GC_5_457 b_5 NI_5 NS_457 0 -1.6006799026690693e-03
GC_5_458 b_5 NI_5 NS_458 0 -1.4593086028127297e-03
GC_5_459 b_5 NI_5 NS_459 0 1.6731670520646303e-04
GC_5_460 b_5 NI_5 NS_460 0 1.2458632753298087e-04
GC_5_461 b_5 NI_5 NS_461 0 -6.7420663220518361e-04
GC_5_462 b_5 NI_5 NS_462 0 9.2119959799569541e-06
GC_5_463 b_5 NI_5 NS_463 0 -4.2469367752487059e-06
GC_5_464 b_5 NI_5 NS_464 0 -1.3434627151044835e-06
GC_5_465 b_5 NI_5 NS_465 0 9.2624482964964814e-03
GC_5_466 b_5 NI_5 NS_466 0 5.1206901426547047e-03
GC_5_467 b_5 NI_5 NS_467 0 -3.7979299271296662e-03
GC_5_468 b_5 NI_5 NS_468 0 -6.8446989339299401e-03
GC_5_469 b_5 NI_5 NS_469 0 -1.1424471249240921e-04
GC_5_470 b_5 NI_5 NS_470 0 3.3269716955616578e-04
GC_5_471 b_5 NI_5 NS_471 0 3.1697470688186859e-07
GC_5_472 b_5 NI_5 NS_472 0 5.6517218515745007e-08
GC_5_473 b_5 NI_5 NS_473 0 9.5350625057421993e-06
GC_5_474 b_5 NI_5 NS_474 0 -8.0270523981653370e-05
GC_5_475 b_5 NI_5 NS_475 0 4.4899288275093137e-07
GC_5_476 b_5 NI_5 NS_476 0 2.4706850582126317e-07
GC_5_477 b_5 NI_5 NS_477 0 1.8223765411241960e-07
GC_5_478 b_5 NI_5 NS_478 0 -2.3335350698957533e-06
GC_5_479 b_5 NI_5 NS_479 0 1.4808791392205892e-04
GC_5_480 b_5 NI_5 NS_480 0 4.5714727759423214e-04
GC_5_481 b_5 NI_5 NS_481 0 -1.4396786532958145e-04
GC_5_482 b_5 NI_5 NS_482 0 6.2618425750418958e-05
GC_5_483 b_5 NI_5 NS_483 0 -1.5086878181414736e-05
GC_5_484 b_5 NI_5 NS_484 0 -5.0400774213453882e-06
GC_5_485 b_5 NI_5 NS_485 0 -4.3958862252502081e-03
GC_5_486 b_5 NI_5 NS_486 0 -9.0777618995771335e-05
GC_5_487 b_5 NI_5 NS_487 0 -3.4404004717977464e-03
GC_5_488 b_5 NI_5 NS_488 0 2.0210165385460980e-03
GC_5_489 b_5 NI_5 NS_489 0 -4.9337974146412096e-04
GC_5_490 b_5 NI_5 NS_490 0 -4.0747012553577948e-03
GC_5_491 b_5 NI_5 NS_491 0 1.3970777582900397e-03
GC_5_492 b_5 NI_5 NS_492 0 -1.1760055933874791e-03
GC_5_493 b_5 NI_5 NS_493 0 1.6563892939223991e-04
GC_5_494 b_5 NI_5 NS_494 0 -1.4757526011808080e-04
GC_5_495 b_5 NI_5 NS_495 0 -9.7312484526983006e-04
GC_5_496 b_5 NI_5 NS_496 0 -2.8312976679026390e-03
GC_5_497 b_5 NI_5 NS_497 0 -1.0726088726844459e-04
GC_5_498 b_5 NI_5 NS_498 0 2.1933156711714948e-04
GC_5_499 b_5 NI_5 NS_499 0 2.0124271079450268e-04
GC_5_500 b_5 NI_5 NS_500 0 -5.4626912225828291e-05
GC_5_501 b_5 NI_5 NS_501 0 -9.9261163484215556e-05
GC_5_502 b_5 NI_5 NS_502 0 -1.6536522588633711e-04
GC_5_503 b_5 NI_5 NS_503 0 -3.2354395029787414e-05
GC_5_504 b_5 NI_5 NS_504 0 -2.5316888210246620e-05
GC_5_505 b_5 NI_5 NS_505 0 -4.7489227179093156e-05
GC_5_506 b_5 NI_5 NS_506 0 -5.6669282189402497e-05
GC_5_507 b_5 NI_5 NS_507 0 1.9670502485342276e-06
GC_5_508 b_5 NI_5 NS_508 0 4.5476291160873383e-07
GC_5_509 b_5 NI_5 NS_509 0 6.3088018014864199e-03
GC_5_510 b_5 NI_5 NS_510 0 2.8314688857696839e-03
GC_5_511 b_5 NI_5 NS_511 0 -3.0528998336207102e-03
GC_5_512 b_5 NI_5 NS_512 0 -2.4994549656510859e-03
GC_5_513 b_5 NI_5 NS_513 0 6.1556831549707216e-05
GC_5_514 b_5 NI_5 NS_514 0 2.1313256518463669e-04
GC_5_515 b_5 NI_5 NS_515 0 4.5412610207979066e-07
GC_5_516 b_5 NI_5 NS_516 0 1.0965892950274096e-06
GC_5_517 b_5 NI_5 NS_517 0 5.0102819824949663e-05
GC_5_518 b_5 NI_5 NS_518 0 4.6042427023939330e-06
GC_5_519 b_5 NI_5 NS_519 0 3.6648195719318533e-07
GC_5_520 b_5 NI_5 NS_520 0 1.9218476246556235e-07
GC_5_521 b_5 NI_5 NS_521 0 3.6178653853462982e-06
GC_5_522 b_5 NI_5 NS_522 0 5.3309154516238464e-07
GC_5_523 b_5 NI_5 NS_523 0 -1.4652616834783018e-04
GC_5_524 b_5 NI_5 NS_524 0 1.0880864250812918e-05
GC_5_525 b_5 NI_5 NS_525 0 -1.4894665965079207e-05
GC_5_526 b_5 NI_5 NS_526 0 -1.5389908727180548e-05
GC_5_527 b_5 NI_5 NS_527 0 -3.3165573412197533e-06
GC_5_528 b_5 NI_5 NS_528 0 7.0127921328692979e-06
GD_5_1 b_5 NI_5 NA_1 0 -2.2869906298709719e-02
GD_5_2 b_5 NI_5 NA_2 0 -3.6721389996634693e-03
GD_5_3 b_5 NI_5 NA_3 0 -3.0752557099579254e-02
GD_5_4 b_5 NI_5 NA_4 0 -1.2057227942289115e-02
GD_5_5 b_5 NI_5 NA_5 0 -1.8337541099106791e-01
GD_5_6 b_5 NI_5 NA_6 0 -1.6162878732128294e-02
GD_5_7 b_5 NI_5 NA_7 0 -2.1416087166423951e-02
GD_5_8 b_5 NI_5 NA_8 0 -2.6693183174679607e-03
GD_5_9 b_5 NI_5 NA_9 0 1.1174945952043472e-02
GD_5_10 b_5 NI_5 NA_10 0 1.3441709675942838e-03
GD_5_11 b_5 NI_5 NA_11 0 3.1059682420072235e-03
GD_5_12 b_5 NI_5 NA_12 0 5.6822052397968968e-03
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 1.4112468708611057e-02
GC_6_2 b_6 NI_6 NS_2 0 -6.0820585627221297e-04
GC_6_3 b_6 NI_6 NS_3 0 -1.5409865371543412e-02
GC_6_4 b_6 NI_6 NS_4 0 6.3372079764282370e-03
GC_6_5 b_6 NI_6 NS_5 0 2.3440157145031950e-03
GC_6_6 b_6 NI_6 NS_6 0 -1.2292674427882599e-02
GC_6_7 b_6 NI_6 NS_7 0 8.6622331958598770e-03
GC_6_8 b_6 NI_6 NS_8 0 9.3590176400118019e-04
GC_6_9 b_6 NI_6 NS_9 0 -4.2273216718258211e-04
GC_6_10 b_6 NI_6 NS_10 0 -6.2490282474033786e-04
GC_6_11 b_6 NI_6 NS_11 0 -7.4366755644204915e-03
GC_6_12 b_6 NI_6 NS_12 0 -2.5616625251924114e-03
GC_6_13 b_6 NI_6 NS_13 0 -2.8290821983852847e-04
GC_6_14 b_6 NI_6 NS_14 0 9.9873141396264594e-05
GC_6_15 b_6 NI_6 NS_15 0 1.4028345289085459e-04
GC_6_16 b_6 NI_6 NS_16 0 3.7184731672336273e-05
GC_6_17 b_6 NI_6 NS_17 0 6.0003137430694059e-04
GC_6_18 b_6 NI_6 NS_18 0 1.3116124746276580e-04
GC_6_19 b_6 NI_6 NS_19 0 2.6151008574502522e-05
GC_6_20 b_6 NI_6 NS_20 0 1.5509521873296917e-05
GC_6_21 b_6 NI_6 NS_21 0 5.2609416930517682e-05
GC_6_22 b_6 NI_6 NS_22 0 -1.6342984312426028e-05
GC_6_23 b_6 NI_6 NS_23 0 7.1935138306258568e-06
GC_6_24 b_6 NI_6 NS_24 0 -5.0563598433835042e-08
GC_6_25 b_6 NI_6 NS_25 0 -3.0349579133228039e-04
GC_6_26 b_6 NI_6 NS_26 0 3.1321499703063039e-03
GC_6_27 b_6 NI_6 NS_27 0 1.9318343152064878e-03
GC_6_28 b_6 NI_6 NS_28 0 -1.7750716646072577e-03
GC_6_29 b_6 NI_6 NS_29 0 1.7999948139529059e-05
GC_6_30 b_6 NI_6 NS_30 0 -2.6283026769945011e-05
GC_6_31 b_6 NI_6 NS_31 0 -1.5737649874535257e-07
GC_6_32 b_6 NI_6 NS_32 0 1.4176124851802802e-08
GC_6_33 b_6 NI_6 NS_33 0 5.8309901270279606e-06
GC_6_34 b_6 NI_6 NS_34 0 -1.3992874588016089e-05
GC_6_35 b_6 NI_6 NS_35 0 9.3550153847118511e-08
GC_6_36 b_6 NI_6 NS_36 0 -6.2686481096073009e-07
GC_6_37 b_6 NI_6 NS_37 0 3.1536238724834728e-06
GC_6_38 b_6 NI_6 NS_38 0 2.3639585707598339e-07
GC_6_39 b_6 NI_6 NS_39 0 -2.5270305902813830e-06
GC_6_40 b_6 NI_6 NS_40 0 2.8776869288140104e-05
GC_6_41 b_6 NI_6 NS_41 0 1.3870237329911900e-05
GC_6_42 b_6 NI_6 NS_42 0 1.4507190030808775e-05
GC_6_43 b_6 NI_6 NS_43 0 6.2453973555453573e-06
GC_6_44 b_6 NI_6 NS_44 0 -1.5536764595718731e-06
GC_6_45 b_6 NI_6 NS_45 0 -1.8304325853742670e-02
GC_6_46 b_6 NI_6 NS_46 0 9.4343763878071990e-05
GC_6_47 b_6 NI_6 NS_47 0 1.0992279551523477e-02
GC_6_48 b_6 NI_6 NS_48 0 -8.8287399600669985e-03
GC_6_49 b_6 NI_6 NS_49 0 -1.4721970915940253e-03
GC_6_50 b_6 NI_6 NS_50 0 7.3804244445370920e-03
GC_6_51 b_6 NI_6 NS_51 0 6.5444475108928186e-03
GC_6_52 b_6 NI_6 NS_52 0 7.2497330727034565e-05
GC_6_53 b_6 NI_6 NS_53 0 -2.1772676130101570e-03
GC_6_54 b_6 NI_6 NS_54 0 -2.0344017971621838e-03
GC_6_55 b_6 NI_6 NS_55 0 -1.0511637422557188e-03
GC_6_56 b_6 NI_6 NS_56 0 4.1364617698711149e-03
GC_6_57 b_6 NI_6 NS_57 0 1.0826425534843945e-04
GC_6_58 b_6 NI_6 NS_58 0 -1.3510495797180289e-04
GC_6_59 b_6 NI_6 NS_59 0 -7.3274034286389581e-06
GC_6_60 b_6 NI_6 NS_60 0 -3.6813368376286995e-05
GC_6_61 b_6 NI_6 NS_61 0 5.9208532565232521e-05
GC_6_62 b_6 NI_6 NS_62 0 -2.3283379809016139e-04
GC_6_63 b_6 NI_6 NS_63 0 -3.4391599992917248e-06
GC_6_64 b_6 NI_6 NS_64 0 -1.1077300717405246e-05
GC_6_65 b_6 NI_6 NS_65 0 -3.5853797609923269e-05
GC_6_66 b_6 NI_6 NS_66 0 -1.2023799108234140e-05
GC_6_67 b_6 NI_6 NS_67 0 -6.5784171957122770e-06
GC_6_68 b_6 NI_6 NS_68 0 -1.1001697587887688e-06
GC_6_69 b_6 NI_6 NS_69 0 5.1981096425168473e-03
GC_6_70 b_6 NI_6 NS_70 0 7.5917200122474120e-03
GC_6_71 b_6 NI_6 NS_71 0 -2.5683500636752444e-03
GC_6_72 b_6 NI_6 NS_72 0 -3.5182470795133143e-03
GC_6_73 b_6 NI_6 NS_73 0 -3.5119961975431553e-04
GC_6_74 b_6 NI_6 NS_74 0 -5.9277701984955511e-05
GC_6_75 b_6 NI_6 NS_75 0 -1.0106058346591284e-08
GC_6_76 b_6 NI_6 NS_76 0 8.7607962482880496e-07
GC_6_77 b_6 NI_6 NS_77 0 -7.8295119980793972e-05
GC_6_78 b_6 NI_6 NS_78 0 1.6659559371619051e-04
GC_6_79 b_6 NI_6 NS_79 0 -4.0090664178988577e-06
GC_6_80 b_6 NI_6 NS_80 0 -3.1648973391936408e-06
GC_6_81 b_6 NI_6 NS_81 0 -7.6632663683458638e-06
GC_6_82 b_6 NI_6 NS_82 0 -2.0112510740782898e-05
GC_6_83 b_6 NI_6 NS_83 0 -3.6834113681124663e-04
GC_6_84 b_6 NI_6 NS_84 0 1.5609629405501956e-04
GC_6_85 b_6 NI_6 NS_85 0 -1.9882963591359121e-04
GC_6_86 b_6 NI_6 NS_86 0 -5.9439222031193308e-05
GC_6_87 b_6 NI_6 NS_87 0 -4.1363970428794943e-05
GC_6_88 b_6 NI_6 NS_88 0 -5.6111904906493818e-06
GC_6_89 b_6 NI_6 NS_89 0 2.1741675366207473e-02
GC_6_90 b_6 NI_6 NS_90 0 -7.0767733721048770e-04
GC_6_91 b_6 NI_6 NS_91 0 -2.4103492833785080e-02
GC_6_92 b_6 NI_6 NS_92 0 2.0857034181942366e-03
GC_6_93 b_6 NI_6 NS_93 0 7.8016341299932653e-03
GC_6_94 b_6 NI_6 NS_94 0 -8.9897627851683211e-03
GC_6_95 b_6 NI_6 NS_95 0 1.0382015344121387e-02
GC_6_96 b_6 NI_6 NS_96 0 1.0956933802609376e-03
GC_6_97 b_6 NI_6 NS_97 0 -2.1120333646929550e-05
GC_6_98 b_6 NI_6 NS_98 0 1.0438424227287204e-03
GC_6_99 b_6 NI_6 NS_99 0 -5.6257911855354713e-03
GC_6_100 b_6 NI_6 NS_100 0 -6.4630736150212420e-03
GC_6_101 b_6 NI_6 NS_101 0 -3.6620978047084484e-04
GC_6_102 b_6 NI_6 NS_102 0 1.7291379601824407e-04
GC_6_103 b_6 NI_6 NS_103 0 2.1628794752744774e-04
GC_6_104 b_6 NI_6 NS_104 0 1.0406288522357281e-04
GC_6_105 b_6 NI_6 NS_105 0 5.1664554234123988e-04
GC_6_106 b_6 NI_6 NS_106 0 3.2572089182549371e-04
GC_6_107 b_6 NI_6 NS_107 0 3.0771089761729666e-05
GC_6_108 b_6 NI_6 NS_108 0 4.4270873586791591e-05
GC_6_109 b_6 NI_6 NS_109 0 7.3720422870431575e-05
GC_6_110 b_6 NI_6 NS_110 0 9.8804042273975063e-06
GC_6_111 b_6 NI_6 NS_111 0 8.8736175996478193e-06
GC_6_112 b_6 NI_6 NS_112 0 -4.4111079801958329e-07
GC_6_113 b_6 NI_6 NS_113 0 -4.0603204597342048e-03
GC_6_114 b_6 NI_6 NS_114 0 6.9355308562895155e-03
GC_6_115 b_6 NI_6 NS_115 0 4.2510532902162021e-03
GC_6_116 b_6 NI_6 NS_116 0 -3.0466215039111782e-03
GC_6_117 b_6 NI_6 NS_117 0 -9.3510920506042000e-05
GC_6_118 b_6 NI_6 NS_118 0 3.0181678768813940e-05
GC_6_119 b_6 NI_6 NS_119 0 -1.2736045548789990e-07
GC_6_120 b_6 NI_6 NS_120 0 -2.3136946862914335e-08
GC_6_121 b_6 NI_6 NS_121 0 6.4282585787549793e-06
GC_6_122 b_6 NI_6 NS_122 0 1.2877456111562950e-05
GC_6_123 b_6 NI_6 NS_123 0 -5.3253719615470932e-07
GC_6_124 b_6 NI_6 NS_124 0 -2.3353212463912596e-07
GC_6_125 b_6 NI_6 NS_125 0 -1.4391840947810239e-06
GC_6_126 b_6 NI_6 NS_126 0 -2.3459791001753782e-06
GC_6_127 b_6 NI_6 NS_127 0 1.8411541441936825e-05
GC_6_128 b_6 NI_6 NS_128 0 5.8513725805753612e-06
GC_6_129 b_6 NI_6 NS_129 0 7.0700508735465627e-06
GC_6_130 b_6 NI_6 NS_130 0 2.3792649206643453e-05
GC_6_131 b_6 NI_6 NS_131 0 1.7612973072130276e-06
GC_6_132 b_6 NI_6 NS_132 0 -4.1088855641264937e-06
GC_6_133 b_6 NI_6 NS_133 0 -1.9416588524809073e-02
GC_6_134 b_6 NI_6 NS_134 0 -7.4615686067070180e-04
GC_6_135 b_6 NI_6 NS_135 0 1.6105158561743358e-02
GC_6_136 b_6 NI_6 NS_136 0 -3.7351583856857899e-03
GC_6_137 b_6 NI_6 NS_137 0 -1.1137222575644999e-02
GC_6_138 b_6 NI_6 NS_138 0 3.9185227344225266e-04
GC_6_139 b_6 NI_6 NS_139 0 9.2206345693901810e-03
GC_6_140 b_6 NI_6 NS_140 0 -6.8232812035264956e-04
GC_6_141 b_6 NI_6 NS_141 0 -2.0524747598416990e-03
GC_6_142 b_6 NI_6 NS_142 0 5.4581271167415987e-05
GC_6_143 b_6 NI_6 NS_143 0 1.6080614885646686e-03
GC_6_144 b_6 NI_6 NS_144 0 1.3979481233104929e-03
GC_6_145 b_6 NI_6 NS_145 0 1.4224350608191874e-04
GC_6_146 b_6 NI_6 NS_146 0 -1.5902372605879829e-04
GC_6_147 b_6 NI_6 NS_147 0 1.9868385411701419e-06
GC_6_148 b_6 NI_6 NS_148 0 -2.8882779192636919e-05
GC_6_149 b_6 NI_6 NS_149 0 1.0048275540928518e-05
GC_6_150 b_6 NI_6 NS_150 0 -1.9636976086257989e-04
GC_6_151 b_6 NI_6 NS_151 0 1.5656797142947321e-06
GC_6_152 b_6 NI_6 NS_152 0 -7.4218636670945531e-06
GC_6_153 b_6 NI_6 NS_153 0 -2.0270584794906362e-05
GC_6_154 b_6 NI_6 NS_154 0 -1.2449759347736102e-05
GC_6_155 b_6 NI_6 NS_155 0 -5.0121853052891173e-06
GC_6_156 b_6 NI_6 NS_156 0 -5.9828597427127702e-07
GC_6_157 b_6 NI_6 NS_157 0 6.5906380909834424e-03
GC_6_158 b_6 NI_6 NS_158 0 9.3893546746954982e-03
GC_6_159 b_6 NI_6 NS_159 0 -2.6109538946935819e-03
GC_6_160 b_6 NI_6 NS_160 0 -4.2191037536823692e-03
GC_6_161 b_6 NI_6 NS_161 0 -3.7390052448463740e-04
GC_6_162 b_6 NI_6 NS_162 0 6.5001597106427789e-05
GC_6_163 b_6 NI_6 NS_163 0 -8.1958710179395253e-07
GC_6_164 b_6 NI_6 NS_164 0 1.8565788423578575e-06
GC_6_165 b_6 NI_6 NS_165 0 -3.5962724070231194e-05
GC_6_166 b_6 NI_6 NS_166 0 1.8810658404863924e-04
GC_6_167 b_6 NI_6 NS_167 0 -4.9033932065431646e-06
GC_6_168 b_6 NI_6 NS_168 0 -2.9326992908920130e-06
GC_6_169 b_6 NI_6 NS_169 0 -9.3865262007800513e-06
GC_6_170 b_6 NI_6 NS_170 0 -2.0049992673940773e-05
GC_6_171 b_6 NI_6 NS_171 0 -3.9349276260890843e-04
GC_6_172 b_6 NI_6 NS_172 0 1.9876592317708626e-04
GC_6_173 b_6 NI_6 NS_173 0 -2.2250355242589876e-04
GC_6_174 b_6 NI_6 NS_174 0 -4.3800112377559726e-05
GC_6_175 b_6 NI_6 NS_175 0 -4.0917490127282586e-05
GC_6_176 b_6 NI_6 NS_176 0 2.1432972345325082e-06
GC_6_177 b_6 NI_6 NS_177 0 4.7547290818107664e-02
GC_6_178 b_6 NI_6 NS_178 0 1.6148575703483766e-02
GC_6_179 b_6 NI_6 NS_179 0 -2.8784676938770175e-02
GC_6_180 b_6 NI_6 NS_180 0 1.3904415597774009e-03
GC_6_181 b_6 NI_6 NS_181 0 -2.8618554001337903e-02
GC_6_182 b_6 NI_6 NS_182 0 -9.2802340156127525e-03
GC_6_183 b_6 NI_6 NS_183 0 9.6204946360267801e-03
GC_6_184 b_6 NI_6 NS_184 0 2.5770766881009401e-03
GC_6_185 b_6 NI_6 NS_185 0 -2.6261267865963791e-03
GC_6_186 b_6 NI_6 NS_186 0 9.3809662928476554e-05
GC_6_187 b_6 NI_6 NS_187 0 1.3380579702192738e-03
GC_6_188 b_6 NI_6 NS_188 0 -2.9466270797785551e-03
GC_6_189 b_6 NI_6 NS_189 0 -5.0555633589762774e-04
GC_6_190 b_6 NI_6 NS_190 0 1.1060588345051277e-04
GC_6_191 b_6 NI_6 NS_191 0 1.3619834283354877e-04
GC_6_192 b_6 NI_6 NS_192 0 4.0475384268710406e-05
GC_6_193 b_6 NI_6 NS_193 0 6.9117352146444357e-04
GC_6_194 b_6 NI_6 NS_194 0 -3.7665960616931244e-04
GC_6_195 b_6 NI_6 NS_195 0 -3.3764247233357185e-06
GC_6_196 b_6 NI_6 NS_196 0 1.0564266413754897e-05
GC_6_197 b_6 NI_6 NS_197 0 -9.0504273426302934e-06
GC_6_198 b_6 NI_6 NS_198 0 -1.2975905285973577e-05
GC_6_199 b_6 NI_6 NS_199 0 7.7709107487828169e-06
GC_6_200 b_6 NI_6 NS_200 0 8.7534026355618751e-07
GC_6_201 b_6 NI_6 NS_201 0 -1.5794618792235573e-03
GC_6_202 b_6 NI_6 NS_202 0 -3.8550470293122795e-03
GC_6_203 b_6 NI_6 NS_203 0 1.4547170328720405e-03
GC_6_204 b_6 NI_6 NS_204 0 5.2850931172190993e-04
GC_6_205 b_6 NI_6 NS_205 0 1.1220256898846258e-04
GC_6_206 b_6 NI_6 NS_206 0 -5.3923010191989334e-05
GC_6_207 b_6 NI_6 NS_207 0 1.3133507411594797e-06
GC_6_208 b_6 NI_6 NS_208 0 1.1915904730954531e-07
GC_6_209 b_6 NI_6 NS_209 0 -8.9935687520718706e-06
GC_6_210 b_6 NI_6 NS_210 0 -5.5497877731408206e-05
GC_6_211 b_6 NI_6 NS_211 0 6.9625767762816229e-07
GC_6_212 b_6 NI_6 NS_212 0 -1.8260244037074301e-06
GC_6_213 b_6 NI_6 NS_213 0 6.6504835290182281e-06
GC_6_214 b_6 NI_6 NS_214 0 -2.9212251284492487e-06
GC_6_215 b_6 NI_6 NS_215 0 5.4536072809944510e-05
GC_6_216 b_6 NI_6 NS_216 0 1.3167163820848756e-04
GC_6_217 b_6 NI_6 NS_217 0 1.9319945599650413e-05
GC_6_218 b_6 NI_6 NS_218 0 2.7113163285906141e-05
GC_6_219 b_6 NI_6 NS_219 0 1.0086511961622308e-05
GC_6_220 b_6 NI_6 NS_220 0 -1.5525391085552296e-06
GC_6_221 b_6 NI_6 NS_221 0 -1.6036979482620947e-01
GC_6_222 b_6 NI_6 NS_222 0 1.8180573520598202e-02
GC_6_223 b_6 NI_6 NS_223 0 1.6103185985543361e-02
GC_6_224 b_6 NI_6 NS_224 0 2.3420820964802354e-03
GC_6_225 b_6 NI_6 NS_225 0 2.0628978578723856e-02
GC_6_226 b_6 NI_6 NS_226 0 -5.6143075882510536e-03
GC_6_227 b_6 NI_6 NS_227 0 6.8412269830907804e-03
GC_6_228 b_6 NI_6 NS_228 0 1.6638614438991991e-03
GC_6_229 b_6 NI_6 NS_229 0 -2.3471875184899738e-03
GC_6_230 b_6 NI_6 NS_230 0 -6.1919328141470391e-04
GC_6_231 b_6 NI_6 NS_231 0 6.6616119731378581e-03
GC_6_232 b_6 NI_6 NS_232 0 6.1516398835021278e-03
GC_6_233 b_6 NI_6 NS_233 0 3.0524911619771507e-05
GC_6_234 b_6 NI_6 NS_234 0 -2.7437074147511651e-04
GC_6_235 b_6 NI_6 NS_235 0 -3.1903054136525899e-05
GC_6_236 b_6 NI_6 NS_236 0 -9.7464419193481550e-05
GC_6_237 b_6 NI_6 NS_237 0 2.6686632079201783e-04
GC_6_238 b_6 NI_6 NS_238 0 -4.6199643468073048e-04
GC_6_239 b_6 NI_6 NS_239 0 5.0988317424300034e-06
GC_6_240 b_6 NI_6 NS_240 0 -2.9519435757094257e-05
GC_6_241 b_6 NI_6 NS_241 0 -3.6614068194187411e-05
GC_6_242 b_6 NI_6 NS_242 0 -4.5405040724007015e-05
GC_6_243 b_6 NI_6 NS_243 0 -8.8640440392632303e-06
GC_6_244 b_6 NI_6 NS_244 0 -4.6261142796860233e-06
GC_6_245 b_6 NI_6 NS_245 0 6.9442178895966298e-03
GC_6_246 b_6 NI_6 NS_246 0 1.3325937100555263e-02
GC_6_247 b_6 NI_6 NS_247 0 -3.1900741482660511e-03
GC_6_248 b_6 NI_6 NS_248 0 -6.2387090453656265e-03
GC_6_249 b_6 NI_6 NS_249 0 -6.2198478071561749e-04
GC_6_250 b_6 NI_6 NS_250 0 -4.4903918916213108e-05
GC_6_251 b_6 NI_6 NS_251 0 -1.0851883511386824e-07
GC_6_252 b_6 NI_6 NS_252 0 5.6520959402104324e-07
GC_6_253 b_6 NI_6 NS_253 0 -1.1446935607342421e-04
GC_6_254 b_6 NI_6 NS_254 0 2.8274520033535149e-04
GC_6_255 b_6 NI_6 NS_255 0 -7.5197961160966510e-06
GC_6_256 b_6 NI_6 NS_256 0 -3.3307551218280824e-06
GC_6_257 b_6 NI_6 NS_257 0 -1.5476577159977199e-05
GC_6_258 b_6 NI_6 NS_258 0 -3.1363472703098145e-05
GC_6_259 b_6 NI_6 NS_259 0 -5.5518129971253590e-04
GC_6_260 b_6 NI_6 NS_260 0 1.8362641922669299e-04
GC_6_261 b_6 NI_6 NS_261 0 -3.2298267639991132e-04
GC_6_262 b_6 NI_6 NS_262 0 -9.2316235180612996e-05
GC_6_263 b_6 NI_6 NS_263 0 -5.8708061017615501e-05
GC_6_264 b_6 NI_6 NS_264 0 -2.5338662126368369e-06
GC_6_265 b_6 NI_6 NS_265 0 6.1507866044296106e-03
GC_6_266 b_6 NI_6 NS_266 0 -3.8636957925102287e-04
GC_6_267 b_6 NI_6 NS_267 0 -2.0319170926007633e-02
GC_6_268 b_6 NI_6 NS_268 0 -2.9799757317841547e-03
GC_6_269 b_6 NI_6 NS_269 0 1.0030808512120916e-02
GC_6_270 b_6 NI_6 NS_270 0 -3.4804738917802737e-03
GC_6_271 b_6 NI_6 NS_271 0 6.1236368894866675e-03
GC_6_272 b_6 NI_6 NS_272 0 6.4978683405598114e-04
GC_6_273 b_6 NI_6 NS_273 0 1.4531255133526193e-03
GC_6_274 b_6 NI_6 NS_274 0 -2.7388354097491698e-05
GC_6_275 b_6 NI_6 NS_275 0 -2.7195649467449951e-04
GC_6_276 b_6 NI_6 NS_276 0 -8.8213910496476172e-03
GC_6_277 b_6 NI_6 NS_277 0 -2.6856746714925596e-04
GC_6_278 b_6 NI_6 NS_278 0 1.0823191844131195e-04
GC_6_279 b_6 NI_6 NS_279 0 2.1792848461554538e-04
GC_6_280 b_6 NI_6 NS_280 0 3.8412687463668644e-05
GC_6_281 b_6 NI_6 NS_281 0 4.6922798432008270e-04
GC_6_282 b_6 NI_6 NS_282 0 4.1093464334406986e-04
GC_6_283 b_6 NI_6 NS_283 0 4.0985501595778674e-05
GC_6_284 b_6 NI_6 NS_284 0 2.7208120908522104e-05
GC_6_285 b_6 NI_6 NS_285 0 8.3515005410065478e-05
GC_6_286 b_6 NI_6 NS_286 0 -1.9874247028458764e-05
GC_6_287 b_6 NI_6 NS_287 0 7.8069488171924485e-06
GC_6_288 b_6 NI_6 NS_288 0 -9.9686667968113612e-07
GC_6_289 b_6 NI_6 NS_289 0 -4.8530597783347064e-03
GC_6_290 b_6 NI_6 NS_290 0 9.8910022813513566e-03
GC_6_291 b_6 NI_6 NS_291 0 3.9529174469969206e-03
GC_6_292 b_6 NI_6 NS_292 0 -4.3989992597532109e-03
GC_6_293 b_6 NI_6 NS_293 0 -2.4430289336018233e-04
GC_6_294 b_6 NI_6 NS_294 0 1.4055318610111325e-04
GC_6_295 b_6 NI_6 NS_295 0 -5.4456124827200396e-07
GC_6_296 b_6 NI_6 NS_296 0 2.8277985714279663e-07
GC_6_297 b_6 NI_6 NS_297 0 -1.4539573798198310e-05
GC_6_298 b_6 NI_6 NS_298 0 5.5277592759158462e-05
GC_6_299 b_6 NI_6 NS_299 0 -8.6591885968592924e-07
GC_6_300 b_6 NI_6 NS_300 0 7.3752165611195587e-07
GC_6_301 b_6 NI_6 NS_301 0 -2.6196530735306848e-06
GC_6_302 b_6 NI_6 NS_302 0 -1.0301308436893354e-06
GC_6_303 b_6 NI_6 NS_303 0 -7.4525893843541889e-05
GC_6_304 b_6 NI_6 NS_304 0 -1.2986853872844846e-04
GC_6_305 b_6 NI_6 NS_305 0 -1.9115744390457456e-05
GC_6_306 b_6 NI_6 NS_306 0 -3.2863758292850780e-05
GC_6_307 b_6 NI_6 NS_307 0 -8.2088450398930087e-06
GC_6_308 b_6 NI_6 NS_308 0 -8.3685220571300952e-06
GC_6_309 b_6 NI_6 NS_309 0 -9.7066265209022947e-03
GC_6_310 b_6 NI_6 NS_310 0 -9.4596811027398519e-04
GC_6_311 b_6 NI_6 NS_311 0 1.3631649729863639e-02
GC_6_312 b_6 NI_6 NS_312 0 2.7905397308381772e-03
GC_6_313 b_6 NI_6 NS_313 0 -1.5667987275341612e-02
GC_6_314 b_6 NI_6 NS_314 0 -3.6561043783437837e-03
GC_6_315 b_6 NI_6 NS_315 0 5.4852631635970124e-03
GC_6_316 b_6 NI_6 NS_316 0 -1.3271597842458836e-03
GC_6_317 b_6 NI_6 NS_317 0 -7.3861607460020534e-04
GC_6_318 b_6 NI_6 NS_318 0 6.8618872769703925e-04
GC_6_319 b_6 NI_6 NS_319 0 1.9224541293903555e-03
GC_6_320 b_6 NI_6 NS_320 0 -3.5056746073897681e-03
GC_6_321 b_6 NI_6 NS_321 0 8.7739258958878410e-05
GC_6_322 b_6 NI_6 NS_322 0 -1.3437037900940755e-04
GC_6_323 b_6 NI_6 NS_323 0 1.4876582476162522e-05
GC_6_324 b_6 NI_6 NS_324 0 -3.8187390179365162e-05
GC_6_325 b_6 NI_6 NS_325 0 7.5485542792309038e-05
GC_6_326 b_6 NI_6 NS_326 0 -7.5105405971183747e-05
GC_6_327 b_6 NI_6 NS_327 0 4.4239403579608258e-06
GC_6_328 b_6 NI_6 NS_328 0 -8.4701318977602430e-06
GC_6_329 b_6 NI_6 NS_329 0 -1.3698030329988629e-05
GC_6_330 b_6 NI_6 NS_330 0 -1.3952994160185997e-05
GC_6_331 b_6 NI_6 NS_331 0 -4.1088225143976469e-06
GC_6_332 b_6 NI_6 NS_332 0 -9.6123718560977532e-07
GC_6_333 b_6 NI_6 NS_333 0 7.4074546445994562e-03
GC_6_334 b_6 NI_6 NS_334 0 6.9523945611948820e-03
GC_6_335 b_6 NI_6 NS_335 0 -2.8837180862516642e-03
GC_6_336 b_6 NI_6 NS_336 0 -3.3439362559328938e-03
GC_6_337 b_6 NI_6 NS_337 0 -2.4770875036417999e-04
GC_6_338 b_6 NI_6 NS_338 0 7.5608802933867247e-05
GC_6_339 b_6 NI_6 NS_339 0 -3.3714632772069532e-07
GC_6_340 b_6 NI_6 NS_340 0 1.5975625822864345e-06
GC_6_341 b_6 NI_6 NS_341 0 -1.1933144619880322e-05
GC_6_342 b_6 NI_6 NS_342 0 1.2769747154881423e-04
GC_6_343 b_6 NI_6 NS_343 0 -2.9501731132763868e-06
GC_6_344 b_6 NI_6 NS_344 0 -7.3138894122136900e-07
GC_6_345 b_6 NI_6 NS_345 0 -7.0394952714519611e-06
GC_6_346 b_6 NI_6 NS_346 0 -1.8912958483678779e-05
GC_6_347 b_6 NI_6 NS_347 0 -3.1588707384847182e-04
GC_6_348 b_6 NI_6 NS_348 0 1.8334380777710799e-04
GC_6_349 b_6 NI_6 NS_349 0 -1.8513841179665865e-04
GC_6_350 b_6 NI_6 NS_350 0 -3.3901960157504569e-05
GC_6_351 b_6 NI_6 NS_351 0 -2.3165393931028059e-05
GC_6_352 b_6 NI_6 NS_352 0 1.0566553169891282e-05
GC_6_353 b_6 NI_6 NS_353 0 -5.2199223672356928e-05
GC_6_354 b_6 NI_6 NS_354 0 -5.2140906564589991e-05
GC_6_355 b_6 NI_6 NS_355 0 -7.0738106743112544e-04
GC_6_356 b_6 NI_6 NS_356 0 2.0717716619665255e-03
GC_6_357 b_6 NI_6 NS_357 0 -2.5928282580306625e-03
GC_6_358 b_6 NI_6 NS_358 0 -1.6990340159135067e-03
GC_6_359 b_6 NI_6 NS_359 0 2.4115312859618532e-04
GC_6_360 b_6 NI_6 NS_360 0 -1.8967101241772779e-03
GC_6_361 b_6 NI_6 NS_361 0 2.3977634774642105e-05
GC_6_362 b_6 NI_6 NS_362 0 6.8445141771105312e-04
GC_6_363 b_6 NI_6 NS_363 0 -8.3743548490737002e-05
GC_6_364 b_6 NI_6 NS_364 0 -1.4351597035106587e-03
GC_6_365 b_6 NI_6 NS_365 0 -5.7653040097257286e-05
GC_6_366 b_6 NI_6 NS_366 0 3.1313225657391075e-04
GC_6_367 b_6 NI_6 NS_367 0 2.7375028563988215e-04
GC_6_368 b_6 NI_6 NS_368 0 -7.1122349996501481e-05
GC_6_369 b_6 NI_6 NS_369 0 -4.8207527221316471e-04
GC_6_370 b_6 NI_6 NS_370 0 -9.0787482154614354e-05
GC_6_371 b_6 NI_6 NS_371 0 -3.7600020720387231e-05
GC_6_372 b_6 NI_6 NS_372 0 -5.4726523660381245e-06
GC_6_373 b_6 NI_6 NS_373 0 -9.0613464194235860e-05
GC_6_374 b_6 NI_6 NS_374 0 -4.4807556787525997e-05
GC_6_375 b_6 NI_6 NS_375 0 4.6109873444846013e-06
GC_6_376 b_6 NI_6 NS_376 0 5.7909092212214392e-06
GC_6_377 b_6 NI_6 NS_377 0 6.2277055389356418e-03
GC_6_378 b_6 NI_6 NS_378 0 1.6826596581070163e-03
GC_6_379 b_6 NI_6 NS_379 0 -3.7003658959584439e-03
GC_6_380 b_6 NI_6 NS_380 0 -2.1166610807514864e-03
GC_6_381 b_6 NI_6 NS_381 0 3.4200685744665795e-05
GC_6_382 b_6 NI_6 NS_382 0 6.3527253615423018e-05
GC_6_383 b_6 NI_6 NS_383 0 2.8980174057699267e-08
GC_6_384 b_6 NI_6 NS_384 0 4.9038390907175583e-07
GC_6_385 b_6 NI_6 NS_385 0 1.5243759811507297e-05
GC_6_386 b_6 NI_6 NS_386 0 -9.4672361167612725e-06
GC_6_387 b_6 NI_6 NS_387 0 -9.6353746656365482e-07
GC_6_388 b_6 NI_6 NS_388 0 6.2614716561419949e-07
GC_6_389 b_6 NI_6 NS_389 0 4.1113230934106040e-06
GC_6_390 b_6 NI_6 NS_390 0 -2.6724157170140923e-07
GC_6_391 b_6 NI_6 NS_391 0 -1.0216090963299474e-04
GC_6_392 b_6 NI_6 NS_392 0 -1.1184956838462202e-05
GC_6_393 b_6 NI_6 NS_393 0 -1.2887820877097823e-05
GC_6_394 b_6 NI_6 NS_394 0 -4.4744706242927303e-05
GC_6_395 b_6 NI_6 NS_395 0 -7.0801867836624319e-06
GC_6_396 b_6 NI_6 NS_396 0 5.7174045974277323e-06
GC_6_397 b_6 NI_6 NS_397 0 -1.0559914108872998e-02
GC_6_398 b_6 NI_6 NS_398 0 2.0843816288909439e-05
GC_6_399 b_6 NI_6 NS_399 0 -3.3160410006659790e-04
GC_6_400 b_6 NI_6 NS_400 0 -1.8547698665160232e-03
GC_6_401 b_6 NI_6 NS_401 0 1.2558829888192104e-03
GC_6_402 b_6 NI_6 NS_402 0 -7.1109852709456498e-05
GC_6_403 b_6 NI_6 NS_403 0 6.1086631612852966e-04
GC_6_404 b_6 NI_6 NS_404 0 -1.1819412533399724e-03
GC_6_405 b_6 NI_6 NS_405 0 7.5931312693843314e-04
GC_6_406 b_6 NI_6 NS_406 0 1.6950600306736511e-04
GC_6_407 b_6 NI_6 NS_407 0 1.0237219393123965e-03
GC_6_408 b_6 NI_6 NS_408 0 5.1774325617669952e-04
GC_6_409 b_6 NI_6 NS_409 0 -1.0576257059065527e-04
GC_6_410 b_6 NI_6 NS_410 0 -8.7955211826900049e-05
GC_6_411 b_6 NI_6 NS_411 0 3.8776716427546895e-05
GC_6_412 b_6 NI_6 NS_412 0 -3.4867364586854898e-05
GC_6_413 b_6 NI_6 NS_413 0 -2.8656566598413743e-04
GC_6_414 b_6 NI_6 NS_414 0 2.5662598428824576e-04
GC_6_415 b_6 NI_6 NS_415 0 -1.5192572833024995e-05
GC_6_416 b_6 NI_6 NS_416 0 3.2850873558218179e-05
GC_6_417 b_6 NI_6 NS_417 0 -9.2917700878562658e-06
GC_6_418 b_6 NI_6 NS_418 0 1.0250305606663257e-04
GC_6_419 b_6 NI_6 NS_419 0 -5.6727872977306927e-07
GC_6_420 b_6 NI_6 NS_420 0 -2.5365804543112824e-07
GC_6_421 b_6 NI_6 NS_421 0 3.9666274569757154e-03
GC_6_422 b_6 NI_6 NS_422 0 -5.4840565659618045e-03
GC_6_423 b_6 NI_6 NS_423 0 -2.7124172157682912e-03
GC_6_424 b_6 NI_6 NS_424 0 3.3085644318646122e-03
GC_6_425 b_6 NI_6 NS_425 0 1.8443797145728619e-04
GC_6_426 b_6 NI_6 NS_426 0 -8.8841184609456139e-06
GC_6_427 b_6 NI_6 NS_427 0 3.4347412548187931e-06
GC_6_428 b_6 NI_6 NS_428 0 -2.7204144181219287e-07
GC_6_429 b_6 NI_6 NS_429 0 -3.4931913086156694e-05
GC_6_430 b_6 NI_6 NS_430 0 -8.6845363855787310e-05
GC_6_431 b_6 NI_6 NS_431 0 5.7021823891697587e-06
GC_6_432 b_6 NI_6 NS_432 0 1.1695718697364809e-05
GC_6_433 b_6 NI_6 NS_433 0 -1.7455794820947887e-05
GC_6_434 b_6 NI_6 NS_434 0 -3.6198380777827585e-05
GC_6_435 b_6 NI_6 NS_435 0 -4.1973154696239698e-05
GC_6_436 b_6 NI_6 NS_436 0 3.7033176494602574e-04
GC_6_437 b_6 NI_6 NS_437 0 -3.0302824596563458e-04
GC_6_438 b_6 NI_6 NS_438 0 3.9296931700078912e-06
GC_6_439 b_6 NI_6 NS_439 0 6.4708976052815927e-05
GC_6_440 b_6 NI_6 NS_440 0 8.3236597939826071e-05
GC_6_441 b_6 NI_6 NS_441 0 -4.6147298263072073e-03
GC_6_442 b_6 NI_6 NS_442 0 -9.1507982483837399e-05
GC_6_443 b_6 NI_6 NS_443 0 -3.4538995597095373e-03
GC_6_444 b_6 NI_6 NS_444 0 2.0673691360280477e-03
GC_6_445 b_6 NI_6 NS_445 0 -5.8284116660255484e-04
GC_6_446 b_6 NI_6 NS_446 0 -4.1404342208974159e-03
GC_6_447 b_6 NI_6 NS_447 0 1.4316771262851851e-03
GC_6_448 b_6 NI_6 NS_448 0 -1.2519594612108056e-03
GC_6_449 b_6 NI_6 NS_449 0 2.6670833434100719e-04
GC_6_450 b_6 NI_6 NS_450 0 -8.4215514876752147e-06
GC_6_451 b_6 NI_6 NS_451 0 -1.0216583821127190e-03
GC_6_452 b_6 NI_6 NS_452 0 -2.8396194224716395e-03
GC_6_453 b_6 NI_6 NS_453 0 -1.0674678049317115e-04
GC_6_454 b_6 NI_6 NS_454 0 2.2366888654651220e-04
GC_6_455 b_6 NI_6 NS_455 0 1.9107917520206469e-04
GC_6_456 b_6 NI_6 NS_456 0 -6.5344362238967788e-05
GC_6_457 b_6 NI_6 NS_457 0 -9.1262700151106750e-05
GC_6_458 b_6 NI_6 NS_458 0 -1.4993492801851786e-04
GC_6_459 b_6 NI_6 NS_459 0 -1.6403030620519296e-05
GC_6_460 b_6 NI_6 NS_460 0 -1.8273693849294730e-05
GC_6_461 b_6 NI_6 NS_461 0 -4.9930957324176615e-05
GC_6_462 b_6 NI_6 NS_462 0 -6.2139820596162265e-05
GC_6_463 b_6 NI_6 NS_463 0 3.5330616217318078e-06
GC_6_464 b_6 NI_6 NS_464 0 1.6964493760107395e-06
GC_6_465 b_6 NI_6 NS_465 0 6.2934678356185055e-03
GC_6_466 b_6 NI_6 NS_466 0 2.1224042927910250e-03
GC_6_467 b_6 NI_6 NS_467 0 -3.0165293495987167e-03
GC_6_468 b_6 NI_6 NS_468 0 -2.0750248415268946e-03
GC_6_469 b_6 NI_6 NS_469 0 7.1025223875465589e-05
GC_6_470 b_6 NI_6 NS_470 0 2.0943215080856920e-04
GC_6_471 b_6 NI_6 NS_471 0 3.3258300127674759e-07
GC_6_472 b_6 NI_6 NS_472 0 8.7719277560942442e-07
GC_6_473 b_6 NI_6 NS_473 0 5.4092566814911349e-05
GC_6_474 b_6 NI_6 NS_474 0 -1.1669013086254587e-06
GC_6_475 b_6 NI_6 NS_475 0 1.8059205099185046e-06
GC_6_476 b_6 NI_6 NS_476 0 -3.4863155656352324e-07
GC_6_477 b_6 NI_6 NS_477 0 -5.1640227808602503e-07
GC_6_478 b_6 NI_6 NS_478 0 -1.6096646465374173e-06
GC_6_479 b_6 NI_6 NS_479 0 -9.3868188881660749e-05
GC_6_480 b_6 NI_6 NS_480 0 4.8865629715452607e-05
GC_6_481 b_6 NI_6 NS_481 0 -3.8746122828526170e-05
GC_6_482 b_6 NI_6 NS_482 0 -1.3114751928981409e-06
GC_6_483 b_6 NI_6 NS_483 0 4.4417562018513674e-06
GC_6_484 b_6 NI_6 NS_484 0 6.8494639327604105e-06
GC_6_485 b_6 NI_6 NS_485 0 -6.5775107440052029e-03
GC_6_486 b_6 NI_6 NS_486 0 1.3709303852555791e-05
GC_6_487 b_6 NI_6 NS_487 0 2.1081904113967212e-03
GC_6_488 b_6 NI_6 NS_488 0 -2.2925817218598685e-03
GC_6_489 b_6 NI_6 NS_489 0 -4.0290652845791070e-04
GC_6_490 b_6 NI_6 NS_490 0 2.3106704686941195e-03
GC_6_491 b_6 NI_6 NS_491 0 7.1393542789883709e-04
GC_6_492 b_6 NI_6 NS_492 0 -6.6889357741712989e-04
GC_6_493 b_6 NI_6 NS_493 0 3.9387720606288572e-04
GC_6_494 b_6 NI_6 NS_494 0 -1.0217273075937490e-04
GC_6_495 b_6 NI_6 NS_495 0 -4.1847632698007446e-04
GC_6_496 b_6 NI_6 NS_496 0 3.8358518306348910e-04
GC_6_497 b_6 NI_6 NS_497 0 -5.4446268966694457e-05
GC_6_498 b_6 NI_6 NS_498 0 -9.6901709719871088e-05
GC_6_499 b_6 NI_6 NS_499 0 2.8557372980684706e-05
GC_6_500 b_6 NI_6 NS_500 0 -4.0820152391292421e-05
GC_6_501 b_6 NI_6 NS_501 0 -1.0444586353167934e-04
GC_6_502 b_6 NI_6 NS_502 0 1.0947178771901545e-04
GC_6_503 b_6 NI_6 NS_503 0 -9.1462794701515412e-06
GC_6_504 b_6 NI_6 NS_504 0 9.6433512051565493e-06
GC_6_505 b_6 NI_6 NS_505 0 -1.0532786818935184e-05
GC_6_506 b_6 NI_6 NS_506 0 4.0942520585255448e-05
GC_6_507 b_6 NI_6 NS_507 0 -1.4333373087439636e-06
GC_6_508 b_6 NI_6 NS_508 0 2.7864853720127531e-07
GC_6_509 b_6 NI_6 NS_509 0 2.8146570081552169e-03
GC_6_510 b_6 NI_6 NS_510 0 -2.0759944606451434e-03
GC_6_511 b_6 NI_6 NS_511 0 -1.7758096632358119e-03
GC_6_512 b_6 NI_6 NS_512 0 1.1015225488893489e-03
GC_6_513 b_6 NI_6 NS_513 0 2.9428568477516061e-05
GC_6_514 b_6 NI_6 NS_514 0 -3.7008624955722896e-05
GC_6_515 b_6 NI_6 NS_515 0 1.6465548220706839e-06
GC_6_516 b_6 NI_6 NS_516 0 -3.3987603491866489e-07
GC_6_517 b_6 NI_6 NS_517 0 -2.3709565226938377e-05
GC_6_518 b_6 NI_6 NS_518 0 -1.3494367349675637e-05
GC_6_519 b_6 NI_6 NS_519 0 7.5996048406742090e-07
GC_6_520 b_6 NI_6 NS_520 0 5.2410059679893349e-06
GC_6_521 b_6 NI_6 NS_521 0 -9.1527659293328630e-06
GC_6_522 b_6 NI_6 NS_522 0 -2.1591622628735276e-05
GC_6_523 b_6 NI_6 NS_523 0 -4.6005615822902157e-05
GC_6_524 b_6 NI_6 NS_524 0 1.8503668660785320e-04
GC_6_525 b_6 NI_6 NS_525 0 -1.5662841441585216e-04
GC_6_526 b_6 NI_6 NS_526 0 -6.5461622154032698e-06
GC_6_527 b_6 NI_6 NS_527 0 2.6304267973395834e-05
GC_6_528 b_6 NI_6 NS_528 0 3.8665299374378454e-05
GD_6_1 b_6 NI_6 NA_1 0 -3.5671852664924475e-03
GD_6_2 b_6 NI_6 NA_2 0 1.3532982709400878e-03
GD_6_3 b_6 NI_6 NA_3 0 -1.3246278655202713e-02
GD_6_4 b_6 NI_6 NA_4 0 8.8946856248933704e-04
GD_6_5 b_6 NI_6 NA_5 0 -1.6162878732134619e-02
GD_6_6 b_6 NI_6 NA_6 0 1.2773641717724929e-01
GD_6_7 b_6 NI_6 NA_7 0 -3.6884604259927816e-03
GD_6_8 b_6 NI_6 NA_8 0 -9.6644532438176805e-05
GD_6_9 b_6 NI_6 NA_9 0 1.3317487238180821e-03
GD_6_10 b_6 NI_6 NA_10 0 7.5521511839722298e-03
GD_6_11 b_6 NI_6 NA_11 0 5.8234355331995315e-03
GD_6_12 b_6 NI_6 NA_12 0 3.7310735701665976e-03
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 8.0678348141416147e-03
GC_7_2 b_7 NI_7 NS_2 0 2.4279265951727863e-04
GC_7_3 b_7 NI_7 NS_3 0 7.0724015355783107e-03
GC_7_4 b_7 NI_7 NS_4 0 -7.0940926046936604e-03
GC_7_5 b_7 NI_7 NS_5 0 3.3452930912150516e-03
GC_7_6 b_7 NI_7 NS_6 0 7.8189965493124791e-03
GC_7_7 b_7 NI_7 NS_7 0 9.6302829097820470e-03
GC_7_8 b_7 NI_7 NS_8 0 7.7632217464526799e-03
GC_7_9 b_7 NI_7 NS_9 0 2.1695161319534653e-05
GC_7_10 b_7 NI_7 NS_10 0 -3.7467283856284423e-03
GC_7_11 b_7 NI_7 NS_11 0 -1.3029598792570016e-02
GC_7_12 b_7 NI_7 NS_12 0 1.1815842226089800e-02
GC_7_13 b_7 NI_7 NS_13 0 4.2549892168000387e-04
GC_7_14 b_7 NI_7 NS_14 0 2.9282716494638186e-04
GC_7_15 b_7 NI_7 NS_15 0 3.6567343485953687e-05
GC_7_16 b_7 NI_7 NS_16 0 2.2547725912695277e-04
GC_7_17 b_7 NI_7 NS_17 0 5.2629767312816302e-04
GC_7_18 b_7 NI_7 NS_18 0 -2.7813714694784319e-04
GC_7_19 b_7 NI_7 NS_19 0 9.5387529800151598e-05
GC_7_20 b_7 NI_7 NS_20 0 1.1274327254585065e-04
GC_7_21 b_7 NI_7 NS_21 0 4.5339081751346355e-05
GC_7_22 b_7 NI_7 NS_22 0 5.4219000620850692e-05
GC_7_23 b_7 NI_7 NS_23 0 -6.6504745767974843e-06
GC_7_24 b_7 NI_7 NS_24 0 2.6857297221467853e-06
GC_7_25 b_7 NI_7 NS_25 0 -1.8209602962112655e-02
GC_7_26 b_7 NI_7 NS_26 0 -7.7990122981954164e-03
GC_7_27 b_7 NI_7 NS_27 0 9.6141322539971836e-03
GC_7_28 b_7 NI_7 NS_28 0 5.1853209234924398e-03
GC_7_29 b_7 NI_7 NS_29 0 -1.6326950250375200e-04
GC_7_30 b_7 NI_7 NS_30 0 -4.4113601250547795e-04
GC_7_31 b_7 NI_7 NS_31 0 7.8930443643316344e-07
GC_7_32 b_7 NI_7 NS_32 0 2.8147367237137539e-08
GC_7_33 b_7 NI_7 NS_33 0 4.8560994068586401e-05
GC_7_34 b_7 NI_7 NS_34 0 -5.4730653968546579e-05
GC_7_35 b_7 NI_7 NS_35 0 1.1114820923336849e-06
GC_7_36 b_7 NI_7 NS_36 0 -1.3801920749524094e-07
GC_7_37 b_7 NI_7 NS_37 0 -8.9165880659144122e-07
GC_7_38 b_7 NI_7 NS_38 0 -2.6989598376235418e-06
GC_7_39 b_7 NI_7 NS_39 0 6.8568315591368303e-05
GC_7_40 b_7 NI_7 NS_40 0 2.0889738559959499e-04
GC_7_41 b_7 NI_7 NS_41 0 1.4083727125750865e-05
GC_7_42 b_7 NI_7 NS_42 0 -2.8696275950915213e-05
GC_7_43 b_7 NI_7 NS_43 0 -3.8665155973581525e-06
GC_7_44 b_7 NI_7 NS_44 0 -1.4059424596533844e-06
GC_7_45 b_7 NI_7 NS_45 0 2.2948301871686332e-02
GC_7_46 b_7 NI_7 NS_46 0 -5.3842917103620158e-04
GC_7_47 b_7 NI_7 NS_47 0 -6.7369915218261729e-03
GC_7_48 b_7 NI_7 NS_48 0 8.1863869839340145e-03
GC_7_49 b_7 NI_7 NS_49 0 -3.3877637453861810e-03
GC_7_50 b_7 NI_7 NS_50 0 -9.1189585495070301e-03
GC_7_51 b_7 NI_7 NS_51 0 6.4574413697185392e-03
GC_7_52 b_7 NI_7 NS_52 0 4.8890777964331845e-04
GC_7_53 b_7 NI_7 NS_53 0 -2.0439170955069796e-03
GC_7_54 b_7 NI_7 NS_54 0 9.0199755405259024e-04
GC_7_55 b_7 NI_7 NS_55 0 -8.2736238464650967e-03
GC_7_56 b_7 NI_7 NS_56 0 2.9338873651041163e-03
GC_7_57 b_7 NI_7 NS_57 0 -1.5612575571939116e-04
GC_7_58 b_7 NI_7 NS_58 0 1.1334855413051254e-04
GC_7_59 b_7 NI_7 NS_59 0 1.0636730255068730e-04
GC_7_60 b_7 NI_7 NS_60 0 6.6658769272087909e-05
GC_7_61 b_7 NI_7 NS_61 0 -6.2653489999532004e-06
GC_7_62 b_7 NI_7 NS_62 0 3.6242976869933858e-05
GC_7_63 b_7 NI_7 NS_63 0 -1.0501946086996858e-05
GC_7_64 b_7 NI_7 NS_64 0 2.5674300525146586e-05
GC_7_65 b_7 NI_7 NS_65 0 -3.6817673478052690e-06
GC_7_66 b_7 NI_7 NS_66 0 4.3958088448507614e-05
GC_7_67 b_7 NI_7 NS_67 0 3.8785826680582748e-06
GC_7_68 b_7 NI_7 NS_68 0 2.6611844246673614e-06
GC_7_69 b_7 NI_7 NS_69 0 1.1590208880779983e-03
GC_7_70 b_7 NI_7 NS_70 0 -3.2210073781254100e-03
GC_7_71 b_7 NI_7 NS_71 0 2.6143654296192958e-04
GC_7_72 b_7 NI_7 NS_72 0 1.2121985100628588e-03
GC_7_73 b_7 NI_7 NS_73 0 2.3177105225123708e-04
GC_7_74 b_7 NI_7 NS_74 0 -3.1244705689381251e-04
GC_7_75 b_7 NI_7 NS_75 0 1.5929202578425777e-06
GC_7_76 b_7 NI_7 NS_76 0 -1.1741403603291267e-06
GC_7_77 b_7 NI_7 NS_77 0 -3.7724423031996653e-05
GC_7_78 b_7 NI_7 NS_78 0 -7.5794675055051246e-05
GC_7_79 b_7 NI_7 NS_79 0 -9.7753472713858331e-07
GC_7_80 b_7 NI_7 NS_80 0 -2.3368512417533961e-06
GC_7_81 b_7 NI_7 NS_81 0 3.3777470673606230e-08
GC_7_82 b_7 NI_7 NS_82 0 -4.4193393432701792e-06
GC_7_83 b_7 NI_7 NS_83 0 1.4335024226088430e-04
GC_7_84 b_7 NI_7 NS_84 0 1.0012941665611746e-04
GC_7_85 b_7 NI_7 NS_85 0 3.2113032995891171e-05
GC_7_86 b_7 NI_7 NS_86 0 3.9293842067923722e-05
GC_7_87 b_7 NI_7 NS_87 0 1.0596578986705207e-05
GC_7_88 b_7 NI_7 NS_88 0 -2.3269419541206455e-06
GC_7_89 b_7 NI_7 NS_89 0 9.9818664266441877e-03
GC_7_90 b_7 NI_7 NS_90 0 1.5045400667294004e-04
GC_7_91 b_7 NI_7 NS_91 0 1.1789443444855904e-02
GC_7_92 b_7 NI_7 NS_92 0 -5.2505934137351273e-03
GC_7_93 b_7 NI_7 NS_93 0 -1.9371351844904069e-03
GC_7_94 b_7 NI_7 NS_94 0 4.9258926213432211e-03
GC_7_95 b_7 NI_7 NS_95 0 1.2517409746386873e-02
GC_7_96 b_7 NI_7 NS_96 0 8.9652562394801003e-03
GC_7_97 b_7 NI_7 NS_97 0 -1.9239124801317552e-03
GC_7_98 b_7 NI_7 NS_98 0 -2.4865856789169616e-03
GC_7_99 b_7 NI_7 NS_99 0 -9.7661868281683269e-03
GC_7_100 b_7 NI_7 NS_100 0 8.8928008328633609e-03
GC_7_101 b_7 NI_7 NS_101 0 5.8049079826565813e-04
GC_7_102 b_7 NI_7 NS_102 0 3.7355971365066697e-04
GC_7_103 b_7 NI_7 NS_103 0 1.2603095789339287e-04
GC_7_104 b_7 NI_7 NS_104 0 2.9540492461345907e-04
GC_7_105 b_7 NI_7 NS_105 0 9.7537432970567887e-04
GC_7_106 b_7 NI_7 NS_106 0 -9.0222303389366721e-05
GC_7_107 b_7 NI_7 NS_107 0 1.9116872871044230e-04
GC_7_108 b_7 NI_7 NS_108 0 1.5172835083544222e-04
GC_7_109 b_7 NI_7 NS_109 0 1.1166578991582868e-04
GC_7_110 b_7 NI_7 NS_110 0 1.4012369637773525e-05
GC_7_111 b_7 NI_7 NS_111 0 -5.6488213994736247e-06
GC_7_112 b_7 NI_7 NS_112 0 2.2481555752384959e-06
GC_7_113 b_7 NI_7 NS_113 0 -2.0697010641678084e-02
GC_7_114 b_7 NI_7 NS_114 0 4.1956786199519384e-04
GC_7_115 b_7 NI_7 NS_115 0 1.3340586991602574e-02
GC_7_116 b_7 NI_7 NS_116 0 2.3195750793349921e-03
GC_7_117 b_7 NI_7 NS_117 0 -3.0587828970174229e-04
GC_7_118 b_7 NI_7 NS_118 0 -4.5083622758745846e-04
GC_7_119 b_7 NI_7 NS_119 0 9.6451887130816307e-07
GC_7_120 b_7 NI_7 NS_120 0 5.6514710221326497e-07
GC_7_121 b_7 NI_7 NS_121 0 9.5799145236906468e-05
GC_7_122 b_7 NI_7 NS_122 0 -6.0553483481342263e-05
GC_7_123 b_7 NI_7 NS_123 0 1.8789972871147877e-06
GC_7_124 b_7 NI_7 NS_124 0 3.9977701151812958e-07
GC_7_125 b_7 NI_7 NS_125 0 -1.2005928945909404e-06
GC_7_126 b_7 NI_7 NS_126 0 -1.9855078906194338e-06
GC_7_127 b_7 NI_7 NS_127 0 -9.4007608696025471e-06
GC_7_128 b_7 NI_7 NS_128 0 2.6929478439756947e-04
GC_7_129 b_7 NI_7 NS_129 0 -7.9152312476600635e-06
GC_7_130 b_7 NI_7 NS_130 0 -5.6596677515228468e-05
GC_7_131 b_7 NI_7 NS_131 0 -1.3865358019714742e-05
GC_7_132 b_7 NI_7 NS_132 0 -1.0496156926868893e-06
GC_7_133 b_7 NI_7 NS_133 0 1.0839454610276017e-02
GC_7_134 b_7 NI_7 NS_134 0 -5.3461293774454180e-04
GC_7_135 b_7 NI_7 NS_135 0 -1.5028118722613422e-02
GC_7_136 b_7 NI_7 NS_136 0 5.6909028619676286e-03
GC_7_137 b_7 NI_7 NS_137 0 2.7206587581655832e-03
GC_7_138 b_7 NI_7 NS_138 0 -1.1950861421298850e-02
GC_7_139 b_7 NI_7 NS_139 0 8.2375395800570895e-03
GC_7_140 b_7 NI_7 NS_140 0 6.6318010624247725e-04
GC_7_141 b_7 NI_7 NS_141 0 -3.8060551260203130e-04
GC_7_142 b_7 NI_7 NS_142 0 -2.9349273032718286e-04
GC_7_143 b_7 NI_7 NS_143 0 -6.5977941874399227e-03
GC_7_144 b_7 NI_7 NS_144 0 -3.1244351094444254e-03
GC_7_145 b_7 NI_7 NS_145 0 -2.5715150274552219e-04
GC_7_146 b_7 NI_7 NS_146 0 9.7651956192425007e-05
GC_7_147 b_7 NI_7 NS_147 0 1.6653327221130258e-04
GC_7_148 b_7 NI_7 NS_148 0 4.3650736593680145e-05
GC_7_149 b_7 NI_7 NS_149 0 4.6034031160150735e-04
GC_7_150 b_7 NI_7 NS_150 0 1.4668897178793248e-04
GC_7_151 b_7 NI_7 NS_151 0 7.0401105503574056e-06
GC_7_152 b_7 NI_7 NS_152 0 1.2265873582749694e-05
GC_7_153 b_7 NI_7 NS_153 0 2.7506507009165545e-06
GC_7_154 b_7 NI_7 NS_154 0 -9.0069109490576210e-06
GC_7_155 b_7 NI_7 NS_155 0 2.6628682629375446e-06
GC_7_156 b_7 NI_7 NS_156 0 -7.2013677696949834e-07
GC_7_157 b_7 NI_7 NS_157 0 2.0783219740401152e-03
GC_7_158 b_7 NI_7 NS_158 0 3.8165485799018014e-03
GC_7_159 b_7 NI_7 NS_159 0 5.8530761632765609e-04
GC_7_160 b_7 NI_7 NS_160 0 -2.3275328653761950e-03
GC_7_161 b_7 NI_7 NS_161 0 2.3189892290253567e-05
GC_7_162 b_7 NI_7 NS_162 0 -7.8370425884858653e-06
GC_7_163 b_7 NI_7 NS_163 0 8.2022390712440437e-07
GC_7_164 b_7 NI_7 NS_164 0 3.7928308725269573e-07
GC_7_165 b_7 NI_7 NS_165 0 1.2016034992935977e-06
GC_7_166 b_7 NI_7 NS_166 0 -7.0171390258925844e-06
GC_7_167 b_7 NI_7 NS_167 0 -4.3696738138045135e-08
GC_7_168 b_7 NI_7 NS_168 0 -2.0550641234003465e-07
GC_7_169 b_7 NI_7 NS_169 0 -1.2705087366532083e-07
GC_7_170 b_7 NI_7 NS_170 0 -1.2096128330752077e-06
GC_7_171 b_7 NI_7 NS_171 0 -6.3494731446081897e-05
GC_7_172 b_7 NI_7 NS_172 0 1.9663962922210394e-05
GC_7_173 b_7 NI_7 NS_173 0 -1.4824933676504345e-05
GC_7_174 b_7 NI_7 NS_174 0 1.9191652089814664e-05
GC_7_175 b_7 NI_7 NS_175 0 -1.1583797214201170e-07
GC_7_176 b_7 NI_7 NS_176 0 3.8801410406707268e-07
GC_7_177 b_7 NI_7 NS_177 0 5.6120539298801205e-03
GC_7_178 b_7 NI_7 NS_178 0 -5.1913700960235236e-04
GC_7_179 b_7 NI_7 NS_179 0 1.1152832382888320e-02
GC_7_180 b_7 NI_7 NS_180 0 3.3286876797509503e-03
GC_7_181 b_7 NI_7 NS_181 0 -8.8802452741731930e-03
GC_7_182 b_7 NI_7 NS_182 0 -8.9204509768649898e-03
GC_7_183 b_7 NI_7 NS_183 0 1.1593344810249741e-02
GC_7_184 b_7 NI_7 NS_184 0 6.5240857665463071e-03
GC_7_185 b_7 NI_7 NS_185 0 -2.6330008472468260e-03
GC_7_186 b_7 NI_7 NS_186 0 -1.1657371882231485e-03
GC_7_187 b_7 NI_7 NS_187 0 2.8837397276921081e-03
GC_7_188 b_7 NI_7 NS_188 0 2.9234219270477938e-03
GC_7_189 b_7 NI_7 NS_189 0 5.7649672114973023e-04
GC_7_190 b_7 NI_7 NS_190 0 3.7833629962890459e-04
GC_7_191 b_7 NI_7 NS_191 0 1.2742624069930948e-04
GC_7_192 b_7 NI_7 NS_192 0 3.4203965796308770e-04
GC_7_193 b_7 NI_7 NS_193 0 7.7293193933660419e-04
GC_7_194 b_7 NI_7 NS_194 0 -6.4517690610893565e-05
GC_7_195 b_7 NI_7 NS_195 0 1.8599392982158832e-04
GC_7_196 b_7 NI_7 NS_196 0 1.6984865408423863e-04
GC_7_197 b_7 NI_7 NS_197 0 8.7402876868479317e-05
GC_7_198 b_7 NI_7 NS_198 0 3.6761398473650177e-05
GC_7_199 b_7 NI_7 NS_199 0 -8.5234104693607557e-06
GC_7_200 b_7 NI_7 NS_200 0 1.9060167792779641e-06
GC_7_201 b_7 NI_7 NS_201 0 -1.7137304426197857e-02
GC_7_202 b_7 NI_7 NS_202 0 9.6737302919323778e-03
GC_7_203 b_7 NI_7 NS_203 0 1.2689828848665674e-02
GC_7_204 b_7 NI_7 NS_204 0 -1.1129100038089303e-03
GC_7_205 b_7 NI_7 NS_205 0 -4.3328715421901465e-04
GC_7_206 b_7 NI_7 NS_206 0 -2.1162014478746413e-05
GC_7_207 b_7 NI_7 NS_207 0 1.2982407320318606e-06
GC_7_208 b_7 NI_7 NS_208 0 2.8962947404359074e-06
GC_7_209 b_7 NI_7 NS_209 0 1.8336278332959665e-04
GC_7_210 b_7 NI_7 NS_210 0 -2.1362352079684109e-05
GC_7_211 b_7 NI_7 NS_211 0 4.3755483143903149e-06
GC_7_212 b_7 NI_7 NS_212 0 1.0716257489376100e-06
GC_7_213 b_7 NI_7 NS_213 0 -4.9215837093277624e-09
GC_7_214 b_7 NI_7 NS_214 0 -8.4765074292317445e-08
GC_7_215 b_7 NI_7 NS_215 0 -1.8712977959643116e-04
GC_7_216 b_7 NI_7 NS_216 0 3.0580470557346127e-04
GC_7_217 b_7 NI_7 NS_217 0 -5.6725967090392505e-05
GC_7_218 b_7 NI_7 NS_218 0 -4.3286565094196980e-05
GC_7_219 b_7 NI_7 NS_219 0 -1.9141010544143624e-05
GC_7_220 b_7 NI_7 NS_220 0 5.9946355818655368e-06
GC_7_221 b_7 NI_7 NS_221 0 6.1507866043792403e-03
GC_7_222 b_7 NI_7 NS_222 0 -3.8636957924981512e-04
GC_7_223 b_7 NI_7 NS_223 0 -2.0319170926007882e-02
GC_7_224 b_7 NI_7 NS_224 0 -2.9799757317896642e-03
GC_7_225 b_7 NI_7 NS_225 0 1.0030808512126590e-02
GC_7_226 b_7 NI_7 NS_226 0 -3.4804738917824695e-03
GC_7_227 b_7 NI_7 NS_227 0 6.1236368894885627e-03
GC_7_228 b_7 NI_7 NS_228 0 6.4978683405443529e-04
GC_7_229 b_7 NI_7 NS_229 0 1.4531255133561139e-03
GC_7_230 b_7 NI_7 NS_230 0 -2.7388354097941564e-05
GC_7_231 b_7 NI_7 NS_231 0 -2.7195649467214261e-04
GC_7_232 b_7 NI_7 NS_232 0 -8.8213910496511335e-03
GC_7_233 b_7 NI_7 NS_233 0 -2.6856746714931353e-04
GC_7_234 b_7 NI_7 NS_234 0 1.0823191844144467e-04
GC_7_235 b_7 NI_7 NS_235 0 2.1792848461543450e-04
GC_7_236 b_7 NI_7 NS_236 0 3.8412687463670989e-05
GC_7_237 b_7 NI_7 NS_237 0 4.6922798432003744e-04
GC_7_238 b_7 NI_7 NS_238 0 4.1093464334346423e-04
GC_7_239 b_7 NI_7 NS_239 0 4.0985501595735408e-05
GC_7_240 b_7 NI_7 NS_240 0 2.7208120908488229e-05
GC_7_241 b_7 NI_7 NS_241 0 8.3515005409951908e-05
GC_7_242 b_7 NI_7 NS_242 0 -1.9874247028491422e-05
GC_7_243 b_7 NI_7 NS_243 0 7.8069488171795804e-06
GC_7_244 b_7 NI_7 NS_244 0 -9.9686667967906915e-07
GC_7_245 b_7 NI_7 NS_245 0 -4.8530597783247916e-03
GC_7_246 b_7 NI_7 NS_246 0 9.8910022813491899e-03
GC_7_247 b_7 NI_7 NS_247 0 3.9529174469917954e-03
GC_7_248 b_7 NI_7 NS_248 0 -4.3989992597534139e-03
GC_7_249 b_7 NI_7 NS_249 0 -2.4430289335984921e-04
GC_7_250 b_7 NI_7 NS_250 0 1.4055318610138758e-04
GC_7_251 b_7 NI_7 NS_251 0 -5.4456124827019449e-07
GC_7_252 b_7 NI_7 NS_252 0 2.8277985714432378e-07
GC_7_253 b_7 NI_7 NS_253 0 -1.4539573798105399e-05
GC_7_254 b_7 NI_7 NS_254 0 5.5277592759103648e-05
GC_7_255 b_7 NI_7 NS_255 0 -8.6591885968278199e-07
GC_7_256 b_7 NI_7 NS_256 0 7.3752165611013496e-07
GC_7_257 b_7 NI_7 NS_257 0 -2.6196530735269443e-06
GC_7_258 b_7 NI_7 NS_258 0 -1.0301308436845626e-06
GC_7_259 b_7 NI_7 NS_259 0 -7.4525893843725770e-05
GC_7_260 b_7 NI_7 NS_260 0 -1.2986853872837061e-04
GC_7_261 b_7 NI_7 NS_261 0 -1.9115744390433140e-05
GC_7_262 b_7 NI_7 NS_262 0 -3.2863758292807561e-05
GC_7_263 b_7 NI_7 NS_263 0 -8.2088450398899763e-06
GC_7_264 b_7 NI_7 NS_264 0 -8.3685220571518301e-06
GC_7_265 b_7 NI_7 NS_265 0 -2.1602519232088883e-02
GC_7_266 b_7 NI_7 NS_266 0 1.3450284115624015e-02
GC_7_267 b_7 NI_7 NS_267 0 4.5213974835390872e-03
GC_7_268 b_7 NI_7 NS_268 0 9.9845169218586872e-03
GC_7_269 b_7 NI_7 NS_269 0 1.6504881593702905e-02
GC_7_270 b_7 NI_7 NS_270 0 -8.9076456318253807e-03
GC_7_271 b_7 NI_7 NS_271 0 5.1437313985785429e-03
GC_7_272 b_7 NI_7 NS_272 0 4.9917189533298899e-03
GC_7_273 b_7 NI_7 NS_273 0 3.3299237405692672e-03
GC_7_274 b_7 NI_7 NS_274 0 4.9943587138322754e-03
GC_7_275 b_7 NI_7 NS_275 0 8.2456656336360838e-03
GC_7_276 b_7 NI_7 NS_276 0 9.5938733082247939e-03
GC_7_277 b_7 NI_7 NS_277 0 3.1638786678116779e-04
GC_7_278 b_7 NI_7 NS_278 0 1.3137167946175796e-04
GC_7_279 b_7 NI_7 NS_279 0 3.5352738176703889e-05
GC_7_280 b_7 NI_7 NS_280 0 2.1097945156722933e-04
GC_7_281 b_7 NI_7 NS_281 0 7.0665597197846119e-04
GC_7_282 b_7 NI_7 NS_282 0 -8.6798196063591292e-04
GC_7_283 b_7 NI_7 NS_283 0 1.2721744269849521e-04
GC_7_284 b_7 NI_7 NS_284 0 6.2231104705610401e-05
GC_7_285 b_7 NI_7 NS_285 0 -8.6570783323473488e-05
GC_7_286 b_7 NI_7 NS_286 0 -8.0591538657770841e-05
GC_7_287 b_7 NI_7 NS_287 0 -8.7153464715979010e-06
GC_7_288 b_7 NI_7 NS_288 0 -1.2768305406428142e-06
GC_7_289 b_7 NI_7 NS_289 0 -1.6026866910917573e-04
GC_7_290 b_7 NI_7 NS_290 0 8.0028415214623318e-03
GC_7_291 b_7 NI_7 NS_291 0 3.2473658389351075e-03
GC_7_292 b_7 NI_7 NS_292 0 -3.1806934000808340e-03
GC_7_293 b_7 NI_7 NS_293 0 -5.0611492434595232e-04
GC_7_294 b_7 NI_7 NS_294 0 6.2773493246689170e-04
GC_7_295 b_7 NI_7 NS_295 0 1.5543907021554829e-06
GC_7_296 b_7 NI_7 NS_296 0 5.2760529937149520e-06
GC_7_297 b_7 NI_7 NS_297 0 2.4274906913631755e-04
GC_7_298 b_7 NI_7 NS_298 0 3.4333801547874384e-05
GC_7_299 b_7 NI_7 NS_299 0 5.4104274580105856e-06
GC_7_300 b_7 NI_7 NS_300 0 1.8636667407238327e-06
GC_7_301 b_7 NI_7 NS_301 0 3.4346222965024605e-06
GC_7_302 b_7 NI_7 NS_302 0 2.4007915336259832e-06
GC_7_303 b_7 NI_7 NS_303 0 -3.4068753547243370e-04
GC_7_304 b_7 NI_7 NS_304 0 3.6175323734042957e-04
GC_7_305 b_7 NI_7 NS_305 0 -1.2101566845695395e-04
GC_7_306 b_7 NI_7 NS_306 0 -1.4533218288905470e-05
GC_7_307 b_7 NI_7 NS_307 0 -2.4865382143977588e-05
GC_7_308 b_7 NI_7 NS_308 0 1.6970170295165842e-05
GC_7_309 b_7 NI_7 NS_309 0 3.0345586105208548e-02
GC_7_310 b_7 NI_7 NS_310 0 1.6567569493163934e-02
GC_7_311 b_7 NI_7 NS_311 0 -1.9639967248424497e-02
GC_7_312 b_7 NI_7 NS_312 0 -6.0010372913804656e-03
GC_7_313 b_7 NI_7 NS_313 0 -2.7653552805386686e-02
GC_7_314 b_7 NI_7 NS_314 0 1.3586390375302741e-03
GC_7_315 b_7 NI_7 NS_315 0 2.3949683403563043e-03
GC_7_316 b_7 NI_7 NS_316 0 1.7316508049602672e-03
GC_7_317 b_7 NI_7 NS_317 0 -1.1942220505414851e-03
GC_7_318 b_7 NI_7 NS_318 0 1.1387796392580997e-03
GC_7_319 b_7 NI_7 NS_319 0 7.9306211588074018e-03
GC_7_320 b_7 NI_7 NS_320 0 -3.8432297545315406e-03
GC_7_321 b_7 NI_7 NS_321 0 -3.1739138430673990e-04
GC_7_322 b_7 NI_7 NS_322 0 5.2908898973899223e-05
GC_7_323 b_7 NI_7 NS_323 0 6.2981587277220912e-05
GC_7_324 b_7 NI_7 NS_324 0 2.0929374550275529e-05
GC_7_325 b_7 NI_7 NS_325 0 1.1905110525430607e-04
GC_7_326 b_7 NI_7 NS_326 0 -4.4050925313760984e-04
GC_7_327 b_7 NI_7 NS_327 0 -4.1805576190874964e-05
GC_7_328 b_7 NI_7 NS_328 0 2.9251233708072179e-07
GC_7_329 b_7 NI_7 NS_329 0 -7.5658259999060164e-05
GC_7_330 b_7 NI_7 NS_330 0 1.8702338408319648e-05
GC_7_331 b_7 NI_7 NS_331 0 4.2147443018672270e-07
GC_7_332 b_7 NI_7 NS_332 0 2.9364603803254640e-06
GC_7_333 b_7 NI_7 NS_333 0 4.0311006347029530e-04
GC_7_334 b_7 NI_7 NS_334 0 -7.8347510415009286e-03
GC_7_335 b_7 NI_7 NS_335 0 -9.5602287718762663e-04
GC_7_336 b_7 NI_7 NS_336 0 2.8189952421668659e-03
GC_7_337 b_7 NI_7 NS_337 0 2.3608923416160269e-04
GC_7_338 b_7 NI_7 NS_338 0 1.5679284374402896e-04
GC_7_339 b_7 NI_7 NS_339 0 2.3456923981426361e-06
GC_7_340 b_7 NI_7 NS_340 0 4.8623968856849969e-07
GC_7_341 b_7 NI_7 NS_341 0 3.9457072116086471e-05
GC_7_342 b_7 NI_7 NS_342 0 -6.2485811107831801e-05
GC_7_343 b_7 NI_7 NS_343 0 8.0395806572731593e-07
GC_7_344 b_7 NI_7 NS_344 0 -1.8006287311656177e-06
GC_7_345 b_7 NI_7 NS_345 0 1.6862245916863339e-06
GC_7_346 b_7 NI_7 NS_346 0 -3.8933125274131063e-06
GC_7_347 b_7 NI_7 NS_347 0 7.2647524476736154e-05
GC_7_348 b_7 NI_7 NS_348 0 1.7115084872874105e-04
GC_7_349 b_7 NI_7 NS_349 0 3.7180883435760076e-06
GC_7_350 b_7 NI_7 NS_350 0 5.2362870108039585e-05
GC_7_351 b_7 NI_7 NS_351 0 1.0282566081291398e-05
GC_7_352 b_7 NI_7 NS_352 0 5.5513726852957736e-06
GC_7_353 b_7 NI_7 NS_353 0 -7.2175652553153457e-03
GC_7_354 b_7 NI_7 NS_354 0 4.0551398261866308e-05
GC_7_355 b_7 NI_7 NS_355 0 1.9335304825858302e-03
GC_7_356 b_7 NI_7 NS_356 0 -1.5459930291885917e-03
GC_7_357 b_7 NI_7 NS_357 0 -1.1753708115920254e-03
GC_7_358 b_7 NI_7 NS_358 0 7.1462146040561026e-04
GC_7_359 b_7 NI_7 NS_359 0 2.4739555043350680e-03
GC_7_360 b_7 NI_7 NS_360 0 -3.4029816455579877e-05
GC_7_361 b_7 NI_7 NS_361 0 1.7508903810365881e-04
GC_7_362 b_7 NI_7 NS_362 0 7.1212522549260709e-04
GC_7_363 b_7 NI_7 NS_363 0 -3.3745137326394144e-03
GC_7_364 b_7 NI_7 NS_364 0 1.8943511562715271e-04
GC_7_365 b_7 NI_7 NS_365 0 4.2453574892510582e-04
GC_7_366 b_7 NI_7 NS_366 0 -1.7728940836727274e-04
GC_7_367 b_7 NI_7 NS_367 0 2.9733426805896349e-04
GC_7_368 b_7 NI_7 NS_368 0 6.0884568735112209e-04
GC_7_369 b_7 NI_7 NS_369 0 -1.5840679109543775e-03
GC_7_370 b_7 NI_7 NS_370 0 -1.4372871478060545e-03
GC_7_371 b_7 NI_7 NS_371 0 1.7043351425808319e-04
GC_7_372 b_7 NI_7 NS_372 0 1.2501332664887615e-04
GC_7_373 b_7 NI_7 NS_373 0 -6.6702467860379545e-04
GC_7_374 b_7 NI_7 NS_374 0 1.0739770262914510e-05
GC_7_375 b_7 NI_7 NS_375 0 -4.0231684304563813e-06
GC_7_376 b_7 NI_7 NS_376 0 -1.6768706567850990e-06
GC_7_377 b_7 NI_7 NS_377 0 8.8095447149813527e-03
GC_7_378 b_7 NI_7 NS_378 0 5.1660340645631672e-03
GC_7_379 b_7 NI_7 NS_379 0 -3.5560662962972503e-03
GC_7_380 b_7 NI_7 NS_380 0 -6.8177765225508396e-03
GC_7_381 b_7 NI_7 NS_381 0 -1.1657069007169432e-04
GC_7_382 b_7 NI_7 NS_382 0 3.0218388354222498e-04
GC_7_383 b_7 NI_7 NS_383 0 2.3041144711677235e-07
GC_7_384 b_7 NI_7 NS_384 0 -1.6325642329087899e-07
GC_7_385 b_7 NI_7 NS_385 0 1.4629907354362692e-06
GC_7_386 b_7 NI_7 NS_386 0 -7.9883577184207825e-05
GC_7_387 b_7 NI_7 NS_387 0 2.0985313971449682e-07
GC_7_388 b_7 NI_7 NS_388 0 3.0768800827040934e-07
GC_7_389 b_7 NI_7 NS_389 0 4.4105782110316373e-09
GC_7_390 b_7 NI_7 NS_390 0 -2.3463716035643938e-06
GC_7_391 b_7 NI_7 NS_391 0 1.5601311942709168e-04
GC_7_392 b_7 NI_7 NS_392 0 4.4744746847381325e-04
GC_7_393 b_7 NI_7 NS_393 0 -1.4084514213392416e-04
GC_7_394 b_7 NI_7 NS_394 0 6.0917700401389494e-05
GC_7_395 b_7 NI_7 NS_395 0 -1.5053221307123436e-05
GC_7_396 b_7 NI_7 NS_396 0 -5.8659903067951298e-06
GC_7_397 b_7 NI_7 NS_397 0 -4.1691162356828635e-03
GC_7_398 b_7 NI_7 NS_398 0 -9.7800668995874586e-05
GC_7_399 b_7 NI_7 NS_399 0 -3.4354452474854558e-03
GC_7_400 b_7 NI_7 NS_400 0 2.1023028694434390e-03
GC_7_401 b_7 NI_7 NS_401 0 -6.1026594135366562e-04
GC_7_402 b_7 NI_7 NS_402 0 -4.1004274608966770e-03
GC_7_403 b_7 NI_7 NS_403 0 1.4299878031195793e-03
GC_7_404 b_7 NI_7 NS_404 0 -1.2193512336292239e-03
GC_7_405 b_7 NI_7 NS_405 0 1.8072629887217446e-04
GC_7_406 b_7 NI_7 NS_406 0 -1.1251587944797828e-04
GC_7_407 b_7 NI_7 NS_407 0 -1.0116146447004298e-03
GC_7_408 b_7 NI_7 NS_408 0 -2.7587722375132457e-03
GC_7_409 b_7 NI_7 NS_409 0 -1.0898185725681590e-04
GC_7_410 b_7 NI_7 NS_410 0 2.2108096524690518e-04
GC_7_411 b_7 NI_7 NS_411 0 1.9213213396477015e-04
GC_7_412 b_7 NI_7 NS_412 0 -6.8711855591089161e-05
GC_7_413 b_7 NI_7 NS_413 0 -7.1607713068507284e-05
GC_7_414 b_7 NI_7 NS_414 0 -1.3686210968904571e-04
GC_7_415 b_7 NI_7 NS_415 0 -1.4114852819097489e-05
GC_7_416 b_7 NI_7 NS_416 0 -1.8759714010636929e-05
GC_7_417 b_7 NI_7 NS_417 0 -4.4744377829930175e-05
GC_7_418 b_7 NI_7 NS_418 0 -6.3879350909429975e-05
GC_7_419 b_7 NI_7 NS_419 0 3.7420373355060911e-06
GC_7_420 b_7 NI_7 NS_420 0 1.5699117063441888e-06
GC_7_421 b_7 NI_7 NS_421 0 5.9046279963274025e-03
GC_7_422 b_7 NI_7 NS_422 0 2.4577989257401024e-03
GC_7_423 b_7 NI_7 NS_423 0 -2.8030277647965551e-03
GC_7_424 b_7 NI_7 NS_424 0 -2.2213267320967340e-03
GC_7_425 b_7 NI_7 NS_425 0 5.2446601353769073e-05
GC_7_426 b_7 NI_7 NS_426 0 1.7578252686970225e-04
GC_7_427 b_7 NI_7 NS_427 0 2.4034225822430473e-07
GC_7_428 b_7 NI_7 NS_428 0 7.0788341607000972e-07
GC_7_429 b_7 NI_7 NS_429 0 4.6067688707350933e-05
GC_7_430 b_7 NI_7 NS_430 0 2.2851957796723199e-06
GC_7_431 b_7 NI_7 NS_431 0 1.3018957438942227e-06
GC_7_432 b_7 NI_7 NS_432 0 -2.1707885484549564e-07
GC_7_433 b_7 NI_7 NS_433 0 -6.8041437939121576e-07
GC_7_434 b_7 NI_7 NS_434 0 -1.3565379716990915e-06
GC_7_435 b_7 NI_7 NS_435 0 -9.4749806933040878e-05
GC_7_436 b_7 NI_7 NS_436 0 2.8698039083336433e-05
GC_7_437 b_7 NI_7 NS_437 0 -3.4791055667476555e-05
GC_7_438 b_7 NI_7 NS_438 0 -8.7737187500790502e-06
GC_7_439 b_7 NI_7 NS_439 0 3.3053766214632694e-06
GC_7_440 b_7 NI_7 NS_440 0 5.5863110921134382e-06
GC_7_441 b_7 NI_7 NS_441 0 -6.0603592032650736e-03
GC_7_442 b_7 NI_7 NS_442 0 -2.1312935981613655e-04
GC_7_443 b_7 NI_7 NS_443 0 2.4418368838900390e-03
GC_7_444 b_7 NI_7 NS_444 0 1.7985969645022747e-03
GC_7_445 b_7 NI_7 NS_445 0 -3.8803098350916050e-03
GC_7_446 b_7 NI_7 NS_446 0 -4.1123799700742781e-03
GC_7_447 b_7 NI_7 NS_447 0 2.4221469032116145e-03
GC_7_448 b_7 NI_7 NS_448 0 3.6138305580558851e-04
GC_7_449 b_7 NI_7 NS_449 0 1.4371147985468448e-04
GC_7_450 b_7 NI_7 NS_450 0 -4.4032904818858045e-04
GC_7_451 b_7 NI_7 NS_451 0 8.5390369759869304e-04
GC_7_452 b_7 NI_7 NS_452 0 -1.4662076137502908e-03
GC_7_453 b_7 NI_7 NS_453 0 2.9759000795817354e-04
GC_7_454 b_7 NI_7 NS_454 0 -5.8796034275011747e-05
GC_7_455 b_7 NI_7 NS_455 0 2.1005013221669154e-04
GC_7_456 b_7 NI_7 NS_456 0 4.4514685835448406e-04
GC_7_457 b_7 NI_7 NS_457 0 -1.0977214127254359e-03
GC_7_458 b_7 NI_7 NS_458 0 -9.2864250975412403e-04
GC_7_459 b_7 NI_7 NS_459 0 1.3465509120811451e-04
GC_7_460 b_7 NI_7 NS_460 0 9.7802956017741476e-05
GC_7_461 b_7 NI_7 NS_461 0 -4.4566627387797401e-04
GC_7_462 b_7 NI_7 NS_462 0 5.5649764901145122e-06
GC_7_463 b_7 NI_7 NS_463 0 -8.0918160373482278e-07
GC_7_464 b_7 NI_7 NS_464 0 -5.0393010720756553e-07
GC_7_465 b_7 NI_7 NS_465 0 4.1119240075792119e-03
GC_7_466 b_7 NI_7 NS_466 0 6.8603493682723770e-03
GC_7_467 b_7 NI_7 NS_467 0 -7.2764908892527526e-04
GC_7_468 b_7 NI_7 NS_468 0 -5.7931892338286082e-03
GC_7_469 b_7 NI_7 NS_469 0 -3.5775308651607012e-04
GC_7_470 b_7 NI_7 NS_470 0 3.8834911402994523e-04
GC_7_471 b_7 NI_7 NS_471 0 9.4512421664228531e-08
GC_7_472 b_7 NI_7 NS_472 0 4.5738255391481510e-07
GC_7_473 b_7 NI_7 NS_473 0 2.6844694184315749e-05
GC_7_474 b_7 NI_7 NS_474 0 -2.2194802683348891e-05
GC_7_475 b_7 NI_7 NS_475 0 3.3931998008711181e-07
GC_7_476 b_7 NI_7 NS_476 0 6.9561053447600165e-07
GC_7_477 b_7 NI_7 NS_477 0 -1.4718253902633587e-06
GC_7_478 b_7 NI_7 NS_478 0 -9.8770241655271839e-07
GC_7_479 b_7 NI_7 NS_479 0 5.9106733586471631e-05
GC_7_480 b_7 NI_7 NS_480 0 2.3858333840164690e-04
GC_7_481 b_7 NI_7 NS_481 0 -1.0408464158216801e-04
GC_7_482 b_7 NI_7 NS_482 0 2.0899988973949210e-05
GC_7_483 b_7 NI_7 NS_483 0 -1.4386399320208944e-05
GC_7_484 b_7 NI_7 NS_484 0 -5.7818104663803490e-06
GC_7_485 b_7 NI_7 NS_485 0 -9.2404038201695615e-04
GC_7_486 b_7 NI_7 NS_486 0 -1.0486435411964030e-04
GC_7_487 b_7 NI_7 NS_487 0 -5.6890150266187545e-03
GC_7_488 b_7 NI_7 NS_488 0 -9.2937909862438333e-04
GC_7_489 b_7 NI_7 NS_489 0 2.1856550581691152e-03
GC_7_490 b_7 NI_7 NS_490 0 -4.4645526662866756e-04
GC_7_491 b_7 NI_7 NS_491 0 6.7367416259125218e-04
GC_7_492 b_7 NI_7 NS_492 0 -4.8131725161458180e-04
GC_7_493 b_7 NI_7 NS_493 0 8.9750050241973784e-04
GC_7_494 b_7 NI_7 NS_494 0 2.8166329620972540e-04
GC_7_495 b_7 NI_7 NS_495 0 6.2080685063446283e-04
GC_7_496 b_7 NI_7 NS_496 0 -4.4931037199533964e-03
GC_7_497 b_7 NI_7 NS_497 0 -1.3699452358760801e-04
GC_7_498 b_7 NI_7 NS_498 0 1.5172652148976633e-04
GC_7_499 b_7 NI_7 NS_499 0 1.5212355527495600e-04
GC_7_500 b_7 NI_7 NS_500 0 -2.6260463575138233e-05
GC_7_501 b_7 NI_7 NS_501 0 -8.1269803623868552e-05
GC_7_502 b_7 NI_7 NS_502 0 -4.0289757989831376e-05
GC_7_503 b_7 NI_7 NS_503 0 -1.9383966378427764e-05
GC_7_504 b_7 NI_7 NS_504 0 -1.0425340580950845e-05
GC_7_505 b_7 NI_7 NS_505 0 -1.8592434584840259e-05
GC_7_506 b_7 NI_7 NS_506 0 -2.7443285999571829e-05
GC_7_507 b_7 NI_7 NS_507 0 1.9958229821025246e-06
GC_7_508 b_7 NI_7 NS_508 0 5.3636260682803701e-07
GC_7_509 b_7 NI_7 NS_509 0 1.6574361944100210e-03
GC_7_510 b_7 NI_7 NS_510 0 3.0647333810401079e-03
GC_7_511 b_7 NI_7 NS_511 0 -7.7998852790826627e-04
GC_7_512 b_7 NI_7 NS_512 0 -1.7043265536214542e-03
GC_7_513 b_7 NI_7 NS_513 0 4.4861243954079224e-05
GC_7_514 b_7 NI_7 NS_514 0 1.9006420059172480e-04
GC_7_515 b_7 NI_7 NS_515 0 3.0979022679617841e-07
GC_7_516 b_7 NI_7 NS_516 0 4.1163530681843359e-07
GC_7_517 b_7 NI_7 NS_517 0 3.9532654428783232e-05
GC_7_518 b_7 NI_7 NS_518 0 1.3984380737778746e-06
GC_7_519 b_7 NI_7 NS_519 0 6.6950162699657955e-07
GC_7_520 b_7 NI_7 NS_520 0 2.0641674768822462e-07
GC_7_521 b_7 NI_7 NS_521 0 -4.6822464253848722e-07
GC_7_522 b_7 NI_7 NS_522 0 -8.9954844251352801e-07
GC_7_523 b_7 NI_7 NS_523 0 -7.3574673989483037e-05
GC_7_524 b_7 NI_7 NS_524 0 -2.1184629916424105e-05
GC_7_525 b_7 NI_7 NS_525 0 -1.2509487085659746e-05
GC_7_526 b_7 NI_7 NS_526 0 -7.5098806214601919e-06
GC_7_527 b_7 NI_7 NS_527 0 2.2524736632329221e-06
GC_7_528 b_7 NI_7 NS_528 0 2.4634424021404142e-06
GD_7_1 b_7 NI_7 NA_1 0 -9.0786133963409038e-03
GD_7_2 b_7 NI_7 NA_2 0 -1.1073250957336118e-02
GD_7_3 b_7 NI_7 NA_3 0 -2.0609250360904677e-02
GD_7_4 b_7 NI_7 NA_4 0 -2.6662571492135595e-03
GD_7_5 b_7 NI_7 NA_5 0 -2.1416087166440473e-02
GD_7_6 b_7 NI_7 NA_6 0 -3.6884604259526214e-03
GD_7_7 b_7 NI_7 NA_7 0 -1.6672114161107437e-01
GD_7_8 b_7 NI_7 NA_8 0 -9.1138840882758511e-03
GD_7_9 b_7 NI_7 NA_9 0 3.1710214399040468e-03
GD_7_10 b_7 NI_7 NA_10 0 5.7785659537107261e-03
GD_7_11 b_7 NI_7 NA_11 0 1.5364429252738832e-03
GD_7_12 b_7 NI_7 NA_12 0 1.4691786521526401e-03
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 2.2701383137622825e-02
GC_8_2 b_8 NI_8 NS_2 0 -5.3164488024111151e-04
GC_8_3 b_8 NI_8 NS_3 0 -6.5503786045687396e-03
GC_8_4 b_8 NI_8 NS_4 0 8.2362773686255122e-03
GC_8_5 b_8 NI_8 NS_5 0 -3.6090198409855540e-03
GC_8_6 b_8 NI_8 NS_6 0 -8.8590221970597204e-03
GC_8_7 b_8 NI_8 NS_7 0 6.1402281782453084e-03
GC_8_8 b_8 NI_8 NS_8 0 4.8129312488712000e-04
GC_8_9 b_8 NI_8 NS_9 0 -1.6902783599212967e-03
GC_8_10 b_8 NI_8 NS_10 0 4.3909960251882707e-04
GC_8_11 b_8 NI_8 NS_11 0 -8.2254729575556504e-03
GC_8_12 b_8 NI_8 NS_12 0 2.8484432460404853e-03
GC_8_13 b_8 NI_8 NS_13 0 -1.6753675302615524e-04
GC_8_14 b_8 NI_8 NS_14 0 1.1463757082214324e-04
GC_8_15 b_8 NI_8 NS_15 0 1.0497005236746672e-04
GC_8_16 b_8 NI_8 NS_16 0 7.3248079189796201e-05
GC_8_17 b_8 NI_8 NS_17 0 4.3404098279567406e-05
GC_8_18 b_8 NI_8 NS_18 0 5.1326448043586284e-05
GC_8_19 b_8 NI_8 NS_19 0 -1.3610507749505152e-05
GC_8_20 b_8 NI_8 NS_20 0 2.9465331777734755e-05
GC_8_21 b_8 NI_8 NS_21 0 -7.8793111362592605e-06
GC_8_22 b_8 NI_8 NS_22 0 4.3639231677379382e-05
GC_8_23 b_8 NI_8 NS_23 0 3.3150395654177417e-06
GC_8_24 b_8 NI_8 NS_24 0 2.7916137086861482e-06
GC_8_25 b_8 NI_8 NS_25 0 -2.6241609617897973e-04
GC_8_26 b_8 NI_8 NS_26 0 -3.6640709710942811e-03
GC_8_27 b_8 NI_8 NS_27 0 1.0167936237770875e-03
GC_8_28 b_8 NI_8 NS_28 0 1.5016845663472780e-03
GC_8_29 b_8 NI_8 NS_29 0 2.3407575291108483e-04
GC_8_30 b_8 NI_8 NS_30 0 -3.3545074027530448e-04
GC_8_31 b_8 NI_8 NS_31 0 1.2063665016274481e-06
GC_8_32 b_8 NI_8 NS_32 0 -1.5445557228348959e-06
GC_8_33 b_8 NI_8 NS_33 0 -3.7386760437213833e-05
GC_8_34 b_8 NI_8 NS_34 0 -8.1394976865917733e-05
GC_8_35 b_8 NI_8 NS_35 0 -5.8536822360965341e-07
GC_8_36 b_8 NI_8 NS_36 0 -2.1526513364171568e-06
GC_8_37 b_8 NI_8 NS_37 0 2.0405916681523366e-06
GC_8_38 b_8 NI_8 NS_38 0 -2.6188172796597336e-06
GC_8_39 b_8 NI_8 NS_39 0 1.4986989963964995e-04
GC_8_40 b_8 NI_8 NS_40 0 9.1312796745943902e-05
GC_8_41 b_8 NI_8 NS_41 0 4.3196311353054962e-05
GC_8_42 b_8 NI_8 NS_42 0 4.3611220708049120e-05
GC_8_43 b_8 NI_8 NS_43 0 1.5167024618446862e-05
GC_8_44 b_8 NI_8 NS_44 0 -9.5060022860345182e-07
GC_8_45 b_8 NI_8 NS_45 0 -1.3893730258818465e-02
GC_8_46 b_8 NI_8 NS_46 0 2.9026102260310259e-04
GC_8_47 b_8 NI_8 NS_47 0 4.8228597249884431e-03
GC_8_48 b_8 NI_8 NS_48 0 -9.7669134193472170e-03
GC_8_49 b_8 NI_8 NS_49 0 5.6062432698940519e-03
GC_8_50 b_8 NI_8 NS_50 0 6.9731523325501097e-03
GC_8_51 b_8 NI_8 NS_51 0 5.5234001046188955e-03
GC_8_52 b_8 NI_8 NS_52 0 7.3380258070906762e-04
GC_8_53 b_8 NI_8 NS_53 0 -1.9106744232109095e-03
GC_8_54 b_8 NI_8 NS_54 0 -1.1727547925268944e-03
GC_8_55 b_8 NI_8 NS_55 0 -8.2268498478375938e-04
GC_8_56 b_8 NI_8 NS_56 0 7.3480383871382888e-03
GC_8_57 b_8 NI_8 NS_57 0 6.9575961953815266e-05
GC_8_58 b_8 NI_8 NS_58 0 -9.5434784510311729e-05
GC_8_59 b_8 NI_8 NS_59 0 1.4706061031806736e-06
GC_8_60 b_8 NI_8 NS_60 0 -1.4718974485807896e-05
GC_8_61 b_8 NI_8 NS_61 0 -8.5476036403115812e-05
GC_8_62 b_8 NI_8 NS_62 0 -8.9163477564232558e-05
GC_8_63 b_8 NI_8 NS_63 0 1.1463293347009888e-06
GC_8_64 b_8 NI_8 NS_64 0 4.7508347406071326e-06
GC_8_65 b_8 NI_8 NS_65 0 3.0264435367831983e-06
GC_8_66 b_8 NI_8 NS_66 0 1.6333030724762291e-05
GC_8_67 b_8 NI_8 NS_67 0 -1.2945820052232606e-06
GC_8_68 b_8 NI_8 NS_68 0 3.6536968317834730e-07
GC_8_69 b_8 NI_8 NS_69 0 -1.3192198976317625e-03
GC_8_70 b_8 NI_8 NS_70 0 3.4185839203156013e-03
GC_8_71 b_8 NI_8 NS_71 0 3.4934756350931030e-04
GC_8_72 b_8 NI_8 NS_72 0 -1.0911559514152076e-03
GC_8_73 b_8 NI_8 NS_73 0 -1.5710296991541535e-04
GC_8_74 b_8 NI_8 NS_74 0 -1.2483946531983051e-04
GC_8_75 b_8 NI_8 NS_75 0 -2.9558702803357790e-07
GC_8_76 b_8 NI_8 NS_76 0 2.2030008635390766e-08
GC_8_77 b_8 NI_8 NS_77 0 -6.0982957870068453e-05
GC_8_78 b_8 NI_8 NS_78 0 6.4431260603480832e-05
GC_8_79 b_8 NI_8 NS_79 0 -3.0538690357745444e-06
GC_8_80 b_8 NI_8 NS_80 0 -1.2068345885271515e-06
GC_8_81 b_8 NI_8 NS_81 0 -5.2754100552009171e-06
GC_8_82 b_8 NI_8 NS_82 0 -1.2386946183512120e-05
GC_8_83 b_8 NI_8 NS_83 0 -1.2300988782441987e-04
GC_8_84 b_8 NI_8 NS_84 0 2.6460789109125649e-05
GC_8_85 b_8 NI_8 NS_85 0 -8.5507141967126700e-05
GC_8_86 b_8 NI_8 NS_86 0 -4.5749619149000487e-05
GC_8_87 b_8 NI_8 NS_87 0 -1.5451556390134291e-05
GC_8_88 b_8 NI_8 NS_88 0 -3.2006998600201073e-06
GC_8_89 b_8 NI_8 NS_89 0 1.0514065926672908e-02
GC_8_90 b_8 NI_8 NS_90 0 -5.4058377238708156e-04
GC_8_91 b_8 NI_8 NS_91 0 -1.5154914903479338e-02
GC_8_92 b_8 NI_8 NS_92 0 5.6633492917467568e-03
GC_8_93 b_8 NI_8 NS_93 0 2.8294697761636505e-03
GC_8_94 b_8 NI_8 NS_94 0 -1.2088446004759322e-02
GC_8_95 b_8 NI_8 NS_95 0 8.3137025276591205e-03
GC_8_96 b_8 NI_8 NS_96 0 6.6309770995790331e-04
GC_8_97 b_8 NI_8 NS_97 0 -3.4484997010405957e-04
GC_8_98 b_8 NI_8 NS_98 0 -2.8598223430459860e-05
GC_8_99 b_8 NI_8 NS_99 0 -6.7348291807609109e-03
GC_8_100 b_8 NI_8 NS_100 0 -3.2229970949944932e-03
GC_8_101 b_8 NI_8 NS_101 0 -2.4894218878713121e-04
GC_8_102 b_8 NI_8 NS_102 0 1.1680764457516718e-04
GC_8_103 b_8 NI_8 NS_103 0 1.7347978838575212e-04
GC_8_104 b_8 NI_8 NS_104 0 4.1149025659733577e-05
GC_8_105 b_8 NI_8 NS_105 0 4.6942272912426085e-04
GC_8_106 b_8 NI_8 NS_106 0 1.4013402084115813e-04
GC_8_107 b_8 NI_8 NS_107 0 1.2727223474938106e-06
GC_8_108 b_8 NI_8 NS_108 0 1.1211335419853672e-05
GC_8_109 b_8 NI_8 NS_109 0 -3.7678167096457141e-07
GC_8_110 b_8 NI_8 NS_110 0 -1.4114224300083362e-05
GC_8_111 b_8 NI_8 NS_111 0 3.0806649660732321e-06
GC_8_112 b_8 NI_8 NS_112 0 -5.3051361946212191e-07
GC_8_113 b_8 NI_8 NS_113 0 2.3954362665779350e-03
GC_8_114 b_8 NI_8 NS_114 0 3.3323572354629120e-03
GC_8_115 b_8 NI_8 NS_115 0 5.1032123515624105e-04
GC_8_116 b_8 NI_8 NS_116 0 -2.1558234051140233e-03
GC_8_117 b_8 NI_8 NS_117 0 6.6241398564926266e-05
GC_8_118 b_8 NI_8 NS_118 0 5.4420217291196535e-05
GC_8_119 b_8 NI_8 NS_119 0 6.4337507987627800e-07
GC_8_120 b_8 NI_8 NS_120 0 4.1806208403149323e-07
GC_8_121 b_8 NI_8 NS_121 0 2.2552325329687113e-05
GC_8_122 b_8 NI_8 NS_122 0 -7.9382844952871129e-06
GC_8_123 b_8 NI_8 NS_123 0 2.1940902841325035e-07
GC_8_124 b_8 NI_8 NS_124 0 -1.4624724365450250e-07
GC_8_125 b_8 NI_8 NS_125 0 2.9189598158366816e-07
GC_8_126 b_8 NI_8 NS_126 0 -1.2057456190519311e-06
GC_8_127 b_8 NI_8 NS_127 0 -4.4287581135871926e-05
GC_8_128 b_8 NI_8 NS_128 0 5.0083392130173806e-05
GC_8_129 b_8 NI_8 NS_129 0 -8.6788980109260580e-06
GC_8_130 b_8 NI_8 NS_130 0 3.3894161815933080e-05
GC_8_131 b_8 NI_8 NS_131 0 3.5248380954709964e-06
GC_8_132 b_8 NI_8 NS_132 0 2.2051796556837772e-06
GC_8_133 b_8 NI_8 NS_133 0 -1.4671280403463148e-02
GC_8_134 b_8 NI_8 NS_134 0 -3.9612008524602078e-05
GC_8_135 b_8 NI_8 NS_135 0 1.0735646632765689e-02
GC_8_136 b_8 NI_8 NS_136 0 -8.0555438698417126e-03
GC_8_137 b_8 NI_8 NS_137 0 -2.2205184117405452e-03
GC_8_138 b_8 NI_8 NS_138 0 7.4174858857309475e-03
GC_8_139 b_8 NI_8 NS_139 0 5.8634918567747234e-03
GC_8_140 b_8 NI_8 NS_140 0 3.2191624985112014e-05
GC_8_141 b_8 NI_8 NS_141 0 -1.0338921838642390e-03
GC_8_142 b_8 NI_8 NS_142 0 -4.5070260359845190e-06
GC_8_143 b_8 NI_8 NS_143 0 -1.3392216981324809e-03
GC_8_144 b_8 NI_8 NS_144 0 3.8124200847916481e-03
GC_8_145 b_8 NI_8 NS_145 0 1.1933038061478903e-04
GC_8_146 b_8 NI_8 NS_146 0 -1.4633060599066020e-04
GC_8_147 b_8 NI_8 NS_147 0 2.3851015762141185e-05
GC_8_148 b_8 NI_8 NS_148 0 -3.7598973388033609e-05
GC_8_149 b_8 NI_8 NS_149 0 6.4637648404614084e-05
GC_8_150 b_8 NI_8 NS_150 0 -6.4426350145507840e-05
GC_8_151 b_8 NI_8 NS_151 0 6.6625356829603700e-06
GC_8_152 b_8 NI_8 NS_152 0 -8.2070104992716462e-07
GC_8_153 b_8 NI_8 NS_153 0 4.4391318304817992e-06
GC_8_154 b_8 NI_8 NS_154 0 1.7479473788167214e-06
GC_8_155 b_8 NI_8 NS_155 0 -1.2042987845890287e-06
GC_8_156 b_8 NI_8 NS_156 0 2.0397137255638690e-07
GC_8_157 b_8 NI_8 NS_157 0 1.4559893821872601e-03
GC_8_158 b_8 NI_8 NS_158 0 3.7260726853052891e-03
GC_8_159 b_8 NI_8 NS_159 0 -5.2046170625081245e-04
GC_8_160 b_8 NI_8 NS_160 0 -1.6075189593958957e-03
GC_8_161 b_8 NI_8 NS_161 0 -2.2441269655397198e-04
GC_8_162 b_8 NI_8 NS_162 0 -5.5430691673778416e-05
GC_8_163 b_8 NI_8 NS_163 0 -1.4782810093874926e-07
GC_8_164 b_8 NI_8 NS_164 0 5.4686732273473771e-07
GC_8_165 b_8 NI_8 NS_165 0 -3.2622666533502071e-05
GC_8_166 b_8 NI_8 NS_166 0 8.0490468727787565e-05
GC_8_167 b_8 NI_8 NS_167 0 -3.0471003588209099e-06
GC_8_168 b_8 NI_8 NS_168 0 1.9903398820918057e-07
GC_8_169 b_8 NI_8 NS_169 0 -6.1210686508460819e-06
GC_8_170 b_8 NI_8 NS_170 0 -1.2557782516335116e-05
GC_8_171 b_8 NI_8 NS_171 0 -1.4722852605906445e-04
GC_8_172 b_8 NI_8 NS_172 0 7.5941640691777311e-05
GC_8_173 b_8 NI_8 NS_173 0 -1.0485339413305144e-04
GC_8_174 b_8 NI_8 NS_174 0 -2.9691151766616629e-05
GC_8_175 b_8 NI_8 NS_175 0 -1.4870896669024282e-05
GC_8_176 b_8 NI_8 NS_176 0 2.6716918566159330e-06
GC_8_177 b_8 NI_8 NS_177 0 5.3117525551164444e-03
GC_8_178 b_8 NI_8 NS_178 0 -3.4365694724904490e-04
GC_8_179 b_8 NI_8 NS_179 0 -1.9971882412578388e-02
GC_8_180 b_8 NI_8 NS_180 0 -3.0245411875640580e-03
GC_8_181 b_8 NI_8 NS_181 0 9.7982095617109004e-03
GC_8_182 b_8 NI_8 NS_182 0 -2.9828054633953224e-03
GC_8_183 b_8 NI_8 NS_183 0 5.6535050806042954e-03
GC_8_184 b_8 NI_8 NS_184 0 5.5762876877719848e-04
GC_8_185 b_8 NI_8 NS_185 0 2.2363204799432240e-03
GC_8_186 b_8 NI_8 NS_186 0 -3.9035827238165520e-04
GC_8_187 b_8 NI_8 NS_187 0 -2.0827490631037559e-04
GC_8_188 b_8 NI_8 NS_188 0 -8.9815090995539245e-03
GC_8_189 b_8 NI_8 NS_189 0 -2.5813605053039319e-04
GC_8_190 b_8 NI_8 NS_190 0 1.0030187056164411e-04
GC_8_191 b_8 NI_8 NS_191 0 2.2578959543765407e-04
GC_8_192 b_8 NI_8 NS_192 0 5.2177047703547898e-05
GC_8_193 b_8 NI_8 NS_193 0 4.3582627497293868e-04
GC_8_194 b_8 NI_8 NS_194 0 4.4577164807080316e-04
GC_8_195 b_8 NI_8 NS_195 0 2.2967443813895806e-05
GC_8_196 b_8 NI_8 NS_196 0 2.7912270853004264e-05
GC_8_197 b_8 NI_8 NS_197 0 5.6546243809255117e-05
GC_8_198 b_8 NI_8 NS_198 0 -6.4920680256287428e-06
GC_8_199 b_8 NI_8 NS_199 0 6.2764557964036020e-06
GC_8_200 b_8 NI_8 NS_200 0 -1.7734222969593341e-06
GC_8_201 b_8 NI_8 NS_201 0 -5.8493308428285672e-03
GC_8_202 b_8 NI_8 NS_202 0 8.9112016487609396e-03
GC_8_203 b_8 NI_8 NS_203 0 4.2883855088155440e-03
GC_8_204 b_8 NI_8 NS_204 0 -3.9254650144776608e-03
GC_8_205 b_8 NI_8 NS_205 0 -2.2543551512393481e-04
GC_8_206 b_8 NI_8 NS_206 0 1.6173885610409623e-04
GC_8_207 b_8 NI_8 NS_207 0 -8.9621890537927558e-07
GC_8_208 b_8 NI_8 NS_208 0 4.5080165508537834e-07
GC_8_209 b_8 NI_8 NS_209 0 -7.1820357024794547e-06
GC_8_210 b_8 NI_8 NS_210 0 5.0950835896463529e-05
GC_8_211 b_8 NI_8 NS_211 0 -1.6752471426257697e-07
GC_8_212 b_8 NI_8 NS_212 0 6.1315702702914363e-07
GC_8_213 b_8 NI_8 NS_213 0 8.9882225359082657e-07
GC_8_214 b_8 NI_8 NS_214 0 8.3013983882002233e-07
GC_8_215 b_8 NI_8 NS_215 0 -7.4655509108434835e-05
GC_8_216 b_8 NI_8 NS_216 0 -1.7674251278363448e-04
GC_8_217 b_8 NI_8 NS_217 0 -2.8288028214657058e-06
GC_8_218 b_8 NI_8 NS_218 0 -2.9368078386252110e-05
GC_8_219 b_8 NI_8 NS_219 0 -2.6804632783537523e-06
GC_8_220 b_8 NI_8 NS_220 0 -7.6383025818860525e-06
GC_8_221 b_8 NI_8 NS_221 0 -9.7066265209055785e-03
GC_8_222 b_8 NI_8 NS_222 0 -9.4596811027393532e-04
GC_8_223 b_8 NI_8 NS_223 0 1.3631649729863426e-02
GC_8_224 b_8 NI_8 NS_224 0 2.7905397308378281e-03
GC_8_225 b_8 NI_8 NS_225 0 -1.5667987275341147e-02
GC_8_226 b_8 NI_8 NS_226 0 -3.6561043783441926e-03
GC_8_227 b_8 NI_8 NS_227 0 5.4852631635972701e-03
GC_8_228 b_8 NI_8 NS_228 0 -1.3271597842460787e-03
GC_8_229 b_8 NI_8 NS_229 0 -7.3861607459965175e-04
GC_8_230 b_8 NI_8 NS_230 0 6.8618872769682664e-04
GC_8_231 b_8 NI_8 NS_231 0 1.9224541293908191e-03
GC_8_232 b_8 NI_8 NS_232 0 -3.5056746073900517e-03
GC_8_233 b_8 NI_8 NS_233 0 8.7739258958870984e-05
GC_8_234 b_8 NI_8 NS_234 0 -1.3437037900939465e-04
GC_8_235 b_8 NI_8 NS_235 0 1.4876582476112849e-05
GC_8_236 b_8 NI_8 NS_236 0 -3.8187390179383173e-05
GC_8_237 b_8 NI_8 NS_237 0 7.5485542792475070e-05
GC_8_238 b_8 NI_8 NS_238 0 -7.5105405971376558e-05
GC_8_239 b_8 NI_8 NS_239 0 4.4239403579659893e-06
GC_8_240 b_8 NI_8 NS_240 0 -8.4701318978033011e-06
GC_8_241 b_8 NI_8 NS_241 0 -1.3698030329947977e-05
GC_8_242 b_8 NI_8 NS_242 0 -1.3952994160285417e-05
GC_8_243 b_8 NI_8 NS_243 0 -4.1088225143861772e-06
GC_8_244 b_8 NI_8 NS_244 0 -9.6123718561603298e-07
GC_8_245 b_8 NI_8 NS_245 0 7.4074546445979262e-03
GC_8_246 b_8 NI_8 NS_246 0 6.9523945611976853e-03
GC_8_247 b_8 NI_8 NS_247 0 -2.8837180862503918e-03
GC_8_248 b_8 NI_8 NS_248 0 -3.3439362559344512e-03
GC_8_249 b_8 NI_8 NS_249 0 -2.4770875036398630e-04
GC_8_250 b_8 NI_8 NS_250 0 7.5608802933518608e-05
GC_8_251 b_8 NI_8 NS_251 0 -3.3714632771410996e-07
GC_8_252 b_8 NI_8 NS_252 0 1.5975625822799488e-06
GC_8_253 b_8 NI_8 NS_253 0 -1.1933144620068720e-05
GC_8_254 b_8 NI_8 NS_254 0 1.2769747154876498e-04
GC_8_255 b_8 NI_8 NS_255 0 -2.9501731132795102e-06
GC_8_256 b_8 NI_8 NS_256 0 -7.3138894121600940e-07
GC_8_257 b_8 NI_8 NS_257 0 -7.0394952714527294e-06
GC_8_258 b_8 NI_8 NS_258 0 -1.8912958483677878e-05
GC_8_259 b_8 NI_8 NS_259 0 -3.1588707384848608e-04
GC_8_260 b_8 NI_8 NS_260 0 1.8334380777699287e-04
GC_8_261 b_8 NI_8 NS_261 0 -1.8513841179665873e-04
GC_8_262 b_8 NI_8 NS_262 0 -3.3901960157555798e-05
GC_8_263 b_8 NI_8 NS_263 0 -2.3165393931035964e-05
GC_8_264 b_8 NI_8 NS_264 0 1.0566553169885876e-05
GC_8_265 b_8 NI_8 NS_265 0 3.0345586105108489e-02
GC_8_266 b_8 NI_8 NS_266 0 1.6567569493169187e-02
GC_8_267 b_8 NI_8 NS_267 0 -1.9639967248414724e-02
GC_8_268 b_8 NI_8 NS_268 0 -6.0010372914104581e-03
GC_8_269 b_8 NI_8 NS_269 0 -2.7653552805349813e-02
GC_8_270 b_8 NI_8 NS_270 0 1.3586390375419000e-03
GC_8_271 b_8 NI_8 NS_271 0 2.3949683403661796e-03
GC_8_272 b_8 NI_8 NS_272 0 1.7316508049722745e-03
GC_8_273 b_8 NI_8 NS_273 0 -1.1942220505416206e-03
GC_8_274 b_8 NI_8 NS_274 0 1.1387796392588780e-03
GC_8_275 b_8 NI_8 NS_275 0 7.9306211588123683e-03
GC_8_276 b_8 NI_8 NS_276 0 -3.8432297545224836e-03
GC_8_277 b_8 NI_8 NS_277 0 -3.1739138430676012e-04
GC_8_278 b_8 NI_8 NS_278 0 5.2908898973599665e-05
GC_8_279 b_8 NI_8 NS_279 0 6.2981587277300221e-05
GC_8_280 b_8 NI_8 NS_280 0 2.0929374550180516e-05
GC_8_281 b_8 NI_8 NS_281 0 1.1905110525494950e-04
GC_8_282 b_8 NI_8 NS_282 0 -4.4050925313729217e-04
GC_8_283 b_8 NI_8 NS_283 0 -4.1805576190820375e-05
GC_8_284 b_8 NI_8 NS_284 0 2.9251233705421564e-07
GC_8_285 b_8 NI_8 NS_285 0 -7.5658259998979648e-05
GC_8_286 b_8 NI_8 NS_286 0 1.8702338408229029e-05
GC_8_287 b_8 NI_8 NS_287 0 4.2147443018835324e-07
GC_8_288 b_8 NI_8 NS_288 0 2.9364603803196664e-06
GC_8_289 b_8 NI_8 NS_289 0 4.0311006346967980e-04
GC_8_290 b_8 NI_8 NS_290 0 -7.8347510414878713e-03
GC_8_291 b_8 NI_8 NS_291 0 -9.5602287718607340e-04
GC_8_292 b_8 NI_8 NS_292 0 2.8189952421607176e-03
GC_8_293 b_8 NI_8 NS_293 0 2.3608923416101009e-04
GC_8_294 b_8 NI_8 NS_294 0 1.5679284374397646e-04
GC_8_295 b_8 NI_8 NS_295 0 2.3456923981379787e-06
GC_8_296 b_8 NI_8 NS_296 0 4.8623968856923491e-07
GC_8_297 b_8 NI_8 NS_297 0 3.9457072116039403e-05
GC_8_298 b_8 NI_8 NS_298 0 -6.2485811107673548e-05
GC_8_299 b_8 NI_8 NS_299 0 8.0395806572695467e-07
GC_8_300 b_8 NI_8 NS_300 0 -1.8006287311613220e-06
GC_8_301 b_8 NI_8 NS_301 0 1.6862245916845824e-06
GC_8_302 b_8 NI_8 NS_302 0 -3.8933125274080267e-06
GC_8_303 b_8 NI_8 NS_303 0 7.2647524476495773e-05
GC_8_304 b_8 NI_8 NS_304 0 1.7115084872844011e-04
GC_8_305 b_8 NI_8 NS_305 0 3.7180883435474291e-06
GC_8_306 b_8 NI_8 NS_306 0 5.2362870107952856e-05
GC_8_307 b_8 NI_8 NS_307 0 1.0282566081272461e-05
GC_8_308 b_8 NI_8 NS_308 0 5.5513726852820152e-06
GC_8_309 b_8 NI_8 NS_309 0 -1.3498871019285411e-01
GC_8_310 b_8 NI_8 NS_310 0 1.7434457226571571e-02
GC_8_311 b_8 NI_8 NS_311 0 9.3838503668210883e-03
GC_8_312 b_8 NI_8 NS_312 0 1.3564129239431597e-02
GC_8_313 b_8 NI_8 NS_313 0 1.5350952531900859e-02
GC_8_314 b_8 NI_8 NS_314 0 -1.2614372714058960e-02
GC_8_315 b_8 NI_8 NS_315 0 8.1955747954231574e-04
GC_8_316 b_8 NI_8 NS_316 0 1.8071449422098326e-03
GC_8_317 b_8 NI_8 NS_317 0 -4.8166459644200356e-04
GC_8_318 b_8 NI_8 NS_318 0 8.2396557054123304e-04
GC_8_319 b_8 NI_8 NS_319 0 5.8465279852721415e-03
GC_8_320 b_8 NI_8 NS_320 0 2.3258646372266876e-03
GC_8_321 b_8 NI_8 NS_321 0 -1.7784439084520480e-05
GC_8_322 b_8 NI_8 NS_322 0 -2.2028093468348734e-04
GC_8_323 b_8 NI_8 NS_323 0 6.1704879066613668e-05
GC_8_324 b_8 NI_8 NS_324 0 -7.5291410151107963e-05
GC_8_325 b_8 NI_8 NS_325 0 1.6895409608898464e-04
GC_8_326 b_8 NI_8 NS_326 0 2.3276318810613433e-04
GC_8_327 b_8 NI_8 NS_327 0 4.3115458961241519e-05
GC_8_328 b_8 NI_8 NS_328 0 1.9503446811346866e-05
GC_8_329 b_8 NI_8 NS_329 0 9.3327039556622581e-05
GC_8_330 b_8 NI_8 NS_330 0 3.0469935515081017e-05
GC_8_331 b_8 NI_8 NS_331 0 4.4182904981139189e-06
GC_8_332 b_8 NI_8 NS_332 0 -3.7257672311095448e-07
GC_8_333 b_8 NI_8 NS_333 0 -7.5974896769242786e-03
GC_8_334 b_8 NI_8 NS_334 0 1.8908993912972168e-03
GC_8_335 b_8 NI_8 NS_335 0 3.9799465921219355e-03
GC_8_336 b_8 NI_8 NS_336 0 -3.4867783615603735e-04
GC_8_337 b_8 NI_8 NS_337 0 1.4647675515051207e-04
GC_8_338 b_8 NI_8 NS_338 0 -4.3295024476761908e-04
GC_8_339 b_8 NI_8 NS_339 0 1.9877769528325788e-06
GC_8_340 b_8 NI_8 NS_340 0 -4.0252535753005299e-06
GC_8_341 b_8 NI_8 NS_341 0 -1.4065495457194385e-04
GC_8_342 b_8 NI_8 NS_342 0 -5.6002758895333426e-05
GC_8_343 b_8 NI_8 NS_343 0 -6.6615125394292038e-06
GC_8_344 b_8 NI_8 NS_344 0 -1.6721155671082020e-06
GC_8_345 b_8 NI_8 NS_345 0 -1.0407931716239219e-05
GC_8_346 b_8 NI_8 NS_346 0 -1.4262571889305074e-05
GC_8_347 b_8 NI_8 NS_347 0 1.7235077957397830e-04
GC_8_348 b_8 NI_8 NS_348 0 -1.5431574844908973e-04
GC_8_349 b_8 NI_8 NS_349 0 1.6786473631244723e-05
GC_8_350 b_8 NI_8 NS_350 0 -4.5881089838307566e-05
GC_8_351 b_8 NI_8 NS_351 0 4.5030897845147346e-06
GC_8_352 b_8 NI_8 NS_352 0 -1.7177901551593523e-05
GC_8_353 b_8 NI_8 NS_353 0 -4.1618362139533164e-03
GC_8_354 b_8 NI_8 NS_354 0 -9.3097685022838116e-05
GC_8_355 b_8 NI_8 NS_355 0 -3.4254422922341413e-03
GC_8_356 b_8 NI_8 NS_356 0 2.0319650507157668e-03
GC_8_357 b_8 NI_8 NS_357 0 -4.9991833770359005e-04
GC_8_358 b_8 NI_8 NS_358 0 -4.0450611884379900e-03
GC_8_359 b_8 NI_8 NS_359 0 1.3964490585492806e-03
GC_8_360 b_8 NI_8 NS_360 0 -1.1547664270375431e-03
GC_8_361 b_8 NI_8 NS_361 0 1.0210927141661200e-04
GC_8_362 b_8 NI_8 NS_362 0 -2.1052225925407298e-04
GC_8_363 b_8 NI_8 NS_363 0 -9.6474519053545323e-04
GC_8_364 b_8 NI_8 NS_364 0 -2.7863777925036639e-03
GC_8_365 b_8 NI_8 NS_365 0 -1.0845047901366903e-04
GC_8_366 b_8 NI_8 NS_366 0 2.1776560376324884e-04
GC_8_367 b_8 NI_8 NS_367 0 2.0328315916884988e-04
GC_8_368 b_8 NI_8 NS_368 0 -5.6948298314745205e-05
GC_8_369 b_8 NI_8 NS_369 0 -9.1897359759624927e-05
GC_8_370 b_8 NI_8 NS_370 0 -1.5687921708736418e-04
GC_8_371 b_8 NI_8 NS_371 0 -3.1204498936372247e-05
GC_8_372 b_8 NI_8 NS_372 0 -2.5658371447840477e-05
GC_8_373 b_8 NI_8 NS_373 0 -4.6427497825901326e-05
GC_8_374 b_8 NI_8 NS_374 0 -5.7913821007369822e-05
GC_8_375 b_8 NI_8 NS_375 0 2.0465184713816032e-06
GC_8_376 b_8 NI_8 NS_376 0 3.6336391204410913e-07
GC_8_377 b_8 NI_8 NS_377 0 6.1605115452973988e-03
GC_8_378 b_8 NI_8 NS_378 0 3.0675404248534772e-03
GC_8_379 b_8 NI_8 NS_379 0 -2.9753533796482239e-03
GC_8_380 b_8 NI_8 NS_380 0 -2.6104651180070644e-03
GC_8_381 b_8 NI_8 NS_381 0 4.3639223105852017e-05
GC_8_382 b_8 NI_8 NS_382 0 1.9023397483743790e-04
GC_8_383 b_8 NI_8 NS_383 0 2.6028249322231284e-07
GC_8_384 b_8 NI_8 NS_384 0 9.6483369795224271e-07
GC_8_385 b_8 NI_8 NS_385 0 4.3188243240466140e-05
GC_8_386 b_8 NI_8 NS_386 0 9.5008043994636516e-06
GC_8_387 b_8 NI_8 NS_387 0 2.2599734396211281e-07
GC_8_388 b_8 NI_8 NS_388 0 3.6287841650171890e-07
GC_8_389 b_8 NI_8 NS_389 0 3.3652251089656273e-06
GC_8_390 b_8 NI_8 NS_390 0 6.6152349714820582e-07
GC_8_391 b_8 NI_8 NS_391 0 -1.5028261652405174e-04
GC_8_392 b_8 NI_8 NS_392 0 -6.0098442395958327e-07
GC_8_393 b_8 NI_8 NS_393 0 -1.5626214077562652e-05
GC_8_394 b_8 NI_8 NS_394 0 -1.8964576528535920e-05
GC_8_395 b_8 NI_8 NS_395 0 -3.8385826151112020e-06
GC_8_396 b_8 NI_8 NS_396 0 6.5804769671178849e-06
GC_8_397 b_8 NI_8 NS_397 0 -6.5654896695792426e-03
GC_8_398 b_8 NI_8 NS_398 0 1.4070739759078426e-05
GC_8_399 b_8 NI_8 NS_399 0 2.1104382165692487e-03
GC_8_400 b_8 NI_8 NS_400 0 -2.2927271862660066e-03
GC_8_401 b_8 NI_8 NS_401 0 -4.0182995272034969e-04
GC_8_402 b_8 NI_8 NS_402 0 2.3103511168937369e-03
GC_8_403 b_8 NI_8 NS_403 0 7.1908537375202179e-04
GC_8_404 b_8 NI_8 NS_404 0 -6.6616716591901893e-04
GC_8_405 b_8 NI_8 NS_405 0 3.8058525062592655e-04
GC_8_406 b_8 NI_8 NS_406 0 -1.0825052297325639e-04
GC_8_407 b_8 NI_8 NS_407 0 -4.1404677224804676e-04
GC_8_408 b_8 NI_8 NS_408 0 3.8833425489222370e-04
GC_8_409 b_8 NI_8 NS_409 0 -5.4546876476851793e-05
GC_8_410 b_8 NI_8 NS_410 0 -9.7045471598222825e-05
GC_8_411 b_8 NI_8 NS_411 0 2.8305771125800490e-05
GC_8_412 b_8 NI_8 NS_412 0 -4.1622894108610652e-05
GC_8_413 b_8 NI_8 NS_413 0 -1.0112047015327693e-04
GC_8_414 b_8 NI_8 NS_414 0 1.1016057188759258e-04
GC_8_415 b_8 NI_8 NS_415 0 -8.8336809976651159e-06
GC_8_416 b_8 NI_8 NS_416 0 9.4572640934447373e-06
GC_8_417 b_8 NI_8 NS_417 0 -9.9977219450211253e-06
GC_8_418 b_8 NI_8 NS_418 0 4.0459777747441157e-05
GC_8_419 b_8 NI_8 NS_419 0 -1.4669081635896448e-06
GC_8_420 b_8 NI_8 NS_420 0 2.0014075069587903e-07
GC_8_421 b_8 NI_8 NS_421 0 2.7811173274871494e-03
GC_8_422 b_8 NI_8 NS_422 0 -2.0345485694487140e-03
GC_8_423 b_8 NI_8 NS_423 0 -1.7534937851623445e-03
GC_8_424 b_8 NI_8 NS_424 0 1.0823793245746374e-03
GC_8_425 b_8 NI_8 NS_425 0 2.7883327216606286e-05
GC_8_426 b_8 NI_8 NS_426 0 -3.5939214159206220e-05
GC_8_427 b_8 NI_8 NS_427 0 1.5361131296352460e-06
GC_8_428 b_8 NI_8 NS_428 0 -2.5906415074307878e-07
GC_8_429 b_8 NI_8 NS_429 0 -2.3407525917555776e-05
GC_8_430 b_8 NI_8 NS_430 0 -1.4251665470824309e-05
GC_8_431 b_8 NI_8 NS_431 0 8.2809318641563421e-07
GC_8_432 b_8 NI_8 NS_432 0 5.2003294970824880e-06
GC_8_433 b_8 NI_8 NS_433 0 -9.2030184331908374e-06
GC_8_434 b_8 NI_8 NS_434 0 -2.1598177008954063e-05
GC_8_435 b_8 NI_8 NS_435 0 -4.5944367057763490e-05
GC_8_436 b_8 NI_8 NS_436 0 1.8296510119918645e-04
GC_8_437 b_8 NI_8 NS_437 0 -1.5583744254588460e-04
GC_8_438 b_8 NI_8 NS_438 0 -7.1629463184886323e-06
GC_8_439 b_8 NI_8 NS_439 0 2.6324116115432645e-05
GC_8_440 b_8 NI_8 NS_440 0 3.8418595726428234e-05
GC_8_441 b_8 NI_8 NS_441 0 -7.2805286979953446e-04
GC_8_442 b_8 NI_8 NS_442 0 -1.0592867708815297e-04
GC_8_443 b_8 NI_8 NS_443 0 -5.6660594162068079e-03
GC_8_444 b_8 NI_8 NS_444 0 -9.1823177327935367e-04
GC_8_445 b_8 NI_8 NS_445 0 2.1705414359744993e-03
GC_8_446 b_8 NI_8 NS_446 0 -4.1311994997430461e-04
GC_8_447 b_8 NI_8 NS_447 0 6.6842937432290059e-04
GC_8_448 b_8 NI_8 NS_448 0 -4.6299382282516481e-04
GC_8_449 b_8 NI_8 NS_449 0 8.4566392280166817e-04
GC_8_450 b_8 NI_8 NS_450 0 2.3034670944396308e-04
GC_8_451 b_8 NI_8 NS_451 0 6.2427406936093504e-04
GC_8_452 b_8 NI_8 NS_452 0 -4.4556831061236049e-03
GC_8_453 b_8 NI_8 NS_453 0 -1.3745598398041256e-04
GC_8_454 b_8 NI_8 NS_454 0 1.5070338868870015e-04
GC_8_455 b_8 NI_8 NS_455 0 1.5406557710496792e-04
GC_8_456 b_8 NI_8 NS_456 0 -2.7668304018819956e-05
GC_8_457 b_8 NI_8 NS_457 0 -7.6293647452307868e-05
GC_8_458 b_8 NI_8 NS_458 0 -3.3923979180487574e-05
GC_8_459 b_8 NI_8 NS_459 0 -1.8395520540958119e-05
GC_8_460 b_8 NI_8 NS_460 0 -1.0688579017044042e-05
GC_8_461 b_8 NI_8 NS_461 0 -1.7353200145267430e-05
GC_8_462 b_8 NI_8 NS_462 0 -2.8379848114266225e-05
GC_8_463 b_8 NI_8 NS_463 0 2.0420192581255030e-06
GC_8_464 b_8 NI_8 NS_464 0 4.1574867662809824e-07
GC_8_465 b_8 NI_8 NS_465 0 1.5056720964588270e-03
GC_8_466 b_8 NI_8 NS_466 0 3.2374092983115444e-03
GC_8_467 b_8 NI_8 NS_467 0 -6.9847109796717646e-04
GC_8_468 b_8 NI_8 NS_468 0 -1.7851805217996551e-03
GC_8_469 b_8 NI_8 NS_469 0 3.3018846141912275e-05
GC_8_470 b_8 NI_8 NS_470 0 1.7319109542166764e-04
GC_8_471 b_8 NI_8 NS_471 0 1.6094935856089560e-07
GC_8_472 b_8 NI_8 NS_472 0 3.1376557243517251e-07
GC_8_473 b_8 NI_8 NS_473 0 3.3999313319914329e-05
GC_8_474 b_8 NI_8 NS_474 0 4.2129591277315830e-06
GC_8_475 b_8 NI_8 NS_475 0 6.5827951778945285e-07
GC_8_476 b_8 NI_8 NS_476 0 3.1769739621215271e-07
GC_8_477 b_8 NI_8 NS_477 0 -6.6327387525926880e-07
GC_8_478 b_8 NI_8 NS_478 0 -8.7826448050231153e-07
GC_8_479 b_8 NI_8 NS_479 0 -7.3533624121265644e-05
GC_8_480 b_8 NI_8 NS_480 0 -3.0345372253579563e-05
GC_8_481 b_8 NI_8 NS_481 0 -1.2848234746741485e-05
GC_8_482 b_8 NI_8 NS_482 0 -8.9770545010869801e-06
GC_8_483 b_8 NI_8 NS_483 0 2.2219855354947344e-06
GC_8_484 b_8 NI_8 NS_484 0 1.9794130799244765e-06
GC_8_485 b_8 NI_8 NS_485 0 -1.5486858777897625e-03
GC_8_486 b_8 NI_8 NS_486 0 -3.5231288951187987e-04
GC_8_487 b_8 NI_8 NS_487 0 3.8115909101870725e-03
GC_8_488 b_8 NI_8 NS_488 0 1.9431288310771844e-03
GC_8_489 b_8 NI_8 NS_489 0 -5.7326668809373127e-03
GC_8_490 b_8 NI_8 NS_490 0 -1.5733240587978115e-03
GC_8_491 b_8 NI_8 NS_491 0 7.8471878613730847e-04
GC_8_492 b_8 NI_8 NS_492 0 -6.0615700562076131e-04
GC_8_493 b_8 NI_8 NS_493 0 2.2348756940763077e-04
GC_8_494 b_8 NI_8 NS_494 0 3.4945715564513004e-04
GC_8_495 b_8 NI_8 NS_495 0 5.4670033154532397e-04
GC_8_496 b_8 NI_8 NS_496 0 -1.9578561260610631e-03
GC_8_497 b_8 NI_8 NS_497 0 -4.4516932215543635e-05
GC_8_498 b_8 NI_8 NS_498 0 -6.0017652261417835e-05
GC_8_499 b_8 NI_8 NS_499 0 1.7366513284304823e-05
GC_8_500 b_8 NI_8 NS_500 0 -2.9323561135619087e-05
GC_8_501 b_8 NI_8 NS_501 0 -7.4360235474980036e-05
GC_8_502 b_8 NI_8 NS_502 0 6.2773929283692400e-05
GC_8_503 b_8 NI_8 NS_503 0 -6.1280135848430101e-06
GC_8_504 b_8 NI_8 NS_504 0 1.2388185532753786e-06
GC_8_505 b_8 NI_8 NS_505 0 -1.0717438370747699e-05
GC_8_506 b_8 NI_8 NS_506 0 1.3690102806513149e-05
GC_8_507 b_8 NI_8 NS_507 0 -1.3302421358625877e-06
GC_8_508 b_8 NI_8 NS_508 0 5.1766192262232493e-07
GC_8_509 b_8 NI_8 NS_509 0 3.0793950464285272e-03
GC_8_510 b_8 NI_8 NS_510 0 3.5657386593729973e-04
GC_8_511 b_8 NI_8 NS_511 0 -1.5595379996991364e-03
GC_8_512 b_8 NI_8 NS_512 0 -2.5251759548984500e-04
GC_8_513 b_8 NI_8 NS_513 0 -4.1907051709867013e-06
GC_8_514 b_8 NI_8 NS_514 0 7.2307595488689931e-05
GC_8_515 b_8 NI_8 NS_515 0 9.3764965681284294e-07
GC_8_516 b_8 NI_8 NS_516 0 1.7017258573198332e-07
GC_8_517 b_8 NI_8 NS_517 0 4.8632805863115321e-06
GC_8_518 b_8 NI_8 NS_518 0 1.3104812675989385e-05
GC_8_519 b_8 NI_8 NS_519 0 -1.3426139828979218e-07
GC_8_520 b_8 NI_8 NS_520 0 3.4906142092922029e-06
GC_8_521 b_8 NI_8 NS_521 0 -4.4742496331481726e-06
GC_8_522 b_8 NI_8 NS_522 0 -1.2432072389930705e-05
GC_8_523 b_8 NI_8 NS_523 0 -7.4957430356572651e-05
GC_8_524 b_8 NI_8 NS_524 0 1.0707737033852531e-04
GC_8_525 b_8 NI_8 NS_525 0 -9.3114093978392359e-05
GC_8_526 b_8 NI_8 NS_526 0 -2.1115771812039443e-06
GC_8_527 b_8 NI_8 NS_527 0 9.5946968373381018e-06
GC_8_528 b_8 NI_8 NS_528 0 2.0479795271432951e-05
GD_8_1 b_8 NI_8 NA_1 0 -9.8904579298574151e-03
GD_8_2 b_8 NI_8 NA_2 0 1.4622702056546722e-03
GD_8_3 b_8 NI_8 NA_3 0 -2.8358596812201697e-03
GD_8_4 b_8 NI_8 NA_4 0 8.7422291379429524e-04
GD_8_5 b_8 NI_8 NA_5 0 -2.6693183174990713e-03
GD_8_6 b_8 NI_8 NA_6 0 -9.6644532436222178e-05
GD_8_7 b_8 NI_8 NA_7 0 -9.1138840882410161e-03
GD_8_8 b_8 NI_8 NA_8 0 1.3163162521421237e-01
GD_8_9 b_8 NI_8 NA_9 0 5.6845931965737954e-03
GD_8_10 b_8 NI_8 NA_10 0 3.7501335521255867e-03
GD_8_11 b_8 NI_8 NA_11 0 1.4948353692688825e-03
GD_8_12 b_8 NI_8 NA_12 0 6.1594338326591616e-04
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 -1.1394110043609230e-02
GC_9_2 b_9 NI_9 NS_2 0 5.3879744221198391e-05
GC_9_3 b_9 NI_9 NS_3 0 -9.8723080462374086e-04
GC_9_4 b_9 NI_9 NS_4 0 -6.7885736986798275e-04
GC_9_5 b_9 NI_9 NS_5 0 2.7015328322822351e-04
GC_9_6 b_9 NI_9 NS_6 0 -1.8137468306987144e-03
GC_9_7 b_9 NI_9 NS_7 0 9.8065716253655844e-04
GC_9_8 b_9 NI_9 NS_8 0 -2.1464622949615665e-03
GC_9_9 b_9 NI_9 NS_9 0 3.6936230799127721e-04
GC_9_10 b_9 NI_9 NS_10 0 1.3125386895622038e-03
GC_9_11 b_9 NI_9 NS_11 0 3.9409123339834162e-04
GC_9_12 b_9 NI_9 NS_12 0 -2.7742375994548876e-04
GC_9_13 b_9 NI_9 NS_13 0 3.4404789774481419e-04
GC_9_14 b_9 NI_9 NS_14 0 -2.7109771613108329e-04
GC_9_15 b_9 NI_9 NS_15 0 2.9707605304675710e-04
GC_9_16 b_9 NI_9 NS_16 0 6.0787934286052228e-04
GC_9_17 b_9 NI_9 NS_17 0 -1.9167768098630569e-03
GC_9_18 b_9 NI_9 NS_18 0 -1.5694669517799153e-03
GC_9_19 b_9 NI_9 NS_19 0 1.4566888759792092e-04
GC_9_20 b_9 NI_9 NS_20 0 9.4418302102694507e-05
GC_9_21 b_9 NI_9 NS_21 0 -7.5079176415204026e-04
GC_9_22 b_9 NI_9 NS_22 0 -2.6223496031895460e-06
GC_9_23 b_9 NI_9 NS_23 0 -1.7724531171804240e-06
GC_9_24 b_9 NI_9 NS_24 0 -4.1820800005522134e-06
GC_9_25 b_9 NI_9 NS_25 0 1.1962236119658774e-02
GC_9_26 b_9 NI_9 NS_26 0 7.5139379540393077e-03
GC_9_27 b_9 NI_9 NS_27 0 -5.7663301145390771e-03
GC_9_28 b_9 NI_9 NS_28 0 -8.4439103321111951e-03
GC_9_29 b_9 NI_9 NS_29 0 5.0316366105045183e-05
GC_9_30 b_9 NI_9 NS_30 0 2.4328749992239812e-04
GC_9_31 b_9 NI_9 NS_31 0 4.7883113125200495e-08
GC_9_32 b_9 NI_9 NS_32 0 -1.9304201918943712e-07
GC_9_33 b_9 NI_9 NS_33 0 -1.6233474382991807e-05
GC_9_34 b_9 NI_9 NS_34 0 -7.3436249902449977e-05
GC_9_35 b_9 NI_9 NS_35 0 -3.9354883776178165e-09
GC_9_36 b_9 NI_9 NS_36 0 1.2088391620990810e-07
GC_9_37 b_9 NI_9 NS_37 0 -6.8269680056082769e-07
GC_9_38 b_9 NI_9 NS_38 0 -3.5484685237741808e-06
GC_9_39 b_9 NI_9 NS_39 0 2.3502666210673716e-04
GC_9_40 b_9 NI_9 NS_40 0 4.0007149268338947e-04
GC_9_41 b_9 NI_9 NS_41 0 -1.4727562969128101e-04
GC_9_42 b_9 NI_9 NS_42 0 8.1879697462761326e-05
GC_9_43 b_9 NI_9 NS_43 0 -1.1231031129478538e-05
GC_9_44 b_9 NI_9 NS_44 0 -7.4139974408346931e-06
GC_9_45 b_9 NI_9 NS_45 0 -3.0548453918608268e-03
GC_9_46 b_9 NI_9 NS_46 0 4.2903336641734222e-05
GC_9_47 b_9 NI_9 NS_47 0 -9.6647408528553249e-06
GC_9_48 b_9 NI_9 NS_48 0 3.6005487693596536e-04
GC_9_49 b_9 NI_9 NS_49 0 -9.9797222235509415e-04
GC_9_50 b_9 NI_9 NS_50 0 -4.1025550018235419e-04
GC_9_51 b_9 NI_9 NS_51 0 -2.4854498401008317e-04
GC_9_52 b_9 NI_9 NS_52 0 -1.4564868200066311e-03
GC_9_53 b_9 NI_9 NS_53 0 3.1072139561258818e-04
GC_9_54 b_9 NI_9 NS_54 0 -4.1918890120018655e-05
GC_9_55 b_9 NI_9 NS_55 0 1.4124705031721863e-03
GC_9_56 b_9 NI_9 NS_56 0 -1.1653485419028079e-03
GC_9_57 b_9 NI_9 NS_57 0 -1.0494437660210654e-05
GC_9_58 b_9 NI_9 NS_58 0 1.8459527648338145e-04
GC_9_59 b_9 NI_9 NS_59 0 2.1211595109364812e-04
GC_9_60 b_9 NI_9 NS_60 0 -8.7597575019115163e-05
GC_9_61 b_9 NI_9 NS_61 0 -1.8971725494102402e-04
GC_9_62 b_9 NI_9 NS_62 0 1.2548583488418197e-04
GC_9_63 b_9 NI_9 NS_63 0 -1.8410270438327116e-05
GC_9_64 b_9 NI_9 NS_64 0 -1.5639364519904848e-05
GC_9_65 b_9 NI_9 NS_65 0 -4.4386195558427800e-06
GC_9_66 b_9 NI_9 NS_66 0 -5.0753899602951689e-05
GC_9_67 b_9 NI_9 NS_67 0 4.7062720113832658e-06
GC_9_68 b_9 NI_9 NS_68 0 2.4035829340758703e-06
GC_9_69 b_9 NI_9 NS_69 0 2.3765047109722843e-03
GC_9_70 b_9 NI_9 NS_70 0 3.0204123580648877e-03
GC_9_71 b_9 NI_9 NS_71 0 -1.4545168383701939e-03
GC_9_72 b_9 NI_9 NS_72 0 -2.2237740734173607e-03
GC_9_73 b_9 NI_9 NS_73 0 -1.4344081759094831e-04
GC_9_74 b_9 NI_9 NS_74 0 4.4317697326561250e-05
GC_9_75 b_9 NI_9 NS_75 0 -7.7608163436788033e-07
GC_9_76 b_9 NI_9 NS_76 0 4.6675061898033908e-07
GC_9_77 b_9 NI_9 NS_77 0 8.0425714866638163e-08
GC_9_78 b_9 NI_9 NS_78 0 2.8073070446819351e-05
GC_9_79 b_9 NI_9 NS_79 0 -9.9666977822783363e-07
GC_9_80 b_9 NI_9 NS_80 0 1.1224869086848839e-06
GC_9_81 b_9 NI_9 NS_81 0 1.7158802719705772e-06
GC_9_82 b_9 NI_9 NS_82 0 6.0925076513487809e-07
GC_9_83 b_9 NI_9 NS_83 0 -1.0052660390033057e-04
GC_9_84 b_9 NI_9 NS_84 0 -8.9327236264791403e-05
GC_9_85 b_9 NI_9 NS_85 0 -4.9561199467064441e-06
GC_9_86 b_9 NI_9 NS_86 0 -5.4431559589160241e-05
GC_9_87 b_9 NI_9 NS_87 0 -6.9059987283781613e-06
GC_9_88 b_9 NI_9 NS_88 0 1.4081668083336577e-06
GC_9_89 b_9 NI_9 NS_89 0 -1.6010149182669655e-02
GC_9_90 b_9 NI_9 NS_90 0 8.4556712492930955e-05
GC_9_91 b_9 NI_9 NS_91 0 -1.0880593474424988e-03
GC_9_92 b_9 NI_9 NS_92 0 -1.3722877455203764e-03
GC_9_93 b_9 NI_9 NS_93 0 7.2095672858119172e-04
GC_9_94 b_9 NI_9 NS_94 0 -2.0089286349000411e-03
GC_9_95 b_9 NI_9 NS_95 0 1.8327073446930959e-03
GC_9_96 b_9 NI_9 NS_96 0 -2.4202876331503092e-03
GC_9_97 b_9 NI_9 NS_97 0 7.5045369873800614e-04
GC_9_98 b_9 NI_9 NS_98 0 9.8520254495127997e-04
GC_9_99 b_9 NI_9 NS_99 0 -6.7278517476774343e-04
GC_9_100 b_9 NI_9 NS_100 0 6.0838331308319684e-04
GC_9_101 b_9 NI_9 NS_101 0 4.6813767728825465e-04
GC_9_102 b_9 NI_9 NS_102 0 -3.4954146280000061e-04
GC_9_103 b_9 NI_9 NS_103 0 4.0783402292010888e-04
GC_9_104 b_9 NI_9 NS_104 0 8.7236767648585570e-04
GC_9_105 b_9 NI_9 NS_105 0 -2.7876297777500586e-03
GC_9_106 b_9 NI_9 NS_106 0 -2.2314859015543022e-03
GC_9_107 b_9 NI_9 NS_107 0 2.0925991794827436e-04
GC_9_108 b_9 NI_9 NS_108 0 1.4856713555087776e-04
GC_9_109 b_9 NI_9 NS_109 0 -1.0575707871659133e-03
GC_9_110 b_9 NI_9 NS_110 0 9.2076646964924510e-07
GC_9_111 b_9 NI_9 NS_111 0 -2.5480238822720166e-06
GC_9_112 b_9 NI_9 NS_112 0 -3.7622174150027566e-06
GC_9_113 b_9 NI_9 NS_113 0 1.5846693001626506e-02
GC_9_114 b_9 NI_9 NS_114 0 8.8977282823699405e-03
GC_9_115 b_9 NI_9 NS_115 0 -7.8134765697858155e-03
GC_9_116 b_9 NI_9 NS_116 0 -1.1117849172031681e-02
GC_9_117 b_9 NI_9 NS_117 0 -2.0510235383857054e-05
GC_9_118 b_9 NI_9 NS_118 0 5.3591418898097905e-04
GC_9_119 b_9 NI_9 NS_119 0 5.5993450234570960e-08
GC_9_120 b_9 NI_9 NS_120 0 4.5085408718905126e-08
GC_9_121 b_9 NI_9 NS_121 0 -1.2243503354691412e-05
GC_9_122 b_9 NI_9 NS_122 0 -9.8372915013667970e-05
GC_9_123 b_9 NI_9 NS_123 0 4.3589435743657952e-07
GC_9_124 b_9 NI_9 NS_124 0 6.3551889308793178e-07
GC_9_125 b_9 NI_9 NS_125 0 -1.5228888850270890e-07
GC_9_126 b_9 NI_9 NS_126 0 -4.7680094947912243e-06
GC_9_127 b_9 NI_9 NS_127 0 3.2025091371577362e-04
GC_9_128 b_9 NI_9 NS_128 0 5.9623175434199947e-04
GC_9_129 b_9 NI_9 NS_129 0 -2.2013619201616773e-04
GC_9_130 b_9 NI_9 NS_130 0 1.1583315698660538e-04
GC_9_131 b_9 NI_9 NS_131 0 -1.8662076386426222e-05
GC_9_132 b_9 NI_9 NS_132 0 -8.2192323719448524e-06
GC_9_133 b_9 NI_9 NS_133 0 -2.7665593770446061e-03
GC_9_134 b_9 NI_9 NS_134 0 2.3848676764869808e-05
GC_9_135 b_9 NI_9 NS_135 0 -1.8665108248710455e-04
GC_9_136 b_9 NI_9 NS_136 0 1.0958629566774237e-03
GC_9_137 b_9 NI_9 NS_137 0 -1.9192392406505874e-03
GC_9_138 b_9 NI_9 NS_138 0 -9.4797577630001525e-04
GC_9_139 b_9 NI_9 NS_139 0 -1.1950401653710780e-04
GC_9_140 b_9 NI_9 NS_140 0 -2.0095925560262864e-03
GC_9_141 b_9 NI_9 NS_141 0 4.0981862017141086e-04
GC_9_142 b_9 NI_9 NS_142 0 4.1401935073116997e-04
GC_9_143 b_9 NI_9 NS_143 0 1.1378844060145803e-03
GC_9_144 b_9 NI_9 NS_144 0 -1.4196426355702540e-03
GC_9_145 b_9 NI_9 NS_145 0 -4.2762759547657756e-05
GC_9_146 b_9 NI_9 NS_146 0 2.8376264063791095e-04
GC_9_147 b_9 NI_9 NS_147 0 2.8615083716652305e-04
GC_9_148 b_9 NI_9 NS_148 0 -5.5018807482893492e-05
GC_9_149 b_9 NI_9 NS_149 0 -4.1482032653995034e-04
GC_9_150 b_9 NI_9 NS_150 0 -8.4882455951506336e-06
GC_9_151 b_9 NI_9 NS_151 0 -3.0721451216136997e-05
GC_9_152 b_9 NI_9 NS_152 0 -5.5385538692325157e-06
GC_9_153 b_9 NI_9 NS_153 0 -4.5921017934898551e-05
GC_9_154 b_9 NI_9 NS_154 0 -3.8872736723803182e-05
GC_9_155 b_9 NI_9 NS_155 0 3.7805612151591879e-06
GC_9_156 b_9 NI_9 NS_156 0 2.6211297484549216e-06
GC_9_157 b_9 NI_9 NS_157 0 4.1537484152293792e-03
GC_9_158 b_9 NI_9 NS_158 0 2.5532816055444060e-03
GC_9_159 b_9 NI_9 NS_159 0 -2.4389329149147473e-03
GC_9_160 b_9 NI_9 NS_160 0 -2.4427823384902958e-03
GC_9_161 b_9 NI_9 NS_161 0 -7.8708910054826574e-05
GC_9_162 b_9 NI_9 NS_162 0 3.4115984232235427e-05
GC_9_163 b_9 NI_9 NS_163 0 -3.5747683842787410e-07
GC_9_164 b_9 NI_9 NS_164 0 4.2833342486016911e-07
GC_9_165 b_9 NI_9 NS_165 0 1.4781630109308610e-06
GC_9_166 b_9 NI_9 NS_166 0 1.8509713307825941e-05
GC_9_167 b_9 NI_9 NS_167 0 -1.0610956312303502e-06
GC_9_168 b_9 NI_9 NS_168 0 5.6424242368557225e-07
GC_9_169 b_9 NI_9 NS_169 0 2.4592730295415037e-06
GC_9_170 b_9 NI_9 NS_170 0 -5.5099077374826148e-07
GC_9_171 b_9 NI_9 NS_171 0 -7.7184383045014922e-05
GC_9_172 b_9 NI_9 NS_172 0 -4.2278010238329049e-05
GC_9_173 b_9 NI_9 NS_173 0 6.1210227458100474e-06
GC_9_174 b_9 NI_9 NS_174 0 -4.0132187195273322e-05
GC_9_175 b_9 NI_9 NS_175 0 -2.5192484268107334e-06
GC_9_176 b_9 NI_9 NS_176 0 3.9560717926350963e-06
GC_9_177 b_9 NI_9 NS_177 0 -1.6158609900312981e-02
GC_9_178 b_9 NI_9 NS_178 0 9.1107310938883386e-05
GC_9_179 b_9 NI_9 NS_179 0 -4.3254019157911881e-04
GC_9_180 b_9 NI_9 NS_180 0 -1.8778414691809754e-03
GC_9_181 b_9 NI_9 NS_181 0 8.0261132070020105e-04
GC_9_182 b_9 NI_9 NS_182 0 -1.0036537689311843e-03
GC_9_183 b_9 NI_9 NS_183 0 2.0572436509999040e-03
GC_9_184 b_9 NI_9 NS_184 0 -1.5296001819547665e-03
GC_9_185 b_9 NI_9 NS_185 0 1.4875913351317105e-03
GC_9_186 b_9 NI_9 NS_186 0 5.0912717544956336e-04
GC_9_187 b_9 NI_9 NS_187 0 -2.8274675581327464e-03
GC_9_188 b_9 NI_9 NS_188 0 9.4844968661059604e-04
GC_9_189 b_9 NI_9 NS_189 0 4.8312754789076804e-04
GC_9_190 b_9 NI_9 NS_190 0 -3.3369915002472216e-04
GC_9_191 b_9 NI_9 NS_191 0 3.9123081488917513e-04
GC_9_192 b_9 NI_9 NS_192 0 8.9631101666165774e-04
GC_9_193 b_9 NI_9 NS_193 0 -2.8039633253659512e-03
GC_9_194 b_9 NI_9 NS_194 0 -2.3539979806315972e-03
GC_9_195 b_9 NI_9 NS_195 0 2.0109589934054514e-04
GC_9_196 b_9 NI_9 NS_196 0 1.4905611231956105e-04
GC_9_197 b_9 NI_9 NS_197 0 -1.0499536289492821e-03
GC_9_198 b_9 NI_9 NS_198 0 2.7558435783096901e-05
GC_9_199 b_9 NI_9 NS_199 0 -5.6646409241988755e-06
GC_9_200 b_9 NI_9 NS_200 0 -1.1322788230996171e-06
GC_9_201 b_9 NI_9 NS_201 0 1.5717068484344694e-02
GC_9_202 b_9 NI_9 NS_202 0 6.6254528864043930e-03
GC_9_203 b_9 NI_9 NS_203 0 -7.9304325621467366e-03
GC_9_204 b_9 NI_9 NS_204 0 -1.0255598463578080e-02
GC_9_205 b_9 NI_9 NS_205 0 -1.0155421041065335e-04
GC_9_206 b_9 NI_9 NS_206 0 5.9377354495707710e-04
GC_9_207 b_9 NI_9 NS_207 0 3.2944058727547605e-07
GC_9_208 b_9 NI_9 NS_208 0 2.3782145447838468e-07
GC_9_209 b_9 NI_9 NS_209 0 4.5743571821407960e-06
GC_9_210 b_9 NI_9 NS_210 0 -1.0484008446771973e-04
GC_9_211 b_9 NI_9 NS_211 0 3.4052897278573002e-07
GC_9_212 b_9 NI_9 NS_212 0 2.3972188554695245e-07
GC_9_213 b_9 NI_9 NS_213 0 -1.4652513307436836e-07
GC_9_214 b_9 NI_9 NS_214 0 -4.4748074803810284e-06
GC_9_215 b_9 NI_9 NS_215 0 3.0142477753231919e-04
GC_9_216 b_9 NI_9 NS_216 0 6.2621930701089047e-04
GC_9_217 b_9 NI_9 NS_217 0 -2.1232441495844113e-04
GC_9_218 b_9 NI_9 NS_218 0 1.0183783725933922e-04
GC_9_219 b_9 NI_9 NS_219 0 -1.9757008162510074e-05
GC_9_220 b_9 NI_9 NS_220 0 -9.2648038572492434e-06
GC_9_221 b_9 NI_9 NS_221 0 -5.2199223667347663e-05
GC_9_222 b_9 NI_9 NS_222 0 -5.2140906564556293e-05
GC_9_223 b_9 NI_9 NS_223 0 -7.0738106743087890e-04
GC_9_224 b_9 NI_9 NS_224 0 2.0717716619663719e-03
GC_9_225 b_9 NI_9 NS_225 0 -2.5928282580302752e-03
GC_9_226 b_9 NI_9 NS_226 0 -1.6990340159133285e-03
GC_9_227 b_9 NI_9 NS_227 0 2.4115312859669110e-04
GC_9_228 b_9 NI_9 NS_228 0 -1.8967101241772534e-03
GC_9_229 b_9 NI_9 NS_229 0 2.3977634773377461e-05
GC_9_230 b_9 NI_9 NS_230 0 6.8445141771082923e-04
GC_9_231 b_9 NI_9 NS_231 0 -8.3743548488997819e-05
GC_9_232 b_9 NI_9 NS_232 0 -1.4351597035105424e-03
GC_9_233 b_9 NI_9 NS_233 0 -5.7653040097293980e-05
GC_9_234 b_9 NI_9 NS_234 0 3.1313225657395803e-04
GC_9_235 b_9 NI_9 NS_235 0 2.7375028563978565e-04
GC_9_236 b_9 NI_9 NS_236 0 -7.1122349996595197e-05
GC_9_237 b_9 NI_9 NS_237 0 -4.8207527221247543e-04
GC_9_238 b_9 NI_9 NS_238 0 -9.0787482155151413e-05
GC_9_239 b_9 NI_9 NS_239 0 -3.7600020720393370e-05
GC_9_240 b_9 NI_9 NS_240 0 -5.4726523661964129e-06
GC_9_241 b_9 NI_9 NS_241 0 -9.0613464194156266e-05
GC_9_242 b_9 NI_9 NS_242 0 -4.4807556788060827e-05
GC_9_243 b_9 NI_9 NS_243 0 4.6109873445416846e-06
GC_9_244 b_9 NI_9 NS_244 0 5.7909092211543169e-06
GC_9_245 b_9 NI_9 NS_245 0 6.2277055389262257e-03
GC_9_246 b_9 NI_9 NS_246 0 1.6826596581216336e-03
GC_9_247 b_9 NI_9 NS_247 0 -3.7003658959505730e-03
GC_9_248 b_9 NI_9 NS_248 0 -2.1166610807594370e-03
GC_9_249 b_9 NI_9 NS_249 0 3.4200685744503009e-05
GC_9_250 b_9 NI_9 NS_250 0 6.3527253614966285e-05
GC_9_251 b_9 NI_9 NS_251 0 2.8980174056735337e-08
GC_9_252 b_9 NI_9 NS_252 0 4.9038390906839872e-07
GC_9_253 b_9 NI_9 NS_253 0 1.5243759811362514e-05
GC_9_254 b_9 NI_9 NS_254 0 -9.4672361167658939e-06
GC_9_255 b_9 NI_9 NS_255 0 -9.6353746656790629e-07
GC_9_256 b_9 NI_9 NS_256 0 6.2614716561377767e-07
GC_9_257 b_9 NI_9 NS_257 0 4.1113230934028740e-06
GC_9_258 b_9 NI_9 NS_258 0 -2.6724157170413053e-07
GC_9_259 b_9 NI_9 NS_259 0 -1.0216090963272538e-04
GC_9_260 b_9 NI_9 NS_260 0 -1.1184956838926862e-05
GC_9_261 b_9 NI_9 NS_261 0 -1.2887820877008131e-05
GC_9_262 b_9 NI_9 NS_262 0 -4.4744706243001300e-05
GC_9_263 b_9 NI_9 NS_263 0 -7.0801867836588557e-06
GC_9_264 b_9 NI_9 NS_264 0 5.7174045974000089e-06
GC_9_265 b_9 NI_9 NS_265 0 -7.2175652553152338e-03
GC_9_266 b_9 NI_9 NS_266 0 4.0551398261913030e-05
GC_9_267 b_9 NI_9 NS_267 0 1.9335304825859043e-03
GC_9_268 b_9 NI_9 NS_268 0 -1.5459930291887895e-03
GC_9_269 b_9 NI_9 NS_269 0 -1.1753708115917504e-03
GC_9_270 b_9 NI_9 NS_270 0 7.1462146040562056e-04
GC_9_271 b_9 NI_9 NS_271 0 2.4739555043352731e-03
GC_9_272 b_9 NI_9 NS_272 0 -3.4029816455556235e-05
GC_9_273 b_9 NI_9 NS_273 0 1.7508903810338564e-04
GC_9_274 b_9 NI_9 NS_274 0 7.1212522549257229e-04
GC_9_275 b_9 NI_9 NS_275 0 -3.3745137326391113e-03
GC_9_276 b_9 NI_9 NS_276 0 1.8943511562717345e-04
GC_9_277 b_9 NI_9 NS_277 0 4.2453574892512154e-04
GC_9_278 b_9 NI_9 NS_278 0 -1.7728940836726865e-04
GC_9_279 b_9 NI_9 NS_279 0 2.9733426805894896e-04
GC_9_280 b_9 NI_9 NS_280 0 6.0884568735111949e-04
GC_9_281 b_9 NI_9 NS_281 0 -1.5840679109543428e-03
GC_9_282 b_9 NI_9 NS_282 0 -1.4372871478061878e-03
GC_9_283 b_9 NI_9 NS_283 0 1.7043351425805386e-04
GC_9_284 b_9 NI_9 NS_284 0 1.2501332664885257e-04
GC_9_285 b_9 NI_9 NS_285 0 -6.6702467860387405e-04
GC_9_286 b_9 NI_9 NS_286 0 1.0739770262798211e-05
GC_9_287 b_9 NI_9 NS_287 0 -4.0231684304593654e-06
GC_9_288 b_9 NI_9 NS_288 0 -1.6768706568130155e-06
GC_9_289 b_9 NI_9 NS_289 0 8.8095447149806327e-03
GC_9_290 b_9 NI_9 NS_290 0 5.1660340645674329e-03
GC_9_291 b_9 NI_9 NS_291 0 -3.5560662962963036e-03
GC_9_292 b_9 NI_9 NS_292 0 -6.8177765225536152e-03
GC_9_293 b_9 NI_9 NS_293 0 -1.1657069007175689e-04
GC_9_294 b_9 NI_9 NS_294 0 3.0218388354212876e-04
GC_9_295 b_9 NI_9 NS_295 0 2.3041144711650662e-07
GC_9_296 b_9 NI_9 NS_296 0 -1.6325642329155786e-07
GC_9_297 b_9 NI_9 NS_297 0 1.4629907354024368e-06
GC_9_298 b_9 NI_9 NS_298 0 -7.9883577184203827e-05
GC_9_299 b_9 NI_9 NS_299 0 2.0985313971337908e-07
GC_9_300 b_9 NI_9 NS_300 0 3.0768800827044502e-07
GC_9_301 b_9 NI_9 NS_301 0 4.4105782084612372e-09
GC_9_302 b_9 NI_9 NS_302 0 -2.3463716035647691e-06
GC_9_303 b_9 NI_9 NS_303 0 1.5601311942713456e-04
GC_9_304 b_9 NI_9 NS_304 0 4.4744746847365902e-04
GC_9_305 b_9 NI_9 NS_305 0 -1.4084514213390256e-04
GC_9_306 b_9 NI_9 NS_306 0 6.0917700401367200e-05
GC_9_307 b_9 NI_9 NS_307 0 -1.5053221307122830e-05
GC_9_308 b_9 NI_9 NS_308 0 -5.8659903068036314e-06
GC_9_309 b_9 NI_9 NS_309 0 -4.1618362139531594e-03
GC_9_310 b_9 NI_9 NS_310 0 -9.3097685022836896e-05
GC_9_311 b_9 NI_9 NS_311 0 -3.4254422922341565e-03
GC_9_312 b_9 NI_9 NS_312 0 2.0319650507158032e-03
GC_9_313 b_9 NI_9 NS_313 0 -4.9991833770366366e-04
GC_9_314 b_9 NI_9 NS_314 0 -4.0450611884380429e-03
GC_9_315 b_9 NI_9 NS_315 0 1.3964490585492216e-03
GC_9_316 b_9 NI_9 NS_316 0 -1.1547664270376351e-03
GC_9_317 b_9 NI_9 NS_317 0 1.0210927141662611e-04
GC_9_318 b_9 NI_9 NS_318 0 -2.1052225925359568e-04
GC_9_319 b_9 NI_9 NS_319 0 -9.6474519053543469e-04
GC_9_320 b_9 NI_9 NS_320 0 -2.7863777925039484e-03
GC_9_321 b_9 NI_9 NS_321 0 -1.0845047901367747e-04
GC_9_322 b_9 NI_9 NS_322 0 2.1776560376325337e-04
GC_9_323 b_9 NI_9 NS_323 0 2.0328315916883381e-04
GC_9_324 b_9 NI_9 NS_324 0 -5.6948298314740732e-05
GC_9_325 b_9 NI_9 NS_325 0 -9.1897359759661641e-05
GC_9_326 b_9 NI_9 NS_326 0 -1.5687921708746615e-04
GC_9_327 b_9 NI_9 NS_327 0 -3.1204498936379680e-05
GC_9_328 b_9 NI_9 NS_328 0 -2.5658371447845664e-05
GC_9_329 b_9 NI_9 NS_329 0 -4.6427497825924982e-05
GC_9_330 b_9 NI_9 NS_330 0 -5.7913821007376585e-05
GC_9_331 b_9 NI_9 NS_331 0 2.0465184713801179e-06
GC_9_332 b_9 NI_9 NS_332 0 3.6336391204387958e-07
GC_9_333 b_9 NI_9 NS_333 0 6.1605115452991674e-03
GC_9_334 b_9 NI_9 NS_334 0 3.0675404248535969e-03
GC_9_335 b_9 NI_9 NS_335 0 -2.9753533796491529e-03
GC_9_336 b_9 NI_9 NS_336 0 -2.6104651180072886e-03
GC_9_337 b_9 NI_9 NS_337 0 4.3639223105848344e-05
GC_9_338 b_9 NI_9 NS_338 0 1.9023397483755044e-04
GC_9_339 b_9 NI_9 NS_339 0 2.6028249322272111e-07
GC_9_340 b_9 NI_9 NS_340 0 9.6483369795285659e-07
GC_9_341 b_9 NI_9 NS_341 0 4.3188243240491680e-05
GC_9_342 b_9 NI_9 NS_342 0 9.5008043994666992e-06
GC_9_343 b_9 NI_9 NS_343 0 2.2599734396259657e-07
GC_9_344 b_9 NI_9 NS_344 0 3.6287841650170429e-07
GC_9_345 b_9 NI_9 NS_345 0 3.3652251089659763e-06
GC_9_346 b_9 NI_9 NS_346 0 6.6152349714925657e-07
GC_9_347 b_9 NI_9 NS_347 0 -1.5028261652409898e-04
GC_9_348 b_9 NI_9 NS_348 0 -6.0098442394116189e-07
GC_9_349 b_9 NI_9 NS_349 0 -1.5626214077572505e-05
GC_9_350 b_9 NI_9 NS_350 0 -1.8964576528530635e-05
GC_9_351 b_9 NI_9 NS_351 0 -3.8385826151117831e-06
GC_9_352 b_9 NI_9 NS_352 0 6.5804769671191902e-06
GC_9_353 b_9 NI_9 NS_353 0 -7.7527667072166179e-04
GC_9_354 b_9 NI_9 NS_354 0 1.3305952547625769e-02
GC_9_355 b_9 NI_9 NS_355 0 1.2996826411509116e-02
GC_9_356 b_9 NI_9 NS_356 0 4.3976287143904788e-03
GC_9_357 b_9 NI_9 NS_357 0 1.6195862944604244e-02
GC_9_358 b_9 NI_9 NS_358 0 4.7096712031957600e-04
GC_9_359 b_9 NI_9 NS_359 0 1.3456158939228009e-02
GC_9_360 b_9 NI_9 NS_360 0 1.2314550568240060e-02
GC_9_361 b_9 NI_9 NS_361 0 2.1449524013703574e-03
GC_9_362 b_9 NI_9 NS_362 0 1.0688788864685282e-03
GC_9_363 b_9 NI_9 NS_363 0 -3.0249190122930330e-03
GC_9_364 b_9 NI_9 NS_364 0 2.0113420119738802e-02
GC_9_365 b_9 NI_9 NS_365 0 7.0377388852215970e-04
GC_9_366 b_9 NI_9 NS_366 0 3.8688464730367506e-04
GC_9_367 b_9 NI_9 NS_367 0 7.6697325049275623e-05
GC_9_368 b_9 NI_9 NS_368 0 3.2199950870826231e-04
GC_9_369 b_9 NI_9 NS_369 0 1.8577676806489649e-03
GC_9_370 b_9 NI_9 NS_370 0 -2.2936875263085494e-04
GC_9_371 b_9 NI_9 NS_371 0 2.1904532649901179e-04
GC_9_372 b_9 NI_9 NS_372 0 1.9383521496494155e-04
GC_9_373 b_9 NI_9 NS_373 0 2.2000521549317870e-04
GC_9_374 b_9 NI_9 NS_374 0 4.9192768325931861e-05
GC_9_375 b_9 NI_9 NS_375 0 -1.5953753512952281e-05
GC_9_376 b_9 NI_9 NS_376 0 6.0041763136611244e-06
GC_9_377 b_9 NI_9 NS_377 0 -2.6659171165114130e-02
GC_9_378 b_9 NI_9 NS_378 0 1.5309075689419107e-03
GC_9_379 b_9 NI_9 NS_379 0 1.8055449941715401e-02
GC_9_380 b_9 NI_9 NS_380 0 3.3674779677797190e-03
GC_9_381 b_9 NI_9 NS_381 0 -5.5701482151924802e-04
GC_9_382 b_9 NI_9 NS_382 0 -3.8147473865200818e-04
GC_9_383 b_9 NI_9 NS_383 0 2.3480419202202051e-06
GC_9_384 b_9 NI_9 NS_384 0 2.0468532400658526e-06
GC_9_385 b_9 NI_9 NS_385 0 1.9994660543287750e-04
GC_9_386 b_9 NI_9 NS_386 0 -6.9178934344280826e-05
GC_9_387 b_9 NI_9 NS_387 0 3.9064351950757742e-06
GC_9_388 b_9 NI_9 NS_388 0 9.0039675910087727e-07
GC_9_389 b_9 NI_9 NS_389 0 -3.6577985772566000e-07
GC_9_390 b_9 NI_9 NS_390 0 4.8832602288814983e-07
GC_9_391 b_9 NI_9 NS_391 0 -2.1265916662441858e-04
GC_9_392 b_9 NI_9 NS_392 0 4.3298846482958583e-04
GC_9_393 b_9 NI_9 NS_393 0 -1.2331674805150498e-05
GC_9_394 b_9 NI_9 NS_394 0 -8.5995123905070576e-05
GC_9_395 b_9 NI_9 NS_395 0 -2.3476857343340883e-05
GC_9_396 b_9 NI_9 NS_396 0 3.1416925225859839e-06
GC_9_397 b_9 NI_9 NS_397 0 5.0036266227609039e-02
GC_9_398 b_9 NI_9 NS_398 0 1.6071584659497134e-02
GC_9_399 b_9 NI_9 NS_399 0 -2.8776424522273119e-02
GC_9_400 b_9 NI_9 NS_400 0 1.7828641248073184e-03
GC_9_401 b_9 NI_9 NS_401 0 -2.9040846883456779e-02
GC_9_402 b_9 NI_9 NS_402 0 -9.1424757304603629e-03
GC_9_403 b_9 NI_9 NS_403 0 9.4344918295574103e-03
GC_9_404 b_9 NI_9 NS_404 0 2.6842595120575249e-03
GC_9_405 b_9 NI_9 NS_405 0 -2.8563734932079057e-03
GC_9_406 b_9 NI_9 NS_406 0 -3.3598973971509275e-04
GC_9_407 b_9 NI_9 NS_407 0 1.0950828795006039e-03
GC_9_408 b_9 NI_9 NS_408 0 -2.6817704714581650e-03
GC_9_409 b_9 NI_9 NS_409 0 -5.0250578372737866e-04
GC_9_410 b_9 NI_9 NS_410 0 9.7861125276343705e-05
GC_9_411 b_9 NI_9 NS_411 0 1.4762414045177400e-04
GC_9_412 b_9 NI_9 NS_412 0 3.6732122271115406e-05
GC_9_413 b_9 NI_9 NS_413 0 7.0511199253420946e-04
GC_9_414 b_9 NI_9 NS_414 0 -3.0702078182155533e-04
GC_9_415 b_9 NI_9 NS_415 0 2.7500133027399067e-06
GC_9_416 b_9 NI_9 NS_416 0 1.4934039353221519e-05
GC_9_417 b_9 NI_9 NS_417 0 4.4996409194623554e-06
GC_9_418 b_9 NI_9 NS_418 0 -8.3039516230941443e-06
GC_9_419 b_9 NI_9 NS_419 0 8.4537840049402721e-06
GC_9_420 b_9 NI_9 NS_420 0 6.3615405589587089e-07
GC_9_421 b_9 NI_9 NS_421 0 -3.1319721579091604e-03
GC_9_422 b_9 NI_9 NS_422 0 -3.6711192177799664e-03
GC_9_423 b_9 NI_9 NS_423 0 2.2340650113115428e-03
GC_9_424 b_9 NI_9 NS_424 0 5.4121741372736680e-04
GC_9_425 b_9 NI_9 NS_425 0 9.4495136852304400e-05
GC_9_426 b_9 NI_9 NS_426 0 -1.6044037374588339e-04
GC_9_427 b_9 NI_9 NS_427 0 9.8972455612949943e-07
GC_9_428 b_9 NI_9 NS_428 0 -6.0340054788681786e-07
GC_9_429 b_9 NI_9 NS_429 0 -3.6274103986946345e-05
GC_9_430 b_9 NI_9 NS_430 0 -5.6085242481036182e-05
GC_9_431 b_9 NI_9 NS_431 0 8.9303607780646928e-10
GC_9_432 b_9 NI_9 NS_432 0 -1.8542850472524777e-06
GC_9_433 b_9 NI_9 NS_433 0 5.5870194966696596e-06
GC_9_434 b_9 NI_9 NS_434 0 -3.0926920090921209e-06
GC_9_435 b_9 NI_9 NS_435 0 8.5765905340609382e-05
GC_9_436 b_9 NI_9 NS_436 0 9.0185910615498077e-05
GC_9_437 b_9 NI_9 NS_437 0 2.9832825597751102e-05
GC_9_438 b_9 NI_9 NS_438 0 1.8953170120870692e-05
GC_9_439 b_9 NI_9 NS_439 0 1.0780351641819062e-05
GC_9_440 b_9 NI_9 NS_440 0 -4.6450942597007735e-06
GC_9_441 b_9 NI_9 NS_441 0 1.1922627028366219e-02
GC_9_442 b_9 NI_9 NS_442 0 -6.5844195732113768e-04
GC_9_443 b_9 NI_9 NS_443 0 1.1369832599582757e-02
GC_9_444 b_9 NI_9 NS_444 0 4.1780408700606659e-03
GC_9_445 b_9 NI_9 NS_445 0 -9.7949700493270581e-03
GC_9_446 b_9 NI_9 NS_446 0 -8.3145698846087777e-03
GC_9_447 b_9 NI_9 NS_447 0 1.1198762804449614e-02
GC_9_448 b_9 NI_9 NS_448 0 6.9171363062514443e-03
GC_9_449 b_9 NI_9 NS_449 0 -3.0683196859481576e-03
GC_9_450 b_9 NI_9 NS_450 0 -2.5359853970917828e-03
GC_9_451 b_9 NI_9 NS_451 0 2.3248066546641835e-03
GC_9_452 b_9 NI_9 NS_452 0 3.8909047096627120e-03
GC_9_453 b_9 NI_9 NS_453 0 5.8142716380972027e-04
GC_9_454 b_9 NI_9 NS_454 0 3.4308214082468176e-04
GC_9_455 b_9 NI_9 NS_455 0 1.6421752533923482e-04
GC_9_456 b_9 NI_9 NS_456 0 3.3136555069081903e-04
GC_9_457 b_9 NI_9 NS_457 0 8.5588573610024133e-04
GC_9_458 b_9 NI_9 NS_458 0 1.6013636999630948e-04
GC_9_459 b_9 NI_9 NS_459 0 2.1246444548422063e-04
GC_9_460 b_9 NI_9 NS_460 0 1.8332738046137359e-04
GC_9_461 b_9 NI_9 NS_461 0 1.4584430503433360e-04
GC_9_462 b_9 NI_9 NS_462 0 4.7664821618550908e-05
GC_9_463 b_9 NI_9 NS_463 0 -5.3882975873412039e-06
GC_9_464 b_9 NI_9 NS_464 0 1.2511407388815709e-06
GC_9_465 b_9 NI_9 NS_465 0 -2.2779904017138111e-02
GC_9_466 b_9 NI_9 NS_466 0 1.0554424335503201e-02
GC_9_467 b_9 NI_9 NS_467 0 1.5573795652923484e-02
GC_9_468 b_9 NI_9 NS_468 0 -1.1837445138570409e-03
GC_9_469 b_9 NI_9 NS_469 0 -4.1324616077250916e-04
GC_9_470 b_9 NI_9 NS_470 0 -4.4059545533350973e-04
GC_9_471 b_9 NI_9 NS_471 0 6.9442206438379790e-07
GC_9_472 b_9 NI_9 NS_472 0 -2.3556084832646371e-07
GC_9_473 b_9 NI_9 NS_473 0 7.0284308372919898e-05
GC_9_474 b_9 NI_9 NS_474 0 -4.3043808869542358e-05
GC_9_475 b_9 NI_9 NS_475 0 1.1118405249021944e-06
GC_9_476 b_9 NI_9 NS_476 0 1.0051844965361363e-06
GC_9_477 b_9 NI_9 NS_477 0 -3.0885202042627007e-06
GC_9_478 b_9 NI_9 NS_478 0 -2.8306337455833390e-07
GC_9_479 b_9 NI_9 NS_479 0 -7.6137090614972035e-05
GC_9_480 b_9 NI_9 NS_480 0 1.4218921465658277e-04
GC_9_481 b_9 NI_9 NS_481 0 -9.1712066797774837e-06
GC_9_482 b_9 NI_9 NS_482 0 -8.2462677603541905e-05
GC_9_483 b_9 NI_9 NS_483 0 -1.8755641146988839e-05
GC_9_484 b_9 NI_9 NS_484 0 -8.2807764409902684e-06
GC_9_485 b_9 NI_9 NS_485 0 7.2221788558346611e-03
GC_9_486 b_9 NI_9 NS_486 0 -3.6221201072844352e-04
GC_9_487 b_9 NI_9 NS_487 0 -1.9882112977590974e-02
GC_9_488 b_9 NI_9 NS_488 0 -2.9310672005078832e-03
GC_9_489 b_9 NI_9 NS_489 0 9.7598244588682544e-03
GC_9_490 b_9 NI_9 NS_490 0 -2.7969796518780140e-03
GC_9_491 b_9 NI_9 NS_491 0 5.7013058624985485e-03
GC_9_492 b_9 NI_9 NS_492 0 6.7618349981701657e-04
GC_9_493 b_9 NI_9 NS_493 0 1.5968830043391513e-03
GC_9_494 b_9 NI_9 NS_494 0 -8.6069402703185761e-04
GC_9_495 b_9 NI_9 NS_495 0 -5.2205901742273725e-05
GC_9_496 b_9 NI_9 NS_496 0 -8.6046019501000055e-03
GC_9_497 b_9 NI_9 NS_497 0 -2.7012461749727754e-04
GC_9_498 b_9 NI_9 NS_498 0 9.0542398599852711e-05
GC_9_499 b_9 NI_9 NS_499 0 2.3050374309889038e-04
GC_9_500 b_9 NI_9 NS_500 0 3.4908456389671164e-05
GC_9_501 b_9 NI_9 NS_501 0 5.3532353537658528e-04
GC_9_502 b_9 NI_9 NS_502 0 4.8342451317561071e-04
GC_9_503 b_9 NI_9 NS_503 0 3.3166282548239424e-05
GC_9_504 b_9 NI_9 NS_504 0 2.3104994189697843e-05
GC_9_505 b_9 NI_9 NS_505 0 7.4281860200917159e-05
GC_9_506 b_9 NI_9 NS_506 0 -2.1860255518730700e-05
GC_9_507 b_9 NI_9 NS_507 0 6.7174860060833674e-06
GC_9_508 b_9 NI_9 NS_508 0 -3.0035187185827824e-06
GC_9_509 b_9 NI_9 NS_509 0 -7.1010896762910810e-03
GC_9_510 b_9 NI_9 NS_510 0 1.1143993545289086e-02
GC_9_511 b_9 NI_9 NS_511 0 5.0151273330537906e-03
GC_9_512 b_9 NI_9 NS_512 0 -4.9722785823224681e-03
GC_9_513 b_9 NI_9 NS_513 0 -3.9017729368488263e-04
GC_9_514 b_9 NI_9 NS_514 0 6.3164745032136471e-06
GC_9_515 b_9 NI_9 NS_515 0 -2.4927630367449831e-06
GC_9_516 b_9 NI_9 NS_516 0 -2.8432544330522360e-07
GC_9_517 b_9 NI_9 NS_517 0 -5.3738301810821695e-05
GC_9_518 b_9 NI_9 NS_518 0 9.0888003668954817e-05
GC_9_519 b_9 NI_9 NS_519 0 -1.1803819706381087e-06
GC_9_520 b_9 NI_9 NS_520 0 1.8404645000086643e-06
GC_9_521 b_9 NI_9 NS_521 0 -2.6448935699970725e-07
GC_9_522 b_9 NI_9 NS_522 0 2.1268368263308317e-06
GC_9_523 b_9 NI_9 NS_523 0 -1.1065874190352067e-04
GC_9_524 b_9 NI_9 NS_524 0 -2.7199021486740827e-04
GC_9_525 b_9 NI_9 NS_525 0 -3.7657372662897387e-06
GC_9_526 b_9 NI_9 NS_526 0 -6.0107678714469310e-05
GC_9_527 b_9 NI_9 NS_527 0 -7.8808636189532053e-06
GC_9_528 b_9 NI_9 NS_528 0 -1.2254870634133747e-05
GD_9_1 b_9 NI_9 NA_1 0 5.9829461827951578e-03
GD_9_2 b_9 NI_9 NA_2 0 1.9149126078420702e-03
GD_9_3 b_9 NI_9 NA_3 0 9.8570499902000848e-03
GD_9_4 b_9 NI_9 NA_4 0 2.1561735887676175e-03
GD_9_5 b_9 NI_9 NA_5 0 1.1174945952043847e-02
GD_9_6 b_9 NI_9 NA_6 0 1.3317487238098647e-03
GD_9_7 b_9 NI_9 NA_7 0 3.1710214399024569e-03
GD_9_8 b_9 NI_9 NA_8 0 5.6845931965721821e-03
GD_9_9 b_9 NI_9 NA_9 0 -1.8334457781461019e-01
GD_9_10 b_9 NI_9 NA_10 0 -1.5985849390849134e-02
GD_9_11 b_9 NI_9 NA_11 0 -2.1286062301483832e-02
GD_9_12 b_9 NI_9 NA_12 0 -2.6100856012958077e-03
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 -3.1343479687051677e-03
GC_10_2 b_10 NI_10 NS_2 0 4.3166440025265953e-05
GC_10_3 b_10 NI_10 NS_3 0 -1.5455853079254559e-05
GC_10_4 b_10 NI_10 NS_4 0 3.6118218363994986e-04
GC_10_5 b_10 NI_10 NS_5 0 -1.0071123414495959e-03
GC_10_6 b_10 NI_10 NS_6 0 -4.2339505591782909e-04
GC_10_7 b_10 NI_10 NS_7 0 -2.5534355234772870e-04
GC_10_8 b_10 NI_10 NS_8 0 -1.4776842959832385e-03
GC_10_9 b_10 NI_10 NS_9 0 2.8524762423575280e-04
GC_10_10 b_10 NI_10 NS_10 0 -5.0422578116646365e-05
GC_10_11 b_10 NI_10 NS_11 0 1.4139041255069678e-03
GC_10_12 b_10 NI_10 NS_12 0 -1.2322107141047958e-03
GC_10_13 b_10 NI_10 NS_13 0 -4.2027475770859668e-06
GC_10_14 b_10 NI_10 NS_14 0 1.8839119023428380e-04
GC_10_15 b_10 NI_10 NS_15 0 2.1091379052458697e-04
GC_10_16 b_10 NI_10 NS_16 0 -7.3898888176858981e-05
GC_10_17 b_10 NI_10 NS_17 0 -2.0294948991869498e-04
GC_10_18 b_10 NI_10 NS_18 0 6.1533548752781315e-05
GC_10_19 b_10 NI_10 NS_19 0 -8.6801400473542218e-06
GC_10_20 b_10 NI_10 NS_20 0 -1.1110998475040167e-05
GC_10_21 b_10 NI_10 NS_21 0 -2.9359761558826341e-05
GC_10_22 b_10 NI_10 NS_22 0 -5.7334880719602936e-05
GC_10_23 b_10 NI_10 NS_23 0 3.5413081315462035e-06
GC_10_24 b_10 NI_10 NS_24 0 3.0127554938967241e-06
GC_10_25 b_10 NI_10 NS_25 0 2.4421199316419324e-03
GC_10_26 b_10 NI_10 NS_26 0 3.7498088124319501e-03
GC_10_27 b_10 NI_10 NS_27 0 -1.4394589167898615e-03
GC_10_28 b_10 NI_10 NS_28 0 -2.8128705914655079e-03
GC_10_29 b_10 NI_10 NS_29 0 -1.4192475295541745e-04
GC_10_30 b_10 NI_10 NS_30 0 2.9433315895309948e-05
GC_10_31 b_10 NI_10 NS_31 0 -6.2237066143714973e-07
GC_10_32 b_10 NI_10 NS_32 0 1.3836169282013703e-07
GC_10_33 b_10 NI_10 NS_33 0 -1.6028860889485160e-05
GC_10_34 b_10 NI_10 NS_34 0 3.0736977570053517e-05
GC_10_35 b_10 NI_10 NS_35 0 -6.8950972062817088e-07
GC_10_36 b_10 NI_10 NS_36 0 7.1768388345752009e-07
GC_10_37 b_10 NI_10 NS_37 0 1.3589709023689366e-06
GC_10_38 b_10 NI_10 NS_38 0 1.0565294902683055e-06
GC_10_39 b_10 NI_10 NS_39 0 -6.0861550190601051e-05
GC_10_40 b_10 NI_10 NS_40 0 -9.6861852872084865e-05
GC_10_41 b_10 NI_10 NS_41 0 -3.3346111761859674e-07
GC_10_42 b_10 NI_10 NS_42 0 -4.3028551479236906e-05
GC_10_43 b_10 NI_10 NS_43 0 -8.2481922745320839e-06
GC_10_44 b_10 NI_10 NS_44 0 -3.2058185792672055e-06
GC_10_45 b_10 NI_10 NS_45 0 -7.4712241648757800e-03
GC_10_46 b_10 NI_10 NS_46 0 -3.7561783335313652e-06
GC_10_47 b_10 NI_10 NS_47 0 -7.0776931132155612e-04
GC_10_48 b_10 NI_10 NS_48 0 -3.6537222418053019e-04
GC_10_49 b_10 NI_10 NS_49 0 1.3974827401092517e-04
GC_10_50 b_10 NI_10 NS_50 0 -9.7990084198339698e-04
GC_10_51 b_10 NI_10 NS_51 0 -5.5936302972056325e-05
GC_10_52 b_10 NI_10 NS_52 0 -1.2390964501962844e-03
GC_10_53 b_10 NI_10 NS_53 0 9.5009474298899201e-04
GC_10_54 b_10 NI_10 NS_54 0 7.0719923835679376e-04
GC_10_55 b_10 NI_10 NS_55 0 1.1643597078637667e-03
GC_10_56 b_10 NI_10 NS_56 0 -8.1019452495916834e-04
GC_10_57 b_10 NI_10 NS_57 0 -6.5949394401339402e-05
GC_10_58 b_10 NI_10 NS_58 0 -7.0904955867127079e-05
GC_10_59 b_10 NI_10 NS_59 0 2.7971431652470190e-05
GC_10_60 b_10 NI_10 NS_60 0 -2.9507957953525018e-05
GC_10_61 b_10 NI_10 NS_61 0 -1.4569953788205381e-04
GC_10_62 b_10 NI_10 NS_62 0 1.9184084497496381e-04
GC_10_63 b_10 NI_10 NS_63 0 -9.9678491836836080e-06
GC_10_64 b_10 NI_10 NS_64 0 1.8883028600055469e-05
GC_10_65 b_10 NI_10 NS_65 0 -4.7106866881902534e-06
GC_10_66 b_10 NI_10 NS_66 0 6.4296425312794649e-05
GC_10_67 b_10 NI_10 NS_67 0 -7.9851578341622355e-07
GC_10_68 b_10 NI_10 NS_68 0 -2.0953949566855504e-07
GC_10_69 b_10 NI_10 NS_69 0 3.4019245258349916e-03
GC_10_70 b_10 NI_10 NS_70 0 -4.2108099289022956e-03
GC_10_71 b_10 NI_10 NS_71 0 -1.9831653689057096e-03
GC_10_72 b_10 NI_10 NS_72 0 2.3988985359620759e-03
GC_10_73 b_10 NI_10 NS_73 0 1.3333553247117378e-04
GC_10_74 b_10 NI_10 NS_74 0 7.1231993320833162e-05
GC_10_75 b_10 NI_10 NS_75 0 2.1726896164720875e-06
GC_10_76 b_10 NI_10 NS_76 0 4.9065804508786726e-07
GC_10_77 b_10 NI_10 NS_77 0 1.8764448668054165e-05
GC_10_78 b_10 NI_10 NS_78 0 -6.6746659652548813e-05
GC_10_79 b_10 NI_10 NS_79 0 3.8683657990555300e-06
GC_10_80 b_10 NI_10 NS_80 0 7.2832691611758826e-06
GC_10_81 b_10 NI_10 NS_81 0 -9.5787296962123863e-06
GC_10_82 b_10 NI_10 NS_82 0 -2.2926818877180186e-05
GC_10_83 b_10 NI_10 NS_83 0 -1.7534704644655432e-05
GC_10_84 b_10 NI_10 NS_84 0 2.5946716169115617e-04
GC_10_85 b_10 NI_10 NS_85 0 -1.8547747699624239e-04
GC_10_86 b_10 NI_10 NS_86 0 1.3937575907495585e-06
GC_10_87 b_10 NI_10 NS_87 0 4.3717681186856205e-05
GC_10_88 b_10 NI_10 NS_88 0 6.0599615467946614e-05
GC_10_89 b_10 NI_10 NS_89 0 -3.2927922961518241e-03
GC_10_90 b_10 NI_10 NS_90 0 2.2446999109578966e-05
GC_10_91 b_10 NI_10 NS_91 0 -2.3649087140538940e-04
GC_10_92 b_10 NI_10 NS_92 0 1.1270724318286779e-03
GC_10_93 b_10 NI_10 NS_93 0 -1.9781904552558351e-03
GC_10_94 b_10 NI_10 NS_94 0 -1.0394287052685352e-03
GC_10_95 b_10 NI_10 NS_95 0 -1.1642155414613576e-04
GC_10_96 b_10 NI_10 NS_96 0 -2.1027193702553614e-03
GC_10_97 b_10 NI_10 NS_97 0 5.4967923160357038e-04
GC_10_98 b_10 NI_10 NS_98 0 4.3256135722342676e-04
GC_10_99 b_10 NI_10 NS_99 0 1.0728716969333404e-03
GC_10_100 b_10 NI_10 NS_100 0 -1.4856778190152564e-03
GC_10_101 b_10 NI_10 NS_101 0 -2.5758262342042431e-05
GC_10_102 b_10 NI_10 NS_102 0 2.8541115645749991e-04
GC_10_103 b_10 NI_10 NS_103 0 2.8697881013274910e-04
GC_10_104 b_10 NI_10 NS_104 0 -8.1332166019953305e-05
GC_10_105 b_10 NI_10 NS_105 0 -4.2960364440372068e-04
GC_10_106 b_10 NI_10 NS_106 0 3.7185475766580182e-05
GC_10_107 b_10 NI_10 NS_107 0 -2.1485800825196973e-05
GC_10_108 b_10 NI_10 NS_108 0 -1.3805957372461017e-06
GC_10_109 b_10 NI_10 NS_109 0 -5.7868421055882179e-05
GC_10_110 b_10 NI_10 NS_110 0 -4.1755665061172945e-05
GC_10_111 b_10 NI_10 NS_111 0 4.8360285741321410e-06
GC_10_112 b_10 NI_10 NS_112 0 4.8951747507593712e-06
GC_10_113 b_10 NI_10 NS_113 0 4.7302599547048617e-03
GC_10_114 b_10 NI_10 NS_114 0 2.0426220108490422e-03
GC_10_115 b_10 NI_10 NS_115 0 -2.8695060019828691e-03
GC_10_116 b_10 NI_10 NS_116 0 -2.1824961772378190e-03
GC_10_117 b_10 NI_10 NS_117 0 -1.0021021831675196e-04
GC_10_118 b_10 NI_10 NS_118 0 1.3801248494058842e-05
GC_10_119 b_10 NI_10 NS_119 0 -6.5732898542652921e-07
GC_10_120 b_10 NI_10 NS_120 0 -3.0161191679797786e-07
GC_10_121 b_10 NI_10 NS_121 0 -1.2367332438258505e-05
GC_10_122 b_10 NI_10 NS_122 0 4.0147865682933249e-05
GC_10_123 b_10 NI_10 NS_123 0 1.0315818908455902e-06
GC_10_124 b_10 NI_10 NS_124 0 4.3900986526991245e-07
GC_10_125 b_10 NI_10 NS_125 0 -1.8678496968802407e-06
GC_10_126 b_10 NI_10 NS_126 0 -1.1860836047632790e-06
GC_10_127 b_10 NI_10 NS_127 0 -5.2268710855028942e-05
GC_10_128 b_10 NI_10 NS_128 0 -2.9095808706721796e-05
GC_10_129 b_10 NI_10 NS_129 0 -1.8127078908019422e-05
GC_10_130 b_10 NI_10 NS_130 0 -1.5549735082452481e-05
GC_10_131 b_10 NI_10 NS_131 0 4.3221708450042545e-06
GC_10_132 b_10 NI_10 NS_132 0 1.7151045972189844e-07
GC_10_133 b_10 NI_10 NS_133 0 -8.5331280581767144e-03
GC_10_134 b_10 NI_10 NS_134 0 -1.0516661592719122e-05
GC_10_135 b_10 NI_10 NS_135 0 -7.3311588018820184e-04
GC_10_136 b_10 NI_10 NS_136 0 -9.8325201273691894e-04
GC_10_137 b_10 NI_10 NS_137 0 7.0731758696430599e-04
GC_10_138 b_10 NI_10 NS_138 0 -7.7756952199129522e-04
GC_10_139 b_10 NI_10 NS_139 0 2.9114187515424787e-04
GC_10_140 b_10 NI_10 NS_140 0 -1.3867303364479000e-03
GC_10_141 b_10 NI_10 NS_141 0 7.7151127018125802e-04
GC_10_142 b_10 NI_10 NS_142 0 5.1468907704980364e-04
GC_10_143 b_10 NI_10 NS_143 0 1.5440900687515439e-03
GC_10_144 b_10 NI_10 NS_144 0 -8.0100793033525169e-05
GC_10_145 b_10 NI_10 NS_145 0 -9.5371414495042204e-05
GC_10_146 b_10 NI_10 NS_146 0 -1.0126519495775106e-04
GC_10_147 b_10 NI_10 NS_147 0 4.9773257698553983e-05
GC_10_148 b_10 NI_10 NS_148 0 -3.2382803585574320e-05
GC_10_149 b_10 NI_10 NS_149 0 -2.3576028298918632e-04
GC_10_150 b_10 NI_10 NS_150 0 2.5376975570770571e-04
GC_10_151 b_10 NI_10 NS_151 0 -1.5147555002122594e-05
GC_10_152 b_10 NI_10 NS_152 0 2.0079655066209039e-05
GC_10_153 b_10 NI_10 NS_153 0 -1.0025987308451503e-05
GC_10_154 b_10 NI_10 NS_154 0 6.4482059525619226e-05
GC_10_155 b_10 NI_10 NS_155 0 -1.0112959989641198e-06
GC_10_156 b_10 NI_10 NS_156 0 8.2034676378789059e-07
GC_10_157 b_10 NI_10 NS_157 0 3.1247846538009095e-03
GC_10_158 b_10 NI_10 NS_158 0 -3.6680387661270344e-03
GC_10_159 b_10 NI_10 NS_159 0 -1.9512084999396848e-03
GC_10_160 b_10 NI_10 NS_160 0 2.0885538930703294e-03
GC_10_161 b_10 NI_10 NS_161 0 1.3427825866401611e-04
GC_10_162 b_10 NI_10 NS_162 0 4.2675392347363664e-05
GC_10_163 b_10 NI_10 NS_163 0 2.6833776912091287e-06
GC_10_164 b_10 NI_10 NS_164 0 -6.4199301991678512e-08
GC_10_165 b_10 NI_10 NS_165 0 4.3939776092113324e-06
GC_10_166 b_10 NI_10 NS_166 0 -6.9435384285648809e-05
GC_10_167 b_10 NI_10 NS_167 0 2.0288190571394275e-06
GC_10_168 b_10 NI_10 NS_168 0 7.7012501325876717e-06
GC_10_169 b_10 NI_10 NS_169 0 -1.2189802455312481e-05
GC_10_170 b_10 NI_10 NS_170 0 -2.3754595997814303e-05
GC_10_171 b_10 NI_10 NS_171 0 -1.7232529037233308e-06
GC_10_172 b_10 NI_10 NS_172 0 2.4439492784718943e-04
GC_10_173 b_10 NI_10 NS_173 0 -1.9289596321363692e-04
GC_10_174 b_10 NI_10 NS_174 0 1.1336651881729845e-05
GC_10_175 b_10 NI_10 NS_175 0 4.5914347452882168e-05
GC_10_176 b_10 NI_10 NS_176 0 5.6879649750137864e-05
GC_10_177 b_10 NI_10 NS_177 0 4.0771973498915411e-05
GC_10_178 b_10 NI_10 NS_178 0 -5.3422053168820784e-05
GC_10_179 b_10 NI_10 NS_179 0 -7.0358329661419840e-04
GC_10_180 b_10 NI_10 NS_180 0 2.0787877769922365e-03
GC_10_181 b_10 NI_10 NS_181 0 -2.5979038424236251e-03
GC_10_182 b_10 NI_10 NS_182 0 -1.6917059050176671e-03
GC_10_183 b_10 NI_10 NS_183 0 2.4394388692881161e-04
GC_10_184 b_10 NI_10 NS_184 0 -1.8902433044394877e-03
GC_10_185 b_10 NI_10 NS_185 0 1.7570369849498278e-06
GC_10_186 b_10 NI_10 NS_186 0 6.5621977445774510e-04
GC_10_187 b_10 NI_10 NS_187 0 -7.5300677771107644e-05
GC_10_188 b_10 NI_10 NS_188 0 -1.4134034929725405e-03
GC_10_189 b_10 NI_10 NS_189 0 -5.8893405805844244e-05
GC_10_190 b_10 NI_10 NS_190 0 3.1286283695235607e-04
GC_10_191 b_10 NI_10 NS_191 0 2.7373746834281405e-04
GC_10_192 b_10 NI_10 NS_192 0 -7.2621914665483688e-05
GC_10_193 b_10 NI_10 NS_193 0 -4.7303299005427242e-04
GC_10_194 b_10 NI_10 NS_194 0 -8.6860354968302505e-05
GC_10_195 b_10 NI_10 NS_195 0 -3.6753425372701478e-05
GC_10_196 b_10 NI_10 NS_196 0 -6.1355427864174982e-06
GC_10_197 b_10 NI_10 NS_197 0 -8.7028929770445904e-05
GC_10_198 b_10 NI_10 NS_198 0 -4.5614640458031845e-05
GC_10_199 b_10 NI_10 NS_199 0 4.9433072544942429e-06
GC_10_200 b_10 NI_10 NS_200 0 5.7013348991328855e-06
GC_10_201 b_10 NI_10 NS_201 0 6.0732001898156874e-03
GC_10_202 b_10 NI_10 NS_202 0 1.7476508141068311e-03
GC_10_203 b_10 NI_10 NS_203 0 -3.6093772074787455e-03
GC_10_204 b_10 NI_10 NS_204 0 -2.1348596486256382e-03
GC_10_205 b_10 NI_10 NS_205 0 3.1621814983588612e-05
GC_10_206 b_10 NI_10 NS_206 0 5.8924596118905005e-05
GC_10_207 b_10 NI_10 NS_207 0 -1.3506942144385507e-08
GC_10_208 b_10 NI_10 NS_208 0 4.8192706716731720e-07
GC_10_209 b_10 NI_10 NS_209 0 1.4552337178345075e-05
GC_10_210 b_10 NI_10 NS_210 0 -1.0268437044772624e-05
GC_10_211 b_10 NI_10 NS_211 0 -9.9978850373308865e-07
GC_10_212 b_10 NI_10 NS_212 0 5.8136052986446978e-07
GC_10_213 b_10 NI_10 NS_213 0 4.2496792251442350e-06
GC_10_214 b_10 NI_10 NS_214 0 -2.6335934198149698e-07
GC_10_215 b_10 NI_10 NS_215 0 -9.9741770372959780e-05
GC_10_216 b_10 NI_10 NS_216 0 -1.5869860359059126e-05
GC_10_217 b_10 NI_10 NS_217 0 -1.0699217883528164e-05
GC_10_218 b_10 NI_10 NS_218 0 -4.5737371146678054e-05
GC_10_219 b_10 NI_10 NS_219 0 -7.2236696280056661e-06
GC_10_220 b_10 NI_10 NS_220 0 5.3444761754227905e-06
GC_10_221 b_10 NI_10 NS_221 0 -1.0559914108875575e-02
GC_10_222 b_10 NI_10 NS_222 0 2.0843816288957808e-05
GC_10_223 b_10 NI_10 NS_223 0 -3.3160410006673983e-04
GC_10_224 b_10 NI_10 NS_224 0 -1.8547698665162826e-03
GC_10_225 b_10 NI_10 NS_225 0 1.2558829888194986e-03
GC_10_226 b_10 NI_10 NS_226 0 -7.1109852709819177e-05
GC_10_227 b_10 NI_10 NS_227 0 6.1086631612878185e-04
GC_10_228 b_10 NI_10 NS_228 0 -1.1819412533401992e-03
GC_10_229 b_10 NI_10 NS_229 0 7.5931312693873953e-04
GC_10_230 b_10 NI_10 NS_230 0 1.6950600306764842e-04
GC_10_231 b_10 NI_10 NS_231 0 1.0237219393127851e-03
GC_10_232 b_10 NI_10 NS_232 0 5.1774325617644429e-04
GC_10_233 b_10 NI_10 NS_233 0 -1.0576257059065674e-04
GC_10_234 b_10 NI_10 NS_234 0 -8.7955211826887689e-05
GC_10_235 b_10 NI_10 NS_235 0 3.8776716427528321e-05
GC_10_236 b_10 NI_10 NS_236 0 -3.4867364586868688e-05
GC_10_237 b_10 NI_10 NS_237 0 -2.8656566598404256e-04
GC_10_238 b_10 NI_10 NS_238 0 2.5662598428814699e-04
GC_10_239 b_10 NI_10 NS_239 0 -1.5192572833023027e-05
GC_10_240 b_10 NI_10 NS_240 0 3.2850873558193242e-05
GC_10_241 b_10 NI_10 NS_241 0 -9.2917700878262672e-06
GC_10_242 b_10 NI_10 NS_242 0 1.0250305606656126e-04
GC_10_243 b_10 NI_10 NS_243 0 -5.6727872976152770e-07
GC_10_244 b_10 NI_10 NS_244 0 -2.5365804543605856e-07
GC_10_245 b_10 NI_10 NS_245 0 3.9666274569746703e-03
GC_10_246 b_10 NI_10 NS_246 0 -5.4840565659614558e-03
GC_10_247 b_10 NI_10 NS_247 0 -2.7124172157672491e-03
GC_10_248 b_10 NI_10 NS_248 0 3.3085644318644135e-03
GC_10_249 b_10 NI_10 NS_249 0 1.8443797145741258e-04
GC_10_250 b_10 NI_10 NS_250 0 -8.8841184608964317e-06
GC_10_251 b_10 NI_10 NS_251 0 3.4347412548200662e-06
GC_10_252 b_10 NI_10 NS_252 0 -2.7204144181210325e-07
GC_10_253 b_10 NI_10 NS_253 0 -3.4931913086142016e-05
GC_10_254 b_10 NI_10 NS_254 0 -8.6845363855826151e-05
GC_10_255 b_10 NI_10 NS_255 0 5.7021823891696486e-06
GC_10_256 b_10 NI_10 NS_256 0 1.1695718697363540e-05
GC_10_257 b_10 NI_10 NS_257 0 -1.7455794820947663e-05
GC_10_258 b_10 NI_10 NS_258 0 -3.6198380777829794e-05
GC_10_259 b_10 NI_10 NS_259 0 -4.1973154696148943e-05
GC_10_260 b_10 NI_10 NS_260 0 3.7033176494604293e-04
GC_10_261 b_10 NI_10 NS_261 0 -3.0302824596561918e-04
GC_10_262 b_10 NI_10 NS_262 0 3.9296931700267174e-06
GC_10_263 b_10 NI_10 NS_263 0 6.4708976052822785e-05
GC_10_264 b_10 NI_10 NS_264 0 8.3236597939825854e-05
GC_10_265 b_10 NI_10 NS_265 0 -4.1691162356842027e-03
GC_10_266 b_10 NI_10 NS_266 0 -9.7800668995835541e-05
GC_10_267 b_10 NI_10 NS_267 0 -3.4354452474853530e-03
GC_10_268 b_10 NI_10 NS_268 0 2.1023028694434243e-03
GC_10_269 b_10 NI_10 NS_269 0 -6.1026594135372590e-04
GC_10_270 b_10 NI_10 NS_270 0 -4.1004274608966067e-03
GC_10_271 b_10 NI_10 NS_271 0 1.4299878031194869e-03
GC_10_272 b_10 NI_10 NS_272 0 -1.2193512336291941e-03
GC_10_273 b_10 NI_10 NS_273 0 1.8072629887254166e-04
GC_10_274 b_10 NI_10 NS_274 0 -1.1251587944811122e-04
GC_10_275 b_10 NI_10 NS_275 0 -1.0116146447007287e-03
GC_10_276 b_10 NI_10 NS_276 0 -2.7587722375132804e-03
GC_10_277 b_10 NI_10 NS_277 0 -1.0898185725681758e-04
GC_10_278 b_10 NI_10 NS_278 0 2.2108096524689640e-04
GC_10_279 b_10 NI_10 NS_279 0 1.9213213396477053e-04
GC_10_280 b_10 NI_10 NS_280 0 -6.8711855591074673e-05
GC_10_281 b_10 NI_10 NS_281 0 -7.1607713068595009e-05
GC_10_282 b_10 NI_10 NS_282 0 -1.3686210968901885e-04
GC_10_283 b_10 NI_10 NS_283 0 -1.4114852819103171e-05
GC_10_284 b_10 NI_10 NS_284 0 -1.8759714010625125e-05
GC_10_285 b_10 NI_10 NS_285 0 -4.4744377829939573e-05
GC_10_286 b_10 NI_10 NS_286 0 -6.3879350909396961e-05
GC_10_287 b_10 NI_10 NS_287 0 3.7420373355024362e-06
GC_10_288 b_10 NI_10 NS_288 0 1.5699117063473696e-06
GC_10_289 b_10 NI_10 NS_289 0 5.9046279963277382e-03
GC_10_290 b_10 NI_10 NS_290 0 2.4577989257384483e-03
GC_10_291 b_10 NI_10 NS_291 0 -2.8030277647969476e-03
GC_10_292 b_10 NI_10 NS_292 0 -2.2213267320959043e-03
GC_10_293 b_10 NI_10 NS_293 0 5.2446601353848369e-05
GC_10_294 b_10 NI_10 NS_294 0 1.7578252686970745e-04
GC_10_295 b_10 NI_10 NS_295 0 2.4034225822471729e-07
GC_10_296 b_10 NI_10 NS_296 0 7.0788341606985493e-07
GC_10_297 b_10 NI_10 NS_297 0 4.6067688707356089e-05
GC_10_298 b_10 NI_10 NS_298 0 2.2851957796547825e-06
GC_10_299 b_10 NI_10 NS_299 0 1.3018957438942949e-06
GC_10_300 b_10 NI_10 NS_300 0 -2.1707885484591784e-07
GC_10_301 b_10 NI_10 NS_301 0 -6.8041437939083809e-07
GC_10_302 b_10 NI_10 NS_302 0 -1.3565379716992319e-06
GC_10_303 b_10 NI_10 NS_303 0 -9.4749806933027068e-05
GC_10_304 b_10 NI_10 NS_304 0 2.8698039083372188e-05
GC_10_305 b_10 NI_10 NS_305 0 -3.4791055667474841e-05
GC_10_306 b_10 NI_10 NS_306 0 -8.7737187500678439e-06
GC_10_307 b_10 NI_10 NS_307 0 3.3053766214657842e-06
GC_10_308 b_10 NI_10 NS_308 0 5.5863110921146749e-06
GC_10_309 b_10 NI_10 NS_309 0 -6.5654896695740757e-03
GC_10_310 b_10 NI_10 NS_310 0 1.4070739758940234e-05
GC_10_311 b_10 NI_10 NS_311 0 2.1104382165692162e-03
GC_10_312 b_10 NI_10 NS_312 0 -2.2927271862654263e-03
GC_10_313 b_10 NI_10 NS_313 0 -4.0182995272094226e-04
GC_10_314 b_10 NI_10 NS_314 0 2.3103511168939264e-03
GC_10_315 b_10 NI_10 NS_315 0 7.1908537375179812e-04
GC_10_316 b_10 NI_10 NS_316 0 -6.6616716591887701e-04
GC_10_317 b_10 NI_10 NS_317 0 3.8058525062556394e-04
GC_10_318 b_10 NI_10 NS_318 0 -1.0825052297319604e-04
GC_10_319 b_10 NI_10 NS_319 0 -4.1404677224828832e-04
GC_10_320 b_10 NI_10 NS_320 0 3.8833425489254045e-04
GC_10_321 b_10 NI_10 NS_321 0 -5.4546876476849035e-05
GC_10_322 b_10 NI_10 NS_322 0 -9.7045471598232650e-05
GC_10_323 b_10 NI_10 NS_323 0 2.8305771125814435e-05
GC_10_324 b_10 NI_10 NS_324 0 -4.1622894108617143e-05
GC_10_325 b_10 NI_10 NS_325 0 -1.0112047015326499e-04
GC_10_326 b_10 NI_10 NS_326 0 1.1016057188768196e-04
GC_10_327 b_10 NI_10 NS_327 0 -8.8336809976569437e-06
GC_10_328 b_10 NI_10 NS_328 0 9.4572640934553066e-06
GC_10_329 b_10 NI_10 NS_329 0 -9.9977219450091246e-06
GC_10_330 b_10 NI_10 NS_330 0 4.0459777747467740e-05
GC_10_331 b_10 NI_10 NS_331 0 -1.4669081635913441e-06
GC_10_332 b_10 NI_10 NS_332 0 2.0014075069861023e-07
GC_10_333 b_10 NI_10 NS_333 0 2.7811173274864165e-03
GC_10_334 b_10 NI_10 NS_334 0 -2.0345485694488108e-03
GC_10_335 b_10 NI_10 NS_335 0 -1.7534937851620732e-03
GC_10_336 b_10 NI_10 NS_336 0 1.0823793245748540e-03
GC_10_337 b_10 NI_10 NS_337 0 2.7883327216573482e-05
GC_10_338 b_10 NI_10 NS_338 0 -3.5939214159219278e-05
GC_10_339 b_10 NI_10 NS_339 0 1.5361131296349735e-06
GC_10_340 b_10 NI_10 NS_340 0 -2.5906415074310170e-07
GC_10_341 b_10 NI_10 NS_341 0 -2.3407525917560543e-05
GC_10_342 b_10 NI_10 NS_342 0 -1.4251665470817962e-05
GC_10_343 b_10 NI_10 NS_343 0 8.2809318641551700e-07
GC_10_344 b_10 NI_10 NS_344 0 5.2003294970826278e-06
GC_10_345 b_10 NI_10 NS_345 0 -9.2030184331909476e-06
GC_10_346 b_10 NI_10 NS_346 0 -2.1598177008953826e-05
GC_10_347 b_10 NI_10 NS_347 0 -4.5944367057763008e-05
GC_10_348 b_10 NI_10 NS_348 0 1.8296510119917783e-04
GC_10_349 b_10 NI_10 NS_349 0 -1.5583744254588430e-04
GC_10_350 b_10 NI_10 NS_350 0 -7.1629463184911996e-06
GC_10_351 b_10 NI_10 NS_351 0 2.6324116115432377e-05
GC_10_352 b_10 NI_10 NS_352 0 3.8418595726427746e-05
GC_10_353 b_10 NI_10 NS_353 0 5.0036266227614569e-02
GC_10_354 b_10 NI_10 NS_354 0 1.6071584659497158e-02
GC_10_355 b_10 NI_10 NS_355 0 -2.8776424522272723e-02
GC_10_356 b_10 NI_10 NS_356 0 1.7828641248069147e-03
GC_10_357 b_10 NI_10 NS_357 0 -2.9040846883456130e-02
GC_10_358 b_10 NI_10 NS_358 0 -9.1424757304597280e-03
GC_10_359 b_10 NI_10 NS_359 0 9.4344918295577260e-03
GC_10_360 b_10 NI_10 NS_360 0 2.6842595120579759e-03
GC_10_361 b_10 NI_10 NS_361 0 -2.8563734932085540e-03
GC_10_362 b_10 NI_10 NS_362 0 -3.3598973971372059e-04
GC_10_363 b_10 NI_10 NS_363 0 1.0950828795011109e-03
GC_10_364 b_10 NI_10 NS_364 0 -2.6817704714575791e-03
GC_10_365 b_10 NI_10 NS_365 0 -5.0250578372737476e-04
GC_10_366 b_10 NI_10 NS_366 0 9.7861125276327347e-05
GC_10_367 b_10 NI_10 NS_367 0 1.4762414045174836e-04
GC_10_368 b_10 NI_10 NS_368 0 3.6732122271088809e-05
GC_10_369 b_10 NI_10 NS_369 0 7.0511199253442999e-04
GC_10_370 b_10 NI_10 NS_370 0 -3.0702078182166380e-04
GC_10_371 b_10 NI_10 NS_371 0 2.7500133027563523e-06
GC_10_372 b_10 NI_10 NS_372 0 1.4934039353182523e-05
GC_10_373 b_10 NI_10 NS_373 0 4.4996409195210879e-06
GC_10_374 b_10 NI_10 NS_374 0 -8.3039516232035640e-06
GC_10_375 b_10 NI_10 NS_375 0 8.4537840049525100e-06
GC_10_376 b_10 NI_10 NS_376 0 6.3615405587470396e-07
GC_10_377 b_10 NI_10 NS_377 0 -3.1319721579107494e-03
GC_10_378 b_10 NI_10 NS_378 0 -3.6711192177777568e-03
GC_10_379 b_10 NI_10 NS_379 0 2.2340650113132849e-03
GC_10_380 b_10 NI_10 NS_380 0 5.4121741372653348e-04
GC_10_381 b_10 NI_10 NS_381 0 9.4495136852261954e-05
GC_10_382 b_10 NI_10 NS_382 0 -1.6044037374566427e-04
GC_10_383 b_10 NI_10 NS_383 0 9.8972455613051503e-07
GC_10_384 b_10 NI_10 NS_384 0 -6.0340054788514592e-07
GC_10_385 b_10 NI_10 NS_385 0 -3.6274103986894791e-05
GC_10_386 b_10 NI_10 NS_386 0 -5.6085242481033329e-05
GC_10_387 b_10 NI_10 NS_387 0 8.9303607888544398e-10
GC_10_388 b_10 NI_10 NS_388 0 -1.8542850472522558e-06
GC_10_389 b_10 NI_10 NS_389 0 5.5870194966708734e-06
GC_10_390 b_10 NI_10 NS_390 0 -3.0926920090944791e-06
GC_10_391 b_10 NI_10 NS_391 0 8.5765905340673756e-05
GC_10_392 b_10 NI_10 NS_392 0 9.0185910615554646e-05
GC_10_393 b_10 NI_10 NS_393 0 2.9832825597743329e-05
GC_10_394 b_10 NI_10 NS_394 0 1.8953170120894327e-05
GC_10_395 b_10 NI_10 NS_395 0 1.0780351641822897e-05
GC_10_396 b_10 NI_10 NS_396 0 -4.6450942596953974e-06
GC_10_397 b_10 NI_10 NS_397 0 -1.6285143664208182e-01
GC_10_398 b_10 NI_10 NS_398 0 1.8237558985346486e-02
GC_10_399 b_10 NI_10 NS_399 0 1.6019965954269490e-02
GC_10_400 b_10 NI_10 NS_400 0 2.0918548904769914e-03
GC_10_401 b_10 NI_10 NS_401 0 2.0892451177833248e-02
GC_10_402 b_10 NI_10 NS_402 0 -5.8848893379503664e-03
GC_10_403 b_10 NI_10 NS_403 0 6.9707216008730657e-03
GC_10_404 b_10 NI_10 NS_404 0 1.4845747421279676e-03
GC_10_405 b_10 NI_10 NS_405 0 -1.9909434367474648e-03
GC_10_406 b_10 NI_10 NS_406 0 -8.7426643319574518e-05
GC_10_407 b_10 NI_10 NS_407 0 6.8105125706824487e-03
GC_10_408 b_10 NI_10 NS_408 0 5.7377609234115787e-03
GC_10_409 b_10 NI_10 NS_409 0 3.3043045630492334e-05
GC_10_410 b_10 NI_10 NS_410 0 -2.6027854915516363e-04
GC_10_411 b_10 NI_10 NS_411 0 -4.5813951836545925e-05
GC_10_412 b_10 NI_10 NS_412 0 -8.9047775677735208e-05
GC_10_413 b_10 NI_10 NS_413 0 2.1492938933389505e-04
GC_10_414 b_10 NI_10 NS_414 0 -5.4471349733023792e-04
GC_10_415 b_10 NI_10 NS_415 0 -5.4512865511624413e-06
GC_10_416 b_10 NI_10 NS_416 0 -3.1757383585698640e-05
GC_10_417 b_10 NI_10 NS_417 0 -5.9117515949932765e-05
GC_10_418 b_10 NI_10 NS_418 0 -4.4120244828797329e-05
GC_10_419 b_10 NI_10 NS_419 0 -9.8847470004144132e-06
GC_10_420 b_10 NI_10 NS_420 0 -4.0079599688344571e-06
GC_10_421 b_10 NI_10 NS_421 0 9.0819937974154132e-03
GC_10_422 b_10 NI_10 NS_422 0 1.2351669653871165e-02
GC_10_423 b_10 NI_10 NS_423 0 -4.3131043626710814e-03
GC_10_424 b_10 NI_10 NS_424 0 -5.8690774809750899e-03
GC_10_425 b_10 NI_10 NS_425 0 -5.8189917816737721e-04
GC_10_426 b_10 NI_10 NS_426 0 1.2354785142631094e-04
GC_10_427 b_10 NI_10 NS_427 0 5.8842349741037418e-07
GC_10_428 b_10 NI_10 NS_428 0 1.9024410084464496e-06
GC_10_429 b_10 NI_10 NS_429 0 -6.6715854409222993e-05
GC_10_430 b_10 NI_10 NS_430 0 2.8039380851372324e-04
GC_10_431 b_10 NI_10 NS_431 0 -5.9815733000079076e-06
GC_10_432 b_10 NI_10 NS_432 0 -3.7208331419945186e-06
GC_10_433 b_10 NI_10 NS_433 0 -1.3951646448004750e-05
GC_10_434 b_10 NI_10 NS_434 0 -3.1580057596213002e-05
GC_10_435 b_10 NI_10 NS_435 0 -5.8765220549857077e-04
GC_10_436 b_10 NI_10 NS_436 0 2.6305254705110895e-04
GC_10_437 b_10 NI_10 NS_437 0 -3.3467466712826043e-04
GC_10_438 b_10 NI_10 NS_438 0 -7.1967089438815279e-05
GC_10_439 b_10 NI_10 NS_439 0 -5.7364050790763673e-05
GC_10_440 b_10 NI_10 NS_440 0 2.4831056354253120e-06
GC_10_441 b_10 NI_10 NS_441 0 7.7423649505788542e-03
GC_10_442 b_10 NI_10 NS_442 0 -4.1421177029182218e-04
GC_10_443 b_10 NI_10 NS_443 0 -2.0219768579471470e-02
GC_10_444 b_10 NI_10 NS_444 0 -2.7823334655723334e-03
GC_10_445 b_10 NI_10 NS_445 0 9.7982195157107470e-03
GC_10_446 b_10 NI_10 NS_446 0 -3.2789151432791566e-03
GC_10_447 b_10 NI_10 NS_447 0 6.0205679263370948e-03
GC_10_448 b_10 NI_10 NS_448 0 7.6929852060689339e-04
GC_10_449 b_10 NI_10 NS_449 0 1.3145505913622268e-03
GC_10_450 b_10 NI_10 NS_450 0 -3.6657908804324664e-04
GC_10_451 b_10 NI_10 NS_451 0 -4.3212047659798030e-04
GC_10_452 b_10 NI_10 NS_452 0 -8.5719794625248903e-03
GC_10_453 b_10 NI_10 NS_453 0 -2.6757163156710707e-04
GC_10_454 b_10 NI_10 NS_454 0 9.7079222657104570e-05
GC_10_455 b_10 NI_10 NS_455 0 2.2861118392615760e-04
GC_10_456 b_10 NI_10 NS_456 0 3.5892678263456658e-05
GC_10_457 b_10 NI_10 NS_457 0 4.8253185983199848e-04
GC_10_458 b_10 NI_10 NS_458 0 4.7333089958962935e-04
GC_10_459 b_10 NI_10 NS_459 0 4.6225701125958112e-05
GC_10_460 b_10 NI_10 NS_460 0 3.1290093999497361e-05
GC_10_461 b_10 NI_10 NS_461 0 9.5013065351021815e-05
GC_10_462 b_10 NI_10 NS_462 0 -1.5162765449756176e-05
GC_10_463 b_10 NI_10 NS_463 0 8.3740366548232160e-06
GC_10_464 b_10 NI_10 NS_464 0 -1.1811460526142630e-06
GC_10_465 b_10 NI_10 NS_465 0 -6.1970677007062089e-03
GC_10_466 b_10 NI_10 NS_466 0 1.0080227723166378e-02
GC_10_467 b_10 NI_10 NS_467 0 4.6325170788556504e-03
GC_10_468 b_10 NI_10 NS_468 0 -4.4066222670871517e-03
GC_10_469 b_10 NI_10 NS_469 0 -2.5058960723425334e-04
GC_10_470 b_10 NI_10 NS_470 0 4.6790434605366632e-05
GC_10_471 b_10 NI_10 NS_471 0 -6.6504500252296160e-07
GC_10_472 b_10 NI_10 NS_472 0 -2.2026185825336876e-07
GC_10_473 b_10 NI_10 NS_473 0 -3.7948828187904381e-05
GC_10_474 b_10 NI_10 NS_474 0 5.1815144498848845e-05
GC_10_475 b_10 NI_10 NS_475 0 -1.6266645378352961e-06
GC_10_476 b_10 NI_10 NS_476 0 9.9565523227367028e-07
GC_10_477 b_10 NI_10 NS_477 0 -3.4631624993037496e-06
GC_10_478 b_10 NI_10 NS_478 0 -1.1988003575533969e-06
GC_10_479 b_10 NI_10 NS_479 0 -4.6950534025452632e-05
GC_10_480 b_10 NI_10 NS_480 0 -1.6846558357179632e-04
GC_10_481 b_10 NI_10 NS_481 0 -8.8715353684078600e-06
GC_10_482 b_10 NI_10 NS_482 0 -3.9401083871149573e-05
GC_10_483 b_10 NI_10 NS_483 0 -7.3300224231212162e-06
GC_10_484 b_10 NI_10 NS_484 0 -1.1822118857012043e-05
GC_10_485 b_10 NI_10 NS_485 0 -9.7443421373240371e-03
GC_10_486 b_10 NI_10 NS_486 0 -9.3917171272317045e-04
GC_10_487 b_10 NI_10 NS_487 0 1.3653746597707867e-02
GC_10_488 b_10 NI_10 NS_488 0 2.7673291230055287e-03
GC_10_489 b_10 NI_10 NS_489 0 -1.5647676844075611e-02
GC_10_490 b_10 NI_10 NS_490 0 -3.6596642560931102e-03
GC_10_491 b_10 NI_10 NS_491 0 5.5280297490402563e-03
GC_10_492 b_10 NI_10 NS_492 0 -1.3324129345129187e-03
GC_10_493 b_10 NI_10 NS_493 0 -8.2810141254378552e-04
GC_10_494 b_10 NI_10 NS_494 0 6.6508459781628143e-04
GC_10_495 b_10 NI_10 NS_495 0 1.9880254564863405e-03
GC_10_496 b_10 NI_10 NS_496 0 -3.4878358547299664e-03
GC_10_497 b_10 NI_10 NS_497 0 8.6027085081741994e-05
GC_10_498 b_10 NI_10 NS_498 0 -1.3374342761635687e-04
GC_10_499 b_10 NI_10 NS_499 0 1.2614452964292485e-05
GC_10_500 b_10 NI_10 NS_500 0 -4.1222658370924556e-05
GC_10_501 b_10 NI_10 NS_501 0 9.4340971347341070e-05
GC_10_502 b_10 NI_10 NS_502 0 -8.2947552189410696e-05
GC_10_503 b_10 NI_10 NS_503 0 5.4963698761735765e-06
GC_10_504 b_10 NI_10 NS_504 0 -1.0735251088344374e-05
GC_10_505 b_10 NI_10 NS_505 0 -1.2131682052749499e-05
GC_10_506 b_10 NI_10 NS_506 0 -1.9429380574433309e-05
GC_10_507 b_10 NI_10 NS_507 0 -4.0447317534849813e-06
GC_10_508 b_10 NI_10 NS_508 0 -1.2811397566794561e-06
GC_10_509 b_10 NI_10 NS_509 0 7.3694096641510852e-03
GC_10_510 b_10 NI_10 NS_510 0 7.3632398657586615e-03
GC_10_511 b_10 NI_10 NS_511 0 -2.8316970022079879e-03
GC_10_512 b_10 NI_10 NS_512 0 -3.5561294446569210e-03
GC_10_513 b_10 NI_10 NS_513 0 -2.7050625177088832e-04
GC_10_514 b_10 NI_10 NS_514 0 6.5144461968653989e-05
GC_10_515 b_10 NI_10 NS_515 0 -3.6858897198832002e-07
GC_10_516 b_10 NI_10 NS_516 0 1.5925358445252273e-06
GC_10_517 b_10 NI_10 NS_517 0 -1.6844486625966736e-05
GC_10_518 b_10 NI_10 NS_518 0 1.3271591819052759e-04
GC_10_519 b_10 NI_10 NS_519 0 -3.0175705031601036e-06
GC_10_520 b_10 NI_10 NS_520 0 -4.7729998784489781e-07
GC_10_521 b_10 NI_10 NS_521 0 -7.0797261048913285e-06
GC_10_522 b_10 NI_10 NS_522 0 -1.8681115657960788e-05
GC_10_523 b_10 NI_10 NS_523 0 -3.2514654921891065e-04
GC_10_524 b_10 NI_10 NS_524 0 1.6915798568128466e-04
GC_10_525 b_10 NI_10 NS_525 0 -1.8429815109946950e-04
GC_10_526 b_10 NI_10 NS_526 0 -3.7599256690343430e-05
GC_10_527 b_10 NI_10 NS_527 0 -2.3736717877287472e-05
GC_10_528 b_10 NI_10 NS_528 0 9.6044429450411431e-06
GD_10_1 b_10 NI_10 NA_1 0 1.9716467045823851e-03
GD_10_2 b_10 NI_10 NA_2 0 5.2730083733370766e-03
GD_10_3 b_10 NI_10 NA_3 0 2.6616533358790632e-03
GD_10_4 b_10 NI_10 NA_4 0 5.7861508507432557e-03
GD_10_5 b_10 NI_10 NA_5 0 1.3441709675939993e-03
GD_10_6 b_10 NI_10 NA_6 0 7.5521511839730937e-03
GD_10_7 b_10 NI_10 NA_7 0 5.7785659537124600e-03
GD_10_8 b_10 NI_10 NA_8 0 3.7501335521216068e-03
GD_10_9 b_10 NI_10 NA_9 0 -1.5985849390861333e-02
GD_10_10 b_10 NI_10 NA_10 0 1.2711021440727771e-01
GD_10_11 b_10 NI_10 NA_11 0 -3.6142134607249693e-03
GD_10_12 b_10 NI_10 NA_12 0 -2.6919946647153093e-05
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 -5.2728379851417701e-03
GC_11_2 b_11 NI_11 NS_2 0 6.6652010760679943e-05
GC_11_3 b_11 NI_11 NS_3 0 -1.8650511765686464e-04
GC_11_4 b_11 NI_11 NS_4 0 -1.6783837526659245e-03
GC_11_5 b_11 NI_11 NS_5 0 1.6669619891632964e-03
GC_11_6 b_11 NI_11 NS_6 0 -3.8660493333066625e-04
GC_11_7 b_11 NI_11 NS_7 0 2.7653820693805823e-03
GC_11_8 b_11 NI_11 NS_8 0 -2.5015957562668809e-04
GC_11_9 b_11 NI_11 NS_9 0 -1.5644520405711160e-05
GC_11_10 b_11 NI_11 NS_10 0 -3.9238276287404365e-04
GC_11_11 b_11 NI_11 NS_11 0 -1.3578920610218307e-03
GC_11_12 b_11 NI_11 NS_12 0 3.8126783621759423e-03
GC_11_13 b_11 NI_11 NS_13 0 3.2378883776582751e-04
GC_11_14 b_11 NI_11 NS_14 0 -1.2353992539099347e-04
GC_11_15 b_11 NI_11 NS_15 0 2.0787701516572203e-04
GC_11_16 b_11 NI_11 NS_16 0 4.4667844758290829e-04
GC_11_17 b_11 NI_11 NS_17 0 -1.2761648388075475e-03
GC_11_18 b_11 NI_11 NS_18 0 -9.8061163894459856e-04
GC_11_19 b_11 NI_11 NS_19 0 1.1216839679869605e-04
GC_11_20 b_11 NI_11 NS_20 0 9.3592020019604580e-05
GC_11_21 b_11 NI_11 NS_21 0 -4.7341479107558955e-04
GC_11_22 b_11 NI_11 NS_22 0 2.2669963689687596e-05
GC_11_23 b_11 NI_11 NS_23 0 -5.5281583023758169e-07
GC_11_24 b_11 NI_11 NS_24 0 -1.7254423011148611e-06
GC_11_25 b_11 NI_11 NS_25 0 2.1479258693227368e-03
GC_11_26 b_11 NI_11 NS_26 0 2.2662692730013195e-03
GC_11_27 b_11 NI_11 NS_27 0 -1.3144167372661801e-03
GC_11_28 b_11 NI_11 NS_28 0 -3.3437514675794685e-03
GC_11_29 b_11 NI_11 NS_29 0 1.6784150063487615e-04
GC_11_30 b_11 NI_11 NS_30 0 -1.5986954132854975e-05
GC_11_31 b_11 NI_11 NS_31 0 2.4682982794887384e-07
GC_11_32 b_11 NI_11 NS_32 0 -6.2979471668040726e-07
GC_11_33 b_11 NI_11 NS_33 0 -1.4337043230955081e-05
GC_11_34 b_11 NI_11 NS_34 0 -7.8788469384514525e-05
GC_11_35 b_11 NI_11 NS_35 0 -2.3683908205130142e-07
GC_11_36 b_11 NI_11 NS_36 0 -2.8911465589717997e-07
GC_11_37 b_11 NI_11 NS_37 0 1.7114269742061901e-07
GC_11_38 b_11 NI_11 NS_38 0 -3.3079790040190286e-06
GC_11_39 b_11 NI_11 NS_39 0 1.9489788625289773e-04
GC_11_40 b_11 NI_11 NS_40 0 3.1959820887117539e-04
GC_11_41 b_11 NI_11 NS_41 0 -8.8378534469247031e-05
GC_11_42 b_11 NI_11 NS_42 0 5.7728659906377122e-05
GC_11_43 b_11 NI_11 NS_43 0 -6.2930208988175095e-06
GC_11_44 b_11 NI_11 NS_44 0 -3.8929526763715744e-06
GC_11_45 b_11 NI_11 NS_45 0 4.7363613247110130e-03
GC_11_46 b_11 NI_11 NS_46 0 -4.3241768768414204e-05
GC_11_47 b_11 NI_11 NS_47 0 -7.5964936883978458e-05
GC_11_48 b_11 NI_11 NS_48 0 1.5091969840032582e-03
GC_11_49 b_11 NI_11 NS_49 0 -1.7719636936819536e-03
GC_11_50 b_11 NI_11 NS_50 0 -7.6151044981315620e-04
GC_11_51 b_11 NI_11 NS_51 0 8.3298023251945821e-04
GC_11_52 b_11 NI_11 NS_52 0 -9.9704595298672686e-04
GC_11_53 b_11 NI_11 NS_53 0 1.1335302015593398e-04
GC_11_54 b_11 NI_11 NS_54 0 1.4084194661349587e-04
GC_11_55 b_11 NI_11 NS_55 0 -3.9469324108981465e-05
GC_11_56 b_11 NI_11 NS_56 0 1.2378843102865550e-03
GC_11_57 b_11 NI_11 NS_57 0 2.5020193867690394e-07
GC_11_58 b_11 NI_11 NS_58 0 1.3294696394776929e-04
GC_11_59 b_11 NI_11 NS_59 0 1.8171066811793754e-04
GC_11_60 b_11 NI_11 NS_60 0 -3.1244219555544793e-05
GC_11_61 b_11 NI_11 NS_61 0 -1.9332152614716359e-04
GC_11_62 b_11 NI_11 NS_62 0 2.7287839375830661e-04
GC_11_63 b_11 NI_11 NS_63 0 -6.9931841373851744e-07
GC_11_64 b_11 NI_11 NS_64 0 7.5432030939707905e-06
GC_11_65 b_11 NI_11 NS_65 0 3.5995035306488056e-05
GC_11_66 b_11 NI_11 NS_66 0 -6.6370412536172835e-06
GC_11_67 b_11 NI_11 NS_67 0 5.4957730258659233e-06
GC_11_68 b_11 NI_11 NS_68 0 1.6960362651073259e-06
GC_11_69 b_11 NI_11 NS_69 0 -1.8441734751117520e-03
GC_11_70 b_11 NI_11 NS_70 0 7.2547656387198455e-04
GC_11_71 b_11 NI_11 NS_71 0 8.8415464303363812e-04
GC_11_72 b_11 NI_11 NS_72 0 -7.2362249586492935e-04
GC_11_73 b_11 NI_11 NS_73 0 -1.7370537981500062e-04
GC_11_74 b_11 NI_11 NS_74 0 -2.5174035245551494e-04
GC_11_75 b_11 NI_11 NS_75 0 -1.1650132152919422e-06
GC_11_76 b_11 NI_11 NS_76 0 -1.1275636457530419e-06
GC_11_77 b_11 NI_11 NS_77 0 -5.4668740162211244e-05
GC_11_78 b_11 NI_11 NS_78 0 1.6240973990118200e-05
GC_11_79 b_11 NI_11 NS_79 0 -1.0587979381138741e-06
GC_11_80 b_11 NI_11 NS_80 0 -3.2037016820337833e-08
GC_11_81 b_11 NI_11 NS_81 0 -2.8400643513653047e-06
GC_11_82 b_11 NI_11 NS_82 0 -1.8549790021034025e-06
GC_11_83 b_11 NI_11 NS_83 0 5.7932958849730484e-05
GC_11_84 b_11 NI_11 NS_84 0 -1.1120971013701847e-04
GC_11_85 b_11 NI_11 NS_85 0 2.0166841556915886e-05
GC_11_86 b_11 NI_11 NS_86 0 -3.6151431612863485e-05
GC_11_87 b_11 NI_11 NS_87 0 5.9349068284471770e-06
GC_11_88 b_11 NI_11 NS_88 0 -6.0312211614387054e-06
GC_11_89 b_11 NI_11 NS_89 0 -8.0348016255976668e-03
GC_11_90 b_11 NI_11 NS_90 0 1.0429383636446338e-04
GC_11_91 b_11 NI_11 NS_91 0 5.9391707802447795e-04
GC_11_92 b_11 NI_11 NS_92 0 -2.3916223286921004e-03
GC_11_93 b_11 NI_11 NS_93 0 1.3647430122108639e-03
GC_11_94 b_11 NI_11 NS_94 0 1.3617959295819974e-04
GC_11_95 b_11 NI_11 NS_95 0 3.5000027138473518e-03
GC_11_96 b_11 NI_11 NS_96 0 -1.1114017620240076e-04
GC_11_97 b_11 NI_11 NS_97 0 1.4459670201111933e-04
GC_11_98 b_11 NI_11 NS_98 0 1.5316438455606867e-04
GC_11_99 b_11 NI_11 NS_99 0 -2.7995810230834312e-03
GC_11_100 b_11 NI_11 NS_100 0 3.3982189247371889e-03
GC_11_101 b_11 NI_11 NS_101 0 4.2530722700842214e-04
GC_11_102 b_11 NI_11 NS_102 0 -1.6037878302586802e-04
GC_11_103 b_11 NI_11 NS_103 0 2.9696162102115328e-04
GC_11_104 b_11 NI_11 NS_104 0 6.1054349855271892e-04
GC_11_105 b_11 NI_11 NS_105 0 -1.7227385516025626e-03
GC_11_106 b_11 NI_11 NS_106 0 -1.3974823703957323e-03
GC_11_107 b_11 NI_11 NS_107 0 1.6234919172521646e-04
GC_11_108 b_11 NI_11 NS_108 0 1.2334858519874633e-04
GC_11_109 b_11 NI_11 NS_109 0 -6.9908029337135600e-04
GC_11_110 b_11 NI_11 NS_110 0 1.9751111344504252e-05
GC_11_111 b_11 NI_11 NS_111 0 -5.8763602407358918e-07
GC_11_112 b_11 NI_11 NS_112 0 -6.5881360556853252e-08
GC_11_113 b_11 NI_11 NS_113 0 6.4245482704106387e-03
GC_11_114 b_11 NI_11 NS_114 0 4.2081817224490373e-03
GC_11_115 b_11 NI_11 NS_115 0 -3.2245895015600707e-03
GC_11_116 b_11 NI_11 NS_116 0 -6.0058478263668473e-03
GC_11_117 b_11 NI_11 NS_117 0 4.7623577950661695e-05
GC_11_118 b_11 NI_11 NS_118 0 1.9860905205647901e-04
GC_11_119 b_11 NI_11 NS_119 0 3.7434772286702537e-07
GC_11_120 b_11 NI_11 NS_120 0 -3.9527667857841418e-07
GC_11_121 b_11 NI_11 NS_121 0 -3.4600673598873627e-06
GC_11_122 b_11 NI_11 NS_122 0 -9.3206189895138664e-05
GC_11_123 b_11 NI_11 NS_123 0 1.5136865834493103e-08
GC_11_124 b_11 NI_11 NS_124 0 -2.5600280302212219e-07
GC_11_125 b_11 NI_11 NS_125 0 -1.1334647212845199e-06
GC_11_126 b_11 NI_11 NS_126 0 -3.8905051214208167e-06
GC_11_127 b_11 NI_11 NS_127 0 2.2688940327509182e-04
GC_11_128 b_11 NI_11 NS_128 0 4.1172440467007276e-04
GC_11_129 b_11 NI_11 NS_129 0 -1.3790953426106692e-04
GC_11_130 b_11 NI_11 NS_130 0 7.5855376296021372e-05
GC_11_131 b_11 NI_11 NS_131 0 -1.2034996968776307e-05
GC_11_132 b_11 NI_11 NS_132 0 -5.7495618201748750e-06
GC_11_133 b_11 NI_11 NS_133 0 1.4921896653376848e-03
GC_11_134 b_11 NI_11 NS_134 0 -7.3701568479689285e-05
GC_11_135 b_11 NI_11 NS_135 0 -1.3799814826982472e-03
GC_11_136 b_11 NI_11 NS_136 0 2.3205548654008034e-03
GC_11_137 b_11 NI_11 NS_137 0 -2.0577647646855602e-03
GC_11_138 b_11 NI_11 NS_138 0 -2.5299259057885650e-03
GC_11_139 b_11 NI_11 NS_139 0 1.2822182235882537e-03
GC_11_140 b_11 NI_11 NS_140 0 -1.4481010212281551e-03
GC_11_141 b_11 NI_11 NS_141 0 7.2089642200661566e-05
GC_11_142 b_11 NI_11 NS_142 0 2.5265585995124228e-04
GC_11_143 b_11 NI_11 NS_143 0 -7.4074317217849876e-04
GC_11_144 b_11 NI_11 NS_144 0 -2.2708897649542322e-04
GC_11_145 b_11 NI_11 NS_145 0 -6.2349947589702772e-05
GC_11_146 b_11 NI_11 NS_146 0 1.9775896212614769e-04
GC_11_147 b_11 NI_11 NS_147 0 2.1171199336411750e-04
GC_11_148 b_11 NI_11 NS_148 0 -2.2826327195561851e-05
GC_11_149 b_11 NI_11 NS_149 0 -2.4338650775554234e-04
GC_11_150 b_11 NI_11 NS_150 0 2.3359700509917591e-05
GC_11_151 b_11 NI_11 NS_151 0 -2.2076438628925655e-05
GC_11_152 b_11 NI_11 NS_152 0 -9.7713130260415342e-07
GC_11_153 b_11 NI_11 NS_153 0 -2.6245403640475611e-05
GC_11_154 b_11 NI_11 NS_154 0 -2.0576384791721053e-05
GC_11_155 b_11 NI_11 NS_155 0 2.7482735030450411e-06
GC_11_156 b_11 NI_11 NS_156 0 1.5709595852626576e-06
GC_11_157 b_11 NI_11 NS_157 0 2.4459695952422861e-03
GC_11_158 b_11 NI_11 NS_158 0 9.3397809426018052e-04
GC_11_159 b_11 NI_11 NS_159 0 -1.2354338004379904e-03
GC_11_160 b_11 NI_11 NS_160 0 -1.3629753273072384e-03
GC_11_161 b_11 NI_11 NS_161 0 -4.6651084354843366e-05
GC_11_162 b_11 NI_11 NS_162 0 -4.6352399645695897e-05
GC_11_163 b_11 NI_11 NS_163 0 -4.4755862498993779e-07
GC_11_164 b_11 NI_11 NS_164 0 -3.9746316546516276e-07
GC_11_165 b_11 NI_11 NS_165 0 -2.9955710982305087e-06
GC_11_166 b_11 NI_11 NS_166 0 -1.0244671923075927e-06
GC_11_167 b_11 NI_11 NS_167 0 -4.4739827057419619e-08
GC_11_168 b_11 NI_11 NS_168 0 1.4190673748532124e-07
GC_11_169 b_11 NI_11 NS_169 0 -1.2784652833569512e-06
GC_11_170 b_11 NI_11 NS_170 0 -1.8597080253315147e-06
GC_11_171 b_11 NI_11 NS_171 0 -7.4426597112023350e-06
GC_11_172 b_11 NI_11 NS_172 0 -2.4977904503347013e-05
GC_11_173 b_11 NI_11 NS_173 0 3.7800083238703306e-06
GC_11_174 b_11 NI_11 NS_174 0 -1.3306520796267974e-05
GC_11_175 b_11 NI_11 NS_175 0 7.0591667677479152e-06
GC_11_176 b_11 NI_11 NS_176 0 7.2630885012150016e-07
GC_11_177 b_11 NI_11 NS_177 0 -7.5740530056826018e-03
GC_11_178 b_11 NI_11 NS_178 0 4.6628792659291687e-05
GC_11_179 b_11 NI_11 NS_179 0 1.9120424654356788e-03
GC_11_180 b_11 NI_11 NS_180 0 -1.5857972592640888e-03
GC_11_181 b_11 NI_11 NS_181 0 -1.1333027495979225e-03
GC_11_182 b_11 NI_11 NS_182 0 6.7014673491507665e-04
GC_11_183 b_11 NI_11 NS_183 0 2.4906704766534905e-03
GC_11_184 b_11 NI_11 NS_184 0 -6.4707425706144099e-05
GC_11_185 b_11 NI_11 NS_185 0 2.1093494274116286e-04
GC_11_186 b_11 NI_11 NS_186 0 8.1204703072573748e-04
GC_11_187 b_11 NI_11 NS_187 0 -3.3539868012668820e-03
GC_11_188 b_11 NI_11 NS_188 0 1.2068615864027568e-04
GC_11_189 b_11 NI_11 NS_189 0 4.2555997092497605e-04
GC_11_190 b_11 NI_11 NS_190 0 -1.7587611308961883e-04
GC_11_191 b_11 NI_11 NS_191 0 2.9436829290275406e-04
GC_11_192 b_11 NI_11 NS_192 0 6.1362507272141821e-04
GC_11_193 b_11 NI_11 NS_193 0 -1.6006799026691363e-03
GC_11_194 b_11 NI_11 NS_194 0 -1.4593086028118845e-03
GC_11_195 b_11 NI_11 NS_195 0 1.6731670520660127e-04
GC_11_196 b_11 NI_11 NS_196 0 1.2458632753310078e-04
GC_11_197 b_11 NI_11 NS_197 0 -6.7420663220479633e-04
GC_11_198 b_11 NI_11 NS_198 0 9.2119959804397002e-06
GC_11_199 b_11 NI_11 NS_199 0 -4.2469367752230399e-06
GC_11_200 b_11 NI_11 NS_200 0 -1.3434627149928545e-06
GC_11_201 b_11 NI_11 NS_201 0 9.2624482964949999e-03
GC_11_202 b_11 NI_11 NS_202 0 5.1206901426344084e-03
GC_11_203 b_11 NI_11 NS_203 0 -3.7979299271310081e-03
GC_11_204 b_11 NI_11 NS_204 0 -6.8446989339165020e-03
GC_11_205 b_11 NI_11 NS_205 0 -1.1424471249193916e-04
GC_11_206 b_11 NI_11 NS_206 0 3.3269716955656038e-04
GC_11_207 b_11 NI_11 NS_207 0 3.1697470688490870e-07
GC_11_208 b_11 NI_11 NS_208 0 5.6517218518678864e-08
GC_11_209 b_11 NI_11 NS_209 0 9.5350625059001557e-06
GC_11_210 b_11 NI_11 NS_210 0 -8.0270523981741502e-05
GC_11_211 b_11 NI_11 NS_211 0 4.4899288275554913e-07
GC_11_212 b_11 NI_11 NS_212 0 2.4706850581858511e-07
GC_11_213 b_11 NI_11 NS_213 0 1.8223765412337158e-07
GC_11_214 b_11 NI_11 NS_214 0 -2.3335350698972771e-06
GC_11_215 b_11 NI_11 NS_215 0 1.4808791392208445e-04
GC_11_216 b_11 NI_11 NS_216 0 4.5714727759493850e-04
GC_11_217 b_11 NI_11 NS_217 0 -1.4396786532963509e-04
GC_11_218 b_11 NI_11 NS_218 0 6.2618425750550160e-05
GC_11_219 b_11 NI_11 NS_219 0 -1.5086878181403018e-05
GC_11_220 b_11 NI_11 NS_220 0 -5.0400774213097849e-06
GC_11_221 b_11 NI_11 NS_221 0 -4.6147298263046286e-03
GC_11_222 b_11 NI_11 NS_222 0 -9.1507982483833008e-05
GC_11_223 b_11 NI_11 NS_223 0 -3.4538995597093386e-03
GC_11_224 b_11 NI_11 NS_224 0 2.0673691360282970e-03
GC_11_225 b_11 NI_11 NS_225 0 -5.8284116660276724e-04
GC_11_226 b_11 NI_11 NS_226 0 -4.1404342208971722e-03
GC_11_227 b_11 NI_11 NS_227 0 1.4316771262851424e-03
GC_11_228 b_11 NI_11 NS_228 0 -1.2519594612106528e-03
GC_11_229 b_11 NI_11 NS_229 0 2.6670833434077338e-04
GC_11_230 b_11 NI_11 NS_230 0 -8.4215514877552441e-06
GC_11_231 b_11 NI_11 NS_231 0 -1.0216583821127216e-03
GC_11_232 b_11 NI_11 NS_232 0 -2.8396194224712340e-03
GC_11_233 b_11 NI_11 NS_233 0 -1.0674678049317883e-04
GC_11_234 b_11 NI_11 NS_234 0 2.2366888654649821e-04
GC_11_235 b_11 NI_11 NS_235 0 1.9107917520208039e-04
GC_11_236 b_11 NI_11 NS_236 0 -6.5344362238989377e-05
GC_11_237 b_11 NI_11 NS_237 0 -9.1262700151008440e-05
GC_11_238 b_11 NI_11 NS_238 0 -1.4993492801840274e-04
GC_11_239 b_11 NI_11 NS_239 0 -1.6403030620490236e-05
GC_11_240 b_11 NI_11 NS_240 0 -1.8273693849286124e-05
GC_11_241 b_11 NI_11 NS_241 0 -4.9930957324118915e-05
GC_11_242 b_11 NI_11 NS_242 0 -6.2139820596125646e-05
GC_11_243 b_11 NI_11 NS_243 0 3.5330616217344916e-06
GC_11_244 b_11 NI_11 NS_244 0 1.6964493760195583e-06
GC_11_245 b_11 NI_11 NS_245 0 6.2934678356170457e-03
GC_11_246 b_11 NI_11 NS_246 0 2.1224042927904720e-03
GC_11_247 b_11 NI_11 NS_247 0 -3.0165293495980185e-03
GC_11_248 b_11 NI_11 NS_248 0 -2.0750248415261981e-03
GC_11_249 b_11 NI_11 NS_249 0 7.1025223875438226e-05
GC_11_250 b_11 NI_11 NS_250 0 2.0943215080853757e-04
GC_11_251 b_11 NI_11 NS_251 0 3.3258300127647924e-07
GC_11_252 b_11 NI_11 NS_252 0 8.7719277560936534e-07
GC_11_253 b_11 NI_11 NS_253 0 5.4092566814904355e-05
GC_11_254 b_11 NI_11 NS_254 0 -1.1669013086196485e-06
GC_11_255 b_11 NI_11 NS_255 0 1.8059205099184407e-06
GC_11_256 b_11 NI_11 NS_256 0 -3.4863155656322392e-07
GC_11_257 b_11 NI_11 NS_257 0 -5.1640227808551417e-07
GC_11_258 b_11 NI_11 NS_258 0 -1.6096646465375310e-06
GC_11_259 b_11 NI_11 NS_259 0 -9.3868188881648864e-05
GC_11_260 b_11 NI_11 NS_260 0 4.8865629715467630e-05
GC_11_261 b_11 NI_11 NS_261 0 -3.8746122828526834e-05
GC_11_262 b_11 NI_11 NS_262 0 -1.3114751928970401e-06
GC_11_263 b_11 NI_11 NS_263 0 4.4417562018517596e-06
GC_11_264 b_11 NI_11 NS_264 0 6.8494639327606731e-06
GC_11_265 b_11 NI_11 NS_265 0 -6.0603592032644526e-03
GC_11_266 b_11 NI_11 NS_266 0 -2.1312935981620138e-04
GC_11_267 b_11 NI_11 NS_267 0 2.4418368838898144e-03
GC_11_268 b_11 NI_11 NS_268 0 1.7985969645023675e-03
GC_11_269 b_11 NI_11 NS_269 0 -3.8803098350916384e-03
GC_11_270 b_11 NI_11 NS_270 0 -4.1123799700745079e-03
GC_11_271 b_11 NI_11 NS_271 0 2.4221469032116535e-03
GC_11_272 b_11 NI_11 NS_272 0 3.6138305580554319e-04
GC_11_273 b_11 NI_11 NS_273 0 1.4371147985464596e-04
GC_11_274 b_11 NI_11 NS_274 0 -4.4032904818843349e-04
GC_11_275 b_11 NI_11 NS_275 0 8.5390369759872264e-04
GC_11_276 b_11 NI_11 NS_276 0 -1.4662076137503450e-03
GC_11_277 b_11 NI_11 NS_277 0 2.9759000795817760e-04
GC_11_278 b_11 NI_11 NS_278 0 -5.8796034275009430e-05
GC_11_279 b_11 NI_11 NS_279 0 2.1005013221668097e-04
GC_11_280 b_11 NI_11 NS_280 0 4.4514685835448043e-04
GC_11_281 b_11 NI_11 NS_281 0 -1.0977214127254002e-03
GC_11_282 b_11 NI_11 NS_282 0 -9.2864250975413932e-04
GC_11_283 b_11 NI_11 NS_283 0 1.3465509120811985e-04
GC_11_284 b_11 NI_11 NS_284 0 9.7802956017739985e-05
GC_11_285 b_11 NI_11 NS_285 0 -4.4566627387795823e-04
GC_11_286 b_11 NI_11 NS_286 0 5.5649764901201103e-06
GC_11_287 b_11 NI_11 NS_287 0 -8.0918160373166493e-07
GC_11_288 b_11 NI_11 NS_288 0 -5.0393010720367458e-07
GC_11_289 b_11 NI_11 NS_289 0 4.1119240075794946e-03
GC_11_290 b_11 NI_11 NS_290 0 6.8603493682720829e-03
GC_11_291 b_11 NI_11 NS_291 0 -7.2764908892541935e-04
GC_11_292 b_11 NI_11 NS_292 0 -5.7931892338283610e-03
GC_11_293 b_11 NI_11 NS_293 0 -3.5775308651608573e-04
GC_11_294 b_11 NI_11 NS_294 0 3.8834911402999028e-04
GC_11_295 b_11 NI_11 NS_295 0 9.4512421664274787e-08
GC_11_296 b_11 NI_11 NS_296 0 4.5738255391522130e-07
GC_11_297 b_11 NI_11 NS_297 0 2.6844694184327686e-05
GC_11_298 b_11 NI_11 NS_298 0 -2.2194802683343514e-05
GC_11_299 b_11 NI_11 NS_299 0 3.3931998008736010e-07
GC_11_300 b_11 NI_11 NS_300 0 6.9561053447628625e-07
GC_11_301 b_11 NI_11 NS_301 0 -1.4718253902625900e-06
GC_11_302 b_11 NI_11 NS_302 0 -9.8770241655272369e-07
GC_11_303 b_11 NI_11 NS_303 0 5.9106733586458546e-05
GC_11_304 b_11 NI_11 NS_304 0 2.3858333840167713e-04
GC_11_305 b_11 NI_11 NS_305 0 -1.0408464158217611e-04
GC_11_306 b_11 NI_11 NS_306 0 2.0899988973954506e-05
GC_11_307 b_11 NI_11 NS_307 0 -1.4386399320209171e-05
GC_11_308 b_11 NI_11 NS_308 0 -5.7818104663779570e-06
GC_11_309 b_11 NI_11 NS_309 0 -7.2805286979607748e-04
GC_11_310 b_11 NI_11 NS_310 0 -1.0592867708821375e-04
GC_11_311 b_11 NI_11 NS_311 0 -5.6660594162066848e-03
GC_11_312 b_11 NI_11 NS_312 0 -9.1823177327914507e-04
GC_11_313 b_11 NI_11 NS_313 0 2.1705414359743276e-03
GC_11_314 b_11 NI_11 NS_314 0 -4.1311994997401459e-04
GC_11_315 b_11 NI_11 NS_315 0 6.6842937432287110e-04
GC_11_316 b_11 NI_11 NS_316 0 -4.6299382282495490e-04
GC_11_317 b_11 NI_11 NS_317 0 8.4566392280101970e-04
GC_11_318 b_11 NI_11 NS_318 0 2.3034670944366948e-04
GC_11_319 b_11 NI_11 NS_319 0 6.2427406936098741e-04
GC_11_320 b_11 NI_11 NS_320 0 -4.4556831061231461e-03
GC_11_321 b_11 NI_11 NS_321 0 -1.3745598398042088e-04
GC_11_322 b_11 NI_11 NS_322 0 1.5070338868868879e-04
GC_11_323 b_11 NI_11 NS_323 0 1.5406557710498082e-04
GC_11_324 b_11 NI_11 NS_324 0 -2.7668304018835477e-05
GC_11_325 b_11 NI_11 NS_325 0 -7.6293647452227664e-05
GC_11_326 b_11 NI_11 NS_326 0 -3.3923979180423810e-05
GC_11_327 b_11 NI_11 NS_327 0 -1.8395520540945986e-05
GC_11_328 b_11 NI_11 NS_328 0 -1.0688579017046462e-05
GC_11_329 b_11 NI_11 NS_329 0 -1.7353200145248270e-05
GC_11_330 b_11 NI_11 NS_330 0 -2.8379848114276000e-05
GC_11_331 b_11 NI_11 NS_331 0 2.0420192581257461e-06
GC_11_332 b_11 NI_11 NS_332 0 4.1574867662730012e-07
GC_11_333 b_11 NI_11 NS_333 0 1.5056720964572634e-03
GC_11_334 b_11 NI_11 NS_334 0 3.2374092983133112e-03
GC_11_335 b_11 NI_11 NS_335 0 -6.9847109796628232e-04
GC_11_336 b_11 NI_11 NS_336 0 -1.7851805218004179e-03
GC_11_337 b_11 NI_11 NS_337 0 3.3018846141791176e-05
GC_11_338 b_11 NI_11 NS_338 0 1.7319109542155009e-04
GC_11_339 b_11 NI_11 NS_339 0 1.6094935855999952e-07
GC_11_340 b_11 NI_11 NS_340 0 3.1376557243468456e-07
GC_11_341 b_11 NI_11 NS_341 0 3.3999313319877446e-05
GC_11_342 b_11 NI_11 NS_342 0 4.2129591277557370e-06
GC_11_343 b_11 NI_11 NS_343 0 6.5827951778850216e-07
GC_11_344 b_11 NI_11 NS_344 0 3.1769739621310123e-07
GC_11_345 b_11 NI_11 NS_345 0 -6.6327387526029011e-07
GC_11_346 b_11 NI_11 NS_346 0 -8.7826448050154624e-07
GC_11_347 b_11 NI_11 NS_347 0 -7.3533624121276011e-05
GC_11_348 b_11 NI_11 NS_348 0 -3.0345372253659465e-05
GC_11_349 b_11 NI_11 NS_349 0 -1.2848234746738474e-05
GC_11_350 b_11 NI_11 NS_350 0 -8.9770545011097992e-06
GC_11_351 b_11 NI_11 NS_351 0 2.2219855354917986e-06
GC_11_352 b_11 NI_11 NS_352 0 1.9794130799202600e-06
GC_11_353 b_11 NI_11 NS_353 0 1.1922627028372230e-02
GC_11_354 b_11 NI_11 NS_354 0 -6.5844195732136178e-04
GC_11_355 b_11 NI_11 NS_355 0 1.1369832599582552e-02
GC_11_356 b_11 NI_11 NS_356 0 4.1780408700608593e-03
GC_11_357 b_11 NI_11 NS_357 0 -9.7949700493272281e-03
GC_11_358 b_11 NI_11 NS_358 0 -8.3145698846085452e-03
GC_11_359 b_11 NI_11 NS_359 0 1.1198762804449413e-02
GC_11_360 b_11 NI_11 NS_360 0 6.9171363062516021e-03
GC_11_361 b_11 NI_11 NS_361 0 -3.0683196859490457e-03
GC_11_362 b_11 NI_11 NS_362 0 -2.5359853970908222e-03
GC_11_363 b_11 NI_11 NS_363 0 2.3248066546639702e-03
GC_11_364 b_11 NI_11 NS_364 0 3.8909047096627224e-03
GC_11_365 b_11 NI_11 NS_365 0 5.8142716380973490e-04
GC_11_366 b_11 NI_11 NS_366 0 3.4308214082466804e-04
GC_11_367 b_11 NI_11 NS_367 0 1.6421752533917855e-04
GC_11_368 b_11 NI_11 NS_368 0 3.3136555069084126e-04
GC_11_369 b_11 NI_11 NS_369 0 8.5588573610017845e-04
GC_11_370 b_11 NI_11 NS_370 0 1.6013636999610644e-04
GC_11_371 b_11 NI_11 NS_371 0 2.1246444548418580e-04
GC_11_372 b_11 NI_11 NS_372 0 1.8332738046135841e-04
GC_11_373 b_11 NI_11 NS_373 0 1.4584430503428172e-04
GC_11_374 b_11 NI_11 NS_374 0 4.7664821618507858e-05
GC_11_375 b_11 NI_11 NS_375 0 -5.3882975873424795e-06
GC_11_376 b_11 NI_11 NS_376 0 1.2511407388761412e-06
GC_11_377 b_11 NI_11 NS_377 0 -2.2779904017134759e-02
GC_11_378 b_11 NI_11 NS_378 0 1.0554424335505526e-02
GC_11_379 b_11 NI_11 NS_379 0 1.5573795652921702e-02
GC_11_380 b_11 NI_11 NS_380 0 -1.1837445138585883e-03
GC_11_381 b_11 NI_11 NS_381 0 -4.1324616077270324e-04
GC_11_382 b_11 NI_11 NS_382 0 -4.4059545533330346e-04
GC_11_383 b_11 NI_11 NS_383 0 6.9442206438359662e-07
GC_11_384 b_11 NI_11 NS_384 0 -2.3556084832419043e-07
GC_11_385 b_11 NI_11 NS_385 0 7.0284308372970707e-05
GC_11_386 b_11 NI_11 NS_386 0 -4.3043808869497377e-05
GC_11_387 b_11 NI_11 NS_387 0 1.1118405249037307e-06
GC_11_388 b_11 NI_11 NS_388 0 1.0051844965364726e-06
GC_11_389 b_11 NI_11 NS_389 0 -3.0885202042634367e-06
GC_11_390 b_11 NI_11 NS_390 0 -2.8306337455314598e-07
GC_11_391 b_11 NI_11 NS_391 0 -7.6137090615126669e-05
GC_11_392 b_11 NI_11 NS_392 0 1.4218921465652766e-04
GC_11_393 b_11 NI_11 NS_393 0 -9.1712066797929844e-06
GC_11_394 b_11 NI_11 NS_394 0 -8.2462677603552571e-05
GC_11_395 b_11 NI_11 NS_395 0 -1.8755641146993362e-05
GC_11_396 b_11 NI_11 NS_396 0 -8.2807764409940292e-06
GC_11_397 b_11 NI_11 NS_397 0 7.7423649505896234e-03
GC_11_398 b_11 NI_11 NS_398 0 -4.1421177029187471e-04
GC_11_399 b_11 NI_11 NS_399 0 -2.0219768579470762e-02
GC_11_400 b_11 NI_11 NS_400 0 -2.7823334655715922e-03
GC_11_401 b_11 NI_11 NS_401 0 9.7982195157099074e-03
GC_11_402 b_11 NI_11 NS_402 0 -3.2789151432782737e-03
GC_11_403 b_11 NI_11 NS_403 0 6.0205679263368875e-03
GC_11_404 b_11 NI_11 NS_404 0 7.6929852060716899e-04
GC_11_405 b_11 NI_11 NS_405 0 1.3145505913615988e-03
GC_11_406 b_11 NI_11 NS_406 0 -3.6657908804202388e-04
GC_11_407 b_11 NI_11 NS_407 0 -4.3212047659777338e-04
GC_11_408 b_11 NI_11 NS_408 0 -8.5719794625244618e-03
GC_11_409 b_11 NI_11 NS_409 0 -2.6757163156709948e-04
GC_11_410 b_11 NI_11 NS_410 0 9.7079222657102239e-05
GC_11_411 b_11 NI_11 NS_411 0 2.2861118392611800e-04
GC_11_412 b_11 NI_11 NS_412 0 3.5892678263436207e-05
GC_11_413 b_11 NI_11 NS_413 0 4.8253185983221039e-04
GC_11_414 b_11 NI_11 NS_414 0 4.7333089958944080e-04
GC_11_415 b_11 NI_11 NS_415 0 4.6225701125957638e-05
GC_11_416 b_11 NI_11 NS_416 0 3.1290093999439397e-05
GC_11_417 b_11 NI_11 NS_417 0 9.5013065351069357e-05
GC_11_418 b_11 NI_11 NS_418 0 -1.5162765449941975e-05
GC_11_419 b_11 NI_11 NS_419 0 8.3740366548445088e-06
GC_11_420 b_11 NI_11 NS_420 0 -1.1811460526317656e-06
GC_11_421 b_11 NI_11 NS_421 0 -6.1970677007095864e-03
GC_11_422 b_11 NI_11 NS_422 0 1.0080227723170868e-02
GC_11_423 b_11 NI_11 NS_423 0 4.6325170788585378e-03
GC_11_424 b_11 NI_11 NS_424 0 -4.4066222670894996e-03
GC_11_425 b_11 NI_11 NS_425 0 -2.5058960723419469e-04
GC_11_426 b_11 NI_11 NS_426 0 4.6790434605361327e-05
GC_11_427 b_11 NI_11 NS_427 0 -6.6504500252201684e-07
GC_11_428 b_11 NI_11 NS_428 0 -2.2026185825413975e-07
GC_11_429 b_11 NI_11 NS_429 0 -3.7948828187924513e-05
GC_11_430 b_11 NI_11 NS_430 0 5.1815144498815892e-05
GC_11_431 b_11 NI_11 NS_431 0 -1.6266645378367460e-06
GC_11_432 b_11 NI_11 NS_432 0 9.9565523227259159e-07
GC_11_433 b_11 NI_11 NS_433 0 -3.4631624993050273e-06
GC_11_434 b_11 NI_11 NS_434 0 -1.1988003575571484e-06
GC_11_435 b_11 NI_11 NS_435 0 -4.6950534025322555e-05
GC_11_436 b_11 NI_11 NS_436 0 -1.6846558357187848e-04
GC_11_437 b_11 NI_11 NS_437 0 -8.8715353683818544e-06
GC_11_438 b_11 NI_11 NS_438 0 -3.9401083871163789e-05
GC_11_439 b_11 NI_11 NS_439 0 -7.3300224231231525e-06
GC_11_440 b_11 NI_11 NS_440 0 -1.1822118857016239e-05
GC_11_441 b_11 NI_11 NS_441 0 -1.4532339503637862e-02
GC_11_442 b_11 NI_11 NS_442 0 1.3254324425956686e-02
GC_11_443 b_11 NI_11 NS_443 0 4.6508562342144405e-03
GC_11_444 b_11 NI_11 NS_444 0 1.0943906627766542e-02
GC_11_445 b_11 NI_11 NS_445 0 1.5396302178797698e-02
GC_11_446 b_11 NI_11 NS_446 0 -8.2779988038482830e-03
GC_11_447 b_11 NI_11 NS_447 0 4.6168368362145872e-03
GC_11_448 b_11 NI_11 NS_448 0 5.3473913877081962e-03
GC_11_449 b_11 NI_11 NS_449 0 2.8763253980888357e-03
GC_11_450 b_11 NI_11 NS_450 0 3.6813361022614540e-03
GC_11_451 b_11 NI_11 NS_451 0 7.5462206187061377e-03
GC_11_452 b_11 NI_11 NS_452 0 1.0423413198144323e-02
GC_11_453 b_11 NI_11 NS_453 0 3.3135833236784133e-04
GC_11_454 b_11 NI_11 NS_454 0 1.0639138259965358e-04
GC_11_455 b_11 NI_11 NS_455 0 6.6283383752329422e-05
GC_11_456 b_11 NI_11 NS_456 0 2.0084392743731537e-04
GC_11_457 b_11 NI_11 NS_457 0 7.7808513345446414e-04
GC_11_458 b_11 NI_11 NS_458 0 -6.6065867055376969e-04
GC_11_459 b_11 NI_11 NS_459 0 1.5059942974481912e-04
GC_11_460 b_11 NI_11 NS_460 0 7.6441776517269860e-05
GC_11_461 b_11 NI_11 NS_461 0 -3.5091679969689604e-05
GC_11_462 b_11 NI_11 NS_462 0 -6.7307417666383031e-05
GC_11_463 b_11 NI_11 NS_463 0 -6.1381264005303898e-06
GC_11_464 b_11 NI_11 NS_464 0 -1.7307987117937475e-06
GC_11_465 b_11 NI_11 NS_465 0 -5.4836899158434132e-03
GC_11_466 b_11 NI_11 NS_466 0 8.6219828262390930e-03
GC_11_467 b_11 NI_11 NS_467 0 5.9454907065339515e-03
GC_11_468 b_11 NI_11 NS_468 0 -3.1620951184483628e-03
GC_11_469 b_11 NI_11 NS_469 0 -4.9322130653768311e-04
GC_11_470 b_11 NI_11 NS_470 0 2.5095536539080992e-04
GC_11_471 b_11 NI_11 NS_471 0 8.5577829005835384e-07
GC_11_472 b_11 NI_11 NS_472 0 2.6051782759537495e-06
GC_11_473 b_11 NI_11 NS_473 0 1.4510373656742510e-04
GC_11_474 b_11 NI_11 NS_474 0 1.5602656448974176e-05
GC_11_475 b_11 NI_11 NS_475 0 2.8317479838257818e-06
GC_11_476 b_11 NI_11 NS_476 0 1.7221576831741541e-06
GC_11_477 b_11 NI_11 NS_477 0 1.5306322801480445e-07
GC_11_478 b_11 NI_11 NS_478 0 1.8737153991071171e-06
GC_11_479 b_11 NI_11 NS_479 0 -2.2253468049318568e-04
GC_11_480 b_11 NI_11 NS_480 0 2.1076576801344173e-04
GC_11_481 b_11 NI_11 NS_481 0 -7.4247080061344282e-05
GC_11_482 b_11 NI_11 NS_482 0 -4.4382564271589045e-05
GC_11_483 b_11 NI_11 NS_483 0 -2.2488891117334205e-05
GC_11_484 b_11 NI_11 NS_484 0 3.9334169342261063e-06
GC_11_485 b_11 NI_11 NS_485 0 3.5289009065834445e-02
GC_11_486 b_11 NI_11 NS_486 0 1.6497220761543814e-02
GC_11_487 b_11 NI_11 NS_487 0 -1.9435780531238289e-02
GC_11_488 b_11 NI_11 NS_488 0 -5.4527637852413036e-03
GC_11_489 b_11 NI_11 NS_489 0 -2.8214541330258500e-02
GC_11_490 b_11 NI_11 NS_490 0 1.8345572205476046e-03
GC_11_491 b_11 NI_11 NS_491 0 2.2404843324811325e-03
GC_11_492 b_11 NI_11 NS_492 0 2.0288883484081968e-03
GC_11_493 b_11 NI_11 NS_493 0 -2.0527313855253013e-03
GC_11_494 b_11 NI_11 NS_494 0 2.8472531335597989e-04
GC_11_495 b_11 NI_11 NS_495 0 7.7524789725776739e-03
GC_11_496 b_11 NI_11 NS_496 0 -3.1287535393299520e-03
GC_11_497 b_11 NI_11 NS_497 0 -3.2243079627035674e-04
GC_11_498 b_11 NI_11 NS_498 0 3.0820890158032158e-05
GC_11_499 b_11 NI_11 NS_499 0 8.3139366925157946e-05
GC_11_500 b_11 NI_11 NS_500 0 4.0063819736194166e-06
GC_11_501 b_11 NI_11 NS_501 0 2.1977055600900738e-04
GC_11_502 b_11 NI_11 NS_502 0 -3.1180510498754103e-04
GC_11_503 b_11 NI_11 NS_503 0 -2.4613569795752457e-05
GC_11_504 b_11 NI_11 NS_504 0 2.3386335034088721e-06
GC_11_505 b_11 NI_11 NS_505 0 -3.9831538056396074e-05
GC_11_506 b_11 NI_11 NS_506 0 1.2518458529314694e-05
GC_11_507 b_11 NI_11 NS_507 0 2.0022389966710403e-06
GC_11_508 b_11 NI_11 NS_508 0 1.7019165922317503e-06
GC_11_509 b_11 NI_11 NS_509 0 -2.9014008520246385e-03
GC_11_510 b_11 NI_11 NS_510 0 -5.7720493218731458e-03
GC_11_511 b_11 NI_11 NS_511 0 8.0019278083641378e-04
GC_11_512 b_11 NI_11 NS_512 0 1.9977889641012649e-03
GC_11_513 b_11 NI_11 NS_513 0 9.8428082168193026e-05
GC_11_514 b_11 NI_11 NS_514 0 -8.8303314472519908e-05
GC_11_515 b_11 NI_11 NS_515 0 9.9704799204156260e-07
GC_11_516 b_11 NI_11 NS_516 0 -7.6665139017412495e-07
GC_11_517 b_11 NI_11 NS_517 0 -2.7720280552699096e-05
GC_11_518 b_11 NI_11 NS_518 0 -3.9678392029073797e-05
GC_11_519 b_11 NI_11 NS_519 0 -9.1732628212781244e-07
GC_11_520 b_11 NI_11 NS_520 0 -9.2002787784369923e-07
GC_11_521 b_11 NI_11 NS_521 0 -5.5606228845199452e-07
GC_11_522 b_11 NI_11 NS_522 0 -3.3394989048881354e-06
GC_11_523 b_11 NI_11 NS_523 0 1.0094568902177828e-04
GC_11_524 b_11 NI_11 NS_524 0 3.5941077296052717e-05
GC_11_525 b_11 NI_11 NS_525 0 2.2153910114390016e-05
GC_11_526 b_11 NI_11 NS_526 0 1.9573523786080400e-05
GC_11_527 b_11 NI_11 NS_527 0 8.1250895541731652e-06
GC_11_528 b_11 NI_11 NS_528 0 -3.1397916808061046e-06
GD_11_1 b_11 NI_11 NA_1 0 2.8504604616419659e-03
GD_11_2 b_11 NI_11 NA_2 0 -3.1761320459139960e-03
GD_11_3 b_11 NI_11 NA_3 0 3.4474710667347242e-03
GD_11_4 b_11 NI_11 NA_4 0 5.7763564577938522e-04
GD_11_5 b_11 NI_11 NA_5 0 3.1059682420099713e-03
GD_11_6 b_11 NI_11 NA_6 0 5.8234355331974541e-03
GD_11_7 b_11 NI_11 NA_7 0 1.5364429252729846e-03
GD_11_8 b_11 NI_11 NA_8 0 1.4948353692672289e-03
GD_11_9 b_11 NI_11 NA_9 0 -2.1286062301490827e-02
GD_11_10 b_11 NI_11 NA_10 0 -3.6142134607399711e-03
GD_11_11 b_11 NI_11 NA_11 0 -1.6684357351320483e-01
GD_11_12 b_11 NI_11 NA_12 0 -9.1444686992623436e-03
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 4.8531323671998083e-03
GC_12_2 b_12 NI_12 NS_2 0 -4.3649876182217649e-05
GC_12_3 b_12 NI_12 NS_3 0 -6.6864802960923950e-05
GC_12_4 b_12 NI_12 NS_4 0 1.5061862253039899e-03
GC_12_5 b_12 NI_12 NS_5 0 -1.7559778821086764e-03
GC_12_6 b_12 NI_12 NS_6 0 -7.3998463627255402e-04
GC_12_7 b_12 NI_12 NS_7 0 8.2701923893396161e-04
GC_12_8 b_12 NI_12 NS_8 0 -9.5862125467594851e-04
GC_12_9 b_12 NI_12 NS_9 0 2.8332973985069090e-05
GC_12_10 b_12 NI_12 NS_10 0 6.3430913104054343e-05
GC_12_11 b_12 NI_12 NS_11 0 -7.5167401952286688e-05
GC_12_12 b_12 NI_12 NS_12 0 1.2237696843840219e-03
GC_12_13 b_12 NI_12 NS_13 0 3.1295802906695642e-06
GC_12_14 b_12 NI_12 NS_14 0 1.3610040821244673e-04
GC_12_15 b_12 NI_12 NS_15 0 1.8544849033467131e-04
GC_12_16 b_12 NI_12 NS_16 0 -1.1512465199294560e-05
GC_12_17 b_12 NI_12 NS_17 0 -2.2096326155143873e-04
GC_12_18 b_12 NI_12 NS_18 0 2.0637401549826443e-04
GC_12_19 b_12 NI_12 NS_19 0 -4.5355204772751033e-06
GC_12_20 b_12 NI_12 NS_20 0 7.2572664302132180e-06
GC_12_21 b_12 NI_12 NS_21 0 2.1469900450834580e-05
GC_12_22 b_12 NI_12 NS_22 0 -6.1794067795413453e-06
GC_12_23 b_12 NI_12 NS_23 0 4.1879283530554900e-06
GC_12_24 b_12 NI_12 NS_24 0 1.3813530524284208e-06
GC_12_25 b_12 NI_12 NS_25 0 -1.7205037505887498e-03
GC_12_26 b_12 NI_12 NS_26 0 1.4659569926855143e-03
GC_12_27 b_12 NI_12 NS_27 0 8.3740845337209897e-04
GC_12_28 b_12 NI_12 NS_28 0 -1.2555801941265075e-03
GC_12_29 b_12 NI_12 NS_29 0 -1.7267001986609289e-04
GC_12_30 b_12 NI_12 NS_30 0 -2.7959000143005228e-04
GC_12_31 b_12 NI_12 NS_31 0 -1.2052302118930189e-06
GC_12_32 b_12 NI_12 NS_32 0 -1.0332950312581274e-06
GC_12_33 b_12 NI_12 NS_33 0 -7.1020870973014232e-05
GC_12_34 b_12 NI_12 NS_34 0 1.4818226572468448e-05
GC_12_35 b_12 NI_12 NS_35 0 -1.8516952569759013e-06
GC_12_36 b_12 NI_12 NS_36 0 4.7519720394391868e-07
GC_12_37 b_12 NI_12 NS_37 0 -4.6311545252998259e-07
GC_12_38 b_12 NI_12 NS_38 0 -2.0724548996706906e-07
GC_12_39 b_12 NI_12 NS_39 0 4.7433695819663435e-05
GC_12_40 b_12 NI_12 NS_40 0 -1.2704949864181996e-04
GC_12_41 b_12 NI_12 NS_41 0 3.5458474176535241e-05
GC_12_42 b_12 NI_12 NS_42 0 -3.7224988754081331e-05
GC_12_43 b_12 NI_12 NS_43 0 9.7157724398932620e-08
GC_12_44 b_12 NI_12 NS_44 0 -7.8350613330000889e-06
GC_12_45 b_12 NI_12 NS_45 0 -7.0009713482045528e-03
GC_12_46 b_12 NI_12 NS_46 0 4.8134337560576913e-05
GC_12_47 b_12 NI_12 NS_47 0 -5.2245231104417660e-04
GC_12_48 b_12 NI_12 NS_48 0 -1.7389684517109907e-03
GC_12_49 b_12 NI_12 NS_49 0 1.7859563375157332e-03
GC_12_50 b_12 NI_12 NS_50 0 -4.9223521168255803e-04
GC_12_51 b_12 NI_12 NS_51 0 1.2938659980306099e-03
GC_12_52 b_12 NI_12 NS_52 0 -9.0056138653113460e-04
GC_12_53 b_12 NI_12 NS_53 0 -2.5114284587946244e-04
GC_12_54 b_12 NI_12 NS_54 0 2.5924648839911849e-04
GC_12_55 b_12 NI_12 NS_55 0 1.7657872136314448e-03
GC_12_56 b_12 NI_12 NS_56 0 1.3062342906827061e-03
GC_12_57 b_12 NI_12 NS_57 0 -2.4702266292376240e-05
GC_12_58 b_12 NI_12 NS_58 0 -6.4663827868776462e-05
GC_12_59 b_12 NI_12 NS_59 0 2.6834901487270061e-05
GC_12_60 b_12 NI_12 NS_60 0 -2.3854992741883493e-05
GC_12_61 b_12 NI_12 NS_61 0 -8.3833893345141739e-05
GC_12_62 b_12 NI_12 NS_62 0 1.5331454558111942e-04
GC_12_63 b_12 NI_12 NS_63 0 -1.8534900343413886e-06
GC_12_64 b_12 NI_12 NS_64 0 1.0180698426838769e-05
GC_12_65 b_12 NI_12 NS_65 0 4.3862392023648088e-06
GC_12_66 b_12 NI_12 NS_66 0 3.0936550171672485e-05
GC_12_67 b_12 NI_12 NS_67 0 -6.2342257390191144e-07
GC_12_68 b_12 NI_12 NS_68 0 2.2712755019806413e-07
GC_12_69 b_12 NI_12 NS_69 0 8.0486074694677788e-04
GC_12_70 b_12 NI_12 NS_70 0 -8.8262624615847776e-05
GC_12_71 b_12 NI_12 NS_71 0 -4.4552090310245456e-04
GC_12_72 b_12 NI_12 NS_72 0 4.3729240434461198e-04
GC_12_73 b_12 NI_12 NS_73 0 1.1171733684972639e-05
GC_12_74 b_12 NI_12 NS_74 0 -2.5726433397829276e-05
GC_12_75 b_12 NI_12 NS_75 0 7.6346496526018443e-07
GC_12_76 b_12 NI_12 NS_76 0 -2.9276901751704534e-08
GC_12_77 b_12 NI_12 NS_77 0 -8.9731485204198246e-06
GC_12_78 b_12 NI_12 NS_78 0 -1.5131074960561316e-05
GC_12_79 b_12 NI_12 NS_79 0 5.3457667862534021e-07
GC_12_80 b_12 NI_12 NS_80 0 3.1692041975584903e-06
GC_12_81 b_12 NI_12 NS_81 0 -5.5403055255166780e-06
GC_12_82 b_12 NI_12 NS_82 0 -1.3507680947908716e-05
GC_12_83 b_12 NI_12 NS_83 0 -2.4375028597632410e-05
GC_12_84 b_12 NI_12 NS_84 0 8.9816869252860740e-05
GC_12_85 b_12 NI_12 NS_85 0 -9.2256127156792127e-05
GC_12_86 b_12 NI_12 NS_86 0 -1.3513340797481907e-05
GC_12_87 b_12 NI_12 NS_87 0 1.6340525871663976e-05
GC_12_88 b_12 NI_12 NS_88 0 2.5546316554647742e-05
GC_12_89 b_12 NI_12 NS_89 0 1.8353629104736328e-03
GC_12_90 b_12 NI_12 NS_90 0 -8.1496573541667562e-05
GC_12_91 b_12 NI_12 NS_91 0 -1.4246904317904096e-03
GC_12_92 b_12 NI_12 NS_92 0 2.3503729805304623e-03
GC_12_93 b_12 NI_12 NS_93 0 -2.0309473490105873e-03
GC_12_94 b_12 NI_12 NS_94 0 -2.5779773943455466e-03
GC_12_95 b_12 NI_12 NS_95 0 1.3478924619194760e-03
GC_12_96 b_12 NI_12 NS_96 0 -1.4137399015676656e-03
GC_12_97 b_12 NI_12 NS_97 0 -1.6671024045083528e-05
GC_12_98 b_12 NI_12 NS_98 0 3.0109292261372016e-04
GC_12_99 b_12 NI_12 NS_99 0 -8.3429487393417467e-04
GC_12_100 b_12 NI_12 NS_100 0 -1.6100691876800034e-04
GC_12_101 b_12 NI_12 NS_101 0 -5.0045096989798652e-05
GC_12_102 b_12 NI_12 NS_102 0 1.9961663943033600e-04
GC_12_103 b_12 NI_12 NS_103 0 2.2201615080165316e-04
GC_12_104 b_12 NI_12 NS_104 0 -3.2028405179757434e-05
GC_12_105 b_12 NI_12 NS_105 0 -2.5660035049358425e-04
GC_12_106 b_12 NI_12 NS_106 0 3.4517837272211383e-05
GC_12_107 b_12 NI_12 NS_107 0 -2.6981829216076552e-05
GC_12_108 b_12 NI_12 NS_108 0 -4.7971095406532196e-06
GC_12_109 b_12 NI_12 NS_109 0 -2.0765423613317498e-05
GC_12_110 b_12 NI_12 NS_110 0 -1.8735738993369651e-05
GC_12_111 b_12 NI_12 NS_111 0 2.9422995686391235e-06
GC_12_112 b_12 NI_12 NS_112 0 1.6729852798690198e-06
GC_12_113 b_12 NI_12 NS_113 0 2.6680134013125937e-03
GC_12_114 b_12 NI_12 NS_114 0 1.0553606427020764e-03
GC_12_115 b_12 NI_12 NS_115 0 -1.3904690700017350e-03
GC_12_116 b_12 NI_12 NS_116 0 -1.4499572984542513e-03
GC_12_117 b_12 NI_12 NS_117 0 -3.5086163313715662e-05
GC_12_118 b_12 NI_12 NS_118 0 -5.9577560389297428e-05
GC_12_119 b_12 NI_12 NS_119 0 -4.1939740353520996e-07
GC_12_120 b_12 NI_12 NS_120 0 -4.0902891029213163e-07
GC_12_121 b_12 NI_12 NS_121 0 -1.1418185354756168e-05
GC_12_122 b_12 NI_12 NS_122 0 1.0428347168328613e-05
GC_12_123 b_12 NI_12 NS_123 0 -2.6985344143699297e-07
GC_12_124 b_12 NI_12 NS_124 0 4.0623754426899130e-07
GC_12_125 b_12 NI_12 NS_125 0 -9.5997446118472446e-07
GC_12_126 b_12 NI_12 NS_126 0 -1.2878619097720091e-06
GC_12_127 b_12 NI_12 NS_127 0 -1.8954257541876173e-05
GC_12_128 b_12 NI_12 NS_128 0 -3.4595309187476067e-05
GC_12_129 b_12 NI_12 NS_129 0 1.1022922227472019e-05
GC_12_130 b_12 NI_12 NS_130 0 -9.1976516587046541e-06
GC_12_131 b_12 NI_12 NS_131 0 5.5940253281930182e-06
GC_12_132 b_12 NI_12 NS_132 0 -8.7726319169471582e-07
GC_12_133 b_12 NI_12 NS_133 0 -7.7201038696604980e-03
GC_12_134 b_12 NI_12 NS_134 0 4.6036720890333272e-05
GC_12_135 b_12 NI_12 NS_135 0 3.5600840642868568e-04
GC_12_136 b_12 NI_12 NS_136 0 -2.5848364737895420e-03
GC_12_137 b_12 NI_12 NS_137 0 1.6943161426997767e-03
GC_12_138 b_12 NI_12 NS_138 0 7.6434861517053331e-04
GC_12_139 b_12 NI_12 NS_139 0 1.4074003772113245e-03
GC_12_140 b_12 NI_12 NS_140 0 -8.6544116223084974e-04
GC_12_141 b_12 NI_12 NS_141 0 -9.6882068985036147e-05
GC_12_142 b_12 NI_12 NS_142 0 1.2011801859381414e-04
GC_12_143 b_12 NI_12 NS_143 0 1.1859183568386129e-03
GC_12_144 b_12 NI_12 NS_144 0 1.5431610557078007e-03
GC_12_145 b_12 NI_12 NS_145 0 -4.1974202777293426e-05
GC_12_146 b_12 NI_12 NS_146 0 -9.4653538199337869e-05
GC_12_147 b_12 NI_12 NS_147 0 3.5520558136251137e-05
GC_12_148 b_12 NI_12 NS_148 0 -3.7570138263593406e-05
GC_12_149 b_12 NI_12 NS_149 0 -9.8097146163083162e-05
GC_12_150 b_12 NI_12 NS_150 0 1.3440293197908136e-04
GC_12_151 b_12 NI_12 NS_151 0 -6.8715956153738578e-06
GC_12_152 b_12 NI_12 NS_152 0 7.5586943959119549e-06
GC_12_153 b_12 NI_12 NS_153 0 -4.8165201091200885e-06
GC_12_154 b_12 NI_12 NS_154 0 2.9354694888476412e-05
GC_12_155 b_12 NI_12 NS_155 0 -6.8688023788069545e-07
GC_12_156 b_12 NI_12 NS_156 0 8.7973206880526479e-07
GC_12_157 b_12 NI_12 NS_157 0 1.4015214406330411e-03
GC_12_158 b_12 NI_12 NS_158 0 -1.1639793123062457e-04
GC_12_159 b_12 NI_12 NS_159 0 -8.8610296437748785e-04
GC_12_160 b_12 NI_12 NS_160 0 2.7449358098781358e-04
GC_12_161 b_12 NI_12 NS_161 0 -5.3103544993893327e-05
GC_12_162 b_12 NI_12 NS_162 0 -2.1662731190091564e-05
GC_12_163 b_12 NI_12 NS_163 0 9.2333175601566430e-07
GC_12_164 b_12 NI_12 NS_164 0 -1.5294455979181771e-07
GC_12_165 b_12 NI_12 NS_165 0 -1.6339952787414514e-05
GC_12_166 b_12 NI_12 NS_166 0 -1.7237379829733060e-07
GC_12_167 b_12 NI_12 NS_167 0 -1.4771839487346266e-08
GC_12_168 b_12 NI_12 NS_168 0 4.6930604172609657e-06
GC_12_169 b_12 NI_12 NS_169 0 -6.8323688717628898e-06
GC_12_170 b_12 NI_12 NS_170 0 -1.3826781834093171e-05
GC_12_171 b_12 NI_12 NS_171 0 -3.6423461675101327e-05
GC_12_172 b_12 NI_12 NS_172 0 9.3394881876893512e-05
GC_12_173 b_12 NI_12 NS_173 0 -1.0377461268375386e-04
GC_12_174 b_12 NI_12 NS_174 0 -5.4861100466000061e-06
GC_12_175 b_12 NI_12 NS_175 0 1.7053330716747981e-05
GC_12_176 b_12 NI_12 NS_176 0 2.5300965507755521e-05
GC_12_177 b_12 NI_12 NS_177 0 -4.3958862252534347e-03
GC_12_178 b_12 NI_12 NS_178 0 -9.0777618995652154e-05
GC_12_179 b_12 NI_12 NS_179 0 -3.4404004717975239e-03
GC_12_180 b_12 NI_12 NS_180 0 2.0210165385456157e-03
GC_12_181 b_12 NI_12 NS_181 0 -4.9337974146362125e-04
GC_12_182 b_12 NI_12 NS_182 0 -4.0747012553577280e-03
GC_12_183 b_12 NI_12 NS_183 0 1.3970777582902731e-03
GC_12_184 b_12 NI_12 NS_184 0 -1.1760055933874582e-03
GC_12_185 b_12 NI_12 NS_185 0 1.6563892939211705e-04
GC_12_186 b_12 NI_12 NS_186 0 -1.4757526011857820e-04
GC_12_187 b_12 NI_12 NS_187 0 -9.7312484526946869e-04
GC_12_188 b_12 NI_12 NS_188 0 -2.8312976679026099e-03
GC_12_189 b_12 NI_12 NS_189 0 -1.0726088726845264e-04
GC_12_190 b_12 NI_12 NS_190 0 2.1933156711715867e-04
GC_12_191 b_12 NI_12 NS_191 0 2.0124271079451184e-04
GC_12_192 b_12 NI_12 NS_192 0 -5.4626912225855118e-05
GC_12_193 b_12 NI_12 NS_193 0 -9.9261163484090168e-05
GC_12_194 b_12 NI_12 NS_194 0 -1.6536522588634056e-04
GC_12_195 b_12 NI_12 NS_195 0 -3.2354395029773109e-05
GC_12_196 b_12 NI_12 NS_196 0 -2.5316888210257283e-05
GC_12_197 b_12 NI_12 NS_197 0 -4.7489227179072543e-05
GC_12_198 b_12 NI_12 NS_198 0 -5.6669282189429107e-05
GC_12_199 b_12 NI_12 NS_199 0 1.9670502485363753e-06
GC_12_200 b_12 NI_12 NS_200 0 4.5476291160612159e-07
GC_12_201 b_12 NI_12 NS_201 0 6.3088018014850504e-03
GC_12_202 b_12 NI_12 NS_202 0 2.8314688857716801e-03
GC_12_203 b_12 NI_12 NS_203 0 -3.0528998336198246e-03
GC_12_204 b_12 NI_12 NS_204 0 -2.4994549656521254e-03
GC_12_205 b_12 NI_12 NS_205 0 6.1556831549677848e-05
GC_12_206 b_12 NI_12 NS_206 0 2.1313256518446563e-04
GC_12_207 b_12 NI_12 NS_207 0 4.5412610207917937e-07
GC_12_208 b_12 NI_12 NS_208 0 1.0965892950260791e-06
GC_12_209 b_12 NI_12 NS_209 0 5.0102819824897967e-05
GC_12_210 b_12 NI_12 NS_210 0 4.6042427023961209e-06
GC_12_211 b_12 NI_12 NS_211 0 3.6648195719169980e-07
GC_12_212 b_12 NI_12 NS_212 0 1.9218476246586410e-07
GC_12_213 b_12 NI_12 NS_213 0 3.6178653853442268e-06
GC_12_214 b_12 NI_12 NS_214 0 5.3309154516297556e-07
GC_12_215 b_12 NI_12 NS_215 0 -1.4652616834782018e-04
GC_12_216 b_12 NI_12 NS_216 0 1.0880864250704987e-05
GC_12_217 b_12 NI_12 NS_217 0 -1.4894665965063044e-05
GC_12_218 b_12 NI_12 NS_218 0 -1.5389908727207599e-05
GC_12_219 b_12 NI_12 NS_219 0 -3.3165573412222516e-06
GC_12_220 b_12 NI_12 NS_220 0 7.0127921328621676e-06
GC_12_221 b_12 NI_12 NS_221 0 -6.5775107440076037e-03
GC_12_222 b_12 NI_12 NS_222 0 1.3709303852559364e-05
GC_12_223 b_12 NI_12 NS_223 0 2.1081904113964575e-03
GC_12_224 b_12 NI_12 NS_224 0 -2.2925817218600372e-03
GC_12_225 b_12 NI_12 NS_225 0 -4.0290652845767158e-04
GC_12_226 b_12 NI_12 NS_226 0 2.3106704686937075e-03
GC_12_227 b_12 NI_12 NS_227 0 7.1393542789899983e-04
GC_12_228 b_12 NI_12 NS_228 0 -6.6889357741732386e-04
GC_12_229 b_12 NI_12 NS_229 0 3.9387720606285167e-04
GC_12_230 b_12 NI_12 NS_230 0 -1.0217273075967349e-04
GC_12_231 b_12 NI_12 NS_231 0 -4.1847632697973613e-04
GC_12_232 b_12 NI_12 NS_232 0 3.8358518306321523e-04
GC_12_233 b_12 NI_12 NS_233 0 -5.4446268966707020e-05
GC_12_234 b_12 NI_12 NS_234 0 -9.6901709719856451e-05
GC_12_235 b_12 NI_12 NS_235 0 2.8557372980666634e-05
GC_12_236 b_12 NI_12 NS_236 0 -4.0820152391300763e-05
GC_12_237 b_12 NI_12 NS_237 0 -1.0444586353162010e-04
GC_12_238 b_12 NI_12 NS_238 0 1.0947178771891059e-04
GC_12_239 b_12 NI_12 NS_239 0 -9.1462794701559001e-06
GC_12_240 b_12 NI_12 NS_240 0 9.6433512051397119e-06
GC_12_241 b_12 NI_12 NS_241 0 -1.0532786818947664e-05
GC_12_242 b_12 NI_12 NS_242 0 4.0942520585208664e-05
GC_12_243 b_12 NI_12 NS_243 0 -1.4333373087430212e-06
GC_12_244 b_12 NI_12 NS_244 0 2.7864853719509981e-07
GC_12_245 b_12 NI_12 NS_245 0 2.8146570081552837e-03
GC_12_246 b_12 NI_12 NS_246 0 -2.0759944606431303e-03
GC_12_247 b_12 NI_12 NS_247 0 -1.7758096632356415e-03
GC_12_248 b_12 NI_12 NS_248 0 1.1015225488881020e-03
GC_12_249 b_12 NI_12 NS_249 0 2.9428568477447997e-05
GC_12_250 b_12 NI_12 NS_250 0 -3.7008624955830266e-05
GC_12_251 b_12 NI_12 NS_251 0 1.6465548220696211e-06
GC_12_252 b_12 NI_12 NS_252 0 -3.3987603491935147e-07
GC_12_253 b_12 NI_12 NS_253 0 -2.3709565226970290e-05
GC_12_254 b_12 NI_12 NS_254 0 -1.3494367349654432e-05
GC_12_255 b_12 NI_12 NS_255 0 7.5996048406688611e-07
GC_12_256 b_12 NI_12 NS_256 0 5.2410059679901151e-06
GC_12_257 b_12 NI_12 NS_257 0 -9.1527659293341115e-06
GC_12_258 b_12 NI_12 NS_258 0 -2.1591622628734808e-05
GC_12_259 b_12 NI_12 NS_259 0 -4.6005615822922798e-05
GC_12_260 b_12 NI_12 NS_260 0 1.8503668660778047e-04
GC_12_261 b_12 NI_12 NS_261 0 -1.5662841441585040e-04
GC_12_262 b_12 NI_12 NS_262 0 -6.5461622154234258e-06
GC_12_263 b_12 NI_12 NS_263 0 2.6304267973392639e-05
GC_12_264 b_12 NI_12 NS_264 0 3.8665299374374876e-05
GC_12_265 b_12 NI_12 NS_265 0 -9.2404038202671148e-04
GC_12_266 b_12 NI_12 NS_266 0 -1.0486435411949298e-04
GC_12_267 b_12 NI_12 NS_267 0 -5.6890150266194076e-03
GC_12_268 b_12 NI_12 NS_268 0 -9.2937909862553854e-04
GC_12_269 b_12 NI_12 NS_269 0 2.1856550581704276e-03
GC_12_270 b_12 NI_12 NS_270 0 -4.4645526662996909e-04
GC_12_271 b_12 NI_12 NS_271 0 6.7367416259189207e-04
GC_12_272 b_12 NI_12 NS_272 0 -4.8131725161539420e-04
GC_12_273 b_12 NI_12 NS_273 0 8.9750050242013433e-04
GC_12_274 b_12 NI_12 NS_274 0 2.8166329621153992e-04
GC_12_275 b_12 NI_12 NS_275 0 6.2080685063564060e-04
GC_12_276 b_12 NI_12 NS_276 0 -4.4931037199550565e-03
GC_12_277 b_12 NI_12 NS_277 0 -1.3699452358763772e-04
GC_12_278 b_12 NI_12 NS_278 0 1.5172652148983198e-04
GC_12_279 b_12 NI_12 NS_279 0 1.5212355527487899e-04
GC_12_280 b_12 NI_12 NS_280 0 -2.6260463575127544e-05
GC_12_281 b_12 NI_12 NS_281 0 -8.1269803623911974e-05
GC_12_282 b_12 NI_12 NS_282 0 -4.0289757990259535e-05
GC_12_283 b_12 NI_12 NS_283 0 -1.9383966378463150e-05
GC_12_284 b_12 NI_12 NS_284 0 -1.0425340580981577e-05
GC_12_285 b_12 NI_12 NS_285 0 -1.8592434584921741e-05
GC_12_286 b_12 NI_12 NS_286 0 -2.7443285999611395e-05
GC_12_287 b_12 NI_12 NS_287 0 1.9958229820974763e-06
GC_12_288 b_12 NI_12 NS_288 0 5.3636260682804199e-07
GC_12_289 b_12 NI_12 NS_289 0 1.6574361944189397e-03
GC_12_290 b_12 NI_12 NS_290 0 3.0647333810407650e-03
GC_12_291 b_12 NI_12 NS_291 0 -7.7998852791277178e-04
GC_12_292 b_12 NI_12 NS_292 0 -1.7043265536223992e-03
GC_12_293 b_12 NI_12 NS_293 0 4.4861243953937031e-05
GC_12_294 b_12 NI_12 NS_294 0 1.9006420059222506e-04
GC_12_295 b_12 NI_12 NS_295 0 3.0979022679603436e-07
GC_12_296 b_12 NI_12 NS_296 0 4.1163530682228621e-07
GC_12_297 b_12 NI_12 NS_297 0 3.9532654428907028e-05
GC_12_298 b_12 NI_12 NS_298 0 1.3984380738417220e-06
GC_12_299 b_12 NI_12 NS_299 0 6.6950162699954343e-07
GC_12_300 b_12 NI_12 NS_300 0 2.0641674768929016e-07
GC_12_301 b_12 NI_12 NS_301 0 -4.6822464253343895e-07
GC_12_302 b_12 NI_12 NS_302 0 -8.9954844251060289e-07
GC_12_303 b_12 NI_12 NS_303 0 -7.3574673989755564e-05
GC_12_304 b_12 NI_12 NS_304 0 -2.1184629916244795e-05
GC_12_305 b_12 NI_12 NS_305 0 -1.2509487085742442e-05
GC_12_306 b_12 NI_12 NS_306 0 -7.5098806214445523e-06
GC_12_307 b_12 NI_12 NS_307 0 2.2524736632212695e-06
GC_12_308 b_12 NI_12 NS_308 0 2.4634424021573379e-06
GC_12_309 b_12 NI_12 NS_309 0 -1.5486858777937565e-03
GC_12_310 b_12 NI_12 NS_310 0 -3.5231288951180587e-04
GC_12_311 b_12 NI_12 NS_311 0 3.8115909101869537e-03
GC_12_312 b_12 NI_12 NS_312 0 1.9431288310767418e-03
GC_12_313 b_12 NI_12 NS_313 0 -5.7326668809368538e-03
GC_12_314 b_12 NI_12 NS_314 0 -1.5733240587980579e-03
GC_12_315 b_12 NI_12 NS_315 0 7.8471878613745299e-04
GC_12_316 b_12 NI_12 NS_316 0 -6.0615700562092231e-04
GC_12_317 b_12 NI_12 NS_317 0 2.2348756940792445e-04
GC_12_318 b_12 NI_12 NS_318 0 3.4945715564520642e-04
GC_12_319 b_12 NI_12 NS_319 0 5.4670033154548823e-04
GC_12_320 b_12 NI_12 NS_320 0 -1.9578561260614321e-03
GC_12_321 b_12 NI_12 NS_321 0 -4.4516932215545953e-05
GC_12_322 b_12 NI_12 NS_322 0 -6.0017652261405035e-05
GC_12_323 b_12 NI_12 NS_323 0 1.7366513284289762e-05
GC_12_324 b_12 NI_12 NS_324 0 -2.9323561135615045e-05
GC_12_325 b_12 NI_12 NS_325 0 -7.4360235474998983e-05
GC_12_326 b_12 NI_12 NS_326 0 6.2773929283612562e-05
GC_12_327 b_12 NI_12 NS_327 0 -6.1280135848502709e-06
GC_12_328 b_12 NI_12 NS_328 0 1.2388185532706647e-06
GC_12_329 b_12 NI_12 NS_329 0 -1.0717438370762434e-05
GC_12_330 b_12 NI_12 NS_330 0 1.3690102806507972e-05
GC_12_331 b_12 NI_12 NS_331 0 -1.3302421358636971e-06
GC_12_332 b_12 NI_12 NS_332 0 5.1766192262235097e-07
GC_12_333 b_12 NI_12 NS_333 0 3.0793950464298413e-03
GC_12_334 b_12 NI_12 NS_334 0 3.5657386593705720e-04
GC_12_335 b_12 NI_12 NS_335 0 -1.5595379996998161e-03
GC_12_336 b_12 NI_12 NS_336 0 -2.5251759548987264e-04
GC_12_337 b_12 NI_12 NS_337 0 -4.1907051709658847e-06
GC_12_338 b_12 NI_12 NS_338 0 7.2307595488740509e-05
GC_12_339 b_12 NI_12 NS_339 0 9.3764965681299880e-07
GC_12_340 b_12 NI_12 NS_340 0 1.7017258573233140e-07
GC_12_341 b_12 NI_12 NS_341 0 4.8632805863255861e-06
GC_12_342 b_12 NI_12 NS_342 0 1.3104812675988972e-05
GC_12_343 b_12 NI_12 NS_343 0 -1.3426139828944773e-07
GC_12_344 b_12 NI_12 NS_344 0 3.4906142092922377e-06
GC_12_345 b_12 NI_12 NS_345 0 -4.4742496331478693e-06
GC_12_346 b_12 NI_12 NS_346 0 -1.2432072389930661e-05
GC_12_347 b_12 NI_12 NS_347 0 -7.4957430356594241e-05
GC_12_348 b_12 NI_12 NS_348 0 1.0707737033855116e-04
GC_12_349 b_12 NI_12 NS_349 0 -9.3114093978399786e-05
GC_12_350 b_12 NI_12 NS_350 0 -2.1115771811984979e-06
GC_12_351 b_12 NI_12 NS_351 0 9.5946968373378443e-06
GC_12_352 b_12 NI_12 NS_352 0 2.0479795271435058e-05
GC_12_353 b_12 NI_12 NS_353 0 7.2221788558421750e-03
GC_12_354 b_12 NI_12 NS_354 0 -3.6221201072865385e-04
GC_12_355 b_12 NI_12 NS_355 0 -1.9882112977590963e-02
GC_12_356 b_12 NI_12 NS_356 0 -2.9310672005069659e-03
GC_12_357 b_12 NI_12 NS_357 0 9.7598244588673194e-03
GC_12_358 b_12 NI_12 NS_358 0 -2.7969796518778340e-03
GC_12_359 b_12 NI_12 NS_359 0 5.7013058624983490e-03
GC_12_360 b_12 NI_12 NS_360 0 6.7618349981718527e-04
GC_12_361 b_12 NI_12 NS_361 0 1.5968830043374706e-03
GC_12_362 b_12 NI_12 NS_362 0 -8.6069402703275078e-04
GC_12_363 b_12 NI_12 NS_363 0 -5.2205901742202866e-05
GC_12_364 b_12 NI_12 NS_364 0 -8.6046019500995562e-03
GC_12_365 b_12 NI_12 NS_365 0 -2.7012461749727619e-04
GC_12_366 b_12 NI_12 NS_366 0 9.0542398599864068e-05
GC_12_367 b_12 NI_12 NS_367 0 2.3050374309891501e-04
GC_12_368 b_12 NI_12 NS_368 0 3.4908456389659773e-05
GC_12_369 b_12 NI_12 NS_369 0 5.3532353537666388e-04
GC_12_370 b_12 NI_12 NS_370 0 4.8342451317561028e-04
GC_12_371 b_12 NI_12 NS_371 0 3.3166282548230622e-05
GC_12_372 b_12 NI_12 NS_372 0 2.3104994189684430e-05
GC_12_373 b_12 NI_12 NS_373 0 7.4281860200873642e-05
GC_12_374 b_12 NI_12 NS_374 0 -2.1860255518790250e-05
GC_12_375 b_12 NI_12 NS_375 0 6.7174860060768698e-06
GC_12_376 b_12 NI_12 NS_376 0 -3.0035187185974060e-06
GC_12_377 b_12 NI_12 NS_377 0 -7.1010896762923881e-03
GC_12_378 b_12 NI_12 NS_378 0 1.1143993545295798e-02
GC_12_379 b_12 NI_12 NS_379 0 5.0151273330545695e-03
GC_12_380 b_12 NI_12 NS_380 0 -4.9722785823262039e-03
GC_12_381 b_12 NI_12 NS_381 0 -3.9017729368529035e-04
GC_12_382 b_12 NI_12 NS_382 0 6.3164745028453487e-06
GC_12_383 b_12 NI_12 NS_383 0 -2.4927630367487045e-06
GC_12_384 b_12 NI_12 NS_384 0 -2.8432544330701852e-07
GC_12_385 b_12 NI_12 NS_385 0 -5.3738301810940158e-05
GC_12_386 b_12 NI_12 NS_386 0 9.0888003669049427e-05
GC_12_387 b_12 NI_12 NS_387 0 -1.1803819706411931e-06
GC_12_388 b_12 NI_12 NS_388 0 1.8404645000118301e-06
GC_12_389 b_12 NI_12 NS_389 0 -2.6448935700382531e-07
GC_12_390 b_12 NI_12 NS_390 0 2.1268368263350893e-06
GC_12_391 b_12 NI_12 NS_391 0 -1.1065874190364190e-04
GC_12_392 b_12 NI_12 NS_392 0 -2.7199021486770886e-04
GC_12_393 b_12 NI_12 NS_393 0 -3.7657372662876076e-06
GC_12_394 b_12 NI_12 NS_394 0 -6.0107678714557062e-05
GC_12_395 b_12 NI_12 NS_395 0 -7.8808636189676150e-06
GC_12_396 b_12 NI_12 NS_396 0 -1.2254870634149081e-05
GC_12_397 b_12 NI_12 NS_397 0 -9.7443421373210569e-03
GC_12_398 b_12 NI_12 NS_398 0 -9.3917171272320894e-04
GC_12_399 b_12 NI_12 NS_399 0 1.3653746597708186e-02
GC_12_400 b_12 NI_12 NS_400 0 2.7673291230059451e-03
GC_12_401 b_12 NI_12 NS_401 0 -1.5647676844076131e-02
GC_12_402 b_12 NI_12 NS_402 0 -3.6596642560925902e-03
GC_12_403 b_12 NI_12 NS_403 0 5.5280297490399675e-03
GC_12_404 b_12 NI_12 NS_404 0 -1.3324129345126080e-03
GC_12_405 b_12 NI_12 NS_405 0 -8.2810141254369238e-04
GC_12_406 b_12 NI_12 NS_406 0 6.6508459781560402e-04
GC_12_407 b_12 NI_12 NS_407 0 1.9880254564857039e-03
GC_12_408 b_12 NI_12 NS_408 0 -3.4878358547294906e-03
GC_12_409 b_12 NI_12 NS_409 0 8.6027085081775008e-05
GC_12_410 b_12 NI_12 NS_410 0 -1.3374342761638249e-04
GC_12_411 b_12 NI_12 NS_411 0 1.2614452964307569e-05
GC_12_412 b_12 NI_12 NS_412 0 -4.1222658370920199e-05
GC_12_413 b_12 NI_12 NS_413 0 9.4340971347328805e-05
GC_12_414 b_12 NI_12 NS_414 0 -8.2947552189313795e-05
GC_12_415 b_12 NI_12 NS_415 0 5.4963698761852063e-06
GC_12_416 b_12 NI_12 NS_416 0 -1.0735251088336974e-05
GC_12_417 b_12 NI_12 NS_417 0 -1.2131682052728064e-05
GC_12_418 b_12 NI_12 NS_418 0 -1.9429380574419946e-05
GC_12_419 b_12 NI_12 NS_419 0 -4.0447317534836989e-06
GC_12_420 b_12 NI_12 NS_420 0 -1.2811397566797350e-06
GC_12_421 b_12 NI_12 NS_421 0 7.3694096641483426e-03
GC_12_422 b_12 NI_12 NS_422 0 7.3632398657584967e-03
GC_12_423 b_12 NI_12 NS_423 0 -2.8316970022066873e-03
GC_12_424 b_12 NI_12 NS_424 0 -3.5561294446567080e-03
GC_12_425 b_12 NI_12 NS_425 0 -2.7050625177076548e-04
GC_12_426 b_12 NI_12 NS_426 0 6.5144461968380716e-05
GC_12_427 b_12 NI_12 NS_427 0 -3.6858897198612891e-07
GC_12_428 b_12 NI_12 NS_428 0 1.5925358445212889e-06
GC_12_429 b_12 NI_12 NS_429 0 -1.6844486626067160e-05
GC_12_430 b_12 NI_12 NS_430 0 1.3271591819048989e-04
GC_12_431 b_12 NI_12 NS_431 0 -3.0175705031636476e-06
GC_12_432 b_12 NI_12 NS_432 0 -4.7729998784314308e-07
GC_12_433 b_12 NI_12 NS_433 0 -7.0797261048928464e-06
GC_12_434 b_12 NI_12 NS_434 0 -1.8681115657960917e-05
GC_12_435 b_12 NI_12 NS_435 0 -3.2514654921884559e-04
GC_12_436 b_12 NI_12 NS_436 0 1.6915798568120608e-04
GC_12_437 b_12 NI_12 NS_437 0 -1.8429815109945093e-04
GC_12_438 b_12 NI_12 NS_438 0 -3.7599256690362281e-05
GC_12_439 b_12 NI_12 NS_439 0 -2.3736717877285243e-05
GC_12_440 b_12 NI_12 NS_440 0 9.6044429450360846e-06
GC_12_441 b_12 NI_12 NS_441 0 3.5289009065899962e-02
GC_12_442 b_12 NI_12 NS_442 0 1.6497220761540046e-02
GC_12_443 b_12 NI_12 NS_443 0 -1.9435780531245280e-02
GC_12_444 b_12 NI_12 NS_444 0 -5.4527637852197766e-03
GC_12_445 b_12 NI_12 NS_445 0 -2.8214541330285624e-02
GC_12_446 b_12 NI_12 NS_446 0 1.8345572205390429e-03
GC_12_447 b_12 NI_12 NS_447 0 2.2404843324733484e-03
GC_12_448 b_12 NI_12 NS_448 0 2.0288883483987512e-03
GC_12_449 b_12 NI_12 NS_449 0 -2.0527313855237929e-03
GC_12_450 b_12 NI_12 NS_450 0 2.8472531335623934e-04
GC_12_451 b_12 NI_12 NS_451 0 7.7524789725735730e-03
GC_12_452 b_12 NI_12 NS_452 0 -3.1287535393384096e-03
GC_12_453 b_12 NI_12 NS_453 0 -3.2243079627031646e-04
GC_12_454 b_12 NI_12 NS_454 0 3.0820890158335456e-05
GC_12_455 b_12 NI_12 NS_455 0 8.3139366925115269e-05
GC_12_456 b_12 NI_12 NS_456 0 4.0063819737582978e-06
GC_12_457 b_12 NI_12 NS_457 0 2.1977055600805589e-04
GC_12_458 b_12 NI_12 NS_458 0 -3.1180510498785192e-04
GC_12_459 b_12 NI_12 NS_459 0 -2.4613569795847345e-05
GC_12_460 b_12 NI_12 NS_460 0 2.3386335034770312e-06
GC_12_461 b_12 NI_12 NS_461 0 -3.9831538056633162e-05
GC_12_462 b_12 NI_12 NS_462 0 1.2518458529547847e-05
GC_12_463 b_12 NI_12 NS_463 0 2.0022389966336227e-06
GC_12_464 b_12 NI_12 NS_464 0 1.7019165922474598e-06
GC_12_465 b_12 NI_12 NS_465 0 -2.9014008520140962e-03
GC_12_466 b_12 NI_12 NS_466 0 -5.7720493218877270e-03
GC_12_467 b_12 NI_12 NS_467 0 8.0019278082879195e-04
GC_12_468 b_12 NI_12 NS_468 0 1.9977889641075845e-03
GC_12_469 b_12 NI_12 NS_469 0 9.8428082168691434e-05
GC_12_470 b_12 NI_12 NS_470 0 -8.8303314472101569e-05
GC_12_471 b_12 NI_12 NS_471 0 9.9704799204547293e-07
GC_12_472 b_12 NI_12 NS_472 0 -7.6665139017212616e-07
GC_12_473 b_12 NI_12 NS_473 0 -2.7720280552560301e-05
GC_12_474 b_12 NI_12 NS_474 0 -3.9678392029173069e-05
GC_12_475 b_12 NI_12 NS_475 0 -9.1732628212465184e-07
GC_12_476 b_12 NI_12 NS_476 0 -9.2002787784670153e-07
GC_12_477 b_12 NI_12 NS_477 0 -5.5606228844583913e-07
GC_12_478 b_12 NI_12 NS_478 0 -3.3394989048878322e-06
GC_12_479 b_12 NI_12 NS_479 0 1.0094568902167450e-04
GC_12_480 b_12 NI_12 NS_480 0 3.5941077296479005e-05
GC_12_481 b_12 NI_12 NS_481 0 2.2153910114354942e-05
GC_12_482 b_12 NI_12 NS_482 0 1.9573523786166113e-05
GC_12_483 b_12 NI_12 NS_483 0 8.1250895541778239e-06
GC_12_484 b_12 NI_12 NS_484 0 -3.1397916807856373e-06
GC_12_485 b_12 NI_12 NS_485 0 -1.3845734641945270e-01
GC_12_486 b_12 NI_12 NS_486 0 1.7548250917139796e-02
GC_12_487 b_12 NI_12 NS_487 0 9.3407566923340065e-03
GC_12_488 b_12 NI_12 NS_488 0 1.3048683820301886e-02
GC_12_489 b_12 NI_12 NS_489 0 1.5988454008662039e-02
GC_12_490 b_12 NI_12 NS_490 0 -1.2931487808525075e-02
GC_12_491 b_12 NI_12 NS_491 0 1.1501307881716623e-03
GC_12_492 b_12 NI_12 NS_492 0 1.6247565364872331e-03
GC_12_493 b_12 NI_12 NS_493 0 -8.0376960535555255e-04
GC_12_494 b_12 NI_12 NS_494 0 1.2910247479092632e-03
GC_12_495 b_12 NI_12 NS_495 0 6.4570434991127702e-03
GC_12_496 b_12 NI_12 NS_496 0 1.9323830748382387e-03
GC_12_497 b_12 NI_12 NS_497 0 -3.2558272433831037e-05
GC_12_498 b_12 NI_12 NS_498 0 -2.0063622956910537e-04
GC_12_499 b_12 NI_12 NS_499 0 3.4487507787755993e-05
GC_12_500 b_12 NI_12 NS_500 0 -8.1759378143015044e-05
GC_12_501 b_12 NI_12 NS_501 0 2.1668245508964603e-04
GC_12_502 b_12 NI_12 NS_502 0 7.6913010063805001e-05
GC_12_503 b_12 NI_12 NS_503 0 3.5181837435084522e-05
GC_12_504 b_12 NI_12 NS_504 0 2.8046296992483823e-06
GC_12_505 b_12 NI_12 NS_505 0 6.8979324111994314e-05
GC_12_506 b_12 NI_12 NS_506 0 1.9958982717123630e-07
GC_12_507 b_12 NI_12 NS_507 0 2.5707845651800845e-06
GC_12_508 b_12 NI_12 NS_508 0 -1.4392022051117192e-06
GC_12_509 b_12 NI_12 NS_509 0 -4.6686783269338965e-03
GC_12_510 b_12 NI_12 NS_510 0 3.8234739101952390e-03
GC_12_511 b_12 NI_12 NS_511 0 2.5926612735620151e-03
GC_12_512 b_12 NI_12 NS_512 0 -1.5289231306136136e-03
GC_12_513 b_12 NI_12 NS_513 0 -4.9540037218678562e-05
GC_12_514 b_12 NI_12 NS_514 0 -3.1679741721227499e-04
GC_12_515 b_12 NI_12 NS_515 0 6.2997191104655607e-07
GC_12_516 b_12 NI_12 NS_516 0 -2.8322669263652216e-06
GC_12_517 b_12 NI_12 NS_517 0 -1.1730679031245074e-04
GC_12_518 b_12 NI_12 NS_518 0 6.8156772743286905e-06
GC_12_519 b_12 NI_12 NS_519 0 -5.7295039492497754e-06
GC_12_520 b_12 NI_12 NS_520 0 4.1832167982717955e-08
GC_12_521 b_12 NI_12 NS_521 0 -9.0285532576718322e-06
GC_12_522 b_12 NI_12 NS_522 0 -1.2382432485693148e-05
GC_12_523 b_12 NI_12 NS_523 0 3.7499556209396115e-05
GC_12_524 b_12 NI_12 NS_524 0 -1.3872036777854620e-04
GC_12_525 b_12 NI_12 NS_525 0 -2.1192399864862596e-05
GC_12_526 b_12 NI_12 NS_526 0 -5.6225567493029068e-05
GC_12_527 b_12 NI_12 NS_527 0 -3.2954566600689946e-06
GC_12_528 b_12 NI_12 NS_528 0 -1.2093632574035077e-05
GD_12_1 b_12 NI_12 NA_1 0 -3.1612752692538998e-03
GD_12_2 b_12 NI_12 NA_2 0 2.9574426789372166e-03
GD_12_3 b_12 NI_12 NA_3 0 2.3832794159780167e-04
GD_12_4 b_12 NI_12 NA_4 0 3.1074003222929555e-03
GD_12_5 b_12 NI_12 NA_5 0 5.6822052398010177e-03
GD_12_6 b_12 NI_12 NA_6 0 3.7310735701693663e-03
GD_12_7 b_12 NI_12 NA_7 0 1.4691786521537848e-03
GD_12_8 b_12 NI_12 NA_8 0 6.1594338326881131e-04
GD_12_9 b_12 NI_12 NA_9 0 -2.6100856012972397e-03
GD_12_10 b_12 NI_12 NA_10 0 -2.6919946647102362e-05
GD_12_11 b_12 NI_12 NA_11 0 -9.1444686992853234e-03
GD_12_12 b_12 NI_12 NA_12 0 1.3327932617766750e-01
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 3.9451851533158515e+00
GS_1_1 0 NS_1 NA_1 0 1.1283794739964070e+00
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 1.8805154767607480e+01
GS_2_1 0 NS_2 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 3/4
CS_3 NS_3 0 9.9999999999999998e-13
CS_4 NS_4 0 9.9999999999999998e-13
RS_3 NS_3 0 1.8483596483142442e+01
RS_4 NS_4 0 1.8483596483142442e+01
GL_3 0 NS_3 NS_4 0 6.9799982353381460e-02
GL_4 0 NS_4 NS_3 0 -6.9799982353381460e-02
GS_3_1 0 NS_3 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 1.9654872352993628e+01
RS_6 NS_6 0 1.9654872352993625e+01
GL_5 0 NS_5 NS_6 0 9.5720932954598423e-02
GL_6 0 NS_6 NS_5 0 -9.5720932954598423e-02
GS_5_1 0 NS_5 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 2.5061544329287912e+01
RS_8 NS_8 0 2.5061544329287909e+01
GL_7 0 NS_7 NS_8 0 1.3536754976539320e-01
GL_8 0 NS_8 NS_7 0 -1.3536754976539320e-01
GS_7_1 0 NS_7 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 7.4239654864745361e+01
RS_10 NS_10 0 7.4239654864745361e+01
GL_9 0 NS_9 NS_10 0 2.8245804011501385e-01
GL_10 0 NS_10 NS_9 0 -2.8245804011501385e-01
GS_9_1 0 NS_9 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 2.8726427419385509e+01
RS_12 NS_12 0 2.8726427419385512e+01
GL_11 0 NS_11 NS_12 0 1.7620265460857126e-01
GL_12 0 NS_12 NS_11 0 -1.7620265460857126e-01
GS_11_1 0 NS_11 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 7.8929016552352451e+01
RS_14 NS_14 0 7.8929016552352465e+01
GL_13 0 NS_13 NS_14 0 1.7267598155977268e-01
GL_14 0 NS_14 NS_13 0 -1.7267598155977268e-01
GS_13_1 0 NS_13 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 1.3876610711235463e+02
RS_16 NS_16 0 1.3876610711235463e+02
GL_15 0 NS_15 NS_16 0 1.9827389109149790e-01
GL_16 0 NS_16 NS_15 0 -1.9827389109149790e-01
GS_15_1 0 NS_15 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 9.4943847388790630e+01
RS_18 NS_18 0 9.4943847388790630e+01
GL_17 0 NS_17 NS_18 0 2.0370912057963636e-01
GL_18 0 NS_18 NS_17 0 -2.0370912057963636e-01
GS_17_1 0 NS_17 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 2.2502148823483816e+02
RS_20 NS_20 0 2.2502148823483816e+02
GL_19 0 NS_19 NS_20 0 2.1140622110318164e-01
GL_20 0 NS_20 NS_19 0 -2.1140622110318164e-01
GS_19_1 0 NS_19 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 2.0359721972446440e+02
RS_22 NS_22 0 2.0359721972446440e+02
GL_21 0 NS_21 NS_22 0 2.1650882528339854e-01
GL_22 0 NS_22 NS_21 0 -2.1650882528339854e-01
GS_21_1 0 NS_21 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 5.4323743269805618e+02
RS_24 NS_24 0 5.4323743269805618e+02
GL_23 0 NS_23 NS_24 0 2.2057741537827197e-01
GL_24 0 NS_24 NS_23 0 -2.2057741537827197e-01
GS_23_1 0 NS_23 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 6.2013592102356057e+01
RS_26 NS_26 0 6.2013592102356057e+01
GL_25 0 NS_25 NS_26 0 2.2721975400227054e-01
GL_26 0 NS_26 NS_25 0 -2.2721975400227054e-01
GS_25_1 0 NS_25 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 8.2527539890421451e+01
RS_28 NS_28 0 8.2527539890421465e+01
GL_27 0 NS_27 NS_28 0 2.2544686857562196e-01
GL_28 0 NS_28 NS_27 0 -2.2544686857562196e-01
GS_27_1 0 NS_27 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 1.5057204740157513e+02
RS_30 NS_30 0 1.5057204740157516e+02
GL_29 0 NS_29 NS_30 0 2.5030962700427895e-01
GL_30 0 NS_30 NS_29 0 -2.5030962700427895e-01
GS_29_1 0 NS_29 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 1.0143406310664166e+03
RS_32 NS_32 0 1.0143406310664167e+03
GL_31 0 NS_31 NS_32 0 2.4802996115452441e-01
GL_32 0 NS_32 NS_31 0 -2.4802996115452441e-01
GS_31_1 0 NS_31 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 2.6049933264405115e+02
RS_34 NS_34 0 2.6049933264405115e+02
GL_33 0 NS_33 NS_34 0 2.4648481498152200e-01
GL_34 0 NS_34 NS_33 0 -2.4648481498152200e-01
GS_33_1 0 NS_33 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 8.6892684135916670e+02
RS_36 NS_36 0 8.6892684135916659e+02
GL_35 0 NS_35 NS_36 0 2.4352824357909131e-01
GL_36 0 NS_36 NS_35 0 -2.4352824357909131e-01
GS_35_1 0 NS_35 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 6.5240189890508168e+02
RS_38 NS_38 0 6.5240189890508168e+02
GL_37 0 NS_37 NS_38 0 2.3166276016037468e-01
GL_38 0 NS_38 NS_37 0 -2.3166276016037468e-01
GS_37_1 0 NS_37 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 1.8572469959933156e+02
RS_40 NS_40 0 1.8572469959933156e+02
GL_39 0 NS_39 NS_40 0 2.3351354491929543e-01
GL_40 0 NS_40 NS_39 0 -2.3351354491929543e-01
GS_39_1 0 NS_39 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 3.0631652744794525e+02
RS_42 NS_42 0 3.0631652744794530e+02
GL_41 0 NS_41 NS_42 0 2.3886925224886552e-01
GL_42 0 NS_42 NS_41 0 -2.3886925224886552e-01
GS_41_1 0 NS_41 NA_1 0 1.1283794739964070e+00
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 5.0301469986378567e+02
RS_44 NS_44 0 5.0301469986378567e+02
GL_43 0 NS_43 NS_44 0 2.3692781195536661e-01
GL_44 0 NS_44 NS_43 0 -2.3692781195536661e-01
GS_43_1 0 NS_43 NA_1 0 1.1283794739964070e+00
*
* Real pole n. 45
CS_45 NS_45 0 9.9999999999999998e-13
RS_45 NS_45 0 3.9451851533158515e+00
GS_45_2 0 NS_45 NA_2 0 1.1283794739964070e+00
*
* Real pole n. 46
CS_46 NS_46 0 9.9999999999999998e-13
RS_46 NS_46 0 1.8805154767607480e+01
GS_46_2 0 NS_46 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 1.8483596483142442e+01
RS_48 NS_48 0 1.8483596483142442e+01
GL_47 0 NS_47 NS_48 0 6.9799982353381460e-02
GL_48 0 NS_48 NS_47 0 -6.9799982353381460e-02
GS_47_2 0 NS_47 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 1.9654872352993628e+01
RS_50 NS_50 0 1.9654872352993625e+01
GL_49 0 NS_49 NS_50 0 9.5720932954598423e-02
GL_50 0 NS_50 NS_49 0 -9.5720932954598423e-02
GS_49_2 0 NS_49 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 2.5061544329287912e+01
RS_52 NS_52 0 2.5061544329287909e+01
GL_51 0 NS_51 NS_52 0 1.3536754976539320e-01
GL_52 0 NS_52 NS_51 0 -1.3536754976539320e-01
GS_51_2 0 NS_51 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 7.4239654864745361e+01
RS_54 NS_54 0 7.4239654864745361e+01
GL_53 0 NS_53 NS_54 0 2.8245804011501385e-01
GL_54 0 NS_54 NS_53 0 -2.8245804011501385e-01
GS_53_2 0 NS_53 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 2.8726427419385509e+01
RS_56 NS_56 0 2.8726427419385512e+01
GL_55 0 NS_55 NS_56 0 1.7620265460857126e-01
GL_56 0 NS_56 NS_55 0 -1.7620265460857126e-01
GS_55_2 0 NS_55 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 7.8929016552352451e+01
RS_58 NS_58 0 7.8929016552352465e+01
GL_57 0 NS_57 NS_58 0 1.7267598155977268e-01
GL_58 0 NS_58 NS_57 0 -1.7267598155977268e-01
GS_57_2 0 NS_57 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 1.3876610711235463e+02
RS_60 NS_60 0 1.3876610711235463e+02
GL_59 0 NS_59 NS_60 0 1.9827389109149790e-01
GL_60 0 NS_60 NS_59 0 -1.9827389109149790e-01
GS_59_2 0 NS_59 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 9.4943847388790630e+01
RS_62 NS_62 0 9.4943847388790630e+01
GL_61 0 NS_61 NS_62 0 2.0370912057963636e-01
GL_62 0 NS_62 NS_61 0 -2.0370912057963636e-01
GS_61_2 0 NS_61 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 2.2502148823483816e+02
RS_64 NS_64 0 2.2502148823483816e+02
GL_63 0 NS_63 NS_64 0 2.1140622110318164e-01
GL_64 0 NS_64 NS_63 0 -2.1140622110318164e-01
GS_63_2 0 NS_63 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 2.0359721972446440e+02
RS_66 NS_66 0 2.0359721972446440e+02
GL_65 0 NS_65 NS_66 0 2.1650882528339854e-01
GL_66 0 NS_66 NS_65 0 -2.1650882528339854e-01
GS_65_2 0 NS_65 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 5.4323743269805618e+02
RS_68 NS_68 0 5.4323743269805618e+02
GL_67 0 NS_67 NS_68 0 2.2057741537827197e-01
GL_68 0 NS_68 NS_67 0 -2.2057741537827197e-01
GS_67_2 0 NS_67 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 6.2013592102356057e+01
RS_70 NS_70 0 6.2013592102356057e+01
GL_69 0 NS_69 NS_70 0 2.2721975400227054e-01
GL_70 0 NS_70 NS_69 0 -2.2721975400227054e-01
GS_69_2 0 NS_69 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 8.2527539890421451e+01
RS_72 NS_72 0 8.2527539890421465e+01
GL_71 0 NS_71 NS_72 0 2.2544686857562196e-01
GL_72 0 NS_72 NS_71 0 -2.2544686857562196e-01
GS_71_2 0 NS_71 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 1.5057204740157513e+02
RS_74 NS_74 0 1.5057204740157516e+02
GL_73 0 NS_73 NS_74 0 2.5030962700427895e-01
GL_74 0 NS_74 NS_73 0 -2.5030962700427895e-01
GS_73_2 0 NS_73 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 1.0143406310664166e+03
RS_76 NS_76 0 1.0143406310664167e+03
GL_75 0 NS_75 NS_76 0 2.4802996115452441e-01
GL_76 0 NS_76 NS_75 0 -2.4802996115452441e-01
GS_75_2 0 NS_75 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 2.6049933264405115e+02
RS_78 NS_78 0 2.6049933264405115e+02
GL_77 0 NS_77 NS_78 0 2.4648481498152200e-01
GL_78 0 NS_78 NS_77 0 -2.4648481498152200e-01
GS_77_2 0 NS_77 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 8.6892684135916670e+02
RS_80 NS_80 0 8.6892684135916659e+02
GL_79 0 NS_79 NS_80 0 2.4352824357909131e-01
GL_80 0 NS_80 NS_79 0 -2.4352824357909131e-01
GS_79_2 0 NS_79 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 6.5240189890508168e+02
RS_82 NS_82 0 6.5240189890508168e+02
GL_81 0 NS_81 NS_82 0 2.3166276016037468e-01
GL_82 0 NS_82 NS_81 0 -2.3166276016037468e-01
GS_81_2 0 NS_81 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 1.8572469959933156e+02
RS_84 NS_84 0 1.8572469959933156e+02
GL_83 0 NS_83 NS_84 0 2.3351354491929543e-01
GL_84 0 NS_84 NS_83 0 -2.3351354491929543e-01
GS_83_2 0 NS_83 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 3.0631652744794525e+02
RS_86 NS_86 0 3.0631652744794530e+02
GL_85 0 NS_85 NS_86 0 2.3886925224886552e-01
GL_86 0 NS_86 NS_85 0 -2.3886925224886552e-01
GS_85_2 0 NS_85 NA_2 0 1.1283794739964070e+00
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 5.0301469986378567e+02
RS_88 NS_88 0 5.0301469986378567e+02
GL_87 0 NS_87 NS_88 0 2.3692781195536661e-01
GL_88 0 NS_88 NS_87 0 -2.3692781195536661e-01
GS_87_2 0 NS_87 NA_2 0 1.1283794739964070e+00
*
* Real pole n. 89
CS_89 NS_89 0 9.9999999999999998e-13
RS_89 NS_89 0 3.9451851533158515e+00
GS_89_3 0 NS_89 NA_3 0 1.1283794739964070e+00
*
* Real pole n. 90
CS_90 NS_90 0 9.9999999999999998e-13
RS_90 NS_90 0 1.8805154767607480e+01
GS_90_3 0 NS_90 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 1.8483596483142442e+01
RS_92 NS_92 0 1.8483596483142442e+01
GL_91 0 NS_91 NS_92 0 6.9799982353381460e-02
GL_92 0 NS_92 NS_91 0 -6.9799982353381460e-02
GS_91_3 0 NS_91 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 1.9654872352993628e+01
RS_94 NS_94 0 1.9654872352993625e+01
GL_93 0 NS_93 NS_94 0 9.5720932954598423e-02
GL_94 0 NS_94 NS_93 0 -9.5720932954598423e-02
GS_93_3 0 NS_93 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 2.5061544329287912e+01
RS_96 NS_96 0 2.5061544329287909e+01
GL_95 0 NS_95 NS_96 0 1.3536754976539320e-01
GL_96 0 NS_96 NS_95 0 -1.3536754976539320e-01
GS_95_3 0 NS_95 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 7.4239654864745361e+01
RS_98 NS_98 0 7.4239654864745361e+01
GL_97 0 NS_97 NS_98 0 2.8245804011501385e-01
GL_98 0 NS_98 NS_97 0 -2.8245804011501385e-01
GS_97_3 0 NS_97 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 2.8726427419385509e+01
RS_100 NS_100 0 2.8726427419385512e+01
GL_99 0 NS_99 NS_100 0 1.7620265460857126e-01
GL_100 0 NS_100 NS_99 0 -1.7620265460857126e-01
GS_99_3 0 NS_99 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 7.8929016552352451e+01
RS_102 NS_102 0 7.8929016552352465e+01
GL_101 0 NS_101 NS_102 0 1.7267598155977268e-01
GL_102 0 NS_102 NS_101 0 -1.7267598155977268e-01
GS_101_3 0 NS_101 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 1.3876610711235463e+02
RS_104 NS_104 0 1.3876610711235463e+02
GL_103 0 NS_103 NS_104 0 1.9827389109149790e-01
GL_104 0 NS_104 NS_103 0 -1.9827389109149790e-01
GS_103_3 0 NS_103 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 9.4943847388790630e+01
RS_106 NS_106 0 9.4943847388790630e+01
GL_105 0 NS_105 NS_106 0 2.0370912057963636e-01
GL_106 0 NS_106 NS_105 0 -2.0370912057963636e-01
GS_105_3 0 NS_105 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 2.2502148823483816e+02
RS_108 NS_108 0 2.2502148823483816e+02
GL_107 0 NS_107 NS_108 0 2.1140622110318164e-01
GL_108 0 NS_108 NS_107 0 -2.1140622110318164e-01
GS_107_3 0 NS_107 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 2.0359721972446440e+02
RS_110 NS_110 0 2.0359721972446440e+02
GL_109 0 NS_109 NS_110 0 2.1650882528339854e-01
GL_110 0 NS_110 NS_109 0 -2.1650882528339854e-01
GS_109_3 0 NS_109 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 5.4323743269805618e+02
RS_112 NS_112 0 5.4323743269805618e+02
GL_111 0 NS_111 NS_112 0 2.2057741537827197e-01
GL_112 0 NS_112 NS_111 0 -2.2057741537827197e-01
GS_111_3 0 NS_111 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 6.2013592102356057e+01
RS_114 NS_114 0 6.2013592102356057e+01
GL_113 0 NS_113 NS_114 0 2.2721975400227054e-01
GL_114 0 NS_114 NS_113 0 -2.2721975400227054e-01
GS_113_3 0 NS_113 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 8.2527539890421451e+01
RS_116 NS_116 0 8.2527539890421465e+01
GL_115 0 NS_115 NS_116 0 2.2544686857562196e-01
GL_116 0 NS_116 NS_115 0 -2.2544686857562196e-01
GS_115_3 0 NS_115 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 1.5057204740157513e+02
RS_118 NS_118 0 1.5057204740157516e+02
GL_117 0 NS_117 NS_118 0 2.5030962700427895e-01
GL_118 0 NS_118 NS_117 0 -2.5030962700427895e-01
GS_117_3 0 NS_117 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 1.0143406310664166e+03
RS_120 NS_120 0 1.0143406310664167e+03
GL_119 0 NS_119 NS_120 0 2.4802996115452441e-01
GL_120 0 NS_120 NS_119 0 -2.4802996115452441e-01
GS_119_3 0 NS_119 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 2.6049933264405115e+02
RS_122 NS_122 0 2.6049933264405115e+02
GL_121 0 NS_121 NS_122 0 2.4648481498152200e-01
GL_122 0 NS_122 NS_121 0 -2.4648481498152200e-01
GS_121_3 0 NS_121 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 8.6892684135916670e+02
RS_124 NS_124 0 8.6892684135916659e+02
GL_123 0 NS_123 NS_124 0 2.4352824357909131e-01
GL_124 0 NS_124 NS_123 0 -2.4352824357909131e-01
GS_123_3 0 NS_123 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 6.5240189890508168e+02
RS_126 NS_126 0 6.5240189890508168e+02
GL_125 0 NS_125 NS_126 0 2.3166276016037468e-01
GL_126 0 NS_126 NS_125 0 -2.3166276016037468e-01
GS_125_3 0 NS_125 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 1.8572469959933156e+02
RS_128 NS_128 0 1.8572469959933156e+02
GL_127 0 NS_127 NS_128 0 2.3351354491929543e-01
GL_128 0 NS_128 NS_127 0 -2.3351354491929543e-01
GS_127_3 0 NS_127 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 3.0631652744794525e+02
RS_130 NS_130 0 3.0631652744794530e+02
GL_129 0 NS_129 NS_130 0 2.3886925224886552e-01
GL_130 0 NS_130 NS_129 0 -2.3886925224886552e-01
GS_129_3 0 NS_129 NA_3 0 1.1283794739964070e+00
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 5.0301469986378567e+02
RS_132 NS_132 0 5.0301469986378567e+02
GL_131 0 NS_131 NS_132 0 2.3692781195536661e-01
GL_132 0 NS_132 NS_131 0 -2.3692781195536661e-01
GS_131_3 0 NS_131 NA_3 0 1.1283794739964070e+00
*
* Real pole n. 133
CS_133 NS_133 0 9.9999999999999998e-13
RS_133 NS_133 0 3.9451851533158515e+00
GS_133_4 0 NS_133 NA_4 0 1.1283794739964070e+00
*
* Real pole n. 134
CS_134 NS_134 0 9.9999999999999998e-13
RS_134 NS_134 0 1.8805154767607480e+01
GS_134_4 0 NS_134 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 1.8483596483142442e+01
RS_136 NS_136 0 1.8483596483142442e+01
GL_135 0 NS_135 NS_136 0 6.9799982353381460e-02
GL_136 0 NS_136 NS_135 0 -6.9799982353381460e-02
GS_135_4 0 NS_135 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 1.9654872352993628e+01
RS_138 NS_138 0 1.9654872352993625e+01
GL_137 0 NS_137 NS_138 0 9.5720932954598423e-02
GL_138 0 NS_138 NS_137 0 -9.5720932954598423e-02
GS_137_4 0 NS_137 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 2.5061544329287912e+01
RS_140 NS_140 0 2.5061544329287909e+01
GL_139 0 NS_139 NS_140 0 1.3536754976539320e-01
GL_140 0 NS_140 NS_139 0 -1.3536754976539320e-01
GS_139_4 0 NS_139 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 7.4239654864745361e+01
RS_142 NS_142 0 7.4239654864745361e+01
GL_141 0 NS_141 NS_142 0 2.8245804011501385e-01
GL_142 0 NS_142 NS_141 0 -2.8245804011501385e-01
GS_141_4 0 NS_141 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 2.8726427419385509e+01
RS_144 NS_144 0 2.8726427419385512e+01
GL_143 0 NS_143 NS_144 0 1.7620265460857126e-01
GL_144 0 NS_144 NS_143 0 -1.7620265460857126e-01
GS_143_4 0 NS_143 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 7.8929016552352451e+01
RS_146 NS_146 0 7.8929016552352465e+01
GL_145 0 NS_145 NS_146 0 1.7267598155977268e-01
GL_146 0 NS_146 NS_145 0 -1.7267598155977268e-01
GS_145_4 0 NS_145 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 1.3876610711235463e+02
RS_148 NS_148 0 1.3876610711235463e+02
GL_147 0 NS_147 NS_148 0 1.9827389109149790e-01
GL_148 0 NS_148 NS_147 0 -1.9827389109149790e-01
GS_147_4 0 NS_147 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 9.4943847388790630e+01
RS_150 NS_150 0 9.4943847388790630e+01
GL_149 0 NS_149 NS_150 0 2.0370912057963636e-01
GL_150 0 NS_150 NS_149 0 -2.0370912057963636e-01
GS_149_4 0 NS_149 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 2.2502148823483816e+02
RS_152 NS_152 0 2.2502148823483816e+02
GL_151 0 NS_151 NS_152 0 2.1140622110318164e-01
GL_152 0 NS_152 NS_151 0 -2.1140622110318164e-01
GS_151_4 0 NS_151 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 2.0359721972446440e+02
RS_154 NS_154 0 2.0359721972446440e+02
GL_153 0 NS_153 NS_154 0 2.1650882528339854e-01
GL_154 0 NS_154 NS_153 0 -2.1650882528339854e-01
GS_153_4 0 NS_153 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 5.4323743269805618e+02
RS_156 NS_156 0 5.4323743269805618e+02
GL_155 0 NS_155 NS_156 0 2.2057741537827197e-01
GL_156 0 NS_156 NS_155 0 -2.2057741537827197e-01
GS_155_4 0 NS_155 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 6.2013592102356057e+01
RS_158 NS_158 0 6.2013592102356057e+01
GL_157 0 NS_157 NS_158 0 2.2721975400227054e-01
GL_158 0 NS_158 NS_157 0 -2.2721975400227054e-01
GS_157_4 0 NS_157 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 8.2527539890421451e+01
RS_160 NS_160 0 8.2527539890421465e+01
GL_159 0 NS_159 NS_160 0 2.2544686857562196e-01
GL_160 0 NS_160 NS_159 0 -2.2544686857562196e-01
GS_159_4 0 NS_159 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 1.5057204740157513e+02
RS_162 NS_162 0 1.5057204740157516e+02
GL_161 0 NS_161 NS_162 0 2.5030962700427895e-01
GL_162 0 NS_162 NS_161 0 -2.5030962700427895e-01
GS_161_4 0 NS_161 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 163/164
CS_163 NS_163 0 9.9999999999999998e-13
CS_164 NS_164 0 9.9999999999999998e-13
RS_163 NS_163 0 1.0143406310664166e+03
RS_164 NS_164 0 1.0143406310664167e+03
GL_163 0 NS_163 NS_164 0 2.4802996115452441e-01
GL_164 0 NS_164 NS_163 0 -2.4802996115452441e-01
GS_163_4 0 NS_163 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 2.6049933264405115e+02
RS_166 NS_166 0 2.6049933264405115e+02
GL_165 0 NS_165 NS_166 0 2.4648481498152200e-01
GL_166 0 NS_166 NS_165 0 -2.4648481498152200e-01
GS_165_4 0 NS_165 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 8.6892684135916670e+02
RS_168 NS_168 0 8.6892684135916659e+02
GL_167 0 NS_167 NS_168 0 2.4352824357909131e-01
GL_168 0 NS_168 NS_167 0 -2.4352824357909131e-01
GS_167_4 0 NS_167 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 6.5240189890508168e+02
RS_170 NS_170 0 6.5240189890508168e+02
GL_169 0 NS_169 NS_170 0 2.3166276016037468e-01
GL_170 0 NS_170 NS_169 0 -2.3166276016037468e-01
GS_169_4 0 NS_169 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 1.8572469959933156e+02
RS_172 NS_172 0 1.8572469959933156e+02
GL_171 0 NS_171 NS_172 0 2.3351354491929543e-01
GL_172 0 NS_172 NS_171 0 -2.3351354491929543e-01
GS_171_4 0 NS_171 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 3.0631652744794525e+02
RS_174 NS_174 0 3.0631652744794530e+02
GL_173 0 NS_173 NS_174 0 2.3886925224886552e-01
GL_174 0 NS_174 NS_173 0 -2.3886925224886552e-01
GS_173_4 0 NS_173 NA_4 0 1.1283794739964070e+00
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 5.0301469986378567e+02
RS_176 NS_176 0 5.0301469986378567e+02
GL_175 0 NS_175 NS_176 0 2.3692781195536661e-01
GL_176 0 NS_176 NS_175 0 -2.3692781195536661e-01
GS_175_4 0 NS_175 NA_4 0 1.1283794739964070e+00
*
* Real pole n. 177
CS_177 NS_177 0 9.9999999999999998e-13
RS_177 NS_177 0 3.9451851533158515e+00
GS_177_5 0 NS_177 NA_5 0 1.1283794739964070e+00
*
* Real pole n. 178
CS_178 NS_178 0 9.9999999999999998e-13
RS_178 NS_178 0 1.8805154767607480e+01
GS_178_5 0 NS_178 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 1.8483596483142442e+01
RS_180 NS_180 0 1.8483596483142442e+01
GL_179 0 NS_179 NS_180 0 6.9799982353381460e-02
GL_180 0 NS_180 NS_179 0 -6.9799982353381460e-02
GS_179_5 0 NS_179 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 181/182
CS_181 NS_181 0 9.9999999999999998e-13
CS_182 NS_182 0 9.9999999999999998e-13
RS_181 NS_181 0 1.9654872352993628e+01
RS_182 NS_182 0 1.9654872352993625e+01
GL_181 0 NS_181 NS_182 0 9.5720932954598423e-02
GL_182 0 NS_182 NS_181 0 -9.5720932954598423e-02
GS_181_5 0 NS_181 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 183/184
CS_183 NS_183 0 9.9999999999999998e-13
CS_184 NS_184 0 9.9999999999999998e-13
RS_183 NS_183 0 2.5061544329287912e+01
RS_184 NS_184 0 2.5061544329287909e+01
GL_183 0 NS_183 NS_184 0 1.3536754976539320e-01
GL_184 0 NS_184 NS_183 0 -1.3536754976539320e-01
GS_183_5 0 NS_183 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 7.4239654864745361e+01
RS_186 NS_186 0 7.4239654864745361e+01
GL_185 0 NS_185 NS_186 0 2.8245804011501385e-01
GL_186 0 NS_186 NS_185 0 -2.8245804011501385e-01
GS_185_5 0 NS_185 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 2.8726427419385509e+01
RS_188 NS_188 0 2.8726427419385512e+01
GL_187 0 NS_187 NS_188 0 1.7620265460857126e-01
GL_188 0 NS_188 NS_187 0 -1.7620265460857126e-01
GS_187_5 0 NS_187 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 7.8929016552352451e+01
RS_190 NS_190 0 7.8929016552352465e+01
GL_189 0 NS_189 NS_190 0 1.7267598155977268e-01
GL_190 0 NS_190 NS_189 0 -1.7267598155977268e-01
GS_189_5 0 NS_189 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 1.3876610711235463e+02
RS_192 NS_192 0 1.3876610711235463e+02
GL_191 0 NS_191 NS_192 0 1.9827389109149790e-01
GL_192 0 NS_192 NS_191 0 -1.9827389109149790e-01
GS_191_5 0 NS_191 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 9.4943847388790630e+01
RS_194 NS_194 0 9.4943847388790630e+01
GL_193 0 NS_193 NS_194 0 2.0370912057963636e-01
GL_194 0 NS_194 NS_193 0 -2.0370912057963636e-01
GS_193_5 0 NS_193 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 2.2502148823483816e+02
RS_196 NS_196 0 2.2502148823483816e+02
GL_195 0 NS_195 NS_196 0 2.1140622110318164e-01
GL_196 0 NS_196 NS_195 0 -2.1140622110318164e-01
GS_195_5 0 NS_195 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 2.0359721972446440e+02
RS_198 NS_198 0 2.0359721972446440e+02
GL_197 0 NS_197 NS_198 0 2.1650882528339854e-01
GL_198 0 NS_198 NS_197 0 -2.1650882528339854e-01
GS_197_5 0 NS_197 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 5.4323743269805618e+02
RS_200 NS_200 0 5.4323743269805618e+02
GL_199 0 NS_199 NS_200 0 2.2057741537827197e-01
GL_200 0 NS_200 NS_199 0 -2.2057741537827197e-01
GS_199_5 0 NS_199 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 201/202
CS_201 NS_201 0 9.9999999999999998e-13
CS_202 NS_202 0 9.9999999999999998e-13
RS_201 NS_201 0 6.2013592102356057e+01
RS_202 NS_202 0 6.2013592102356057e+01
GL_201 0 NS_201 NS_202 0 2.2721975400227054e-01
GL_202 0 NS_202 NS_201 0 -2.2721975400227054e-01
GS_201_5 0 NS_201 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 203/204
CS_203 NS_203 0 9.9999999999999998e-13
CS_204 NS_204 0 9.9999999999999998e-13
RS_203 NS_203 0 8.2527539890421451e+01
RS_204 NS_204 0 8.2527539890421465e+01
GL_203 0 NS_203 NS_204 0 2.2544686857562196e-01
GL_204 0 NS_204 NS_203 0 -2.2544686857562196e-01
GS_203_5 0 NS_203 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 1.5057204740157513e+02
RS_206 NS_206 0 1.5057204740157516e+02
GL_205 0 NS_205 NS_206 0 2.5030962700427895e-01
GL_206 0 NS_206 NS_205 0 -2.5030962700427895e-01
GS_205_5 0 NS_205 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 1.0143406310664166e+03
RS_208 NS_208 0 1.0143406310664167e+03
GL_207 0 NS_207 NS_208 0 2.4802996115452441e-01
GL_208 0 NS_208 NS_207 0 -2.4802996115452441e-01
GS_207_5 0 NS_207 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 2.6049933264405115e+02
RS_210 NS_210 0 2.6049933264405115e+02
GL_209 0 NS_209 NS_210 0 2.4648481498152200e-01
GL_210 0 NS_210 NS_209 0 -2.4648481498152200e-01
GS_209_5 0 NS_209 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 8.6892684135916670e+02
RS_212 NS_212 0 8.6892684135916659e+02
GL_211 0 NS_211 NS_212 0 2.4352824357909131e-01
GL_212 0 NS_212 NS_211 0 -2.4352824357909131e-01
GS_211_5 0 NS_211 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 6.5240189890508168e+02
RS_214 NS_214 0 6.5240189890508168e+02
GL_213 0 NS_213 NS_214 0 2.3166276016037468e-01
GL_214 0 NS_214 NS_213 0 -2.3166276016037468e-01
GS_213_5 0 NS_213 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 1.8572469959933156e+02
RS_216 NS_216 0 1.8572469959933156e+02
GL_215 0 NS_215 NS_216 0 2.3351354491929543e-01
GL_216 0 NS_216 NS_215 0 -2.3351354491929543e-01
GS_215_5 0 NS_215 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 3.0631652744794525e+02
RS_218 NS_218 0 3.0631652744794530e+02
GL_217 0 NS_217 NS_218 0 2.3886925224886552e-01
GL_218 0 NS_218 NS_217 0 -2.3886925224886552e-01
GS_217_5 0 NS_217 NA_5 0 1.1283794739964070e+00
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 5.0301469986378567e+02
RS_220 NS_220 0 5.0301469986378567e+02
GL_219 0 NS_219 NS_220 0 2.3692781195536661e-01
GL_220 0 NS_220 NS_219 0 -2.3692781195536661e-01
GS_219_5 0 NS_219 NA_5 0 1.1283794739964070e+00
*
* Real pole n. 221
CS_221 NS_221 0 9.9999999999999998e-13
RS_221 NS_221 0 3.9451851533158515e+00
GS_221_6 0 NS_221 NA_6 0 1.1283794739964070e+00
*
* Real pole n. 222
CS_222 NS_222 0 9.9999999999999998e-13
RS_222 NS_222 0 1.8805154767607480e+01
GS_222_6 0 NS_222 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 223/224
CS_223 NS_223 0 9.9999999999999998e-13
CS_224 NS_224 0 9.9999999999999998e-13
RS_223 NS_223 0 1.8483596483142442e+01
RS_224 NS_224 0 1.8483596483142442e+01
GL_223 0 NS_223 NS_224 0 6.9799982353381460e-02
GL_224 0 NS_224 NS_223 0 -6.9799982353381460e-02
GS_223_6 0 NS_223 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 225/226
CS_225 NS_225 0 9.9999999999999998e-13
CS_226 NS_226 0 9.9999999999999998e-13
RS_225 NS_225 0 1.9654872352993628e+01
RS_226 NS_226 0 1.9654872352993625e+01
GL_225 0 NS_225 NS_226 0 9.5720932954598423e-02
GL_226 0 NS_226 NS_225 0 -9.5720932954598423e-02
GS_225_6 0 NS_225 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 2.5061544329287912e+01
RS_228 NS_228 0 2.5061544329287909e+01
GL_227 0 NS_227 NS_228 0 1.3536754976539320e-01
GL_228 0 NS_228 NS_227 0 -1.3536754976539320e-01
GS_227_6 0 NS_227 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 229/230
CS_229 NS_229 0 9.9999999999999998e-13
CS_230 NS_230 0 9.9999999999999998e-13
RS_229 NS_229 0 7.4239654864745361e+01
RS_230 NS_230 0 7.4239654864745361e+01
GL_229 0 NS_229 NS_230 0 2.8245804011501385e-01
GL_230 0 NS_230 NS_229 0 -2.8245804011501385e-01
GS_229_6 0 NS_229 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 2.8726427419385509e+01
RS_232 NS_232 0 2.8726427419385512e+01
GL_231 0 NS_231 NS_232 0 1.7620265460857126e-01
GL_232 0 NS_232 NS_231 0 -1.7620265460857126e-01
GS_231_6 0 NS_231 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 7.8929016552352451e+01
RS_234 NS_234 0 7.8929016552352465e+01
GL_233 0 NS_233 NS_234 0 1.7267598155977268e-01
GL_234 0 NS_234 NS_233 0 -1.7267598155977268e-01
GS_233_6 0 NS_233 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 1.3876610711235463e+02
RS_236 NS_236 0 1.3876610711235463e+02
GL_235 0 NS_235 NS_236 0 1.9827389109149790e-01
GL_236 0 NS_236 NS_235 0 -1.9827389109149790e-01
GS_235_6 0 NS_235 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 9.4943847388790630e+01
RS_238 NS_238 0 9.4943847388790630e+01
GL_237 0 NS_237 NS_238 0 2.0370912057963636e-01
GL_238 0 NS_238 NS_237 0 -2.0370912057963636e-01
GS_237_6 0 NS_237 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 2.2502148823483816e+02
RS_240 NS_240 0 2.2502148823483816e+02
GL_239 0 NS_239 NS_240 0 2.1140622110318164e-01
GL_240 0 NS_240 NS_239 0 -2.1140622110318164e-01
GS_239_6 0 NS_239 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 241/242
CS_241 NS_241 0 9.9999999999999998e-13
CS_242 NS_242 0 9.9999999999999998e-13
RS_241 NS_241 0 2.0359721972446440e+02
RS_242 NS_242 0 2.0359721972446440e+02
GL_241 0 NS_241 NS_242 0 2.1650882528339854e-01
GL_242 0 NS_242 NS_241 0 -2.1650882528339854e-01
GS_241_6 0 NS_241 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 243/244
CS_243 NS_243 0 9.9999999999999998e-13
CS_244 NS_244 0 9.9999999999999998e-13
RS_243 NS_243 0 5.4323743269805618e+02
RS_244 NS_244 0 5.4323743269805618e+02
GL_243 0 NS_243 NS_244 0 2.2057741537827197e-01
GL_244 0 NS_244 NS_243 0 -2.2057741537827197e-01
GS_243_6 0 NS_243 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 245/246
CS_245 NS_245 0 9.9999999999999998e-13
CS_246 NS_246 0 9.9999999999999998e-13
RS_245 NS_245 0 6.2013592102356057e+01
RS_246 NS_246 0 6.2013592102356057e+01
GL_245 0 NS_245 NS_246 0 2.2721975400227054e-01
GL_246 0 NS_246 NS_245 0 -2.2721975400227054e-01
GS_245_6 0 NS_245 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 247/248
CS_247 NS_247 0 9.9999999999999998e-13
CS_248 NS_248 0 9.9999999999999998e-13
RS_247 NS_247 0 8.2527539890421451e+01
RS_248 NS_248 0 8.2527539890421465e+01
GL_247 0 NS_247 NS_248 0 2.2544686857562196e-01
GL_248 0 NS_248 NS_247 0 -2.2544686857562196e-01
GS_247_6 0 NS_247 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 249/250
CS_249 NS_249 0 9.9999999999999998e-13
CS_250 NS_250 0 9.9999999999999998e-13
RS_249 NS_249 0 1.5057204740157513e+02
RS_250 NS_250 0 1.5057204740157516e+02
GL_249 0 NS_249 NS_250 0 2.5030962700427895e-01
GL_250 0 NS_250 NS_249 0 -2.5030962700427895e-01
GS_249_6 0 NS_249 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 251/252
CS_251 NS_251 0 9.9999999999999998e-13
CS_252 NS_252 0 9.9999999999999998e-13
RS_251 NS_251 0 1.0143406310664166e+03
RS_252 NS_252 0 1.0143406310664167e+03
GL_251 0 NS_251 NS_252 0 2.4802996115452441e-01
GL_252 0 NS_252 NS_251 0 -2.4802996115452441e-01
GS_251_6 0 NS_251 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 253/254
CS_253 NS_253 0 9.9999999999999998e-13
CS_254 NS_254 0 9.9999999999999998e-13
RS_253 NS_253 0 2.6049933264405115e+02
RS_254 NS_254 0 2.6049933264405115e+02
GL_253 0 NS_253 NS_254 0 2.4648481498152200e-01
GL_254 0 NS_254 NS_253 0 -2.4648481498152200e-01
GS_253_6 0 NS_253 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 255/256
CS_255 NS_255 0 9.9999999999999998e-13
CS_256 NS_256 0 9.9999999999999998e-13
RS_255 NS_255 0 8.6892684135916670e+02
RS_256 NS_256 0 8.6892684135916659e+02
GL_255 0 NS_255 NS_256 0 2.4352824357909131e-01
GL_256 0 NS_256 NS_255 0 -2.4352824357909131e-01
GS_255_6 0 NS_255 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 257/258
CS_257 NS_257 0 9.9999999999999998e-13
CS_258 NS_258 0 9.9999999999999998e-13
RS_257 NS_257 0 6.5240189890508168e+02
RS_258 NS_258 0 6.5240189890508168e+02
GL_257 0 NS_257 NS_258 0 2.3166276016037468e-01
GL_258 0 NS_258 NS_257 0 -2.3166276016037468e-01
GS_257_6 0 NS_257 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 259/260
CS_259 NS_259 0 9.9999999999999998e-13
CS_260 NS_260 0 9.9999999999999998e-13
RS_259 NS_259 0 1.8572469959933156e+02
RS_260 NS_260 0 1.8572469959933156e+02
GL_259 0 NS_259 NS_260 0 2.3351354491929543e-01
GL_260 0 NS_260 NS_259 0 -2.3351354491929543e-01
GS_259_6 0 NS_259 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 261/262
CS_261 NS_261 0 9.9999999999999998e-13
CS_262 NS_262 0 9.9999999999999998e-13
RS_261 NS_261 0 3.0631652744794525e+02
RS_262 NS_262 0 3.0631652744794530e+02
GL_261 0 NS_261 NS_262 0 2.3886925224886552e-01
GL_262 0 NS_262 NS_261 0 -2.3886925224886552e-01
GS_261_6 0 NS_261 NA_6 0 1.1283794739964070e+00
*
* Complex pair n. 263/264
CS_263 NS_263 0 9.9999999999999998e-13
CS_264 NS_264 0 9.9999999999999998e-13
RS_263 NS_263 0 5.0301469986378567e+02
RS_264 NS_264 0 5.0301469986378567e+02
GL_263 0 NS_263 NS_264 0 2.3692781195536661e-01
GL_264 0 NS_264 NS_263 0 -2.3692781195536661e-01
GS_263_6 0 NS_263 NA_6 0 1.1283794739964070e+00
*
* Real pole n. 265
CS_265 NS_265 0 9.9999999999999998e-13
RS_265 NS_265 0 3.9451851533158515e+00
GS_265_7 0 NS_265 NA_7 0 1.1283794739964070e+00
*
* Real pole n. 266
CS_266 NS_266 0 9.9999999999999998e-13
RS_266 NS_266 0 1.8805154767607480e+01
GS_266_7 0 NS_266 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 267/268
CS_267 NS_267 0 9.9999999999999998e-13
CS_268 NS_268 0 9.9999999999999998e-13
RS_267 NS_267 0 1.8483596483142442e+01
RS_268 NS_268 0 1.8483596483142442e+01
GL_267 0 NS_267 NS_268 0 6.9799982353381460e-02
GL_268 0 NS_268 NS_267 0 -6.9799982353381460e-02
GS_267_7 0 NS_267 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 269/270
CS_269 NS_269 0 9.9999999999999998e-13
CS_270 NS_270 0 9.9999999999999998e-13
RS_269 NS_269 0 1.9654872352993628e+01
RS_270 NS_270 0 1.9654872352993625e+01
GL_269 0 NS_269 NS_270 0 9.5720932954598423e-02
GL_270 0 NS_270 NS_269 0 -9.5720932954598423e-02
GS_269_7 0 NS_269 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 271/272
CS_271 NS_271 0 9.9999999999999998e-13
CS_272 NS_272 0 9.9999999999999998e-13
RS_271 NS_271 0 2.5061544329287912e+01
RS_272 NS_272 0 2.5061544329287909e+01
GL_271 0 NS_271 NS_272 0 1.3536754976539320e-01
GL_272 0 NS_272 NS_271 0 -1.3536754976539320e-01
GS_271_7 0 NS_271 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 273/274
CS_273 NS_273 0 9.9999999999999998e-13
CS_274 NS_274 0 9.9999999999999998e-13
RS_273 NS_273 0 7.4239654864745361e+01
RS_274 NS_274 0 7.4239654864745361e+01
GL_273 0 NS_273 NS_274 0 2.8245804011501385e-01
GL_274 0 NS_274 NS_273 0 -2.8245804011501385e-01
GS_273_7 0 NS_273 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 275/276
CS_275 NS_275 0 9.9999999999999998e-13
CS_276 NS_276 0 9.9999999999999998e-13
RS_275 NS_275 0 2.8726427419385509e+01
RS_276 NS_276 0 2.8726427419385512e+01
GL_275 0 NS_275 NS_276 0 1.7620265460857126e-01
GL_276 0 NS_276 NS_275 0 -1.7620265460857126e-01
GS_275_7 0 NS_275 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 277/278
CS_277 NS_277 0 9.9999999999999998e-13
CS_278 NS_278 0 9.9999999999999998e-13
RS_277 NS_277 0 7.8929016552352451e+01
RS_278 NS_278 0 7.8929016552352465e+01
GL_277 0 NS_277 NS_278 0 1.7267598155977268e-01
GL_278 0 NS_278 NS_277 0 -1.7267598155977268e-01
GS_277_7 0 NS_277 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 279/280
CS_279 NS_279 0 9.9999999999999998e-13
CS_280 NS_280 0 9.9999999999999998e-13
RS_279 NS_279 0 1.3876610711235463e+02
RS_280 NS_280 0 1.3876610711235463e+02
GL_279 0 NS_279 NS_280 0 1.9827389109149790e-01
GL_280 0 NS_280 NS_279 0 -1.9827389109149790e-01
GS_279_7 0 NS_279 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 281/282
CS_281 NS_281 0 9.9999999999999998e-13
CS_282 NS_282 0 9.9999999999999998e-13
RS_281 NS_281 0 9.4943847388790630e+01
RS_282 NS_282 0 9.4943847388790630e+01
GL_281 0 NS_281 NS_282 0 2.0370912057963636e-01
GL_282 0 NS_282 NS_281 0 -2.0370912057963636e-01
GS_281_7 0 NS_281 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 283/284
CS_283 NS_283 0 9.9999999999999998e-13
CS_284 NS_284 0 9.9999999999999998e-13
RS_283 NS_283 0 2.2502148823483816e+02
RS_284 NS_284 0 2.2502148823483816e+02
GL_283 0 NS_283 NS_284 0 2.1140622110318164e-01
GL_284 0 NS_284 NS_283 0 -2.1140622110318164e-01
GS_283_7 0 NS_283 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 285/286
CS_285 NS_285 0 9.9999999999999998e-13
CS_286 NS_286 0 9.9999999999999998e-13
RS_285 NS_285 0 2.0359721972446440e+02
RS_286 NS_286 0 2.0359721972446440e+02
GL_285 0 NS_285 NS_286 0 2.1650882528339854e-01
GL_286 0 NS_286 NS_285 0 -2.1650882528339854e-01
GS_285_7 0 NS_285 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 287/288
CS_287 NS_287 0 9.9999999999999998e-13
CS_288 NS_288 0 9.9999999999999998e-13
RS_287 NS_287 0 5.4323743269805618e+02
RS_288 NS_288 0 5.4323743269805618e+02
GL_287 0 NS_287 NS_288 0 2.2057741537827197e-01
GL_288 0 NS_288 NS_287 0 -2.2057741537827197e-01
GS_287_7 0 NS_287 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 289/290
CS_289 NS_289 0 9.9999999999999998e-13
CS_290 NS_290 0 9.9999999999999998e-13
RS_289 NS_289 0 6.2013592102356057e+01
RS_290 NS_290 0 6.2013592102356057e+01
GL_289 0 NS_289 NS_290 0 2.2721975400227054e-01
GL_290 0 NS_290 NS_289 0 -2.2721975400227054e-01
GS_289_7 0 NS_289 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 291/292
CS_291 NS_291 0 9.9999999999999998e-13
CS_292 NS_292 0 9.9999999999999998e-13
RS_291 NS_291 0 8.2527539890421451e+01
RS_292 NS_292 0 8.2527539890421465e+01
GL_291 0 NS_291 NS_292 0 2.2544686857562196e-01
GL_292 0 NS_292 NS_291 0 -2.2544686857562196e-01
GS_291_7 0 NS_291 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 293/294
CS_293 NS_293 0 9.9999999999999998e-13
CS_294 NS_294 0 9.9999999999999998e-13
RS_293 NS_293 0 1.5057204740157513e+02
RS_294 NS_294 0 1.5057204740157516e+02
GL_293 0 NS_293 NS_294 0 2.5030962700427895e-01
GL_294 0 NS_294 NS_293 0 -2.5030962700427895e-01
GS_293_7 0 NS_293 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 295/296
CS_295 NS_295 0 9.9999999999999998e-13
CS_296 NS_296 0 9.9999999999999998e-13
RS_295 NS_295 0 1.0143406310664166e+03
RS_296 NS_296 0 1.0143406310664167e+03
GL_295 0 NS_295 NS_296 0 2.4802996115452441e-01
GL_296 0 NS_296 NS_295 0 -2.4802996115452441e-01
GS_295_7 0 NS_295 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 297/298
CS_297 NS_297 0 9.9999999999999998e-13
CS_298 NS_298 0 9.9999999999999998e-13
RS_297 NS_297 0 2.6049933264405115e+02
RS_298 NS_298 0 2.6049933264405115e+02
GL_297 0 NS_297 NS_298 0 2.4648481498152200e-01
GL_298 0 NS_298 NS_297 0 -2.4648481498152200e-01
GS_297_7 0 NS_297 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 299/300
CS_299 NS_299 0 9.9999999999999998e-13
CS_300 NS_300 0 9.9999999999999998e-13
RS_299 NS_299 0 8.6892684135916670e+02
RS_300 NS_300 0 8.6892684135916659e+02
GL_299 0 NS_299 NS_300 0 2.4352824357909131e-01
GL_300 0 NS_300 NS_299 0 -2.4352824357909131e-01
GS_299_7 0 NS_299 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 301/302
CS_301 NS_301 0 9.9999999999999998e-13
CS_302 NS_302 0 9.9999999999999998e-13
RS_301 NS_301 0 6.5240189890508168e+02
RS_302 NS_302 0 6.5240189890508168e+02
GL_301 0 NS_301 NS_302 0 2.3166276016037468e-01
GL_302 0 NS_302 NS_301 0 -2.3166276016037468e-01
GS_301_7 0 NS_301 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 303/304
CS_303 NS_303 0 9.9999999999999998e-13
CS_304 NS_304 0 9.9999999999999998e-13
RS_303 NS_303 0 1.8572469959933156e+02
RS_304 NS_304 0 1.8572469959933156e+02
GL_303 0 NS_303 NS_304 0 2.3351354491929543e-01
GL_304 0 NS_304 NS_303 0 -2.3351354491929543e-01
GS_303_7 0 NS_303 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 305/306
CS_305 NS_305 0 9.9999999999999998e-13
CS_306 NS_306 0 9.9999999999999998e-13
RS_305 NS_305 0 3.0631652744794525e+02
RS_306 NS_306 0 3.0631652744794530e+02
GL_305 0 NS_305 NS_306 0 2.3886925224886552e-01
GL_306 0 NS_306 NS_305 0 -2.3886925224886552e-01
GS_305_7 0 NS_305 NA_7 0 1.1283794739964070e+00
*
* Complex pair n. 307/308
CS_307 NS_307 0 9.9999999999999998e-13
CS_308 NS_308 0 9.9999999999999998e-13
RS_307 NS_307 0 5.0301469986378567e+02
RS_308 NS_308 0 5.0301469986378567e+02
GL_307 0 NS_307 NS_308 0 2.3692781195536661e-01
GL_308 0 NS_308 NS_307 0 -2.3692781195536661e-01
GS_307_7 0 NS_307 NA_7 0 1.1283794739964070e+00
*
* Real pole n. 309
CS_309 NS_309 0 9.9999999999999998e-13
RS_309 NS_309 0 3.9451851533158515e+00
GS_309_8 0 NS_309 NA_8 0 1.1283794739964070e+00
*
* Real pole n. 310
CS_310 NS_310 0 9.9999999999999998e-13
RS_310 NS_310 0 1.8805154767607480e+01
GS_310_8 0 NS_310 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 311/312
CS_311 NS_311 0 9.9999999999999998e-13
CS_312 NS_312 0 9.9999999999999998e-13
RS_311 NS_311 0 1.8483596483142442e+01
RS_312 NS_312 0 1.8483596483142442e+01
GL_311 0 NS_311 NS_312 0 6.9799982353381460e-02
GL_312 0 NS_312 NS_311 0 -6.9799982353381460e-02
GS_311_8 0 NS_311 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 313/314
CS_313 NS_313 0 9.9999999999999998e-13
CS_314 NS_314 0 9.9999999999999998e-13
RS_313 NS_313 0 1.9654872352993628e+01
RS_314 NS_314 0 1.9654872352993625e+01
GL_313 0 NS_313 NS_314 0 9.5720932954598423e-02
GL_314 0 NS_314 NS_313 0 -9.5720932954598423e-02
GS_313_8 0 NS_313 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 315/316
CS_315 NS_315 0 9.9999999999999998e-13
CS_316 NS_316 0 9.9999999999999998e-13
RS_315 NS_315 0 2.5061544329287912e+01
RS_316 NS_316 0 2.5061544329287909e+01
GL_315 0 NS_315 NS_316 0 1.3536754976539320e-01
GL_316 0 NS_316 NS_315 0 -1.3536754976539320e-01
GS_315_8 0 NS_315 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 317/318
CS_317 NS_317 0 9.9999999999999998e-13
CS_318 NS_318 0 9.9999999999999998e-13
RS_317 NS_317 0 7.4239654864745361e+01
RS_318 NS_318 0 7.4239654864745361e+01
GL_317 0 NS_317 NS_318 0 2.8245804011501385e-01
GL_318 0 NS_318 NS_317 0 -2.8245804011501385e-01
GS_317_8 0 NS_317 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 319/320
CS_319 NS_319 0 9.9999999999999998e-13
CS_320 NS_320 0 9.9999999999999998e-13
RS_319 NS_319 0 2.8726427419385509e+01
RS_320 NS_320 0 2.8726427419385512e+01
GL_319 0 NS_319 NS_320 0 1.7620265460857126e-01
GL_320 0 NS_320 NS_319 0 -1.7620265460857126e-01
GS_319_8 0 NS_319 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 321/322
CS_321 NS_321 0 9.9999999999999998e-13
CS_322 NS_322 0 9.9999999999999998e-13
RS_321 NS_321 0 7.8929016552352451e+01
RS_322 NS_322 0 7.8929016552352465e+01
GL_321 0 NS_321 NS_322 0 1.7267598155977268e-01
GL_322 0 NS_322 NS_321 0 -1.7267598155977268e-01
GS_321_8 0 NS_321 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 323/324
CS_323 NS_323 0 9.9999999999999998e-13
CS_324 NS_324 0 9.9999999999999998e-13
RS_323 NS_323 0 1.3876610711235463e+02
RS_324 NS_324 0 1.3876610711235463e+02
GL_323 0 NS_323 NS_324 0 1.9827389109149790e-01
GL_324 0 NS_324 NS_323 0 -1.9827389109149790e-01
GS_323_8 0 NS_323 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 325/326
CS_325 NS_325 0 9.9999999999999998e-13
CS_326 NS_326 0 9.9999999999999998e-13
RS_325 NS_325 0 9.4943847388790630e+01
RS_326 NS_326 0 9.4943847388790630e+01
GL_325 0 NS_325 NS_326 0 2.0370912057963636e-01
GL_326 0 NS_326 NS_325 0 -2.0370912057963636e-01
GS_325_8 0 NS_325 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 327/328
CS_327 NS_327 0 9.9999999999999998e-13
CS_328 NS_328 0 9.9999999999999998e-13
RS_327 NS_327 0 2.2502148823483816e+02
RS_328 NS_328 0 2.2502148823483816e+02
GL_327 0 NS_327 NS_328 0 2.1140622110318164e-01
GL_328 0 NS_328 NS_327 0 -2.1140622110318164e-01
GS_327_8 0 NS_327 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 329/330
CS_329 NS_329 0 9.9999999999999998e-13
CS_330 NS_330 0 9.9999999999999998e-13
RS_329 NS_329 0 2.0359721972446440e+02
RS_330 NS_330 0 2.0359721972446440e+02
GL_329 0 NS_329 NS_330 0 2.1650882528339854e-01
GL_330 0 NS_330 NS_329 0 -2.1650882528339854e-01
GS_329_8 0 NS_329 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 331/332
CS_331 NS_331 0 9.9999999999999998e-13
CS_332 NS_332 0 9.9999999999999998e-13
RS_331 NS_331 0 5.4323743269805618e+02
RS_332 NS_332 0 5.4323743269805618e+02
GL_331 0 NS_331 NS_332 0 2.2057741537827197e-01
GL_332 0 NS_332 NS_331 0 -2.2057741537827197e-01
GS_331_8 0 NS_331 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 333/334
CS_333 NS_333 0 9.9999999999999998e-13
CS_334 NS_334 0 9.9999999999999998e-13
RS_333 NS_333 0 6.2013592102356057e+01
RS_334 NS_334 0 6.2013592102356057e+01
GL_333 0 NS_333 NS_334 0 2.2721975400227054e-01
GL_334 0 NS_334 NS_333 0 -2.2721975400227054e-01
GS_333_8 0 NS_333 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 335/336
CS_335 NS_335 0 9.9999999999999998e-13
CS_336 NS_336 0 9.9999999999999998e-13
RS_335 NS_335 0 8.2527539890421451e+01
RS_336 NS_336 0 8.2527539890421465e+01
GL_335 0 NS_335 NS_336 0 2.2544686857562196e-01
GL_336 0 NS_336 NS_335 0 -2.2544686857562196e-01
GS_335_8 0 NS_335 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 337/338
CS_337 NS_337 0 9.9999999999999998e-13
CS_338 NS_338 0 9.9999999999999998e-13
RS_337 NS_337 0 1.5057204740157513e+02
RS_338 NS_338 0 1.5057204740157516e+02
GL_337 0 NS_337 NS_338 0 2.5030962700427895e-01
GL_338 0 NS_338 NS_337 0 -2.5030962700427895e-01
GS_337_8 0 NS_337 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 339/340
CS_339 NS_339 0 9.9999999999999998e-13
CS_340 NS_340 0 9.9999999999999998e-13
RS_339 NS_339 0 1.0143406310664166e+03
RS_340 NS_340 0 1.0143406310664167e+03
GL_339 0 NS_339 NS_340 0 2.4802996115452441e-01
GL_340 0 NS_340 NS_339 0 -2.4802996115452441e-01
GS_339_8 0 NS_339 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 341/342
CS_341 NS_341 0 9.9999999999999998e-13
CS_342 NS_342 0 9.9999999999999998e-13
RS_341 NS_341 0 2.6049933264405115e+02
RS_342 NS_342 0 2.6049933264405115e+02
GL_341 0 NS_341 NS_342 0 2.4648481498152200e-01
GL_342 0 NS_342 NS_341 0 -2.4648481498152200e-01
GS_341_8 0 NS_341 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 343/344
CS_343 NS_343 0 9.9999999999999998e-13
CS_344 NS_344 0 9.9999999999999998e-13
RS_343 NS_343 0 8.6892684135916670e+02
RS_344 NS_344 0 8.6892684135916659e+02
GL_343 0 NS_343 NS_344 0 2.4352824357909131e-01
GL_344 0 NS_344 NS_343 0 -2.4352824357909131e-01
GS_343_8 0 NS_343 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 345/346
CS_345 NS_345 0 9.9999999999999998e-13
CS_346 NS_346 0 9.9999999999999998e-13
RS_345 NS_345 0 6.5240189890508168e+02
RS_346 NS_346 0 6.5240189890508168e+02
GL_345 0 NS_345 NS_346 0 2.3166276016037468e-01
GL_346 0 NS_346 NS_345 0 -2.3166276016037468e-01
GS_345_8 0 NS_345 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 347/348
CS_347 NS_347 0 9.9999999999999998e-13
CS_348 NS_348 0 9.9999999999999998e-13
RS_347 NS_347 0 1.8572469959933156e+02
RS_348 NS_348 0 1.8572469959933156e+02
GL_347 0 NS_347 NS_348 0 2.3351354491929543e-01
GL_348 0 NS_348 NS_347 0 -2.3351354491929543e-01
GS_347_8 0 NS_347 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 349/350
CS_349 NS_349 0 9.9999999999999998e-13
CS_350 NS_350 0 9.9999999999999998e-13
RS_349 NS_349 0 3.0631652744794525e+02
RS_350 NS_350 0 3.0631652744794530e+02
GL_349 0 NS_349 NS_350 0 2.3886925224886552e-01
GL_350 0 NS_350 NS_349 0 -2.3886925224886552e-01
GS_349_8 0 NS_349 NA_8 0 1.1283794739964070e+00
*
* Complex pair n. 351/352
CS_351 NS_351 0 9.9999999999999998e-13
CS_352 NS_352 0 9.9999999999999998e-13
RS_351 NS_351 0 5.0301469986378567e+02
RS_352 NS_352 0 5.0301469986378567e+02
GL_351 0 NS_351 NS_352 0 2.3692781195536661e-01
GL_352 0 NS_352 NS_351 0 -2.3692781195536661e-01
GS_351_8 0 NS_351 NA_8 0 1.1283794739964070e+00
*
* Real pole n. 353
CS_353 NS_353 0 9.9999999999999998e-13
RS_353 NS_353 0 3.9451851533158515e+00
GS_353_9 0 NS_353 NA_9 0 1.1283794739964070e+00
*
* Real pole n. 354
CS_354 NS_354 0 9.9999999999999998e-13
RS_354 NS_354 0 1.8805154767607480e+01
GS_354_9 0 NS_354 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 355/356
CS_355 NS_355 0 9.9999999999999998e-13
CS_356 NS_356 0 9.9999999999999998e-13
RS_355 NS_355 0 1.8483596483142442e+01
RS_356 NS_356 0 1.8483596483142442e+01
GL_355 0 NS_355 NS_356 0 6.9799982353381460e-02
GL_356 0 NS_356 NS_355 0 -6.9799982353381460e-02
GS_355_9 0 NS_355 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 357/358
CS_357 NS_357 0 9.9999999999999998e-13
CS_358 NS_358 0 9.9999999999999998e-13
RS_357 NS_357 0 1.9654872352993628e+01
RS_358 NS_358 0 1.9654872352993625e+01
GL_357 0 NS_357 NS_358 0 9.5720932954598423e-02
GL_358 0 NS_358 NS_357 0 -9.5720932954598423e-02
GS_357_9 0 NS_357 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 359/360
CS_359 NS_359 0 9.9999999999999998e-13
CS_360 NS_360 0 9.9999999999999998e-13
RS_359 NS_359 0 2.5061544329287912e+01
RS_360 NS_360 0 2.5061544329287909e+01
GL_359 0 NS_359 NS_360 0 1.3536754976539320e-01
GL_360 0 NS_360 NS_359 0 -1.3536754976539320e-01
GS_359_9 0 NS_359 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 361/362
CS_361 NS_361 0 9.9999999999999998e-13
CS_362 NS_362 0 9.9999999999999998e-13
RS_361 NS_361 0 7.4239654864745361e+01
RS_362 NS_362 0 7.4239654864745361e+01
GL_361 0 NS_361 NS_362 0 2.8245804011501385e-01
GL_362 0 NS_362 NS_361 0 -2.8245804011501385e-01
GS_361_9 0 NS_361 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 363/364
CS_363 NS_363 0 9.9999999999999998e-13
CS_364 NS_364 0 9.9999999999999998e-13
RS_363 NS_363 0 2.8726427419385509e+01
RS_364 NS_364 0 2.8726427419385512e+01
GL_363 0 NS_363 NS_364 0 1.7620265460857126e-01
GL_364 0 NS_364 NS_363 0 -1.7620265460857126e-01
GS_363_9 0 NS_363 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 365/366
CS_365 NS_365 0 9.9999999999999998e-13
CS_366 NS_366 0 9.9999999999999998e-13
RS_365 NS_365 0 7.8929016552352451e+01
RS_366 NS_366 0 7.8929016552352465e+01
GL_365 0 NS_365 NS_366 0 1.7267598155977268e-01
GL_366 0 NS_366 NS_365 0 -1.7267598155977268e-01
GS_365_9 0 NS_365 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 367/368
CS_367 NS_367 0 9.9999999999999998e-13
CS_368 NS_368 0 9.9999999999999998e-13
RS_367 NS_367 0 1.3876610711235463e+02
RS_368 NS_368 0 1.3876610711235463e+02
GL_367 0 NS_367 NS_368 0 1.9827389109149790e-01
GL_368 0 NS_368 NS_367 0 -1.9827389109149790e-01
GS_367_9 0 NS_367 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 369/370
CS_369 NS_369 0 9.9999999999999998e-13
CS_370 NS_370 0 9.9999999999999998e-13
RS_369 NS_369 0 9.4943847388790630e+01
RS_370 NS_370 0 9.4943847388790630e+01
GL_369 0 NS_369 NS_370 0 2.0370912057963636e-01
GL_370 0 NS_370 NS_369 0 -2.0370912057963636e-01
GS_369_9 0 NS_369 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 371/372
CS_371 NS_371 0 9.9999999999999998e-13
CS_372 NS_372 0 9.9999999999999998e-13
RS_371 NS_371 0 2.2502148823483816e+02
RS_372 NS_372 0 2.2502148823483816e+02
GL_371 0 NS_371 NS_372 0 2.1140622110318164e-01
GL_372 0 NS_372 NS_371 0 -2.1140622110318164e-01
GS_371_9 0 NS_371 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 373/374
CS_373 NS_373 0 9.9999999999999998e-13
CS_374 NS_374 0 9.9999999999999998e-13
RS_373 NS_373 0 2.0359721972446440e+02
RS_374 NS_374 0 2.0359721972446440e+02
GL_373 0 NS_373 NS_374 0 2.1650882528339854e-01
GL_374 0 NS_374 NS_373 0 -2.1650882528339854e-01
GS_373_9 0 NS_373 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 375/376
CS_375 NS_375 0 9.9999999999999998e-13
CS_376 NS_376 0 9.9999999999999998e-13
RS_375 NS_375 0 5.4323743269805618e+02
RS_376 NS_376 0 5.4323743269805618e+02
GL_375 0 NS_375 NS_376 0 2.2057741537827197e-01
GL_376 0 NS_376 NS_375 0 -2.2057741537827197e-01
GS_375_9 0 NS_375 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 377/378
CS_377 NS_377 0 9.9999999999999998e-13
CS_378 NS_378 0 9.9999999999999998e-13
RS_377 NS_377 0 6.2013592102356057e+01
RS_378 NS_378 0 6.2013592102356057e+01
GL_377 0 NS_377 NS_378 0 2.2721975400227054e-01
GL_378 0 NS_378 NS_377 0 -2.2721975400227054e-01
GS_377_9 0 NS_377 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 379/380
CS_379 NS_379 0 9.9999999999999998e-13
CS_380 NS_380 0 9.9999999999999998e-13
RS_379 NS_379 0 8.2527539890421451e+01
RS_380 NS_380 0 8.2527539890421465e+01
GL_379 0 NS_379 NS_380 0 2.2544686857562196e-01
GL_380 0 NS_380 NS_379 0 -2.2544686857562196e-01
GS_379_9 0 NS_379 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 381/382
CS_381 NS_381 0 9.9999999999999998e-13
CS_382 NS_382 0 9.9999999999999998e-13
RS_381 NS_381 0 1.5057204740157513e+02
RS_382 NS_382 0 1.5057204740157516e+02
GL_381 0 NS_381 NS_382 0 2.5030962700427895e-01
GL_382 0 NS_382 NS_381 0 -2.5030962700427895e-01
GS_381_9 0 NS_381 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 383/384
CS_383 NS_383 0 9.9999999999999998e-13
CS_384 NS_384 0 9.9999999999999998e-13
RS_383 NS_383 0 1.0143406310664166e+03
RS_384 NS_384 0 1.0143406310664167e+03
GL_383 0 NS_383 NS_384 0 2.4802996115452441e-01
GL_384 0 NS_384 NS_383 0 -2.4802996115452441e-01
GS_383_9 0 NS_383 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 385/386
CS_385 NS_385 0 9.9999999999999998e-13
CS_386 NS_386 0 9.9999999999999998e-13
RS_385 NS_385 0 2.6049933264405115e+02
RS_386 NS_386 0 2.6049933264405115e+02
GL_385 0 NS_385 NS_386 0 2.4648481498152200e-01
GL_386 0 NS_386 NS_385 0 -2.4648481498152200e-01
GS_385_9 0 NS_385 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 387/388
CS_387 NS_387 0 9.9999999999999998e-13
CS_388 NS_388 0 9.9999999999999998e-13
RS_387 NS_387 0 8.6892684135916670e+02
RS_388 NS_388 0 8.6892684135916659e+02
GL_387 0 NS_387 NS_388 0 2.4352824357909131e-01
GL_388 0 NS_388 NS_387 0 -2.4352824357909131e-01
GS_387_9 0 NS_387 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 389/390
CS_389 NS_389 0 9.9999999999999998e-13
CS_390 NS_390 0 9.9999999999999998e-13
RS_389 NS_389 0 6.5240189890508168e+02
RS_390 NS_390 0 6.5240189890508168e+02
GL_389 0 NS_389 NS_390 0 2.3166276016037468e-01
GL_390 0 NS_390 NS_389 0 -2.3166276016037468e-01
GS_389_9 0 NS_389 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 391/392
CS_391 NS_391 0 9.9999999999999998e-13
CS_392 NS_392 0 9.9999999999999998e-13
RS_391 NS_391 0 1.8572469959933156e+02
RS_392 NS_392 0 1.8572469959933156e+02
GL_391 0 NS_391 NS_392 0 2.3351354491929543e-01
GL_392 0 NS_392 NS_391 0 -2.3351354491929543e-01
GS_391_9 0 NS_391 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 393/394
CS_393 NS_393 0 9.9999999999999998e-13
CS_394 NS_394 0 9.9999999999999998e-13
RS_393 NS_393 0 3.0631652744794525e+02
RS_394 NS_394 0 3.0631652744794530e+02
GL_393 0 NS_393 NS_394 0 2.3886925224886552e-01
GL_394 0 NS_394 NS_393 0 -2.3886925224886552e-01
GS_393_9 0 NS_393 NA_9 0 1.1283794739964070e+00
*
* Complex pair n. 395/396
CS_395 NS_395 0 9.9999999999999998e-13
CS_396 NS_396 0 9.9999999999999998e-13
RS_395 NS_395 0 5.0301469986378567e+02
RS_396 NS_396 0 5.0301469986378567e+02
GL_395 0 NS_395 NS_396 0 2.3692781195536661e-01
GL_396 0 NS_396 NS_395 0 -2.3692781195536661e-01
GS_395_9 0 NS_395 NA_9 0 1.1283794739964070e+00
*
* Real pole n. 397
CS_397 NS_397 0 9.9999999999999998e-13
RS_397 NS_397 0 3.9451851533158515e+00
GS_397_10 0 NS_397 NA_10 0 1.1283794739964070e+00
*
* Real pole n. 398
CS_398 NS_398 0 9.9999999999999998e-13
RS_398 NS_398 0 1.8805154767607480e+01
GS_398_10 0 NS_398 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 399/400
CS_399 NS_399 0 9.9999999999999998e-13
CS_400 NS_400 0 9.9999999999999998e-13
RS_399 NS_399 0 1.8483596483142442e+01
RS_400 NS_400 0 1.8483596483142442e+01
GL_399 0 NS_399 NS_400 0 6.9799982353381460e-02
GL_400 0 NS_400 NS_399 0 -6.9799982353381460e-02
GS_399_10 0 NS_399 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 401/402
CS_401 NS_401 0 9.9999999999999998e-13
CS_402 NS_402 0 9.9999999999999998e-13
RS_401 NS_401 0 1.9654872352993628e+01
RS_402 NS_402 0 1.9654872352993625e+01
GL_401 0 NS_401 NS_402 0 9.5720932954598423e-02
GL_402 0 NS_402 NS_401 0 -9.5720932954598423e-02
GS_401_10 0 NS_401 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 403/404
CS_403 NS_403 0 9.9999999999999998e-13
CS_404 NS_404 0 9.9999999999999998e-13
RS_403 NS_403 0 2.5061544329287912e+01
RS_404 NS_404 0 2.5061544329287909e+01
GL_403 0 NS_403 NS_404 0 1.3536754976539320e-01
GL_404 0 NS_404 NS_403 0 -1.3536754976539320e-01
GS_403_10 0 NS_403 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 405/406
CS_405 NS_405 0 9.9999999999999998e-13
CS_406 NS_406 0 9.9999999999999998e-13
RS_405 NS_405 0 7.4239654864745361e+01
RS_406 NS_406 0 7.4239654864745361e+01
GL_405 0 NS_405 NS_406 0 2.8245804011501385e-01
GL_406 0 NS_406 NS_405 0 -2.8245804011501385e-01
GS_405_10 0 NS_405 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 407/408
CS_407 NS_407 0 9.9999999999999998e-13
CS_408 NS_408 0 9.9999999999999998e-13
RS_407 NS_407 0 2.8726427419385509e+01
RS_408 NS_408 0 2.8726427419385512e+01
GL_407 0 NS_407 NS_408 0 1.7620265460857126e-01
GL_408 0 NS_408 NS_407 0 -1.7620265460857126e-01
GS_407_10 0 NS_407 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 409/410
CS_409 NS_409 0 9.9999999999999998e-13
CS_410 NS_410 0 9.9999999999999998e-13
RS_409 NS_409 0 7.8929016552352451e+01
RS_410 NS_410 0 7.8929016552352465e+01
GL_409 0 NS_409 NS_410 0 1.7267598155977268e-01
GL_410 0 NS_410 NS_409 0 -1.7267598155977268e-01
GS_409_10 0 NS_409 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 411/412
CS_411 NS_411 0 9.9999999999999998e-13
CS_412 NS_412 0 9.9999999999999998e-13
RS_411 NS_411 0 1.3876610711235463e+02
RS_412 NS_412 0 1.3876610711235463e+02
GL_411 0 NS_411 NS_412 0 1.9827389109149790e-01
GL_412 0 NS_412 NS_411 0 -1.9827389109149790e-01
GS_411_10 0 NS_411 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 413/414
CS_413 NS_413 0 9.9999999999999998e-13
CS_414 NS_414 0 9.9999999999999998e-13
RS_413 NS_413 0 9.4943847388790630e+01
RS_414 NS_414 0 9.4943847388790630e+01
GL_413 0 NS_413 NS_414 0 2.0370912057963636e-01
GL_414 0 NS_414 NS_413 0 -2.0370912057963636e-01
GS_413_10 0 NS_413 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 415/416
CS_415 NS_415 0 9.9999999999999998e-13
CS_416 NS_416 0 9.9999999999999998e-13
RS_415 NS_415 0 2.2502148823483816e+02
RS_416 NS_416 0 2.2502148823483816e+02
GL_415 0 NS_415 NS_416 0 2.1140622110318164e-01
GL_416 0 NS_416 NS_415 0 -2.1140622110318164e-01
GS_415_10 0 NS_415 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 417/418
CS_417 NS_417 0 9.9999999999999998e-13
CS_418 NS_418 0 9.9999999999999998e-13
RS_417 NS_417 0 2.0359721972446440e+02
RS_418 NS_418 0 2.0359721972446440e+02
GL_417 0 NS_417 NS_418 0 2.1650882528339854e-01
GL_418 0 NS_418 NS_417 0 -2.1650882528339854e-01
GS_417_10 0 NS_417 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 419/420
CS_419 NS_419 0 9.9999999999999998e-13
CS_420 NS_420 0 9.9999999999999998e-13
RS_419 NS_419 0 5.4323743269805618e+02
RS_420 NS_420 0 5.4323743269805618e+02
GL_419 0 NS_419 NS_420 0 2.2057741537827197e-01
GL_420 0 NS_420 NS_419 0 -2.2057741537827197e-01
GS_419_10 0 NS_419 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 421/422
CS_421 NS_421 0 9.9999999999999998e-13
CS_422 NS_422 0 9.9999999999999998e-13
RS_421 NS_421 0 6.2013592102356057e+01
RS_422 NS_422 0 6.2013592102356057e+01
GL_421 0 NS_421 NS_422 0 2.2721975400227054e-01
GL_422 0 NS_422 NS_421 0 -2.2721975400227054e-01
GS_421_10 0 NS_421 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 423/424
CS_423 NS_423 0 9.9999999999999998e-13
CS_424 NS_424 0 9.9999999999999998e-13
RS_423 NS_423 0 8.2527539890421451e+01
RS_424 NS_424 0 8.2527539890421465e+01
GL_423 0 NS_423 NS_424 0 2.2544686857562196e-01
GL_424 0 NS_424 NS_423 0 -2.2544686857562196e-01
GS_423_10 0 NS_423 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 425/426
CS_425 NS_425 0 9.9999999999999998e-13
CS_426 NS_426 0 9.9999999999999998e-13
RS_425 NS_425 0 1.5057204740157513e+02
RS_426 NS_426 0 1.5057204740157516e+02
GL_425 0 NS_425 NS_426 0 2.5030962700427895e-01
GL_426 0 NS_426 NS_425 0 -2.5030962700427895e-01
GS_425_10 0 NS_425 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 427/428
CS_427 NS_427 0 9.9999999999999998e-13
CS_428 NS_428 0 9.9999999999999998e-13
RS_427 NS_427 0 1.0143406310664166e+03
RS_428 NS_428 0 1.0143406310664167e+03
GL_427 0 NS_427 NS_428 0 2.4802996115452441e-01
GL_428 0 NS_428 NS_427 0 -2.4802996115452441e-01
GS_427_10 0 NS_427 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 429/430
CS_429 NS_429 0 9.9999999999999998e-13
CS_430 NS_430 0 9.9999999999999998e-13
RS_429 NS_429 0 2.6049933264405115e+02
RS_430 NS_430 0 2.6049933264405115e+02
GL_429 0 NS_429 NS_430 0 2.4648481498152200e-01
GL_430 0 NS_430 NS_429 0 -2.4648481498152200e-01
GS_429_10 0 NS_429 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 431/432
CS_431 NS_431 0 9.9999999999999998e-13
CS_432 NS_432 0 9.9999999999999998e-13
RS_431 NS_431 0 8.6892684135916670e+02
RS_432 NS_432 0 8.6892684135916659e+02
GL_431 0 NS_431 NS_432 0 2.4352824357909131e-01
GL_432 0 NS_432 NS_431 0 -2.4352824357909131e-01
GS_431_10 0 NS_431 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 433/434
CS_433 NS_433 0 9.9999999999999998e-13
CS_434 NS_434 0 9.9999999999999998e-13
RS_433 NS_433 0 6.5240189890508168e+02
RS_434 NS_434 0 6.5240189890508168e+02
GL_433 0 NS_433 NS_434 0 2.3166276016037468e-01
GL_434 0 NS_434 NS_433 0 -2.3166276016037468e-01
GS_433_10 0 NS_433 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 435/436
CS_435 NS_435 0 9.9999999999999998e-13
CS_436 NS_436 0 9.9999999999999998e-13
RS_435 NS_435 0 1.8572469959933156e+02
RS_436 NS_436 0 1.8572469959933156e+02
GL_435 0 NS_435 NS_436 0 2.3351354491929543e-01
GL_436 0 NS_436 NS_435 0 -2.3351354491929543e-01
GS_435_10 0 NS_435 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 437/438
CS_437 NS_437 0 9.9999999999999998e-13
CS_438 NS_438 0 9.9999999999999998e-13
RS_437 NS_437 0 3.0631652744794525e+02
RS_438 NS_438 0 3.0631652744794530e+02
GL_437 0 NS_437 NS_438 0 2.3886925224886552e-01
GL_438 0 NS_438 NS_437 0 -2.3886925224886552e-01
GS_437_10 0 NS_437 NA_10 0 1.1283794739964070e+00
*
* Complex pair n. 439/440
CS_439 NS_439 0 9.9999999999999998e-13
CS_440 NS_440 0 9.9999999999999998e-13
RS_439 NS_439 0 5.0301469986378567e+02
RS_440 NS_440 0 5.0301469986378567e+02
GL_439 0 NS_439 NS_440 0 2.3692781195536661e-01
GL_440 0 NS_440 NS_439 0 -2.3692781195536661e-01
GS_439_10 0 NS_439 NA_10 0 1.1283794739964070e+00
*
* Real pole n. 441
CS_441 NS_441 0 9.9999999999999998e-13
RS_441 NS_441 0 3.9451851533158515e+00
GS_441_11 0 NS_441 NA_11 0 1.1283794739964070e+00
*
* Real pole n. 442
CS_442 NS_442 0 9.9999999999999998e-13
RS_442 NS_442 0 1.8805154767607480e+01
GS_442_11 0 NS_442 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 443/444
CS_443 NS_443 0 9.9999999999999998e-13
CS_444 NS_444 0 9.9999999999999998e-13
RS_443 NS_443 0 1.8483596483142442e+01
RS_444 NS_444 0 1.8483596483142442e+01
GL_443 0 NS_443 NS_444 0 6.9799982353381460e-02
GL_444 0 NS_444 NS_443 0 -6.9799982353381460e-02
GS_443_11 0 NS_443 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 445/446
CS_445 NS_445 0 9.9999999999999998e-13
CS_446 NS_446 0 9.9999999999999998e-13
RS_445 NS_445 0 1.9654872352993628e+01
RS_446 NS_446 0 1.9654872352993625e+01
GL_445 0 NS_445 NS_446 0 9.5720932954598423e-02
GL_446 0 NS_446 NS_445 0 -9.5720932954598423e-02
GS_445_11 0 NS_445 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 447/448
CS_447 NS_447 0 9.9999999999999998e-13
CS_448 NS_448 0 9.9999999999999998e-13
RS_447 NS_447 0 2.5061544329287912e+01
RS_448 NS_448 0 2.5061544329287909e+01
GL_447 0 NS_447 NS_448 0 1.3536754976539320e-01
GL_448 0 NS_448 NS_447 0 -1.3536754976539320e-01
GS_447_11 0 NS_447 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 449/450
CS_449 NS_449 0 9.9999999999999998e-13
CS_450 NS_450 0 9.9999999999999998e-13
RS_449 NS_449 0 7.4239654864745361e+01
RS_450 NS_450 0 7.4239654864745361e+01
GL_449 0 NS_449 NS_450 0 2.8245804011501385e-01
GL_450 0 NS_450 NS_449 0 -2.8245804011501385e-01
GS_449_11 0 NS_449 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 451/452
CS_451 NS_451 0 9.9999999999999998e-13
CS_452 NS_452 0 9.9999999999999998e-13
RS_451 NS_451 0 2.8726427419385509e+01
RS_452 NS_452 0 2.8726427419385512e+01
GL_451 0 NS_451 NS_452 0 1.7620265460857126e-01
GL_452 0 NS_452 NS_451 0 -1.7620265460857126e-01
GS_451_11 0 NS_451 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 453/454
CS_453 NS_453 0 9.9999999999999998e-13
CS_454 NS_454 0 9.9999999999999998e-13
RS_453 NS_453 0 7.8929016552352451e+01
RS_454 NS_454 0 7.8929016552352465e+01
GL_453 0 NS_453 NS_454 0 1.7267598155977268e-01
GL_454 0 NS_454 NS_453 0 -1.7267598155977268e-01
GS_453_11 0 NS_453 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 455/456
CS_455 NS_455 0 9.9999999999999998e-13
CS_456 NS_456 0 9.9999999999999998e-13
RS_455 NS_455 0 1.3876610711235463e+02
RS_456 NS_456 0 1.3876610711235463e+02
GL_455 0 NS_455 NS_456 0 1.9827389109149790e-01
GL_456 0 NS_456 NS_455 0 -1.9827389109149790e-01
GS_455_11 0 NS_455 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 457/458
CS_457 NS_457 0 9.9999999999999998e-13
CS_458 NS_458 0 9.9999999999999998e-13
RS_457 NS_457 0 9.4943847388790630e+01
RS_458 NS_458 0 9.4943847388790630e+01
GL_457 0 NS_457 NS_458 0 2.0370912057963636e-01
GL_458 0 NS_458 NS_457 0 -2.0370912057963636e-01
GS_457_11 0 NS_457 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 459/460
CS_459 NS_459 0 9.9999999999999998e-13
CS_460 NS_460 0 9.9999999999999998e-13
RS_459 NS_459 0 2.2502148823483816e+02
RS_460 NS_460 0 2.2502148823483816e+02
GL_459 0 NS_459 NS_460 0 2.1140622110318164e-01
GL_460 0 NS_460 NS_459 0 -2.1140622110318164e-01
GS_459_11 0 NS_459 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 461/462
CS_461 NS_461 0 9.9999999999999998e-13
CS_462 NS_462 0 9.9999999999999998e-13
RS_461 NS_461 0 2.0359721972446440e+02
RS_462 NS_462 0 2.0359721972446440e+02
GL_461 0 NS_461 NS_462 0 2.1650882528339854e-01
GL_462 0 NS_462 NS_461 0 -2.1650882528339854e-01
GS_461_11 0 NS_461 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 463/464
CS_463 NS_463 0 9.9999999999999998e-13
CS_464 NS_464 0 9.9999999999999998e-13
RS_463 NS_463 0 5.4323743269805618e+02
RS_464 NS_464 0 5.4323743269805618e+02
GL_463 0 NS_463 NS_464 0 2.2057741537827197e-01
GL_464 0 NS_464 NS_463 0 -2.2057741537827197e-01
GS_463_11 0 NS_463 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 465/466
CS_465 NS_465 0 9.9999999999999998e-13
CS_466 NS_466 0 9.9999999999999998e-13
RS_465 NS_465 0 6.2013592102356057e+01
RS_466 NS_466 0 6.2013592102356057e+01
GL_465 0 NS_465 NS_466 0 2.2721975400227054e-01
GL_466 0 NS_466 NS_465 0 -2.2721975400227054e-01
GS_465_11 0 NS_465 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 467/468
CS_467 NS_467 0 9.9999999999999998e-13
CS_468 NS_468 0 9.9999999999999998e-13
RS_467 NS_467 0 8.2527539890421451e+01
RS_468 NS_468 0 8.2527539890421465e+01
GL_467 0 NS_467 NS_468 0 2.2544686857562196e-01
GL_468 0 NS_468 NS_467 0 -2.2544686857562196e-01
GS_467_11 0 NS_467 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 469/470
CS_469 NS_469 0 9.9999999999999998e-13
CS_470 NS_470 0 9.9999999999999998e-13
RS_469 NS_469 0 1.5057204740157513e+02
RS_470 NS_470 0 1.5057204740157516e+02
GL_469 0 NS_469 NS_470 0 2.5030962700427895e-01
GL_470 0 NS_470 NS_469 0 -2.5030962700427895e-01
GS_469_11 0 NS_469 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 471/472
CS_471 NS_471 0 9.9999999999999998e-13
CS_472 NS_472 0 9.9999999999999998e-13
RS_471 NS_471 0 1.0143406310664166e+03
RS_472 NS_472 0 1.0143406310664167e+03
GL_471 0 NS_471 NS_472 0 2.4802996115452441e-01
GL_472 0 NS_472 NS_471 0 -2.4802996115452441e-01
GS_471_11 0 NS_471 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 473/474
CS_473 NS_473 0 9.9999999999999998e-13
CS_474 NS_474 0 9.9999999999999998e-13
RS_473 NS_473 0 2.6049933264405115e+02
RS_474 NS_474 0 2.6049933264405115e+02
GL_473 0 NS_473 NS_474 0 2.4648481498152200e-01
GL_474 0 NS_474 NS_473 0 -2.4648481498152200e-01
GS_473_11 0 NS_473 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 475/476
CS_475 NS_475 0 9.9999999999999998e-13
CS_476 NS_476 0 9.9999999999999998e-13
RS_475 NS_475 0 8.6892684135916670e+02
RS_476 NS_476 0 8.6892684135916659e+02
GL_475 0 NS_475 NS_476 0 2.4352824357909131e-01
GL_476 0 NS_476 NS_475 0 -2.4352824357909131e-01
GS_475_11 0 NS_475 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 477/478
CS_477 NS_477 0 9.9999999999999998e-13
CS_478 NS_478 0 9.9999999999999998e-13
RS_477 NS_477 0 6.5240189890508168e+02
RS_478 NS_478 0 6.5240189890508168e+02
GL_477 0 NS_477 NS_478 0 2.3166276016037468e-01
GL_478 0 NS_478 NS_477 0 -2.3166276016037468e-01
GS_477_11 0 NS_477 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 479/480
CS_479 NS_479 0 9.9999999999999998e-13
CS_480 NS_480 0 9.9999999999999998e-13
RS_479 NS_479 0 1.8572469959933156e+02
RS_480 NS_480 0 1.8572469959933156e+02
GL_479 0 NS_479 NS_480 0 2.3351354491929543e-01
GL_480 0 NS_480 NS_479 0 -2.3351354491929543e-01
GS_479_11 0 NS_479 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 481/482
CS_481 NS_481 0 9.9999999999999998e-13
CS_482 NS_482 0 9.9999999999999998e-13
RS_481 NS_481 0 3.0631652744794525e+02
RS_482 NS_482 0 3.0631652744794530e+02
GL_481 0 NS_481 NS_482 0 2.3886925224886552e-01
GL_482 0 NS_482 NS_481 0 -2.3886925224886552e-01
GS_481_11 0 NS_481 NA_11 0 1.1283794739964070e+00
*
* Complex pair n. 483/484
CS_483 NS_483 0 9.9999999999999998e-13
CS_484 NS_484 0 9.9999999999999998e-13
RS_483 NS_483 0 5.0301469986378567e+02
RS_484 NS_484 0 5.0301469986378567e+02
GL_483 0 NS_483 NS_484 0 2.3692781195536661e-01
GL_484 0 NS_484 NS_483 0 -2.3692781195536661e-01
GS_483_11 0 NS_483 NA_11 0 1.1283794739964070e+00
*
* Real pole n. 485
CS_485 NS_485 0 9.9999999999999998e-13
RS_485 NS_485 0 3.9451851533158515e+00
GS_485_12 0 NS_485 NA_12 0 1.1283794739964070e+00
*
* Real pole n. 486
CS_486 NS_486 0 9.9999999999999998e-13
RS_486 NS_486 0 1.8805154767607480e+01
GS_486_12 0 NS_486 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 487/488
CS_487 NS_487 0 9.9999999999999998e-13
CS_488 NS_488 0 9.9999999999999998e-13
RS_487 NS_487 0 1.8483596483142442e+01
RS_488 NS_488 0 1.8483596483142442e+01
GL_487 0 NS_487 NS_488 0 6.9799982353381460e-02
GL_488 0 NS_488 NS_487 0 -6.9799982353381460e-02
GS_487_12 0 NS_487 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 489/490
CS_489 NS_489 0 9.9999999999999998e-13
CS_490 NS_490 0 9.9999999999999998e-13
RS_489 NS_489 0 1.9654872352993628e+01
RS_490 NS_490 0 1.9654872352993625e+01
GL_489 0 NS_489 NS_490 0 9.5720932954598423e-02
GL_490 0 NS_490 NS_489 0 -9.5720932954598423e-02
GS_489_12 0 NS_489 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 491/492
CS_491 NS_491 0 9.9999999999999998e-13
CS_492 NS_492 0 9.9999999999999998e-13
RS_491 NS_491 0 2.5061544329287912e+01
RS_492 NS_492 0 2.5061544329287909e+01
GL_491 0 NS_491 NS_492 0 1.3536754976539320e-01
GL_492 0 NS_492 NS_491 0 -1.3536754976539320e-01
GS_491_12 0 NS_491 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 493/494
CS_493 NS_493 0 9.9999999999999998e-13
CS_494 NS_494 0 9.9999999999999998e-13
RS_493 NS_493 0 7.4239654864745361e+01
RS_494 NS_494 0 7.4239654864745361e+01
GL_493 0 NS_493 NS_494 0 2.8245804011501385e-01
GL_494 0 NS_494 NS_493 0 -2.8245804011501385e-01
GS_493_12 0 NS_493 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 495/496
CS_495 NS_495 0 9.9999999999999998e-13
CS_496 NS_496 0 9.9999999999999998e-13
RS_495 NS_495 0 2.8726427419385509e+01
RS_496 NS_496 0 2.8726427419385512e+01
GL_495 0 NS_495 NS_496 0 1.7620265460857126e-01
GL_496 0 NS_496 NS_495 0 -1.7620265460857126e-01
GS_495_12 0 NS_495 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 497/498
CS_497 NS_497 0 9.9999999999999998e-13
CS_498 NS_498 0 9.9999999999999998e-13
RS_497 NS_497 0 7.8929016552352451e+01
RS_498 NS_498 0 7.8929016552352465e+01
GL_497 0 NS_497 NS_498 0 1.7267598155977268e-01
GL_498 0 NS_498 NS_497 0 -1.7267598155977268e-01
GS_497_12 0 NS_497 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 499/500
CS_499 NS_499 0 9.9999999999999998e-13
CS_500 NS_500 0 9.9999999999999998e-13
RS_499 NS_499 0 1.3876610711235463e+02
RS_500 NS_500 0 1.3876610711235463e+02
GL_499 0 NS_499 NS_500 0 1.9827389109149790e-01
GL_500 0 NS_500 NS_499 0 -1.9827389109149790e-01
GS_499_12 0 NS_499 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 501/502
CS_501 NS_501 0 9.9999999999999998e-13
CS_502 NS_502 0 9.9999999999999998e-13
RS_501 NS_501 0 9.4943847388790630e+01
RS_502 NS_502 0 9.4943847388790630e+01
GL_501 0 NS_501 NS_502 0 2.0370912057963636e-01
GL_502 0 NS_502 NS_501 0 -2.0370912057963636e-01
GS_501_12 0 NS_501 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 503/504
CS_503 NS_503 0 9.9999999999999998e-13
CS_504 NS_504 0 9.9999999999999998e-13
RS_503 NS_503 0 2.2502148823483816e+02
RS_504 NS_504 0 2.2502148823483816e+02
GL_503 0 NS_503 NS_504 0 2.1140622110318164e-01
GL_504 0 NS_504 NS_503 0 -2.1140622110318164e-01
GS_503_12 0 NS_503 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 505/506
CS_505 NS_505 0 9.9999999999999998e-13
CS_506 NS_506 0 9.9999999999999998e-13
RS_505 NS_505 0 2.0359721972446440e+02
RS_506 NS_506 0 2.0359721972446440e+02
GL_505 0 NS_505 NS_506 0 2.1650882528339854e-01
GL_506 0 NS_506 NS_505 0 -2.1650882528339854e-01
GS_505_12 0 NS_505 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 507/508
CS_507 NS_507 0 9.9999999999999998e-13
CS_508 NS_508 0 9.9999999999999998e-13
RS_507 NS_507 0 5.4323743269805618e+02
RS_508 NS_508 0 5.4323743269805618e+02
GL_507 0 NS_507 NS_508 0 2.2057741537827197e-01
GL_508 0 NS_508 NS_507 0 -2.2057741537827197e-01
GS_507_12 0 NS_507 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 509/510
CS_509 NS_509 0 9.9999999999999998e-13
CS_510 NS_510 0 9.9999999999999998e-13
RS_509 NS_509 0 6.2013592102356057e+01
RS_510 NS_510 0 6.2013592102356057e+01
GL_509 0 NS_509 NS_510 0 2.2721975400227054e-01
GL_510 0 NS_510 NS_509 0 -2.2721975400227054e-01
GS_509_12 0 NS_509 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 511/512
CS_511 NS_511 0 9.9999999999999998e-13
CS_512 NS_512 0 9.9999999999999998e-13
RS_511 NS_511 0 8.2527539890421451e+01
RS_512 NS_512 0 8.2527539890421465e+01
GL_511 0 NS_511 NS_512 0 2.2544686857562196e-01
GL_512 0 NS_512 NS_511 0 -2.2544686857562196e-01
GS_511_12 0 NS_511 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 513/514
CS_513 NS_513 0 9.9999999999999998e-13
CS_514 NS_514 0 9.9999999999999998e-13
RS_513 NS_513 0 1.5057204740157513e+02
RS_514 NS_514 0 1.5057204740157516e+02
GL_513 0 NS_513 NS_514 0 2.5030962700427895e-01
GL_514 0 NS_514 NS_513 0 -2.5030962700427895e-01
GS_513_12 0 NS_513 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 515/516
CS_515 NS_515 0 9.9999999999999998e-13
CS_516 NS_516 0 9.9999999999999998e-13
RS_515 NS_515 0 1.0143406310664166e+03
RS_516 NS_516 0 1.0143406310664167e+03
GL_515 0 NS_515 NS_516 0 2.4802996115452441e-01
GL_516 0 NS_516 NS_515 0 -2.4802996115452441e-01
GS_515_12 0 NS_515 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 517/518
CS_517 NS_517 0 9.9999999999999998e-13
CS_518 NS_518 0 9.9999999999999998e-13
RS_517 NS_517 0 2.6049933264405115e+02
RS_518 NS_518 0 2.6049933264405115e+02
GL_517 0 NS_517 NS_518 0 2.4648481498152200e-01
GL_518 0 NS_518 NS_517 0 -2.4648481498152200e-01
GS_517_12 0 NS_517 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 519/520
CS_519 NS_519 0 9.9999999999999998e-13
CS_520 NS_520 0 9.9999999999999998e-13
RS_519 NS_519 0 8.6892684135916670e+02
RS_520 NS_520 0 8.6892684135916659e+02
GL_519 0 NS_519 NS_520 0 2.4352824357909131e-01
GL_520 0 NS_520 NS_519 0 -2.4352824357909131e-01
GS_519_12 0 NS_519 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 521/522
CS_521 NS_521 0 9.9999999999999998e-13
CS_522 NS_522 0 9.9999999999999998e-13
RS_521 NS_521 0 6.5240189890508168e+02
RS_522 NS_522 0 6.5240189890508168e+02
GL_521 0 NS_521 NS_522 0 2.3166276016037468e-01
GL_522 0 NS_522 NS_521 0 -2.3166276016037468e-01
GS_521_12 0 NS_521 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 523/524
CS_523 NS_523 0 9.9999999999999998e-13
CS_524 NS_524 0 9.9999999999999998e-13
RS_523 NS_523 0 1.8572469959933156e+02
RS_524 NS_524 0 1.8572469959933156e+02
GL_523 0 NS_523 NS_524 0 2.3351354491929543e-01
GL_524 0 NS_524 NS_523 0 -2.3351354491929543e-01
GS_523_12 0 NS_523 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 525/526
CS_525 NS_525 0 9.9999999999999998e-13
CS_526 NS_526 0 9.9999999999999998e-13
RS_525 NS_525 0 3.0631652744794525e+02
RS_526 NS_526 0 3.0631652744794530e+02
GL_525 0 NS_525 NS_526 0 2.3886925224886552e-01
GL_526 0 NS_526 NS_525 0 -2.3886925224886552e-01
GS_525_12 0 NS_525 NA_12 0 1.1283794739964070e+00
*
* Complex pair n. 527/528
CS_527 NS_527 0 9.9999999999999998e-13
CS_528 NS_528 0 9.9999999999999998e-13
RS_527 NS_527 0 5.0301469986378567e+02
RS_528 NS_528 0 5.0301469986378567e+02
GL_527 0 NS_527 NS_528 0 2.3692781195536661e-01
GL_528 0 NS_528 NS_527 0 -2.3692781195536661e-01
GS_527_12 0 NS_527 NA_12 0 1.1283794739964070e+00
*
******************************


.ends
*******************
* End of subcircuit
*******************
