**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 15-Feb-2023 by IdEM MP 12 (12.3.0)
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 4.0000e+10 Hz
** Order: [8 4 42] 
** SplitType: none 
** tol: 1.0000e-04 
** Weights: relative 
**    Alpha: 0.5
**    RelThreshold: 1e-06
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Data based
** Weights: relative
**    Alpha: 0.5
**    Relative threshold: 1e-06
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: separate (floating)
** Resistor synthesis: standard
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt subckt_1_BoardVia_backdrill
+  a_1 b_1
+  a_2 b_2
+  a_3 b_3
+  a_4 b_4
+  a_5 b_5
+  a_6 b_6
+  a_7 b_7
+  a_8 b_8
+  a_9 b_9
+  a_10 b_10
+  a_11 b_11
+  a_12 b_12
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+01
GC_1_1 b_1 NI_1 NS_1 0 -7.1969660995340398e-02
GC_1_2 b_1 NI_1 NS_2 0 9.5312628270231969e-03
GC_1_3 b_1 NI_1 NS_3 0 3.2250982195424203e-03
GC_1_4 b_1 NI_1 NS_4 0 6.2763081918353137e-03
GC_1_5 b_1 NI_1 NS_5 0 1.1246624936333971e-02
GC_1_6 b_1 NI_1 NS_6 0 -2.3693677175052053e-03
GC_1_7 b_1 NI_1 NS_7 0 1.1394212751562342e-03
GC_1_8 b_1 NI_1 NS_8 0 1.0197078746025114e-03
GC_1_9 b_1 NI_1 NS_9 0 4.2462360838533322e-04
GC_1_10 b_1 NI_1 NS_10 0 3.3292872122667812e-03
GC_1_11 b_1 NI_1 NS_11 0 3.3728878823981643e-03
GC_1_12 b_1 NI_1 NS_12 0 2.3655016827033642e-03
GC_1_13 b_1 NI_1 NS_13 0 5.0394906765831304e-04
GC_1_14 b_1 NI_1 NS_14 0 3.3428139556481009e-04
GC_1_15 b_1 NI_1 NS_15 0 4.7678607552763992e-03
GC_1_16 b_1 NI_1 NS_16 0 8.4549757278073610e-04
GC_1_17 b_1 NI_1 NS_17 0 -6.1335695525057912e-05
GC_1_18 b_1 NI_1 NS_18 0 1.2680551275062789e-04
GC_1_19 b_1 NI_1 NS_19 0 -1.7615567362194002e-04
GC_1_20 b_1 NI_1 NS_20 0 -1.4766092863784527e-03
GC_1_21 b_1 NI_1 NS_21 0 -1.1202662682435437e-03
GC_1_22 b_1 NI_1 NS_22 0 1.2447359492185860e-04
GC_1_23 b_1 NI_1 NS_23 0 1.5680561618548750e-04
GC_1_24 b_1 NI_1 NS_24 0 3.6310398802851822e-05
GC_1_25 b_1 NI_1 NS_25 0 5.7419160365947403e-05
GC_1_26 b_1 NI_1 NS_26 0 -8.8452644571021665e-05
GC_1_27 b_1 NI_1 NS_27 0 3.9879753238560873e-03
GC_1_28 b_1 NI_1 NS_28 0 1.3979555693077435e-02
GC_1_29 b_1 NI_1 NS_29 0 -9.9542720660413994e-06
GC_1_30 b_1 NI_1 NS_30 0 -2.3722553064329456e-05
GC_1_31 b_1 NI_1 NS_31 0 3.4976243030679188e-03
GC_1_32 b_1 NI_1 NS_32 0 -4.5619812781798772e-03
GC_1_33 b_1 NI_1 NS_33 0 4.3171973477329331e-06
GC_1_34 b_1 NI_1 NS_34 0 -2.6821184099461346e-05
GC_1_35 b_1 NI_1 NS_35 0 -2.5734512650576304e-03
GC_1_36 b_1 NI_1 NS_36 0 1.1700663539822489e-03
GC_1_37 b_1 NI_1 NS_37 0 2.7196313482785237e-05
GC_1_38 b_1 NI_1 NS_38 0 3.7092155904566583e-05
GC_1_39 b_1 NI_1 NS_39 0 -7.1041285663088731e-06
GC_1_40 b_1 NI_1 NS_40 0 5.4001318526767396e-06
GC_1_41 b_1 NI_1 NS_41 0 -2.1228074839564005e-06
GC_1_42 b_1 NI_1 NS_42 0 -1.3826419507325876e-05
GC_1_43 b_1 NI_1 NS_43 0 -3.9169331785920795e-04
GC_1_44 b_1 NI_1 NS_44 0 -4.7958591843307189e-05
GC_1_45 b_1 NI_1 NS_45 0 1.4058402996183497e-03
GC_1_46 b_1 NI_1 NS_46 0 1.0834322596834561e-02
GC_1_47 b_1 NI_1 NS_47 0 -6.4869261954459845e-03
GC_1_48 b_1 NI_1 NS_48 0 -5.6190407803363221e-03
GC_1_49 b_1 NI_1 NS_49 0 -1.0866853919043729e-02
GC_1_50 b_1 NI_1 NS_50 0 1.8212815213589897e-03
GC_1_51 b_1 NI_1 NS_51 0 1.1492372185410180e-05
GC_1_52 b_1 NI_1 NS_52 0 2.6773245782678936e-04
GC_1_53 b_1 NI_1 NS_53 0 1.4706217189955938e-03
GC_1_54 b_1 NI_1 NS_54 0 1.5313483725568249e-03
GC_1_55 b_1 NI_1 NS_55 0 3.6979373772631210e-03
GC_1_56 b_1 NI_1 NS_56 0 -1.5576417364613587e-03
GC_1_57 b_1 NI_1 NS_57 0 8.9090973336950968e-06
GC_1_58 b_1 NI_1 NS_58 0 1.7982064842082847e-04
GC_1_59 b_1 NI_1 NS_59 0 3.7662360748474751e-03
GC_1_60 b_1 NI_1 NS_60 0 -9.6566071387888203e-04
GC_1_61 b_1 NI_1 NS_61 0 -1.2923373991674011e-05
GC_1_62 b_1 NI_1 NS_62 0 -1.8248740659875532e-05
GC_1_63 b_1 NI_1 NS_63 0 7.1094157626784148e-04
GC_1_64 b_1 NI_1 NS_64 0 7.8789453803976815e-04
GC_1_65 b_1 NI_1 NS_65 0 6.9875439836003537e-06
GC_1_66 b_1 NI_1 NS_66 0 -1.6667512570323851e-04
GC_1_67 b_1 NI_1 NS_67 0 1.0603608875771069e-05
GC_1_68 b_1 NI_1 NS_68 0 8.5927254266119775e-06
GC_1_69 b_1 NI_1 NS_69 0 -1.4703864252303207e-05
GC_1_70 b_1 NI_1 NS_70 0 4.2781098711767963e-05
GC_1_71 b_1 NI_1 NS_71 0 -3.2539133291888179e-03
GC_1_72 b_1 NI_1 NS_72 0 4.8648781222129724e-04
GC_1_73 b_1 NI_1 NS_73 0 1.2987898314872627e-05
GC_1_74 b_1 NI_1 NS_74 0 2.0804772805273408e-05
GC_1_75 b_1 NI_1 NS_75 0 6.0614633942236652e-04
GC_1_76 b_1 NI_1 NS_76 0 1.2521698098069936e-03
GC_1_77 b_1 NI_1 NS_77 0 3.4036488361297422e-06
GC_1_78 b_1 NI_1 NS_78 0 -8.9213045439782156e-07
GC_1_79 b_1 NI_1 NS_79 0 -1.3308613259046257e-04
GC_1_80 b_1 NI_1 NS_80 0 -6.3314922668327670e-04
GC_1_81 b_1 NI_1 NS_81 0 -3.7984225504397801e-06
GC_1_82 b_1 NI_1 NS_82 0 5.3450663379809049e-06
GC_1_83 b_1 NI_1 NS_83 0 -1.0293960352943536e-06
GC_1_84 b_1 NI_1 NS_84 0 -2.9364902467235754e-07
GC_1_85 b_1 NI_1 NS_85 0 1.9991216132128086e-06
GC_1_86 b_1 NI_1 NS_86 0 -2.1966949780688022e-06
GC_1_87 b_1 NI_1 NS_87 0 2.3950603489111473e-06
GC_1_88 b_1 NI_1 NS_88 0 -1.8509803733067500e-04
GC_1_89 b_1 NI_1 NS_89 0 1.6697373819334945e-03
GC_1_90 b_1 NI_1 NS_90 0 -5.0120088894000953e-05
GC_1_91 b_1 NI_1 NS_91 0 5.0844969784760562e-03
GC_1_92 b_1 NI_1 NS_92 0 4.8276131715846516e-03
GC_1_93 b_1 NI_1 NS_93 0 -5.5576302552346347e-03
GC_1_94 b_1 NI_1 NS_94 0 -4.8354387995109020e-03
GC_1_95 b_1 NI_1 NS_95 0 -3.1164530503589058e-04
GC_1_96 b_1 NI_1 NS_96 0 2.5189387951675537e-04
GC_1_97 b_1 NI_1 NS_97 0 1.4815451307419731e-03
GC_1_98 b_1 NI_1 NS_98 0 5.4309255497519658e-03
GC_1_99 b_1 NI_1 NS_99 0 -3.0290115909179212e-03
GC_1_100 b_1 NI_1 NS_100 0 -1.0501070390127047e-03
GC_1_101 b_1 NI_1 NS_101 0 8.7340228414929395e-04
GC_1_102 b_1 NI_1 NS_102 0 2.8128318091006206e-04
GC_1_103 b_1 NI_1 NS_103 0 -5.4787229084373255e-03
GC_1_104 b_1 NI_1 NS_104 0 -2.2171752965860947e-03
GC_1_105 b_1 NI_1 NS_105 0 -1.0992863609807997e-04
GC_1_106 b_1 NI_1 NS_106 0 9.7725631757524566e-05
GC_1_107 b_1 NI_1 NS_107 0 -1.9544070003646077e-03
GC_1_108 b_1 NI_1 NS_108 0 -3.2931014996275616e-03
GC_1_109 b_1 NI_1 NS_109 0 -2.1733802054046847e-04
GC_1_110 b_1 NI_1 NS_110 0 4.2382574280200124e-04
GC_1_111 b_1 NI_1 NS_111 0 1.6775058785315053e-04
GC_1_112 b_1 NI_1 NS_112 0 -6.0504504543195670e-05
GC_1_113 b_1 NI_1 NS_113 0 1.2085079702516062e-05
GC_1_114 b_1 NI_1 NS_114 0 -1.1186492330431959e-04
GC_1_115 b_1 NI_1 NS_115 0 7.2947654497897332e-03
GC_1_116 b_1 NI_1 NS_116 0 2.0806936961779458e-03
GC_1_117 b_1 NI_1 NS_117 0 -1.4267197436467143e-05
GC_1_118 b_1 NI_1 NS_118 0 -9.5877947873880992e-06
GC_1_119 b_1 NI_1 NS_119 0 6.7126821598653534e-04
GC_1_120 b_1 NI_1 NS_120 0 -3.8047555250349543e-03
GC_1_121 b_1 NI_1 NS_121 0 5.2078306130550098e-07
GC_1_122 b_1 NI_1 NS_122 0 -1.1131565179263749e-05
GC_1_123 b_1 NI_1 NS_123 0 8.3907073796223204e-04
GC_1_124 b_1 NI_1 NS_124 0 1.1031860659254759e-03
GC_1_125 b_1 NI_1 NS_125 0 1.5777727547449042e-05
GC_1_126 b_1 NI_1 NS_126 0 9.4458341171161437e-06
GC_1_127 b_1 NI_1 NS_127 0 8.1870871110488924e-08
GC_1_128 b_1 NI_1 NS_128 0 4.9826430716174011e-06
GC_1_129 b_1 NI_1 NS_129 0 -1.6793242351356264e-06
GC_1_130 b_1 NI_1 NS_130 0 -3.2297986071230524e-06
GC_1_131 b_1 NI_1 NS_131 0 2.1471902395387210e-05
GC_1_132 b_1 NI_1 NS_132 0 1.4413908645220596e-04
GC_1_133 b_1 NI_1 NS_133 0 5.8037900906121216e-02
GC_1_134 b_1 NI_1 NS_134 0 -4.5391613495295567e-05
GC_1_135 b_1 NI_1 NS_135 0 -6.3536055289223712e-03
GC_1_136 b_1 NI_1 NS_136 0 -2.8143303563142067e-03
GC_1_137 b_1 NI_1 NS_137 0 4.5439174102081233e-03
GC_1_138 b_1 NI_1 NS_138 0 2.6349731676868372e-03
GC_1_139 b_1 NI_1 NS_139 0 -4.5415304332687467e-05
GC_1_140 b_1 NI_1 NS_140 0 -1.7645941422076472e-04
GC_1_141 b_1 NI_1 NS_141 0 1.4094138612822024e-03
GC_1_142 b_1 NI_1 NS_142 0 1.6567426435881026e-03
GC_1_143 b_1 NI_1 NS_143 0 -3.2810119539541509e-04
GC_1_144 b_1 NI_1 NS_144 0 -6.3409302635688159e-04
GC_1_145 b_1 NI_1 NS_145 0 -7.6751548956815942e-05
GC_1_146 b_1 NI_1 NS_146 0 6.6003546610050718e-05
GC_1_147 b_1 NI_1 NS_147 0 -3.9096021769548361e-03
GC_1_148 b_1 NI_1 NS_148 0 7.7685266607894815e-04
GC_1_149 b_1 NI_1 NS_149 0 -4.9588475767236331e-05
GC_1_150 b_1 NI_1 NS_150 0 -6.0471268019264827e-05
GC_1_151 b_1 NI_1 NS_151 0 -1.7887581782519916e-04
GC_1_152 b_1 NI_1 NS_152 0 8.0545532402763193e-04
GC_1_153 b_1 NI_1 NS_153 0 3.3912111260390131e-04
GC_1_154 b_1 NI_1 NS_154 0 1.0742553045665405e-04
GC_1_155 b_1 NI_1 NS_155 0 -2.2963037655245031e-05
GC_1_156 b_1 NI_1 NS_156 0 -2.3066274517281786e-05
GC_1_157 b_1 NI_1 NS_157 0 -4.0039232481966269e-05
GC_1_158 b_1 NI_1 NS_158 0 5.7029416419148864e-05
GC_1_159 b_1 NI_1 NS_159 0 -2.9145374628041184e-03
GC_1_160 b_1 NI_1 NS_160 0 -3.6207520560060371e-03
GC_1_161 b_1 NI_1 NS_161 0 1.3068746771748823e-05
GC_1_162 b_1 NI_1 NS_162 0 3.1587675462647662e-05
GC_1_163 b_1 NI_1 NS_163 0 -4.5771698857901790e-04
GC_1_164 b_1 NI_1 NS_164 0 1.9610214189121032e-03
GC_1_165 b_1 NI_1 NS_165 0 -2.2807158662638967e-07
GC_1_166 b_1 NI_1 NS_166 0 6.2996816325074340e-06
GC_1_167 b_1 NI_1 NS_167 0 8.8143137151351593e-04
GC_1_168 b_1 NI_1 NS_168 0 -3.5786971009416844e-04
GC_1_169 b_1 NI_1 NS_169 0 -7.6419218427490811e-06
GC_1_170 b_1 NI_1 NS_170 0 -7.5620559026666551e-06
GC_1_171 b_1 NI_1 NS_171 0 1.6426148471316235e-06
GC_1_172 b_1 NI_1 NS_172 0 -1.8962551749925845e-07
GC_1_173 b_1 NI_1 NS_173 0 1.4166606020935609e-06
GC_1_174 b_1 NI_1 NS_174 0 2.3011833010093542e-06
GC_1_175 b_1 NI_1 NS_175 0 1.4619905505239847e-04
GC_1_176 b_1 NI_1 NS_176 0 -9.6902802604472359e-05
GC_1_177 b_1 NI_1 NS_177 0 3.2244365381018311e-02
GC_1_178 b_1 NI_1 NS_178 0 9.9828524789883093e-05
GC_1_179 b_1 NI_1 NS_179 0 6.0074318997944878e-03
GC_1_180 b_1 NI_1 NS_180 0 1.1808748036717923e-03
GC_1_181 b_1 NI_1 NS_181 0 -4.3858387871981439e-03
GC_1_182 b_1 NI_1 NS_182 0 2.6167250205408215e-03
GC_1_183 b_1 NI_1 NS_183 0 -1.9520787425790704e-04
GC_1_184 b_1 NI_1 NS_184 0 -9.2904559743261844e-04
GC_1_185 b_1 NI_1 NS_185 0 1.2072633119759133e-03
GC_1_186 b_1 NI_1 NS_186 0 6.0278955275660968e-03
GC_1_187 b_1 NI_1 NS_187 0 -1.0133194922044588e-02
GC_1_188 b_1 NI_1 NS_188 0 -1.2931473172068770e-03
GC_1_189 b_1 NI_1 NS_189 0 8.6808542154881343e-04
GC_1_190 b_1 NI_1 NS_190 0 2.4012285397753946e-04
GC_1_191 b_1 NI_1 NS_191 0 -2.6165023295719367e-03
GC_1_192 b_1 NI_1 NS_192 0 3.6605151018870085e-04
GC_1_193 b_1 NI_1 NS_193 0 -7.6933221237117253e-05
GC_1_194 b_1 NI_1 NS_194 0 1.2695582223971649e-04
GC_1_195 b_1 NI_1 NS_195 0 -1.9995731939127601e-03
GC_1_196 b_1 NI_1 NS_196 0 -3.7551143656492378e-03
GC_1_197 b_1 NI_1 NS_197 0 -9.6756900529073423e-05
GC_1_198 b_1 NI_1 NS_198 0 6.2460712247690037e-04
GC_1_199 b_1 NI_1 NS_199 0 1.5201611792864758e-04
GC_1_200 b_1 NI_1 NS_200 0 -7.2212052149634782e-05
GC_1_201 b_1 NI_1 NS_201 0 -4.6513391131842514e-06
GC_1_202 b_1 NI_1 NS_202 0 -1.0029132993858410e-04
GC_1_203 b_1 NI_1 NS_203 0 3.3711763004230580e-03
GC_1_204 b_1 NI_1 NS_204 0 -2.1823934856325337e-03
GC_1_205 b_1 NI_1 NS_205 0 -1.4940585946518276e-05
GC_1_206 b_1 NI_1 NS_206 0 -2.1910509333569713e-06
GC_1_207 b_1 NI_1 NS_207 0 -4.3001084136361548e-04
GC_1_208 b_1 NI_1 NS_208 0 -2.5085607215778504e-03
GC_1_209 b_1 NI_1 NS_209 0 -4.7110668039431212e-07
GC_1_210 b_1 NI_1 NS_210 0 -6.5528040241115868e-06
GC_1_211 b_1 NI_1 NS_211 0 1.4780811372272541e-03
GC_1_212 b_1 NI_1 NS_212 0 8.3287926240553460e-04
GC_1_213 b_1 NI_1 NS_213 0 8.6742405901321320e-06
GC_1_214 b_1 NI_1 NS_214 0 2.8103872213186546e-06
GC_1_215 b_1 NI_1 NS_215 0 1.7339333176097825e-06
GC_1_216 b_1 NI_1 NS_216 0 3.7347143986822790e-06
GC_1_217 b_1 NI_1 NS_217 0 3.9892378281140207e-07
GC_1_218 b_1 NI_1 NS_218 0 9.7631192673859712e-08
GC_1_219 b_1 NI_1 NS_219 0 1.6077375853778324e-04
GC_1_220 b_1 NI_1 NS_220 0 1.1337143098284064e-04
GC_1_221 b_1 NI_1 NS_221 0 3.9830603413155523e-02
GC_1_222 b_1 NI_1 NS_222 0 -2.4322542858021167e-04
GC_1_223 b_1 NI_1 NS_223 0 -5.7110893755188321e-03
GC_1_224 b_1 NI_1 NS_224 0 7.2542276915758179e-04
GC_1_225 b_1 NI_1 NS_225 0 2.5474744465967744e-03
GC_1_226 b_1 NI_1 NS_226 0 -2.5373687858313574e-03
GC_1_227 b_1 NI_1 NS_227 0 -1.4254927955505018e-04
GC_1_228 b_1 NI_1 NS_228 0 -9.8480191357938954e-05
GC_1_229 b_1 NI_1 NS_229 0 2.2444319477639644e-03
GC_1_230 b_1 NI_1 NS_230 0 1.5038716766531536e-03
GC_1_231 b_1 NI_1 NS_231 0 -3.9323770329182869e-03
GC_1_232 b_1 NI_1 NS_232 0 -2.6470139829315816e-04
GC_1_233 b_1 NI_1 NS_233 0 4.0227174841897206e-05
GC_1_234 b_1 NI_1 NS_234 0 4.4920581907517977e-05
GC_1_235 b_1 NI_1 NS_235 0 -5.2289784564181366e-04
GC_1_236 b_1 NI_1 NS_236 0 4.9940666810009111e-05
GC_1_237 b_1 NI_1 NS_237 0 -3.9921698107531255e-05
GC_1_238 b_1 NI_1 NS_238 0 -6.7229226929192793e-05
GC_1_239 b_1 NI_1 NS_239 0 3.7977461228863298e-04
GC_1_240 b_1 NI_1 NS_240 0 6.0672558288453449e-04
GC_1_241 b_1 NI_1 NS_241 0 2.6790942013859567e-04
GC_1_242 b_1 NI_1 NS_242 0 9.6544193118335508e-05
GC_1_243 b_1 NI_1 NS_243 0 6.6752439797879249e-06
GC_1_244 b_1 NI_1 NS_244 0 -4.0602730927203883e-05
GC_1_245 b_1 NI_1 NS_245 0 -4.8598436738465764e-05
GC_1_246 b_1 NI_1 NS_246 0 6.2512102460201036e-05
GC_1_247 b_1 NI_1 NS_247 0 -1.3971105494407123e-03
GC_1_248 b_1 NI_1 NS_248 0 -3.7813793889459961e-03
GC_1_249 b_1 NI_1 NS_249 0 1.2454946637459335e-05
GC_1_250 b_1 NI_1 NS_250 0 3.7793609042421377e-05
GC_1_251 b_1 NI_1 NS_251 0 -7.5664292325685234e-04
GC_1_252 b_1 NI_1 NS_252 0 1.7285494986425504e-03
GC_1_253 b_1 NI_1 NS_253 0 -2.0679609809084274e-06
GC_1_254 b_1 NI_1 NS_254 0 4.9619035889870845e-06
GC_1_255 b_1 NI_1 NS_255 0 8.0168064261095591e-04
GC_1_256 b_1 NI_1 NS_256 0 -1.1023020684585917e-04
GC_1_257 b_1 NI_1 NS_257 0 -3.9683682383379087e-06
GC_1_258 b_1 NI_1 NS_258 0 -7.6300296422107490e-06
GC_1_259 b_1 NI_1 NS_259 0 1.5154235565014082e-06
GC_1_260 b_1 NI_1 NS_260 0 1.3076496067110403e-06
GC_1_261 b_1 NI_1 NS_261 0 3.0137216686272537e-07
GC_1_262 b_1 NI_1 NS_262 0 4.8592073808610220e-07
GC_1_263 b_1 NI_1 NS_263 0 8.3304624356564415e-05
GC_1_264 b_1 NI_1 NS_264 0 -1.1370974196743040e-04
GC_1_265 b_1 NI_1 NS_265 0 5.9439141075038277e-03
GC_1_266 b_1 NI_1 NS_266 0 2.1847207595827707e-04
GC_1_267 b_1 NI_1 NS_267 0 3.9291690159792246e-03
GC_1_268 b_1 NI_1 NS_268 0 -1.0764521587493950e-03
GC_1_269 b_1 NI_1 NS_269 0 -1.1873467967318211e-03
GC_1_270 b_1 NI_1 NS_270 0 3.8898348437263626e-03
GC_1_271 b_1 NI_1 NS_271 0 -5.8511401980053447e-05
GC_1_272 b_1 NI_1 NS_272 0 9.3949177498926003e-05
GC_1_273 b_1 NI_1 NS_273 0 1.0192425276668016e-03
GC_1_274 b_1 NI_1 NS_274 0 4.4797091585926313e-03
GC_1_275 b_1 NI_1 NS_275 0 -1.1924405994036094e-02
GC_1_276 b_1 NI_1 NS_276 0 -9.9346967045963819e-04
GC_1_277 b_1 NI_1 NS_277 0 6.9198140464818805e-04
GC_1_278 b_1 NI_1 NS_278 0 8.6915782298134980e-05
GC_1_279 b_1 NI_1 NS_279 0 2.5020735855891155e-03
GC_1_280 b_1 NI_1 NS_280 0 -2.0610917870754458e-03
GC_1_281 b_1 NI_1 NS_281 0 -1.3573399584812669e-05
GC_1_282 b_1 NI_1 NS_282 0 9.8333464698855075e-05
GC_1_283 b_1 NI_1 NS_283 0 -1.0167624825651426e-03
GC_1_284 b_1 NI_1 NS_284 0 -3.1477886591752329e-03
GC_1_285 b_1 NI_1 NS_285 0 -1.5179162226960585e-04
GC_1_286 b_1 NI_1 NS_286 0 1.1321621590843058e-03
GC_1_287 b_1 NI_1 NS_287 0 1.3200640895543001e-04
GC_1_288 b_1 NI_1 NS_288 0 -8.2116949274852312e-05
GC_1_289 b_1 NI_1 NS_289 0 -1.0844656256587999e-05
GC_1_290 b_1 NI_1 NS_290 0 -6.6003135291765514e-05
GC_1_291 b_1 NI_1 NS_291 0 4.3543271228872089e-03
GC_1_292 b_1 NI_1 NS_292 0 -1.1807794080609722e-03
GC_1_293 b_1 NI_1 NS_293 0 -1.2831524221951114e-05
GC_1_294 b_1 NI_1 NS_294 0 1.3708259122505064e-06
GC_1_295 b_1 NI_1 NS_295 0 -9.4374339325577488e-04
GC_1_296 b_1 NI_1 NS_296 0 -2.1709858007473068e-03
GC_1_297 b_1 NI_1 NS_297 0 -8.8601880366951639e-06
GC_1_298 b_1 NI_1 NS_298 0 -3.6726130159209824e-06
GC_1_299 b_1 NI_1 NS_299 0 1.2863760193726514e-03
GC_1_300 b_1 NI_1 NS_300 0 1.6432059899656487e-03
GC_1_301 b_1 NI_1 NS_301 0 1.4652244934737856e-05
GC_1_302 b_1 NI_1 NS_302 0 -6.3341415224213071e-06
GC_1_303 b_1 NI_1 NS_303 0 2.6462469594757966e-06
GC_1_304 b_1 NI_1 NS_304 0 5.0865518989540508e-06
GC_1_305 b_1 NI_1 NS_305 0 -4.2435176385800989e-06
GC_1_306 b_1 NI_1 NS_306 0 1.4705365649890285e-06
GC_1_307 b_1 NI_1 NS_307 0 6.4674498450183537e-05
GC_1_308 b_1 NI_1 NS_308 0 2.0173185710046343e-04
GC_1_309 b_1 NI_1 NS_309 0 2.4593395635430306e-02
GC_1_310 b_1 NI_1 NS_310 0 -2.7114935220220673e-04
GC_1_311 b_1 NI_1 NS_311 0 -3.1075014061223358e-03
GC_1_312 b_1 NI_1 NS_312 0 2.1556221558190055e-03
GC_1_313 b_1 NI_1 NS_313 0 -1.6908285275136971e-04
GC_1_314 b_1 NI_1 NS_314 0 -2.9744396168019599e-03
GC_1_315 b_1 NI_1 NS_315 0 7.5991706639915376e-05
GC_1_316 b_1 NI_1 NS_316 0 -2.4659598432703747e-04
GC_1_317 b_1 NI_1 NS_317 0 1.4466916131030448e-03
GC_1_318 b_1 NI_1 NS_318 0 9.0058273376340749e-04
GC_1_319 b_1 NI_1 NS_319 0 -5.0460613125761812e-03
GC_1_320 b_1 NI_1 NS_320 0 8.7682714817568055e-04
GC_1_321 b_1 NI_1 NS_321 0 3.0130002307541898e-05
GC_1_322 b_1 NI_1 NS_322 0 4.0039849902530651e-07
GC_1_323 b_1 NI_1 NS_323 0 1.8645445605347554e-04
GC_1_324 b_1 NI_1 NS_324 0 -1.9818018239620618e-03
GC_1_325 b_1 NI_1 NS_325 0 -2.0176917700360823e-05
GC_1_326 b_1 NI_1 NS_326 0 -3.9507402812617429e-05
GC_1_327 b_1 NI_1 NS_327 0 2.8860100231298833e-04
GC_1_328 b_1 NI_1 NS_328 0 -4.9452534854412775e-06
GC_1_329 b_1 NI_1 NS_329 0 7.1942322667059179e-05
GC_1_330 b_1 NI_1 NS_330 0 3.7908808386443627e-06
GC_1_331 b_1 NI_1 NS_331 0 1.1194651046383540e-05
GC_1_332 b_1 NI_1 NS_332 0 -4.4453585841238168e-05
GC_1_333 b_1 NI_1 NS_333 0 -3.1554967382992325e-05
GC_1_334 b_1 NI_1 NS_334 0 3.3040657505891118e-05
GC_1_335 b_1 NI_1 NS_335 0 9.3944094759640156e-04
GC_1_336 b_1 NI_1 NS_336 0 -2.6364004920619018e-03
GC_1_337 b_1 NI_1 NS_337 0 -1.2270495979963039e-07
GC_1_338 b_1 NI_1 NS_338 0 1.9316389584396044e-05
GC_1_339 b_1 NI_1 NS_339 0 -8.6168010287738606e-04
GC_1_340 b_1 NI_1 NS_340 0 4.2423950698938496e-04
GC_1_341 b_1 NI_1 NS_341 0 -1.8533796821895697e-06
GC_1_342 b_1 NI_1 NS_342 0 6.8712208339130478e-07
GC_1_343 b_1 NI_1 NS_343 0 3.4391126458477008e-04
GC_1_344 b_1 NI_1 NS_344 0 1.6790993975083265e-04
GC_1_345 b_1 NI_1 NS_345 0 8.0359013802303584e-07
GC_1_346 b_1 NI_1 NS_346 0 -5.0402799792679988e-06
GC_1_347 b_1 NI_1 NS_347 0 5.9990434538679998e-07
GC_1_348 b_1 NI_1 NS_348 0 1.8242004974385361e-06
GC_1_349 b_1 NI_1 NS_349 0 -1.2684532561972118e-06
GC_1_350 b_1 NI_1 NS_350 0 3.3700601046523444e-07
GC_1_351 b_1 NI_1 NS_351 0 1.1952390348898651e-05
GC_1_352 b_1 NI_1 NS_352 0 -4.1352774710926037e-06
GC_1_353 b_1 NI_1 NS_353 0 1.2161754773318831e-02
GC_1_354 b_1 NI_1 NS_354 0 2.9743901560526829e-05
GC_1_355 b_1 NI_1 NS_355 0 -8.0268601602778903e-05
GC_1_356 b_1 NI_1 NS_356 0 -3.8275723532711897e-04
GC_1_357 b_1 NI_1 NS_357 0 5.0603859991711056e-04
GC_1_358 b_1 NI_1 NS_358 0 -3.1256005231616223e-04
GC_1_359 b_1 NI_1 NS_359 0 -6.7844626113888794e-04
GC_1_360 b_1 NI_1 NS_360 0 -7.6615536974570898e-05
GC_1_361 b_1 NI_1 NS_361 0 8.2391435273082862e-04
GC_1_362 b_1 NI_1 NS_362 0 -3.4301927393208309e-04
GC_1_363 b_1 NI_1 NS_363 0 -3.8630160292228244e-04
GC_1_364 b_1 NI_1 NS_364 0 7.9971579165249841e-05
GC_1_365 b_1 NI_1 NS_365 0 4.1339530172847537e-04
GC_1_366 b_1 NI_1 NS_366 0 -5.0204318453818853e-04
GC_1_367 b_1 NI_1 NS_367 0 4.5638961828215977e-03
GC_1_368 b_1 NI_1 NS_368 0 -3.0340001917996290e-04
GC_1_369 b_1 NI_1 NS_369 0 3.0315089964361332e-04
GC_1_370 b_1 NI_1 NS_370 0 2.6717916448789529e-04
GC_1_371 b_1 NI_1 NS_371 0 -1.1764918184446032e-04
GC_1_372 b_1 NI_1 NS_372 0 2.6577146495062494e-03
GC_1_373 b_1 NI_1 NS_373 0 3.7125976346917252e-04
GC_1_374 b_1 NI_1 NS_374 0 -3.2361049430442660e-04
GC_1_375 b_1 NI_1 NS_375 0 1.2111192952154360e-04
GC_1_376 b_1 NI_1 NS_376 0 -2.2611626581933857e-05
GC_1_377 b_1 NI_1 NS_377 0 2.2635844586056694e-05
GC_1_378 b_1 NI_1 NS_378 0 1.1332281423413358e-04
GC_1_379 b_1 NI_1 NS_379 0 -6.9718390861099929e-03
GC_1_380 b_1 NI_1 NS_380 0 5.8338761727879541e-03
GC_1_381 b_1 NI_1 NS_381 0 1.3223443970589110e-05
GC_1_382 b_1 NI_1 NS_382 0 -1.0943210253338501e-05
GC_1_383 b_1 NI_1 NS_383 0 1.9431588743779613e-03
GC_1_384 b_1 NI_1 NS_384 0 -1.5744097608636569e-04
GC_1_385 b_1 NI_1 NS_385 0 4.6981066949268674e-06
GC_1_386 b_1 NI_1 NS_386 0 8.4502206083166101e-06
GC_1_387 b_1 NI_1 NS_387 0 -3.6496771315986596e-05
GC_1_388 b_1 NI_1 NS_388 0 -2.6828697374517915e-03
GC_1_389 b_1 NI_1 NS_389 0 -2.5651202033680220e-05
GC_1_390 b_1 NI_1 NS_390 0 5.1753396875528456e-06
GC_1_391 b_1 NI_1 NS_391 0 -1.6607257808640483e-06
GC_1_392 b_1 NI_1 NS_392 0 -2.6004079991518493e-06
GC_1_393 b_1 NI_1 NS_393 0 4.4174125241373036e-06
GC_1_394 b_1 NI_1 NS_394 0 1.8743929860939114e-06
GC_1_395 b_1 NI_1 NS_395 0 -5.3721009394822115e-05
GC_1_396 b_1 NI_1 NS_396 0 -6.8479971902531600e-04
GC_1_397 b_1 NI_1 NS_397 0 1.0445798345799338e-02
GC_1_398 b_1 NI_1 NS_398 0 1.1156105787391245e-05
GC_1_399 b_1 NI_1 NS_399 0 5.2714340756271368e-05
GC_1_400 b_1 NI_1 NS_400 0 1.2181908853533330e-04
GC_1_401 b_1 NI_1 NS_401 0 -1.6323517217964767e-04
GC_1_402 b_1 NI_1 NS_402 0 -3.8764789147163845e-05
GC_1_403 b_1 NI_1 NS_403 0 -5.0431481608023438e-04
GC_1_404 b_1 NI_1 NS_404 0 -1.4340181293234010e-04
GC_1_405 b_1 NI_1 NS_405 0 1.8245941052613744e-04
GC_1_406 b_1 NI_1 NS_406 0 -2.8130670806088590e-04
GC_1_407 b_1 NI_1 NS_407 0 9.4346780596149429e-04
GC_1_408 b_1 NI_1 NS_408 0 6.3595592619178980e-05
GC_1_409 b_1 NI_1 NS_409 0 9.3702367669502176e-05
GC_1_410 b_1 NI_1 NS_410 0 6.1330313913267068e-05
GC_1_411 b_1 NI_1 NS_411 0 -1.2731414047403253e-04
GC_1_412 b_1 NI_1 NS_412 0 1.7312365815718067e-03
GC_1_413 b_1 NI_1 NS_413 0 -1.3386865054418418e-04
GC_1_414 b_1 NI_1 NS_414 0 6.5364885657300027e-05
GC_1_415 b_1 NI_1 NS_415 0 -5.9194929116048540e-04
GC_1_416 b_1 NI_1 NS_416 0 -7.9692111308655078e-05
GC_1_417 b_1 NI_1 NS_417 0 2.6351458290963873e-05
GC_1_418 b_1 NI_1 NS_418 0 -1.3989659762915805e-04
GC_1_419 b_1 NI_1 NS_419 0 -3.3709172043436306e-05
GC_1_420 b_1 NI_1 NS_420 0 -1.0934840339605252e-04
GC_1_421 b_1 NI_1 NS_421 0 -5.2985295735444861e-06
GC_1_422 b_1 NI_1 NS_422 0 1.0607258538616541e-04
GC_1_423 b_1 NI_1 NS_423 0 -2.3076863553969540e-04
GC_1_424 b_1 NI_1 NS_424 0 5.7415774006542566e-04
GC_1_425 b_1 NI_1 NS_425 0 -2.2802594025869045e-05
GC_1_426 b_1 NI_1 NS_426 0 -1.2185415449016612e-05
GC_1_427 b_1 NI_1 NS_427 0 -1.6734881734388918e-04
GC_1_428 b_1 NI_1 NS_428 0 -1.8254091194523051e-04
GC_1_429 b_1 NI_1 NS_429 0 1.4834463486013979e-06
GC_1_430 b_1 NI_1 NS_430 0 1.1010844429528562e-06
GC_1_431 b_1 NI_1 NS_431 0 -1.1480178823947508e-04
GC_1_432 b_1 NI_1 NS_432 0 -3.8368668689656475e-04
GC_1_433 b_1 NI_1 NS_433 0 -9.8078584141059137e-06
GC_1_434 b_1 NI_1 NS_434 0 -8.7495988507300288e-06
GC_1_435 b_1 NI_1 NS_435 0 -1.0728586460534463e-06
GC_1_436 b_1 NI_1 NS_436 0 1.2891761205058786e-06
GC_1_437 b_1 NI_1 NS_437 0 2.1697494960313980e-06
GC_1_438 b_1 NI_1 NS_438 0 -2.0403189742074284e-06
GC_1_439 b_1 NI_1 NS_439 0 -2.2730625127760854e-04
GC_1_440 b_1 NI_1 NS_440 0 -7.0817492632299452e-05
GC_1_441 b_1 NI_1 NS_441 0 -4.8473916815966744e-03
GC_1_442 b_1 NI_1 NS_442 0 5.8193002899354805e-05
GC_1_443 b_1 NI_1 NS_443 0 2.5851860320962462e-04
GC_1_444 b_1 NI_1 NS_444 0 -6.1696650161298307e-04
GC_1_445 b_1 NI_1 NS_445 0 6.0893005021074066e-04
GC_1_446 b_1 NI_1 NS_446 0 2.5700322186621345e-04
GC_1_447 b_1 NI_1 NS_447 0 -1.7215809551212569e-04
GC_1_448 b_1 NI_1 NS_448 0 3.9989942726323299e-04
GC_1_449 b_1 NI_1 NS_449 0 8.3994807589333478e-04
GC_1_450 b_1 NI_1 NS_450 0 4.8884773325162168e-04
GC_1_451 b_1 NI_1 NS_451 0 -3.1212609639162934e-03
GC_1_452 b_1 NI_1 NS_452 0 9.1896700909249089e-04
GC_1_453 b_1 NI_1 NS_453 0 4.3581395274903625e-04
GC_1_454 b_1 NI_1 NS_454 0 -3.5686710409483195e-04
GC_1_455 b_1 NI_1 NS_455 0 3.0565703427524200e-03
GC_1_456 b_1 NI_1 NS_456 0 -2.4852298295441099e-03
GC_1_457 b_1 NI_1 NS_457 0 1.9537278461188187e-04
GC_1_458 b_1 NI_1 NS_458 0 1.9681133655354317e-04
GC_1_459 b_1 NI_1 NS_459 0 -2.6528209068734504e-04
GC_1_460 b_1 NI_1 NS_460 0 5.8143462088452525e-04
GC_1_461 b_1 NI_1 NS_461 0 1.9205127423270568e-04
GC_1_462 b_1 NI_1 NS_462 0 2.1095558442975064e-04
GC_1_463 b_1 NI_1 NS_463 0 1.0190831681283976e-04
GC_1_464 b_1 NI_1 NS_464 0 -5.0656230314723996e-05
GC_1_465 b_1 NI_1 NS_465 0 9.5731218470539933e-06
GC_1_466 b_1 NI_1 NS_466 0 6.0035205395878281e-05
GC_1_467 b_1 NI_1 NS_467 0 -1.7194347522206880e-03
GC_1_468 b_1 NI_1 NS_468 0 3.4195686875029985e-03
GC_1_469 b_1 NI_1 NS_469 0 2.2758905213513674e-06
GC_1_470 b_1 NI_1 NS_470 0 -4.2636900078676000e-06
GC_1_471 b_1 NI_1 NS_471 0 7.5314323528875523e-04
GC_1_472 b_1 NI_1 NS_472 0 -8.1751453313269509e-04
GC_1_473 b_1 NI_1 NS_473 0 -2.9690206858981618e-06
GC_1_474 b_1 NI_1 NS_474 0 4.5026133948528741e-06
GC_1_475 b_1 NI_1 NS_475 0 6.2327514251190653e-04
GC_1_476 b_1 NI_1 NS_476 0 -1.0591643280832223e-03
GC_1_477 b_1 NI_1 NS_477 0 -1.0813235041668274e-05
GC_1_478 b_1 NI_1 NS_478 0 -4.9049726031546414e-06
GC_1_479 b_1 NI_1 NS_479 0 1.1004026911296968e-06
GC_1_480 b_1 NI_1 NS_480 0 -1.0385899983451548e-07
GC_1_481 b_1 NI_1 NS_481 0 2.0437311008098350e-07
GC_1_482 b_1 NI_1 NS_482 0 3.5235791937134921e-06
GC_1_483 b_1 NI_1 NS_483 0 1.3478051518594475e-05
GC_1_484 b_1 NI_1 NS_484 0 -3.0832416697572894e-04
GC_1_485 b_1 NI_1 NS_485 0 1.6296100570224542e-02
GC_1_486 b_1 NI_1 NS_486 0 -4.1214930759864766e-05
GC_1_487 b_1 NI_1 NS_487 0 -1.2942858890983497e-04
GC_1_488 b_1 NI_1 NS_488 0 5.5166694215232992e-04
GC_1_489 b_1 NI_1 NS_489 0 -4.9372937055256470e-04
GC_1_490 b_1 NI_1 NS_490 0 -2.2001000782586537e-04
GC_1_491 b_1 NI_1 NS_491 0 -2.9651335720361595e-04
GC_1_492 b_1 NI_1 NS_492 0 -2.6444772323873215e-04
GC_1_493 b_1 NI_1 NS_493 0 3.1164403721717137e-04
GC_1_494 b_1 NI_1 NS_494 0 -1.7842808431383875e-05
GC_1_495 b_1 NI_1 NS_495 0 -2.9608771828721709e-04
GC_1_496 b_1 NI_1 NS_496 0 1.0793521325186579e-03
GC_1_497 b_1 NI_1 NS_497 0 6.5206642067170114e-05
GC_1_498 b_1 NI_1 NS_498 0 3.2526449929976082e-05
GC_1_499 b_1 NI_1 NS_499 0 -8.6557103879074176e-04
GC_1_500 b_1 NI_1 NS_500 0 3.8880528829984969e-04
GC_1_501 b_1 NI_1 NS_501 0 -7.9355488105477235e-05
GC_1_502 b_1 NI_1 NS_502 0 1.9610232945007817e-05
GC_1_503 b_1 NI_1 NS_503 0 -3.6832062914757372e-04
GC_1_504 b_1 NI_1 NS_504 0 -1.0776770031783321e-04
GC_1_505 b_1 NI_1 NS_505 0 3.4176600060913799e-05
GC_1_506 b_1 NI_1 NS_506 0 -1.0181431009055039e-04
GC_1_507 b_1 NI_1 NS_507 0 -1.9440086224947945e-05
GC_1_508 b_1 NI_1 NS_508 0 -7.0944857015246696e-05
GC_1_509 b_1 NI_1 NS_509 0 -1.2758381870427810e-05
GC_1_510 b_1 NI_1 NS_510 0 5.8006996866279153e-05
GC_1_511 b_1 NI_1 NS_511 0 -2.6139701436804388e-04
GC_1_512 b_1 NI_1 NS_512 0 -8.9675752226575211e-04
GC_1_513 b_1 NI_1 NS_513 0 -1.2869092278264391e-05
GC_1_514 b_1 NI_1 NS_514 0 -1.3641917638211865e-06
GC_1_515 b_1 NI_1 NS_515 0 -3.7957515310975534e-04
GC_1_516 b_1 NI_1 NS_516 0 1.4095067303047156e-04
GC_1_517 b_1 NI_1 NS_517 0 -7.3520098505045047e-08
GC_1_518 b_1 NI_1 NS_518 0 1.2107210602289666e-06
GC_1_519 b_1 NI_1 NS_519 0 1.2449040022568297e-04
GC_1_520 b_1 NI_1 NS_520 0 -1.0300443840577027e-04
GC_1_521 b_1 NI_1 NS_521 0 -4.9067850407212953e-06
GC_1_522 b_1 NI_1 NS_522 0 -6.2409973311675107e-06
GC_1_523 b_1 NI_1 NS_523 0 -2.0865144614751249e-07
GC_1_524 b_1 NI_1 NS_524 0 4.1086273005358835e-07
GC_1_525 b_1 NI_1 NS_525 0 1.0466101576849394e-06
GC_1_526 b_1 NI_1 NS_526 0 -1.1962861358791947e-07
GC_1_527 b_1 NI_1 NS_527 0 -7.0941532992741831e-05
GC_1_528 b_1 NI_1 NS_528 0 -2.8922823971479749e-05
GD_1_1 b_1 NI_1 NA_1 0 -1.0100667137732340e-01
GD_1_2 b_1 NI_1 NA_2 0 -4.2054647073772027e-03
GD_1_3 b_1 NI_1 NA_3 0 1.4295396546490033e-03
GD_1_4 b_1 NI_1 NA_4 0 -6.1519775667041386e-02
GD_1_5 b_1 NI_1 NA_5 0 -2.7144956678962173e-02
GD_1_6 b_1 NI_1 NA_6 0 -3.8611709331086236e-02
GD_1_7 b_1 NI_1 NA_7 0 -7.3137574927988709e-03
GD_1_8 b_1 NI_1 NA_8 0 -1.8618147620688572e-02
GD_1_9 b_1 NI_1 NA_9 0 -1.6578067018809286e-02
GD_1_10 b_1 NI_1 NA_10 0 -1.0469193834719726e-02
GD_1_11 b_1 NI_1 NA_11 0 1.6877265313405155e-03
GD_1_12 b_1 NI_1 NA_12 0 -1.4221113416621084e-02
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+01
GC_2_1 b_2 NI_2 NS_1 0 1.4058402975212405e-03
GC_2_2 b_2 NI_2 NS_2 0 1.0834322596881258e-02
GC_2_3 b_2 NI_2 NS_3 0 -6.4869261953688405e-03
GC_2_4 b_2 NI_2 NS_4 0 -5.6190407804785365e-03
GC_2_5 b_2 NI_2 NS_5 0 -1.0866853918875303e-02
GC_2_6 b_2 NI_2 NS_6 0 1.8212815213829120e-03
GC_2_7 b_2 NI_2 NS_7 0 1.1492372158718833e-05
GC_2_8 b_2 NI_2 NS_8 0 2.6773245806776446e-04
GC_2_9 b_2 NI_2 NS_9 0 1.4706217190605111e-03
GC_2_10 b_2 NI_2 NS_10 0 1.5313483725415908e-03
GC_2_11 b_2 NI_2 NS_11 0 3.6979373773191023e-03
GC_2_12 b_2 NI_2 NS_12 0 -1.5576417366394027e-03
GC_2_13 b_2 NI_2 NS_13 0 8.9090973468283019e-06
GC_2_14 b_2 NI_2 NS_14 0 1.7982064842492052e-04
GC_2_15 b_2 NI_2 NS_15 0 3.7662360751606143e-03
GC_2_16 b_2 NI_2 NS_16 0 -9.6566071399317363e-04
GC_2_17 b_2 NI_2 NS_17 0 -1.2923373986944569e-05
GC_2_18 b_2 NI_2 NS_18 0 -1.8248740656974027e-05
GC_2_19 b_2 NI_2 NS_19 0 7.1094157640879730e-04
GC_2_20 b_2 NI_2 NS_20 0 7.8789453802377487e-04
GC_2_21 b_2 NI_2 NS_21 0 6.9875439484755668e-06
GC_2_22 b_2 NI_2 NS_22 0 -1.6667512571381617e-04
GC_2_23 b_2 NI_2 NS_23 0 1.0603608882941899e-05
GC_2_24 b_2 NI_2 NS_24 0 8.5927254291963919e-06
GC_2_25 b_2 NI_2 NS_25 0 -1.4703864248740010e-05
GC_2_26 b_2 NI_2 NS_26 0 4.2781098708692474e-05
GC_2_27 b_2 NI_2 NS_27 0 -3.2539133289059248e-03
GC_2_28 b_2 NI_2 NS_28 0 4.8648781301922954e-04
GC_2_29 b_2 NI_2 NS_29 0 1.2987898314229245e-05
GC_2_30 b_2 NI_2 NS_30 0 2.0804772803695941e-05
GC_2_31 b_2 NI_2 NS_31 0 6.0614633956061835e-04
GC_2_32 b_2 NI_2 NS_32 0 1.2521698095847341e-03
GC_2_33 b_2 NI_2 NS_33 0 3.4036488367886915e-06
GC_2_34 b_2 NI_2 NS_34 0 -8.9213045563448183e-07
GC_2_35 b_2 NI_2 NS_35 0 -1.3308613274863723e-04
GC_2_36 b_2 NI_2 NS_36 0 -6.3314922665237737e-04
GC_2_37 b_2 NI_2 NS_37 0 -3.7984225492094529e-06
GC_2_38 b_2 NI_2 NS_38 0 5.3450663401339889e-06
GC_2_39 b_2 NI_2 NS_39 0 -1.0293960357746952e-06
GC_2_40 b_2 NI_2 NS_40 0 -2.9364902438912153e-07
GC_2_41 b_2 NI_2 NS_41 0 1.9991216129817346e-06
GC_2_42 b_2 NI_2 NS_42 0 -2.1966949788894641e-06
GC_2_43 b_2 NI_2 NS_43 0 2.3950603178843309e-06
GC_2_44 b_2 NI_2 NS_44 0 -1.8509803733382786e-04
GC_2_45 b_2 NI_2 NS_45 0 -2.2001127553199096e-01
GC_2_46 b_2 NI_2 NS_46 0 8.6776004812808439e-03
GC_2_47 b_2 NI_2 NS_47 0 4.1287540551673586e-03
GC_2_48 b_2 NI_2 NS_48 0 6.0575340134017552e-03
GC_2_49 b_2 NI_2 NS_49 0 6.8346783401236552e-03
GC_2_50 b_2 NI_2 NS_50 0 -1.9621000288993738e-03
GC_2_51 b_2 NI_2 NS_51 0 1.2246461149757746e-03
GC_2_52 b_2 NI_2 NS_52 0 -1.0786783028566162e-04
GC_2_53 b_2 NI_2 NS_53 0 3.8411590336271501e-04
GC_2_54 b_2 NI_2 NS_54 0 1.3264045829367681e-03
GC_2_55 b_2 NI_2 NS_55 0 5.2349361556080359e-03
GC_2_56 b_2 NI_2 NS_56 0 1.2154742595105682e-03
GC_2_57 b_2 NI_2 NS_57 0 -1.4363020765269165e-04
GC_2_58 b_2 NI_2 NS_58 0 3.0662137637170906e-04
GC_2_59 b_2 NI_2 NS_59 0 2.7666525253714816e-03
GC_2_60 b_2 NI_2 NS_60 0 7.1763483728655405e-03
GC_2_61 b_2 NI_2 NS_61 0 -5.3418004796635774e-05
GC_2_62 b_2 NI_2 NS_62 0 1.1067716016956187e-04
GC_2_63 b_2 NI_2 NS_63 0 1.1993860530529138e-04
GC_2_64 b_2 NI_2 NS_64 0 3.4692618782689003e-03
GC_2_65 b_2 NI_2 NS_65 0 6.6544117773241680e-04
GC_2_66 b_2 NI_2 NS_66 0 -3.9442377442099123e-04
GC_2_67 b_2 NI_2 NS_67 0 -8.5818206827495638e-05
GC_2_68 b_2 NI_2 NS_68 0 1.5883890125604339e-04
GC_2_69 b_2 NI_2 NS_69 0 3.7994419532440881e-05
GC_2_70 b_2 NI_2 NS_70 0 2.9757036850694510e-05
GC_2_71 b_2 NI_2 NS_71 0 -1.7575594545693539e-02
GC_2_72 b_2 NI_2 NS_72 0 2.6455701825043366e-03
GC_2_73 b_2 NI_2 NS_73 0 1.4353643927555864e-05
GC_2_74 b_2 NI_2 NS_74 0 -4.7573627166124203e-05
GC_2_75 b_2 NI_2 NS_75 0 5.0567764071091795e-03
GC_2_76 b_2 NI_2 NS_76 0 4.1359723107699982e-03
GC_2_77 b_2 NI_2 NS_77 0 -2.5016663078765796e-06
GC_2_78 b_2 NI_2 NS_78 0 3.9399324406717892e-05
GC_2_79 b_2 NI_2 NS_79 0 1.0324850793571577e-03
GC_2_80 b_2 NI_2 NS_80 0 -2.7131626074668683e-03
GC_2_81 b_2 NI_2 NS_81 0 -5.5258007880177276e-05
GC_2_82 b_2 NI_2 NS_82 0 -1.2894103312298068e-05
GC_2_83 b_2 NI_2 NS_83 0 1.4977403051059307e-05
GC_2_84 b_2 NI_2 NS_84 0 -1.5205905818172141e-05
GC_2_85 b_2 NI_2 NS_85 0 4.6166792103562786e-05
GC_2_86 b_2 NI_2 NS_86 0 -5.9782340225934370e-06
GC_2_87 b_2 NI_2 NS_87 0 1.8588492924885271e-04
GC_2_88 b_2 NI_2 NS_88 0 -5.6239918868666958e-04
GC_2_89 b_2 NI_2 NS_89 0 5.8822982993476276e-02
GC_2_90 b_2 NI_2 NS_90 0 -2.0743972438092671e-05
GC_2_91 b_2 NI_2 NS_91 0 -6.4253479494355550e-03
GC_2_92 b_2 NI_2 NS_92 0 -2.9556840752267169e-03
GC_2_93 b_2 NI_2 NS_93 0 4.8501814027708491e-03
GC_2_94 b_2 NI_2 NS_94 0 2.5544219366961363e-03
GC_2_95 b_2 NI_2 NS_95 0 -1.1777984066523793e-04
GC_2_96 b_2 NI_2 NS_96 0 -1.0482802430901682e-04
GC_2_97 b_2 NI_2 NS_97 0 1.6246303186501379e-03
GC_2_98 b_2 NI_2 NS_98 0 1.6016138331532486e-03
GC_2_99 b_2 NI_2 NS_99 0 -3.1790549529395109e-04
GC_2_100 b_2 NI_2 NS_100 0 -7.7117063514732021e-04
GC_2_101 b_2 NI_2 NS_101 0 -2.6956419841883970e-05
GC_2_102 b_2 NI_2 NS_102 0 6.6565596268967304e-05
GC_2_103 b_2 NI_2 NS_103 0 -3.2915211789542789e-03
GC_2_104 b_2 NI_2 NS_104 0 1.1532590937596040e-03
GC_2_105 b_2 NI_2 NS_105 0 -4.8040738315665625e-05
GC_2_106 b_2 NI_2 NS_106 0 -7.1932092230862354e-05
GC_2_107 b_2 NI_2 NS_107 0 7.8901572706784268e-05
GC_2_108 b_2 NI_2 NS_108 0 1.1148674095202333e-03
GC_2_109 b_2 NI_2 NS_109 0 3.2507030977643226e-04
GC_2_110 b_2 NI_2 NS_110 0 6.9320459497553295e-05
GC_2_111 b_2 NI_2 NS_111 0 -2.1473022745161151e-05
GC_2_112 b_2 NI_2 NS_112 0 -2.3815535506497823e-05
GC_2_113 b_2 NI_2 NS_113 0 -4.9121302110090362e-05
GC_2_114 b_2 NI_2 NS_114 0 6.9075315037400083e-05
GC_2_115 b_2 NI_2 NS_115 0 -3.8810926570470566e-03
GC_2_116 b_2 NI_2 NS_116 0 -3.5079993583827175e-03
GC_2_117 b_2 NI_2 NS_117 0 1.4624435922295197e-05
GC_2_118 b_2 NI_2 NS_118 0 3.8510511261582809e-05
GC_2_119 b_2 NI_2 NS_119 0 -2.5984647498068336e-04
GC_2_120 b_2 NI_2 NS_120 0 2.3947784806132894e-03
GC_2_121 b_2 NI_2 NS_121 0 2.0090779392228769e-06
GC_2_122 b_2 NI_2 NS_122 0 9.9947949816447224e-06
GC_2_123 b_2 NI_2 NS_123 0 9.0676155276280879e-04
GC_2_124 b_2 NI_2 NS_124 0 -5.4484277564635403e-04
GC_2_125 b_2 NI_2 NS_125 0 -1.1759195875378817e-05
GC_2_126 b_2 NI_2 NS_126 0 -5.0239537945320735e-06
GC_2_127 b_2 NI_2 NS_127 0 2.0059892893832328e-06
GC_2_128 b_2 NI_2 NS_128 0 -1.7978369556616921e-06
GC_2_129 b_2 NI_2 NS_129 0 2.4366121628434648e-06
GC_2_130 b_2 NI_2 NS_130 0 -4.5690842062221068e-07
GC_2_131 b_2 NI_2 NS_131 0 1.4765342009750664e-04
GC_2_132 b_2 NI_2 NS_132 0 -1.5970040653064875e-04
GC_2_133 b_2 NI_2 NS_133 0 8.7751625046887886e-03
GC_2_134 b_2 NI_2 NS_134 0 -8.8798500392520878e-04
GC_2_135 b_2 NI_2 NS_135 0 4.0914945985620595e-03
GC_2_136 b_2 NI_2 NS_136 0 1.6307259179175616e-03
GC_2_137 b_2 NI_2 NS_137 0 -5.3014703535108620e-03
GC_2_138 b_2 NI_2 NS_138 0 -2.1301209067059856e-03
GC_2_139 b_2 NI_2 NS_139 0 2.8460769626067312e-04
GC_2_140 b_2 NI_2 NS_140 0 -2.7857758521860411e-04
GC_2_141 b_2 NI_2 NS_141 0 1.2238021832174327e-03
GC_2_142 b_2 NI_2 NS_142 0 1.5352189565951638e-04
GC_2_143 b_2 NI_2 NS_143 0 -1.1202117110782689e-04
GC_2_144 b_2 NI_2 NS_144 0 -5.2488576626504957e-04
GC_2_145 b_2 NI_2 NS_145 0 -1.8818100180628142e-05
GC_2_146 b_2 NI_2 NS_146 0 -3.7427298985640742e-05
GC_2_147 b_2 NI_2 NS_147 0 -1.1719674759323828e-03
GC_2_148 b_2 NI_2 NS_148 0 7.9808056929939523e-04
GC_2_149 b_2 NI_2 NS_149 0 2.2581156956849196e-05
GC_2_150 b_2 NI_2 NS_150 0 -1.1119962763800029e-05
GC_2_151 b_2 NI_2 NS_151 0 -3.3838560937798249e-05
GC_2_152 b_2 NI_2 NS_152 0 -6.9917908934367335e-05
GC_2_153 b_2 NI_2 NS_153 0 3.5064736468603446e-04
GC_2_154 b_2 NI_2 NS_154 0 -1.1489355420430048e-04
GC_2_155 b_2 NI_2 NS_155 0 -9.7941340582002348e-06
GC_2_156 b_2 NI_2 NS_156 0 -2.4824519250572327e-05
GC_2_157 b_2 NI_2 NS_157 0 -4.2367230515585613e-05
GC_2_158 b_2 NI_2 NS_158 0 -7.9066594821469361e-05
GC_2_159 b_2 NI_2 NS_159 0 9.9007343473547370e-04
GC_2_160 b_2 NI_2 NS_160 0 -9.7965342306983441e-04
GC_2_161 b_2 NI_2 NS_161 0 -3.3535994706684618e-05
GC_2_162 b_2 NI_2 NS_162 0 -3.7480040636434769e-05
GC_2_163 b_2 NI_2 NS_163 0 2.8908942326769013e-04
GC_2_164 b_2 NI_2 NS_164 0 -1.1664426970746394e-04
GC_2_165 b_2 NI_2 NS_165 0 -1.0500935039992515e-05
GC_2_166 b_2 NI_2 NS_166 0 1.2001480741592045e-05
GC_2_167 b_2 NI_2 NS_167 0 4.3994234634063420e-04
GC_2_168 b_2 NI_2 NS_168 0 6.7489705339294191e-05
GC_2_169 b_2 NI_2 NS_169 0 -1.8378090190189464e-07
GC_2_170 b_2 NI_2 NS_170 0 -9.7233119663194222e-06
GC_2_171 b_2 NI_2 NS_171 0 1.9425684177483119e-05
GC_2_172 b_2 NI_2 NS_172 0 2.9634541921464538e-07
GC_2_173 b_2 NI_2 NS_173 0 2.7196986586220121e-05
GC_2_174 b_2 NI_2 NS_174 0 -8.8295382135156994e-06
GC_2_175 b_2 NI_2 NS_175 0 -1.4646195799778239e-04
GC_2_176 b_2 NI_2 NS_176 0 8.9473388724064956e-05
GC_2_177 b_2 NI_2 NS_177 0 3.9622292483376273e-02
GC_2_178 b_2 NI_2 NS_178 0 -2.3691614670392602e-04
GC_2_179 b_2 NI_2 NS_179 0 -5.6773487281091091e-03
GC_2_180 b_2 NI_2 NS_180 0 6.9768052856374453e-04
GC_2_181 b_2 NI_2 NS_181 0 2.5618358951758997e-03
GC_2_182 b_2 NI_2 NS_182 0 -2.4925754830115656e-03
GC_2_183 b_2 NI_2 NS_183 0 -9.2175038542939894e-05
GC_2_184 b_2 NI_2 NS_184 0 -2.7688128249419995e-05
GC_2_185 b_2 NI_2 NS_185 0 2.2172444865325488e-03
GC_2_186 b_2 NI_2 NS_186 0 1.5253139973653328e-03
GC_2_187 b_2 NI_2 NS_187 0 -3.9397653556183026e-03
GC_2_188 b_2 NI_2 NS_188 0 -2.6243794844541332e-04
GC_2_189 b_2 NI_2 NS_189 0 3.7947450824796962e-05
GC_2_190 b_2 NI_2 NS_190 0 2.6486134502808498e-05
GC_2_191 b_2 NI_2 NS_191 0 -5.9147239085280466e-04
GC_2_192 b_2 NI_2 NS_192 0 -3.0435858891708229e-05
GC_2_193 b_2 NI_2 NS_193 0 -3.5906261591978308e-05
GC_2_194 b_2 NI_2 NS_194 0 -6.8523126878391820e-05
GC_2_195 b_2 NI_2 NS_195 0 3.9647464962658111e-04
GC_2_196 b_2 NI_2 NS_196 0 5.8710706304085185e-04
GC_2_197 b_2 NI_2 NS_197 0 2.6985515070225216e-04
GC_2_198 b_2 NI_2 NS_198 0 9.9496333014702481e-05
GC_2_199 b_2 NI_2 NS_199 0 1.6862576870972010e-06
GC_2_200 b_2 NI_2 NS_200 0 -3.9011134412972583e-05
GC_2_201 b_2 NI_2 NS_201 0 -4.0921664144193867e-05
GC_2_202 b_2 NI_2 NS_202 0 5.9107831721073261e-05
GC_2_203 b_2 NI_2 NS_203 0 -1.1821912787583939e-03
GC_2_204 b_2 NI_2 NS_204 0 -3.6957213809411834e-03
GC_2_205 b_2 NI_2 NS_205 0 1.2454417973425652e-05
GC_2_206 b_2 NI_2 NS_206 0 3.5707535556032961e-05
GC_2_207 b_2 NI_2 NS_207 0 -7.7345298232948327e-04
GC_2_208 b_2 NI_2 NS_208 0 1.6500640224596580e-03
GC_2_209 b_2 NI_2 NS_209 0 -3.2939445411258653e-06
GC_2_210 b_2 NI_2 NS_210 0 6.0222030231706096e-06
GC_2_211 b_2 NI_2 NS_211 0 7.5502075952894280e-04
GC_2_212 b_2 NI_2 NS_212 0 -1.1755906205145573e-04
GC_2_213 b_2 NI_2 NS_213 0 -3.7668355133041891e-06
GC_2_214 b_2 NI_2 NS_214 0 -5.7648358654874508e-06
GC_2_215 b_2 NI_2 NS_215 0 1.8659211073840687e-06
GC_2_216 b_2 NI_2 NS_216 0 1.1002313747246817e-06
GC_2_217 b_2 NI_2 NS_217 0 1.6261228557864982e-06
GC_2_218 b_2 NI_2 NS_218 0 9.8172636406247311e-07
GC_2_219 b_2 NI_2 NS_219 0 7.5333039514158877e-05
GC_2_220 b_2 NI_2 NS_220 0 -9.8976170960829473e-05
GC_2_221 b_2 NI_2 NS_221 0 1.0174600217514049e-02
GC_2_222 b_2 NI_2 NS_222 0 -2.8650416274140188e-04
GC_2_223 b_2 NI_2 NS_223 0 3.9837980473647529e-03
GC_2_224 b_2 NI_2 NS_224 0 -1.4862491485396927e-03
GC_2_225 b_2 NI_2 NS_225 0 -1.9750021259840791e-03
GC_2_226 b_2 NI_2 NS_226 0 2.5692173911277057e-03
GC_2_227 b_2 NI_2 NS_227 0 -4.0285519020060058e-04
GC_2_228 b_2 NI_2 NS_228 0 5.4624486785869429e-04
GC_2_229 b_2 NI_2 NS_229 0 1.0533751763607553e-03
GC_2_230 b_2 NI_2 NS_230 0 3.9215571415191609e-04
GC_2_231 b_2 NI_2 NS_231 0 -8.0041842156533625e-04
GC_2_232 b_2 NI_2 NS_232 0 1.5810096051280015e-03
GC_2_233 b_2 NI_2 NS_233 0 -7.2381194507423633e-05
GC_2_234 b_2 NI_2 NS_234 0 -1.1174353925629420e-05
GC_2_235 b_2 NI_2 NS_235 0 -8.1638383092287939e-04
GC_2_236 b_2 NI_2 NS_236 0 1.6523830353573422e-03
GC_2_237 b_2 NI_2 NS_237 0 5.3324304202860453e-06
GC_2_238 b_2 NI_2 NS_238 0 -9.9047558842280247e-06
GC_2_239 b_2 NI_2 NS_239 0 -5.7076756902267568e-04
GC_2_240 b_2 NI_2 NS_240 0 3.5892225163082194e-04
GC_2_241 b_2 NI_2 NS_241 0 8.0492513272587452e-04
GC_2_242 b_2 NI_2 NS_242 0 -2.5425679855862842e-04
GC_2_243 b_2 NI_2 NS_243 0 -5.0150945575030886e-05
GC_2_244 b_2 NI_2 NS_244 0 -2.0214685125658327e-05
GC_2_245 b_2 NI_2 NS_245 0 -6.4779125502897243e-05
GC_2_246 b_2 NI_2 NS_246 0 -8.3375408564636028e-05
GC_2_247 b_2 NI_2 NS_247 0 -1.9983725863938983e-03
GC_2_248 b_2 NI_2 NS_248 0 -4.0871062309706324e-03
GC_2_249 b_2 NI_2 NS_249 0 -3.7151760291130797e-05
GC_2_250 b_2 NI_2 NS_250 0 -4.0640124262322217e-05
GC_2_251 b_2 NI_2 NS_251 0 4.6431047538323593e-04
GC_2_252 b_2 NI_2 NS_252 0 1.1400822471267587e-03
GC_2_253 b_2 NI_2 NS_253 0 -1.1854253226335043e-05
GC_2_254 b_2 NI_2 NS_254 0 2.8311009773873334e-05
GC_2_255 b_2 NI_2 NS_255 0 1.3271215911634117e-03
GC_2_256 b_2 NI_2 NS_256 0 -5.6138040432383363e-04
GC_2_257 b_2 NI_2 NS_257 0 -1.6263062675046617e-05
GC_2_258 b_2 NI_2 NS_258 0 -2.1206591787451017e-05
GC_2_259 b_2 NI_2 NS_259 0 2.8840060827824208e-05
GC_2_260 b_2 NI_2 NS_260 0 -5.1580401549091257e-06
GC_2_261 b_2 NI_2 NS_261 0 3.6899101272514538e-05
GC_2_262 b_2 NI_2 NS_262 0 -1.3010675945555084e-05
GC_2_263 b_2 NI_2 NS_263 0 -2.4542530470495523e-05
GC_2_264 b_2 NI_2 NS_264 0 1.0909947824194106e-04
GC_2_265 b_2 NI_2 NS_265 0 2.3421754060701194e-02
GC_2_266 b_2 NI_2 NS_266 0 -2.5744160039830753e-04
GC_2_267 b_2 NI_2 NS_267 0 -3.1492332532563404e-03
GC_2_268 b_2 NI_2 NS_268 0 2.0868689764460303e-03
GC_2_269 b_2 NI_2 NS_269 0 -4.7099148742947230e-05
GC_2_270 b_2 NI_2 NS_270 0 -3.0612636009167806e-03
GC_2_271 b_2 NI_2 NS_271 0 1.8864770728500277e-04
GC_2_272 b_2 NI_2 NS_272 0 6.7951159675567053e-05
GC_2_273 b_2 NI_2 NS_273 0 1.5603791899446507e-03
GC_2_274 b_2 NI_2 NS_274 0 8.3668656894354235e-04
GC_2_275 b_2 NI_2 NS_275 0 -5.1453057171476184e-03
GC_2_276 b_2 NI_2 NS_276 0 8.9095471939097876e-04
GC_2_277 b_2 NI_2 NS_277 0 5.5190051676671750e-05
GC_2_278 b_2 NI_2 NS_278 0 -1.6637660310671270e-05
GC_2_279 b_2 NI_2 NS_279 0 4.4096880984075660e-04
GC_2_280 b_2 NI_2 NS_280 0 -2.0968202350977929e-03
GC_2_281 b_2 NI_2 NS_281 0 -1.8612084073678738e-05
GC_2_282 b_2 NI_2 NS_282 0 -4.8223265365245900e-05
GC_2_283 b_2 NI_2 NS_283 0 4.1823346917757554e-04
GC_2_284 b_2 NI_2 NS_284 0 9.3471779330581737e-06
GC_2_285 b_2 NI_2 NS_285 0 2.4959788696287627e-05
GC_2_286 b_2 NI_2 NS_286 0 4.9544013233657312e-05
GC_2_287 b_2 NI_2 NS_287 0 1.4606028204939783e-05
GC_2_288 b_2 NI_2 NS_288 0 -5.2036211392615490e-05
GC_2_289 b_2 NI_2 NS_289 0 -4.0054349092238765e-05
GC_2_290 b_2 NI_2 NS_290 0 3.5301421247469943e-05
GC_2_291 b_2 NI_2 NS_291 0 1.2943919319335780e-03
GC_2_292 b_2 NI_2 NS_292 0 -2.6457135430012716e-03
GC_2_293 b_2 NI_2 NS_293 0 -3.0503865605488646e-06
GC_2_294 b_2 NI_2 NS_294 0 2.3441240391273414e-05
GC_2_295 b_2 NI_2 NS_295 0 -9.6046850696390848e-04
GC_2_296 b_2 NI_2 NS_296 0 4.3628075600917669e-04
GC_2_297 b_2 NI_2 NS_297 0 -3.6554029444506027e-06
GC_2_298 b_2 NI_2 NS_298 0 2.1266828987161705e-06
GC_2_299 b_2 NI_2 NS_299 0 3.3213154647212064e-04
GC_2_300 b_2 NI_2 NS_300 0 2.8075420755081418e-04
GC_2_301 b_2 NI_2 NS_301 0 1.7568629392998689e-06
GC_2_302 b_2 NI_2 NS_302 0 -4.7935201512217311e-06
GC_2_303 b_2 NI_2 NS_303 0 1.4472919116464806e-06
GC_2_304 b_2 NI_2 NS_304 0 9.2826859779193354e-07
GC_2_305 b_2 NI_2 NS_305 0 -1.2266856703596844e-06
GC_2_306 b_2 NI_2 NS_306 0 -1.4451505815800557e-06
GC_2_307 b_2 NI_2 NS_307 0 -2.2064618497229544e-06
GC_2_308 b_2 NI_2 NS_308 0 -1.2790581526204861e-06
GC_2_309 b_2 NI_2 NS_309 0 8.6673466842748480e-03
GC_2_310 b_2 NI_2 NS_310 0 -2.9984941045278235e-05
GC_2_311 b_2 NI_2 NS_311 0 2.1816743945567685e-03
GC_2_312 b_2 NI_2 NS_312 0 -2.1543335272967120e-03
GC_2_313 b_2 NI_2 NS_313 0 4.7628283030937970e-04
GC_2_314 b_2 NI_2 NS_314 0 2.8951595499750711e-03
GC_2_315 b_2 NI_2 NS_315 0 -6.1397029162077411e-04
GC_2_316 b_2 NI_2 NS_316 0 1.0765340971984046e-03
GC_2_317 b_2 NI_2 NS_317 0 8.2212247299277461e-04
GC_2_318 b_2 NI_2 NS_318 0 5.1234698844731716e-04
GC_2_319 b_2 NI_2 NS_319 0 -7.4259407375248704e-04
GC_2_320 b_2 NI_2 NS_320 0 2.1129567375385199e-03
GC_2_321 b_2 NI_2 NS_321 0 -6.1191759666043996e-05
GC_2_322 b_2 NI_2 NS_322 0 1.4744946931973188e-05
GC_2_323 b_2 NI_2 NS_323 0 -2.2804571884143314e-04
GC_2_324 b_2 NI_2 NS_324 0 6.5316934884589628e-04
GC_2_325 b_2 NI_2 NS_325 0 -1.5995759587598118e-06
GC_2_326 b_2 NI_2 NS_326 0 -1.2931702820064241e-06
GC_2_327 b_2 NI_2 NS_327 0 -2.8228159295444889e-04
GC_2_328 b_2 NI_2 NS_328 0 4.2644225250386192e-04
GC_2_329 b_2 NI_2 NS_329 0 3.8310011441909794e-04
GC_2_330 b_2 NI_2 NS_330 0 -1.1535321345794987e-04
GC_2_331 b_2 NI_2 NS_331 0 -3.4956354085518470e-05
GC_2_332 b_2 NI_2 NS_332 0 1.4524546447094819e-08
GC_2_333 b_2 NI_2 NS_333 0 -3.1199052874815309e-05
GC_2_334 b_2 NI_2 NS_334 0 -5.2999155688372945e-05
GC_2_335 b_2 NI_2 NS_335 0 -3.2585180286899551e-03
GC_2_336 b_2 NI_2 NS_336 0 -2.4625876746099569e-03
GC_2_337 b_2 NI_2 NS_337 0 -1.2474920980920529e-05
GC_2_338 b_2 NI_2 NS_338 0 -2.2356700288472807e-05
GC_2_339 b_2 NI_2 NS_339 0 8.9320177555247211e-04
GC_2_340 b_2 NI_2 NS_340 0 1.1299644971558666e-03
GC_2_341 b_2 NI_2 NS_341 0 -6.0030462614792080e-06
GC_2_342 b_2 NI_2 NS_342 0 1.6306029806294771e-05
GC_2_343 b_2 NI_2 NS_343 0 8.9863476514840594e-04
GC_2_344 b_2 NI_2 NS_344 0 -5.2531439804427758e-04
GC_2_345 b_2 NI_2 NS_345 0 -1.6778739698919485e-05
GC_2_346 b_2 NI_2 NS_346 0 -1.4778186089422897e-05
GC_2_347 b_2 NI_2 NS_347 0 1.8946097026053893e-05
GC_2_348 b_2 NI_2 NS_348 0 -2.7209500094450393e-06
GC_2_349 b_2 NI_2 NS_349 0 1.9862635422973987e-05
GC_2_350 b_2 NI_2 NS_350 0 -1.9588298806423391e-06
GC_2_351 b_2 NI_2 NS_351 0 9.0585069224960061e-05
GC_2_352 b_2 NI_2 NS_352 0 7.8226262058151502e-06
GC_2_353 b_2 NI_2 NS_353 0 1.0870601563714907e-02
GC_2_354 b_2 NI_2 NS_354 0 1.2683920774152757e-05
GC_2_355 b_2 NI_2 NS_355 0 5.2885786626707009e-05
GC_2_356 b_2 NI_2 NS_356 0 1.1568908028762091e-04
GC_2_357 b_2 NI_2 NS_357 0 -1.5750037883532954e-04
GC_2_358 b_2 NI_2 NS_358 0 -4.0872092965699806e-05
GC_2_359 b_2 NI_2 NS_359 0 -4.8227685775480139e-04
GC_2_360 b_2 NI_2 NS_360 0 4.6562153168842036e-05
GC_2_361 b_2 NI_2 NS_361 0 1.8156450060305917e-04
GC_2_362 b_2 NI_2 NS_362 0 -2.7879076984466518e-04
GC_2_363 b_2 NI_2 NS_363 0 9.2224055981692573e-04
GC_2_364 b_2 NI_2 NS_364 0 8.0881795339263850e-05
GC_2_365 b_2 NI_2 NS_365 0 8.6181904774627893e-05
GC_2_366 b_2 NI_2 NS_366 0 6.4647132228726252e-05
GC_2_367 b_2 NI_2 NS_367 0 -2.1132938271754638e-04
GC_2_368 b_2 NI_2 NS_368 0 1.6262901390331835e-03
GC_2_369 b_2 NI_2 NS_369 0 -1.3064987932619060e-04
GC_2_370 b_2 NI_2 NS_370 0 6.0058879274983234e-05
GC_2_371 b_2 NI_2 NS_371 0 -5.6746966413376016e-04
GC_2_372 b_2 NI_2 NS_372 0 -1.3590971366137119e-04
GC_2_373 b_2 NI_2 NS_373 0 4.7008698406114655e-06
GC_2_374 b_2 NI_2 NS_374 0 -9.8943493808445473e-05
GC_2_375 b_2 NI_2 NS_375 0 -3.1885075065227977e-05
GC_2_376 b_2 NI_2 NS_376 0 -1.0495393744103823e-04
GC_2_377 b_2 NI_2 NS_377 0 -3.1288021049432834e-06
GC_2_378 b_2 NI_2 NS_378 0 9.4842169186961259e-05
GC_2_379 b_2 NI_2 NS_379 0 6.0029511818771546e-05
GC_2_380 b_2 NI_2 NS_380 0 3.8375889880457980e-04
GC_2_381 b_2 NI_2 NS_381 0 -2.2343874718889361e-05
GC_2_382 b_2 NI_2 NS_382 0 -1.1997769890331521e-05
GC_2_383 b_2 NI_2 NS_383 0 -2.2102137088552426e-04
GC_2_384 b_2 NI_2 NS_384 0 -1.8404117036573196e-04
GC_2_385 b_2 NI_2 NS_385 0 4.5603143309998562e-07
GC_2_386 b_2 NI_2 NS_386 0 2.4999756912231468e-06
GC_2_387 b_2 NI_2 NS_387 0 -6.2589325104402105e-05
GC_2_388 b_2 NI_2 NS_388 0 -2.4324721598342037e-04
GC_2_389 b_2 NI_2 NS_389 0 -1.0946832818777369e-05
GC_2_390 b_2 NI_2 NS_390 0 -1.6208402772433096e-05
GC_2_391 b_2 NI_2 NS_391 0 -2.3535191890995672e-07
GC_2_392 b_2 NI_2 NS_392 0 1.2084763953029411e-06
GC_2_393 b_2 NI_2 NS_393 0 -4.9809921931546235e-07
GC_2_394 b_2 NI_2 NS_394 0 -1.3863858257978143e-06
GC_2_395 b_2 NI_2 NS_395 0 -2.1116633730242554e-04
GC_2_396 b_2 NI_2 NS_396 0 -4.4890192148491981e-05
GC_2_397 b_2 NI_2 NS_397 0 3.1392042271330082e-03
GC_2_398 b_2 NI_2 NS_398 0 -1.4727048154883592e-05
GC_2_399 b_2 NI_2 NS_399 0 -1.1665231639286008e-04
GC_2_400 b_2 NI_2 NS_400 0 -1.2814012631517493e-04
GC_2_401 b_2 NI_2 NS_401 0 1.4448570205746722e-04
GC_2_402 b_2 NI_2 NS_402 0 -1.4445975474241816e-04
GC_2_403 b_2 NI_2 NS_403 0 -3.9538377910831261e-04
GC_2_404 b_2 NI_2 NS_404 0 -2.4173288853534340e-04
GC_2_405 b_2 NI_2 NS_405 0 7.3811167201124028e-05
GC_2_406 b_2 NI_2 NS_406 0 -2.2448948768474908e-04
GC_2_407 b_2 NI_2 NS_407 0 4.2540236479495397e-04
GC_2_408 b_2 NI_2 NS_408 0 -3.9300490848393843e-04
GC_2_409 b_2 NI_2 NS_409 0 1.4198989477816041e-05
GC_2_410 b_2 NI_2 NS_410 0 1.9463010675101719e-05
GC_2_411 b_2 NI_2 NS_411 0 5.4659502947640480e-04
GC_2_412 b_2 NI_2 NS_412 0 -1.8602978415976833e-04
GC_2_413 b_2 NI_2 NS_413 0 1.3269887275672601e-05
GC_2_414 b_2 NI_2 NS_414 0 -4.7731187553006411e-05
GC_2_415 b_2 NI_2 NS_415 0 6.8516055778878020e-04
GC_2_416 b_2 NI_2 NS_416 0 -2.9954464364919872e-04
GC_2_417 b_2 NI_2 NS_417 0 -2.9310255715611302e-04
GC_2_418 b_2 NI_2 NS_418 0 -3.4750843297431450e-04
GC_2_419 b_2 NI_2 NS_419 0 9.3111115450827301e-06
GC_2_420 b_2 NI_2 NS_420 0 -2.3233505323610497e-05
GC_2_421 b_2 NI_2 NS_421 0 -4.3855666995742667e-05
GC_2_422 b_2 NI_2 NS_422 0 -1.5810115206186729e-04
GC_2_423 b_2 NI_2 NS_423 0 -3.9515666256355391e-03
GC_2_424 b_2 NI_2 NS_424 0 4.6472531506230458e-03
GC_2_425 b_2 NI_2 NS_425 0 2.0019926850336466e-05
GC_2_426 b_2 NI_2 NS_426 0 2.0213601388572663e-05
GC_2_427 b_2 NI_2 NS_427 0 3.3768989065631832e-03
GC_2_428 b_2 NI_2 NS_428 0 -1.3815276327076335e-03
GC_2_429 b_2 NI_2 NS_429 0 2.2583083982773844e-05
GC_2_430 b_2 NI_2 NS_430 0 9.3600499649308565e-07
GC_2_431 b_2 NI_2 NS_431 0 -4.3990879309831020e-04
GC_2_432 b_2 NI_2 NS_432 0 -3.0573733420169051e-04
GC_2_433 b_2 NI_2 NS_433 0 -5.3083223841606214e-05
GC_2_434 b_2 NI_2 NS_434 0 1.0412448028675841e-05
GC_2_435 b_2 NI_2 NS_435 0 2.8754363054836546e-05
GC_2_436 b_2 NI_2 NS_436 0 -6.5451805270149169e-06
GC_2_437 b_2 NI_2 NS_437 0 -2.2397670208464243e-05
GC_2_438 b_2 NI_2 NS_438 0 1.6570121379780317e-05
GC_2_439 b_2 NI_2 NS_439 0 4.1369151991612084e-04
GC_2_440 b_2 NI_2 NS_440 0 1.6392327745152528e-04
GC_2_441 b_2 NI_2 NS_441 0 1.5906152990694398e-02
GC_2_442 b_2 NI_2 NS_442 0 -4.0320958787586285e-05
GC_2_443 b_2 NI_2 NS_443 0 -1.3164639886855339e-04
GC_2_444 b_2 NI_2 NS_444 0 5.5101531540962829e-04
GC_2_445 b_2 NI_2 NS_445 0 -4.9856300340315183e-04
GC_2_446 b_2 NI_2 NS_446 0 -2.2826786249437468e-04
GC_2_447 b_2 NI_2 NS_447 0 -2.8765696167797555e-04
GC_2_448 b_2 NI_2 NS_448 0 -2.4519609639307141e-04
GC_2_449 b_2 NI_2 NS_449 0 3.1290750932164949e-04
GC_2_450 b_2 NI_2 NS_450 0 -3.7855692011843651e-05
GC_2_451 b_2 NI_2 NS_451 0 -2.9433566055447858e-04
GC_2_452 b_2 NI_2 NS_452 0 1.1003663910515344e-03
GC_2_453 b_2 NI_2 NS_453 0 6.2766487938688791e-05
GC_2_454 b_2 NI_2 NS_454 0 2.4802187765279457e-05
GC_2_455 b_2 NI_2 NS_455 0 -8.8249458765867405e-04
GC_2_456 b_2 NI_2 NS_456 0 3.7653877625063727e-04
GC_2_457 b_2 NI_2 NS_457 0 -9.2341021478101919e-05
GC_2_458 b_2 NI_2 NS_458 0 2.0573036701235263e-05
GC_2_459 b_2 NI_2 NS_459 0 -3.9481746081860712e-04
GC_2_460 b_2 NI_2 NS_460 0 -1.7241590939246908e-04
GC_2_461 b_2 NI_2 NS_461 0 2.6955932893908707e-05
GC_2_462 b_2 NI_2 NS_462 0 -7.4548020936684181e-05
GC_2_463 b_2 NI_2 NS_463 0 -2.3087067414931348e-05
GC_2_464 b_2 NI_2 NS_464 0 -8.4196444768609032e-05
GC_2_465 b_2 NI_2 NS_465 0 -2.3650398469970587e-05
GC_2_466 b_2 NI_2 NS_466 0 6.6120774689864935e-05
GC_2_467 b_2 NI_2 NS_467 0 -9.0195343951839530e-05
GC_2_468 b_2 NI_2 NS_468 0 -6.9243516557707444e-04
GC_2_469 b_2 NI_2 NS_469 0 -1.2485816604892127e-05
GC_2_470 b_2 NI_2 NS_470 0 -4.1085535298028477e-06
GC_2_471 b_2 NI_2 NS_471 0 -3.9465721507362587e-04
GC_2_472 b_2 NI_2 NS_472 0 -3.0741204985492321e-05
GC_2_473 b_2 NI_2 NS_473 0 -1.3312791493469533e-06
GC_2_474 b_2 NI_2 NS_474 0 4.3627742556709074e-07
GC_2_475 b_2 NI_2 NS_475 0 1.6509918591009427e-04
GC_2_476 b_2 NI_2 NS_476 0 -9.4789060458620901e-05
GC_2_477 b_2 NI_2 NS_477 0 -6.6463075016063377e-06
GC_2_478 b_2 NI_2 NS_478 0 -1.1071355173283538e-05
GC_2_479 b_2 NI_2 NS_479 0 7.2949670909183096e-07
GC_2_480 b_2 NI_2 NS_480 0 -8.3041486990541921e-07
GC_2_481 b_2 NI_2 NS_481 0 -2.1488601104114804e-07
GC_2_482 b_2 NI_2 NS_482 0 6.2332904529867857e-07
GC_2_483 b_2 NI_2 NS_483 0 -9.0268000834495108e-05
GC_2_484 b_2 NI_2 NS_484 0 -4.7819389246511390e-05
GC_2_485 b_2 NI_2 NS_485 0 3.5220261804268921e-04
GC_2_486 b_2 NI_2 NS_486 0 -8.7579771939140887e-07
GC_2_487 b_2 NI_2 NS_487 0 2.2948473626658778e-05
GC_2_488 b_2 NI_2 NS_488 0 -4.6155101834811750e-04
GC_2_489 b_2 NI_2 NS_489 0 4.6433028186834441e-04
GC_2_490 b_2 NI_2 NS_490 0 1.2267897826735745e-04
GC_2_491 b_2 NI_2 NS_491 0 -1.0891672109593519e-04
GC_2_492 b_2 NI_2 NS_492 0 4.1163610800533227e-04
GC_2_493 b_2 NI_2 NS_493 0 2.6657530170351559e-04
GC_2_494 b_2 NI_2 NS_494 0 -8.3139522777805940e-05
GC_2_495 b_2 NI_2 NS_495 0 3.1627686206168434e-04
GC_2_496 b_2 NI_2 NS_496 0 2.9248871819290834e-04
GC_2_497 b_2 NI_2 NS_497 0 6.4677128968528039e-06
GC_2_498 b_2 NI_2 NS_498 0 8.6588215472158032e-06
GC_2_499 b_2 NI_2 NS_499 0 7.4413225126459040e-05
GC_2_500 b_2 NI_2 NS_500 0 -2.1320762985365413e-04
GC_2_501 b_2 NI_2 NS_501 0 1.1842537556931905e-05
GC_2_502 b_2 NI_2 NS_502 0 -2.6766013678128197e-05
GC_2_503 b_2 NI_2 NS_503 0 3.7253633749375156e-04
GC_2_504 b_2 NI_2 NS_504 0 -1.5572727544771974e-04
GC_2_505 b_2 NI_2 NS_505 0 -7.4389146665418385e-05
GC_2_506 b_2 NI_2 NS_506 0 -1.3788867617316509e-04
GC_2_507 b_2 NI_2 NS_507 0 3.4360858482206164e-06
GC_2_508 b_2 NI_2 NS_508 0 -1.3216125935904048e-05
GC_2_509 b_2 NI_2 NS_509 0 -2.5993779587109962e-05
GC_2_510 b_2 NI_2 NS_510 0 -9.7663551509354478e-05
GC_2_511 b_2 NI_2 NS_511 0 -2.1904077919706901e-03
GC_2_512 b_2 NI_2 NS_512 0 2.0228372329643609e-03
GC_2_513 b_2 NI_2 NS_513 0 7.2443997936740680e-06
GC_2_514 b_2 NI_2 NS_514 0 4.9913088758708821e-06
GC_2_515 b_2 NI_2 NS_515 0 1.8971031711093041e-03
GC_2_516 b_2 NI_2 NS_516 0 -5.9841340003978461e-04
GC_2_517 b_2 NI_2 NS_517 0 7.5215563614554383e-06
GC_2_518 b_2 NI_2 NS_518 0 2.6488480219568198e-06
GC_2_519 b_2 NI_2 NS_519 0 -6.5665550047507896e-05
GC_2_520 b_2 NI_2 NS_520 0 -1.6379777743826909e-04
GC_2_521 b_2 NI_2 NS_521 0 -2.3493216193444779e-05
GC_2_522 b_2 NI_2 NS_522 0 1.7814404444711093e-07
GC_2_523 b_2 NI_2 NS_523 0 1.7964554907164197e-05
GC_2_524 b_2 NI_2 NS_524 0 -1.4685968394562758e-06
GC_2_525 b_2 NI_2 NS_525 0 -9.4303416140760345e-06
GC_2_526 b_2 NI_2 NS_526 0 5.6555931641704060e-06
GC_2_527 b_2 NI_2 NS_527 0 1.9716278086594541e-04
GC_2_528 b_2 NI_2 NS_528 0 9.8075526295261209e-05
GD_2_1 b_2 NI_2 NA_1 0 -4.2054647074284985e-03
GD_2_2 b_2 NI_2 NA_2 0 2.6541420089927270e-01
GD_2_3 b_2 NI_2 NA_3 0 -6.4005299132231325e-02
GD_2_4 b_2 NI_2 NA_4 0 -1.5790005140188620e-02
GD_2_5 b_2 NI_2 NA_5 0 -3.8919846984812934e-02
GD_2_6 b_2 NI_2 NA_6 0 -1.9402984504259455e-02
GD_2_7 b_2 NI_2 NA_7 0 -1.9300869900889587e-02
GD_2_8 b_2 NI_2 NA_8 0 -1.1805446344193763e-02
GD_2_9 b_2 NI_2 NA_9 0 -1.1751497739138013e-02
GD_2_10 b_2 NI_2 NA_10 0 -4.5743763923083046e-03
GD_2_11 b_2 NI_2 NA_11 0 -1.4025804121709841e-02
GD_2_12 b_2 NI_2 NA_12 0 -2.9557136715318458e-03
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+01
GC_3_1 b_3 NI_3 NS_1 0 1.6697373826330768e-03
GC_3_2 b_3 NI_3 NS_2 0 -5.0120088912037097e-05
GC_3_3 b_3 NI_3 NS_3 0 5.0844969784566447e-03
GC_3_4 b_3 NI_3 NS_4 0 4.8276131716655356e-03
GC_3_5 b_3 NI_3 NS_5 0 -5.5576302553340812e-03
GC_3_6 b_3 NI_3 NS_6 0 -4.8354387994992021e-03
GC_3_7 b_3 NI_3 NS_7 0 -3.1164530487497383e-04
GC_3_8 b_3 NI_3 NS_8 0 2.5189387947428083e-04
GC_3_9 b_3 NI_3 NS_9 0 1.4815451306979149e-03
GC_3_10 b_3 NI_3 NS_10 0 5.4309255497730713e-03
GC_3_11 b_3 NI_3 NS_11 0 -3.0290115909591179e-03
GC_3_12 b_3 NI_3 NS_12 0 -1.0501070388557708e-03
GC_3_13 b_3 NI_3 NS_13 0 8.7340228413658168e-04
GC_3_14 b_3 NI_3 NS_14 0 2.8128318090735459e-04
GC_3_15 b_3 NI_3 NS_15 0 -5.4787229087480786e-03
GC_3_16 b_3 NI_3 NS_16 0 -2.2171752964961424e-03
GC_3_17 b_3 NI_3 NS_17 0 -1.0992863610316397e-04
GC_3_18 b_3 NI_3 NS_18 0 9.7725631754450650e-05
GC_3_19 b_3 NI_3 NS_19 0 -1.9544070005312717e-03
GC_3_20 b_3 NI_3 NS_20 0 -3.2931014996272863e-03
GC_3_21 b_3 NI_3 NS_21 0 -2.1733802052923635e-04
GC_3_22 b_3 NI_3 NS_22 0 4.2382574285442268e-04
GC_3_23 b_3 NI_3 NS_23 0 1.6775058784348836e-04
GC_3_24 b_3 NI_3 NS_24 0 -6.0504504547231125e-05
GC_3_25 b_3 NI_3 NS_25 0 1.2085079696477738e-05
GC_3_26 b_3 NI_3 NS_26 0 -1.1186492330023307e-04
GC_3_27 b_3 NI_3 NS_27 0 7.2947654499706683e-03
GC_3_28 b_3 NI_3 NS_28 0 2.0806936950625186e-03
GC_3_29 b_3 NI_3 NS_29 0 -1.4267197435995281e-05
GC_3_30 b_3 NI_3 NS_30 0 -9.5877947844583292e-06
GC_3_31 b_3 NI_3 NS_31 0 6.7126821568138924e-04
GC_3_32 b_3 NI_3 NS_32 0 -3.8047555248101454e-03
GC_3_33 b_3 NI_3 NS_33 0 5.2078305872094003e-07
GC_3_34 b_3 NI_3 NS_34 0 -1.1131565178775968e-05
GC_3_35 b_3 NI_3 NS_35 0 8.3907073816453159e-04
GC_3_36 b_3 NI_3 NS_36 0 1.1031860660603654e-03
GC_3_37 b_3 NI_3 NS_37 0 1.5777727548355984e-05
GC_3_38 b_3 NI_3 NS_38 0 9.4458341126459036e-06
GC_3_39 b_3 NI_3 NS_39 0 8.1870872074220420e-08
GC_3_40 b_3 NI_3 NS_40 0 4.9826430716133226e-06
GC_3_41 b_3 NI_3 NS_41 0 -1.6793242355999360e-06
GC_3_42 b_3 NI_3 NS_42 0 -3.2297986056757899e-06
GC_3_43 b_3 NI_3 NS_43 0 2.1471902435505831e-05
GC_3_44 b_3 NI_3 NS_44 0 1.4413908648412140e-04
GC_3_45 b_3 NI_3 NS_45 0 5.8822982995212207e-02
GC_3_46 b_3 NI_3 NS_46 0 -2.0743972462068616e-05
GC_3_47 b_3 NI_3 NS_47 0 -6.4253479494493018e-03
GC_3_48 b_3 NI_3 NS_48 0 -2.9556840751187212e-03
GC_3_49 b_3 NI_3 NS_49 0 4.8501814026438829e-03
GC_3_50 b_3 NI_3 NS_50 0 2.5544219367301135e-03
GC_3_51 b_3 NI_3 NS_51 0 -1.1777984058970646e-04
GC_3_52 b_3 NI_3 NS_52 0 -1.0482802453540824e-04
GC_3_53 b_3 NI_3 NS_53 0 1.6246303186001074e-03
GC_3_54 b_3 NI_3 NS_54 0 1.6016138331904220e-03
GC_3_55 b_3 NI_3 NS_55 0 -3.1790549529455922e-04
GC_3_56 b_3 NI_3 NS_56 0 -7.7117063494307279e-04
GC_3_57 b_3 NI_3 NS_57 0 -2.6956419858134053e-05
GC_3_58 b_3 NI_3 NS_58 0 6.6565596269392189e-05
GC_3_59 b_3 NI_3 NS_59 0 -3.2915211792845403e-03
GC_3_60 b_3 NI_3 NS_60 0 1.1532590939654314e-03
GC_3_61 b_3 NI_3 NS_61 0 -4.8040738322351669e-05
GC_3_62 b_3 NI_3 NS_62 0 -7.1932092233284936e-05
GC_3_63 b_3 NI_3 NS_63 0 7.8901572536778399e-05
GC_3_64 b_3 NI_3 NS_64 0 1.1148674095655673e-03
GC_3_65 b_3 NI_3 NS_65 0 3.2507030982101141e-04
GC_3_66 b_3 NI_3 NS_66 0 6.9320459517763583e-05
GC_3_67 b_3 NI_3 NS_67 0 -2.1473022754481272e-05
GC_3_68 b_3 NI_3 NS_68 0 -2.3815535508117540e-05
GC_3_69 b_3 NI_3 NS_69 0 -4.9121302113917501e-05
GC_3_70 b_3 NI_3 NS_70 0 6.9075315042488758e-05
GC_3_71 b_3 NI_3 NS_71 0 -3.8810926574099659e-03
GC_3_72 b_3 NI_3 NS_72 0 -3.5079993593994854e-03
GC_3_73 b_3 NI_3 NS_73 0 1.4624435923628045e-05
GC_3_74 b_3 NI_3 NS_74 0 3.8510511263810099e-05
GC_3_75 b_3 NI_3 NS_75 0 -2.5984647515243795e-04
GC_3_76 b_3 NI_3 NS_76 0 2.3947784809197196e-03
GC_3_77 b_3 NI_3 NS_77 0 2.0090779382554700e-06
GC_3_78 b_3 NI_3 NS_78 0 9.9947949831887517e-06
GC_3_79 b_3 NI_3 NS_79 0 9.0676155296782991e-04
GC_3_80 b_3 NI_3 NS_80 0 -5.4484277567099317e-04
GC_3_81 b_3 NI_3 NS_81 0 -1.1759195876801402e-05
GC_3_82 b_3 NI_3 NS_82 0 -5.0239537974276268e-06
GC_3_83 b_3 NI_3 NS_83 0 2.0059892901133951e-06
GC_3_84 b_3 NI_3 NS_84 0 -1.7978369559478067e-06
GC_3_85 b_3 NI_3 NS_85 0 2.4366121630486865e-06
GC_3_86 b_3 NI_3 NS_86 0 -4.5690841956521753e-07
GC_3_87 b_3 NI_3 NS_87 0 1.4765342013792183e-04
GC_3_88 b_3 NI_3 NS_88 0 -1.5970040652347155e-04
GC_3_89 b_3 NI_3 NS_89 0 -2.7813104327690644e-02
GC_3_90 b_3 NI_3 NS_90 0 9.6538579712003372e-03
GC_3_91 b_3 NI_3 NS_91 0 7.8752686850444079e-03
GC_3_92 b_3 NI_3 NS_92 0 6.1519676468109394e-03
GC_3_93 b_3 NI_3 NS_93 0 8.2829979337408748e-03
GC_3_94 b_3 NI_3 NS_94 0 2.0449185388556881e-03
GC_3_95 b_3 NI_3 NS_95 0 7.1053369598405138e-04
GC_3_96 b_3 NI_3 NS_96 0 2.0741246033059404e-04
GC_3_97 b_3 NI_3 NS_97 0 1.1023432736495730e-03
GC_3_98 b_3 NI_3 NS_98 0 7.9110017201479699e-03
GC_3_99 b_3 NI_3 NS_99 0 -6.8340661601968304e-03
GC_3_100 b_3 NI_3 NS_100 0 1.0647814635740495e-03
GC_3_101 b_3 NI_3 NS_101 0 1.1189789758399645e-03
GC_3_102 b_3 NI_3 NS_102 0 4.4758910855571197e-04
GC_3_103 b_3 NI_3 NS_103 0 5.0354480370335165e-03
GC_3_104 b_3 NI_3 NS_104 0 2.4688826113652270e-03
GC_3_105 b_3 NI_3 NS_105 0 -1.4970618927056880e-04
GC_3_106 b_3 NI_3 NS_106 0 1.8229105698711436e-04
GC_3_107 b_3 NI_3 NS_107 0 -1.9258006899604174e-03
GC_3_108 b_3 NI_3 NS_108 0 -4.0632535310363331e-03
GC_3_109 b_3 NI_3 NS_109 0 -1.1839145718317754e-03
GC_3_110 b_3 NI_3 NS_110 0 8.4206522190378118e-04
GC_3_111 b_3 NI_3 NS_111 0 2.4353562312994033e-04
GC_3_112 b_3 NI_3 NS_112 0 -6.5159242668895006e-05
GC_3_113 b_3 NI_3 NS_113 0 3.1437609174515116e-05
GC_3_114 b_3 NI_3 NS_114 0 -1.3396086425438114e-04
GC_3_115 b_3 NI_3 NS_115 0 4.5083017075787137e-03
GC_3_116 b_3 NI_3 NS_116 0 1.0673757271343280e-02
GC_3_117 b_3 NI_3 NS_117 0 -1.4503006225397461e-05
GC_3_118 b_3 NI_3 NS_118 0 -1.7258518224225833e-05
GC_3_119 b_3 NI_3 NS_119 0 2.7877448746857964e-03
GC_3_120 b_3 NI_3 NS_120 0 -5.6236496332293271e-03
GC_3_121 b_3 NI_3 NS_121 0 2.3030820530859464e-06
GC_3_122 b_3 NI_3 NS_122 0 -2.7756264012735332e-05
GC_3_123 b_3 NI_3 NS_123 0 -1.1520329115536081e-03
GC_3_124 b_3 NI_3 NS_124 0 1.5921083575454499e-03
GC_3_125 b_3 NI_3 NS_125 0 2.9159028741754128e-05
GC_3_126 b_3 NI_3 NS_126 0 3.4968342871342105e-05
GC_3_127 b_3 NI_3 NS_127 0 -4.7168380153889548e-06
GC_3_128 b_3 NI_3 NS_128 0 7.7073176631086566e-06
GC_3_129 b_3 NI_3 NS_129 0 -1.7510130353752674e-06
GC_3_130 b_3 NI_3 NS_130 0 -1.2625622834726441e-05
GC_3_131 b_3 NI_3 NS_131 0 -2.4484793536580588e-04
GC_3_132 b_3 NI_3 NS_132 0 3.0458847943203702e-05
GC_3_133 b_3 NI_3 NS_133 0 3.5592756495924686e-02
GC_3_134 b_3 NI_3 NS_134 0 1.0566342780604204e-02
GC_3_135 b_3 NI_3 NS_135 0 -1.0030245333905813e-02
GC_3_136 b_3 NI_3 NS_136 0 -3.9402786534513158e-03
GC_3_137 b_3 NI_3 NS_137 0 -9.6876630065494632e-03
GC_3_138 b_3 NI_3 NS_138 0 -1.5121362878166415e-03
GC_3_139 b_3 NI_3 NS_139 0 1.0311872853682791e-04
GC_3_140 b_3 NI_3 NS_140 0 1.2871602691894745e-04
GC_3_141 b_3 NI_3 NS_141 0 3.1272239934004207e-03
GC_3_142 b_3 NI_3 NS_142 0 2.8101416701915450e-03
GC_3_143 b_3 NI_3 NS_143 0 -2.3553740039813534e-05
GC_3_144 b_3 NI_3 NS_144 0 -1.3694868968736173e-03
GC_3_145 b_3 NI_3 NS_145 0 -3.0695225980546811e-06
GC_3_146 b_3 NI_3 NS_146 0 2.1713712331328271e-04
GC_3_147 b_3 NI_3 NS_147 0 3.8553268809377044e-03
GC_3_148 b_3 NI_3 NS_148 0 -6.7826699451358603e-04
GC_3_149 b_3 NI_3 NS_149 0 -2.0010021924324542e-05
GC_3_150 b_3 NI_3 NS_150 0 -3.8245690479485515e-05
GC_3_151 b_3 NI_3 NS_151 0 9.2898787957249496e-04
GC_3_152 b_3 NI_3 NS_152 0 8.1451531256195400e-04
GC_3_153 b_3 NI_3 NS_153 0 1.0575758960818454e-04
GC_3_154 b_3 NI_3 NS_154 0 -3.4831406201477441e-04
GC_3_155 b_3 NI_3 NS_155 0 1.9680245504233894e-05
GC_3_156 b_3 NI_3 NS_156 0 -1.2167884847204299e-05
GC_3_157 b_3 NI_3 NS_157 0 -3.1699702503668995e-05
GC_3_158 b_3 NI_3 NS_158 0 6.2682040356698012e-05
GC_3_159 b_3 NI_3 NS_159 0 -3.7150273355134908e-03
GC_3_160 b_3 NI_3 NS_160 0 -8.4011822875825523e-04
GC_3_161 b_3 NI_3 NS_161 0 1.2136870851590749e-05
GC_3_162 b_3 NI_3 NS_162 0 3.1614162040219620e-05
GC_3_163 b_3 NI_3 NS_163 0 3.2005310122932017e-04
GC_3_164 b_3 NI_3 NS_164 0 1.4242989290049887e-03
GC_3_165 b_3 NI_3 NS_165 0 7.8628303361070483e-06
GC_3_166 b_3 NI_3 NS_166 0 1.1551604587429456e-06
GC_3_167 b_3 NI_3 NS_167 0 4.2314713160320845e-06
GC_3_168 b_3 NI_3 NS_168 0 -9.4246059433054767e-04
GC_3_169 b_3 NI_3 NS_169 0 -7.4444313934079905e-06
GC_3_170 b_3 NI_3 NS_170 0 8.3986347871685795e-06
GC_3_171 b_3 NI_3 NS_171 0 -6.2998892640875551e-07
GC_3_172 b_3 NI_3 NS_172 0 -1.1435436800126161e-06
GC_3_173 b_3 NI_3 NS_173 0 2.3364262781697297e-06
GC_3_174 b_3 NI_3 NS_174 0 -4.2027290172871308e-06
GC_3_175 b_3 NI_3 NS_175 0 1.4553374968741205e-05
GC_3_176 b_3 NI_3 NS_176 0 -2.0877287916715965e-04
GC_3_177 b_3 NI_3 NS_177 0 2.6042158902624879e-03
GC_3_178 b_3 NI_3 NS_178 0 8.9383988543734509e-05
GC_3_179 b_3 NI_3 NS_179 0 7.3168842305533603e-03
GC_3_180 b_3 NI_3 NS_180 0 3.7799779023695132e-03
GC_3_181 b_3 NI_3 NS_181 0 -5.6738793868173010e-03
GC_3_182 b_3 NI_3 NS_182 0 -2.2607660269795102e-03
GC_3_183 b_3 NI_3 NS_183 0 -5.6491115080521667e-06
GC_3_184 b_3 NI_3 NS_184 0 3.1195551145224009e-04
GC_3_185 b_3 NI_3 NS_185 0 2.1334644263346432e-03
GC_3_186 b_3 NI_3 NS_186 0 8.2163653387993512e-03
GC_3_187 b_3 NI_3 NS_187 0 -1.0559431133147267e-02
GC_3_188 b_3 NI_3 NS_188 0 -1.3285589993006759e-03
GC_3_189 b_3 NI_3 NS_189 0 1.2038340771644478e-03
GC_3_190 b_3 NI_3 NS_190 0 3.3587979404143934e-04
GC_3_191 b_3 NI_3 NS_191 0 -3.1080656924231623e-03
GC_3_192 b_3 NI_3 NS_192 0 -3.7438129827699683e-03
GC_3_193 b_3 NI_3 NS_193 0 -1.0879779738903608e-04
GC_3_194 b_3 NI_3 NS_194 0 1.6956704232885464e-04
GC_3_195 b_3 NI_3 NS_195 0 -2.8483499053675448e-03
GC_3_196 b_3 NI_3 NS_196 0 -4.7724640016720424e-03
GC_3_197 b_3 NI_3 NS_197 0 -2.0528968081745216e-04
GC_3_198 b_3 NI_3 NS_198 0 1.3525004221957610e-03
GC_3_199 b_3 NI_3 NS_199 0 2.3453680791593964e-04
GC_3_200 b_3 NI_3 NS_200 0 -1.0747945072964575e-04
GC_3_201 b_3 NI_3 NS_201 0 3.5790555302533272e-06
GC_3_202 b_3 NI_3 NS_202 0 -1.3549743493972654e-04
GC_3_203 b_3 NI_3 NS_203 0 9.4726475675990605e-03
GC_3_204 b_3 NI_3 NS_204 0 -4.0329155887249333e-04
GC_3_205 b_3 NI_3 NS_205 0 -1.8693687614625173e-05
GC_3_206 b_3 NI_3 NS_206 0 -7.4224207518019258e-06
GC_3_207 b_3 NI_3 NS_207 0 -2.5277859540045132e-04
GC_3_208 b_3 NI_3 NS_208 0 -4.4868851112336416e-03
GC_3_209 b_3 NI_3 NS_209 0 -9.9295665740361995e-06
GC_3_210 b_3 NI_3 NS_210 0 -1.0716933609802776e-05
GC_3_211 b_3 NI_3 NS_211 0 2.0753773614150240e-03
GC_3_212 b_3 NI_3 NS_212 0 2.4612096181939077e-03
GC_3_213 b_3 NI_3 NS_213 0 2.4869002602177156e-05
GC_3_214 b_3 NI_3 NS_214 0 -4.5088540072844606e-06
GC_3_215 b_3 NI_3 NS_215 0 4.0935831709417132e-06
GC_3_216 b_3 NI_3 NS_216 0 6.6436021457229467e-06
GC_3_217 b_3 NI_3 NS_217 0 -4.0065427052048209e-06
GC_3_218 b_3 NI_3 NS_218 0 1.5010664251672653e-06
GC_3_219 b_3 NI_3 NS_219 0 1.6970189879687942e-04
GC_3_220 b_3 NI_3 NS_220 0 2.9856672132072825e-04
GC_3_221 b_3 NI_3 NS_221 0 8.1634989490941307e-02
GC_3_222 b_3 NI_3 NS_222 0 -1.7855520853916228e-04
GC_3_223 b_3 NI_3 NS_223 0 -8.1217039939237463e-03
GC_3_224 b_3 NI_3 NS_224 0 -1.4130427044683716e-03
GC_3_225 b_3 NI_3 NS_225 0 4.3646354926537966e-03
GC_3_226 b_3 NI_3 NS_226 0 7.2119099465149422e-04
GC_3_227 b_3 NI_3 NS_227 0 -1.8113522897682797e-04
GC_3_228 b_3 NI_3 NS_228 0 -1.6145934146914276e-04
GC_3_229 b_3 NI_3 NS_229 0 2.5751373574904590e-03
GC_3_230 b_3 NI_3 NS_230 0 2.0530627791780611e-03
GC_3_231 b_3 NI_3 NS_231 0 -3.6491066352081943e-03
GC_3_232 b_3 NI_3 NS_232 0 7.0375492097906426e-05
GC_3_233 b_3 NI_3 NS_233 0 2.6301012027688776e-06
GC_3_234 b_3 NI_3 NS_234 0 8.5417228931486031e-05
GC_3_235 b_3 NI_3 NS_235 0 -2.8536830700692452e-03
GC_3_236 b_3 NI_3 NS_236 0 -4.3976365258547668e-04
GC_3_237 b_3 NI_3 NS_237 0 -7.1372657817288482e-05
GC_3_238 b_3 NI_3 NS_238 0 -9.3882816997135343e-05
GC_3_239 b_3 NI_3 NS_239 0 3.2933766667055618e-04
GC_3_240 b_3 NI_3 NS_240 0 1.1937540403010925e-03
GC_3_241 b_3 NI_3 NS_241 0 2.9779979147040550e-04
GC_3_242 b_3 NI_3 NS_242 0 6.9897393722915394e-05
GC_3_243 b_3 NI_3 NS_243 0 -1.0138278241485231e-05
GC_3_244 b_3 NI_3 NS_244 0 -5.8810761897973491e-05
GC_3_245 b_3 NI_3 NS_245 0 -7.3616762330699443e-05
GC_3_246 b_3 NI_3 NS_246 0 9.6077852797422030e-05
GC_3_247 b_3 NI_3 NS_247 0 -3.5047392222259687e-03
GC_3_248 b_3 NI_3 NS_248 0 -4.6442490872359533e-03
GC_3_249 b_3 NI_3 NS_249 0 1.5227540024704298e-05
GC_3_250 b_3 NI_3 NS_250 0 5.2820572144558862e-05
GC_3_251 b_3 NI_3 NS_251 0 -6.9522072591016897e-04
GC_3_252 b_3 NI_3 NS_252 0 2.6562085577577855e-03
GC_3_253 b_3 NI_3 NS_253 0 1.6594180220010803e-06
GC_3_254 b_3 NI_3 NS_254 0 1.0312508177949698e-05
GC_3_255 b_3 NI_3 NS_255 0 9.8502296587803261e-04
GC_3_256 b_3 NI_3 NS_256 0 -5.1952539210635483e-04
GC_3_257 b_3 NI_3 NS_257 0 -1.1041367161835178e-05
GC_3_258 b_3 NI_3 NS_258 0 -6.1479352959576096e-06
GC_3_259 b_3 NI_3 NS_259 0 2.4642040319624094e-06
GC_3_260 b_3 NI_3 NS_260 0 -1.0710691391096471e-06
GC_3_261 b_3 NI_3 NS_261 0 1.5538657267531779e-06
GC_3_262 b_3 NI_3 NS_262 0 -1.9821850085522444e-06
GC_3_263 b_3 NI_3 NS_263 0 1.2731390762932539e-04
GC_3_264 b_3 NI_3 NS_264 0 -1.9349184096920674e-04
GC_3_265 b_3 NI_3 NS_265 0 3.6231626107201986e-02
GC_3_266 b_3 NI_3 NS_266 0 1.5138667923376503e-04
GC_3_267 b_3 NI_3 NS_267 0 5.9839007046566016e-03
GC_3_268 b_3 NI_3 NS_268 0 1.2391252333337648e-03
GC_3_269 b_3 NI_3 NS_269 0 -4.2692852410106917e-03
GC_3_270 b_3 NI_3 NS_270 0 2.4099803366221394e-03
GC_3_271 b_3 NI_3 NS_271 0 -1.8580069002237218e-04
GC_3_272 b_3 NI_3 NS_272 0 -8.7100542158822993e-04
GC_3_273 b_3 NI_3 NS_273 0 1.3876197649314605e-03
GC_3_274 b_3 NI_3 NS_274 0 6.0150671935160624e-03
GC_3_275 b_3 NI_3 NS_275 0 -1.0172212263085746e-02
GC_3_276 b_3 NI_3 NS_276 0 -1.3505052452540505e-03
GC_3_277 b_3 NI_3 NS_277 0 9.3708588828209777e-04
GC_3_278 b_3 NI_3 NS_278 0 1.5662942157225061e-04
GC_3_279 b_3 NI_3 NS_279 0 -1.4485518766771486e-03
GC_3_280 b_3 NI_3 NS_280 0 3.5854117444563668e-04
GC_3_281 b_3 NI_3 NS_281 0 -4.7419853035017922e-05
GC_3_282 b_3 NI_3 NS_282 0 1.3954276661550156e-04
GC_3_283 b_3 NI_3 NS_283 0 -1.9605622258669292e-03
GC_3_284 b_3 NI_3 NS_284 0 -3.0129734996712644e-03
GC_3_285 b_3 NI_3 NS_285 0 -9.1329852592065083e-05
GC_3_286 b_3 NI_3 NS_286 0 5.5448636410118169e-04
GC_3_287 b_3 NI_3 NS_287 0 1.5028063213266669e-04
GC_3_288 b_3 NI_3 NS_288 0 -9.0394723586656429e-05
GC_3_289 b_3 NI_3 NS_289 0 -6.3512238781921696e-06
GC_3_290 b_3 NI_3 NS_290 0 -5.3563262496847638e-05
GC_3_291 b_3 NI_3 NS_291 0 1.5528939192375928e-03
GC_3_292 b_3 NI_3 NS_292 0 -1.7847901804861949e-03
GC_3_293 b_3 NI_3 NS_293 0 -5.4102261695552342e-06
GC_3_294 b_3 NI_3 NS_294 0 1.0647019428326802e-07
GC_3_295 b_3 NI_3 NS_295 0 9.8253138908344594e-05
GC_3_296 b_3 NI_3 NS_296 0 -1.9582777913704540e-03
GC_3_297 b_3 NI_3 NS_297 0 3.9378267290370911e-07
GC_3_298 b_3 NI_3 NS_298 0 -4.4113111955376758e-06
GC_3_299 b_3 NI_3 NS_299 0 1.5333070809374751e-03
GC_3_300 b_3 NI_3 NS_300 0 3.4475709704128354e-04
GC_3_301 b_3 NI_3 NS_301 0 2.5739790550274864e-06
GC_3_302 b_3 NI_3 NS_302 0 2.1758756787208977e-06
GC_3_303 b_3 NI_3 NS_303 0 1.8069203401081262e-06
GC_3_304 b_3 NI_3 NS_304 0 2.7659732114236420e-06
GC_3_305 b_3 NI_3 NS_305 0 1.1298204583907870e-06
GC_3_306 b_3 NI_3 NS_306 0 9.3955426981398902e-07
GC_3_307 b_3 NI_3 NS_307 0 1.4884658142249148e-04
GC_3_308 b_3 NI_3 NS_308 0 1.9234487329115774e-05
GC_3_309 b_3 NI_3 NS_309 0 3.9278846319671573e-02
GC_3_310 b_3 NI_3 NS_310 0 -2.3265152078646759e-04
GC_3_311 b_3 NI_3 NS_311 0 -5.5253451610476605e-03
GC_3_312 b_3 NI_3 NS_312 0 6.2104283213495028e-04
GC_3_313 b_3 NI_3 NS_313 0 2.5852580645971388e-03
GC_3_314 b_3 NI_3 NS_314 0 -2.3322111819097913e-03
GC_3_315 b_3 NI_3 NS_315 0 -1.2110043352646215e-04
GC_3_316 b_3 NI_3 NS_316 0 -1.0841748006731438e-04
GC_3_317 b_3 NI_3 NS_317 0 2.1251555571569812e-03
GC_3_318 b_3 NI_3 NS_318 0 1.5334216510420455e-03
GC_3_319 b_3 NI_3 NS_319 0 -3.5719108323410231e-03
GC_3_320 b_3 NI_3 NS_320 0 -2.5194945382941530e-04
GC_3_321 b_3 NI_3 NS_321 0 2.5534493265226119e-05
GC_3_322 b_3 NI_3 NS_322 0 5.0696215896596042e-05
GC_3_323 b_3 NI_3 NS_323 0 -1.1603657125566437e-03
GC_3_324 b_3 NI_3 NS_324 0 4.3393020799918923e-04
GC_3_325 b_3 NI_3 NS_325 0 -4.0767606302257895e-05
GC_3_326 b_3 NI_3 NS_326 0 -4.9184528497440732e-05
GC_3_327 b_3 NI_3 NS_327 0 1.6115967672843787e-04
GC_3_328 b_3 NI_3 NS_328 0 3.2723857605888829e-04
GC_3_329 b_3 NI_3 NS_329 0 1.7364231066550759e-04
GC_3_330 b_3 NI_3 NS_330 0 2.0402195858405807e-05
GC_3_331 b_3 NI_3 NS_331 0 -1.9107067360143412e-06
GC_3_332 b_3 NI_3 NS_332 0 -5.3476859265268545e-05
GC_3_333 b_3 NI_3 NS_333 0 -4.4206306562920479e-05
GC_3_334 b_3 NI_3 NS_334 0 5.9070667225463250e-05
GC_3_335 b_3 NI_3 NS_335 0 -4.5025573543699959e-04
GC_3_336 b_3 NI_3 NS_336 0 -3.1591330051792843e-03
GC_3_337 b_3 NI_3 NS_337 0 1.9145429702667331e-06
GC_3_338 b_3 NI_3 NS_338 0 2.6495128073807286e-05
GC_3_339 b_3 NI_3 NS_339 0 -8.6230308380936930e-04
GC_3_340 b_3 NI_3 NS_340 0 1.0286235614388336e-03
GC_3_341 b_3 NI_3 NS_341 0 2.6847870840379067e-07
GC_3_342 b_3 NI_3 NS_342 0 5.0567698572762927e-06
GC_3_343 b_3 NI_3 NS_343 0 5.7311274989870647e-04
GC_3_344 b_3 NI_3 NS_344 0 -1.0736585789356332e-04
GC_3_345 b_3 NI_3 NS_345 0 -4.3512627387778442e-06
GC_3_346 b_3 NI_3 NS_346 0 -4.8626484671159753e-06
GC_3_347 b_3 NI_3 NS_347 0 1.4331945475448505e-06
GC_3_348 b_3 NI_3 NS_348 0 2.7487829690398908e-07
GC_3_349 b_3 NI_3 NS_349 0 -2.4890050212962990e-07
GC_3_350 b_3 NI_3 NS_350 0 -5.5507407334394552e-07
GC_3_351 b_3 NI_3 NS_351 0 4.3337950653775354e-05
GC_3_352 b_3 NI_3 NS_352 0 -4.9008439767990072e-05
GC_3_353 b_3 NI_3 NS_353 0 6.6558836821005206e-03
GC_3_354 b_3 NI_3 NS_354 0 7.2037377053801513e-05
GC_3_355 b_3 NI_3 NS_355 0 7.7325136206700394e-06
GC_3_356 b_3 NI_3 NS_356 0 -7.3280918763181813e-04
GC_3_357 b_3 NI_3 NS_357 0 7.9624033450129855e-04
GC_3_358 b_3 NI_3 NS_358 0 -3.2506063197656001e-04
GC_3_359 b_3 NI_3 NS_359 0 -1.1197732186616755e-03
GC_3_360 b_3 NI_3 NS_360 0 1.8635816206653803e-04
GC_3_361 b_3 NI_3 NS_361 0 1.1683215654292537e-03
GC_3_362 b_3 NI_3 NS_362 0 -3.2146532527671241e-04
GC_3_363 b_3 NI_3 NS_363 0 -1.7507408033528796e-03
GC_3_364 b_3 NI_3 NS_364 0 -2.5742536918941871e-04
GC_3_365 b_3 NI_3 NS_365 0 5.7845458146531237e-04
GC_3_366 b_3 NI_3 NS_366 0 -6.8230827729786052e-04
GC_3_367 b_3 NI_3 NS_367 0 7.2709872965023752e-03
GC_3_368 b_3 NI_3 NS_368 0 -1.6936100436036933e-03
GC_3_369 b_3 NI_3 NS_369 0 4.0505317000308794e-04
GC_3_370 b_3 NI_3 NS_370 0 3.9573834929369263e-04
GC_3_371 b_3 NI_3 NS_371 0 -1.6840727730758007e-05
GC_3_372 b_3 NI_3 NS_372 0 3.4144445070558279e-03
GC_3_373 b_3 NI_3 NS_373 0 4.6607954033359416e-04
GC_3_374 b_3 NI_3 NS_374 0 -3.4889675087111405e-04
GC_3_375 b_3 NI_3 NS_375 0 2.0083092384186576e-04
GC_3_376 b_3 NI_3 NS_376 0 -7.4041779310533035e-05
GC_3_377 b_3 NI_3 NS_377 0 3.7699005102849681e-05
GC_3_378 b_3 NI_3 NS_378 0 1.3194479967427802e-04
GC_3_379 b_3 NI_3 NS_379 0 -7.2294081533545171e-03
GC_3_380 b_3 NI_3 NS_380 0 8.8351753125818170e-03
GC_3_381 b_3 NI_3 NS_381 0 9.4168030265317799e-06
GC_3_382 b_3 NI_3 NS_382 0 -1.8238204867832124e-05
GC_3_383 b_3 NI_3 NS_383 0 2.3124639190475155e-03
GC_3_384 b_3 NI_3 NS_384 0 -1.0858815280901605e-03
GC_3_385 b_3 NI_3 NS_385 0 -2.2710860780182424e-06
GC_3_386 b_3 NI_3 NS_386 0 6.2393270381985824e-06
GC_3_387 b_3 NI_3 NS_387 0 -2.9346244137102261e-04
GC_3_388 b_3 NI_3 NS_388 0 -2.7375782709812327e-03
GC_3_389 b_3 NI_3 NS_389 0 -2.3823606197419470e-05
GC_3_390 b_3 NI_3 NS_390 0 7.0564506277769330e-07
GC_3_391 b_3 NI_3 NS_391 0 -4.5845482414722577e-07
GC_3_392 b_3 NI_3 NS_392 0 -2.3108276893463953e-06
GC_3_393 b_3 NI_3 NS_393 0 2.5409493166158059e-06
GC_3_394 b_3 NI_3 NS_394 0 3.3613287522651328e-06
GC_3_395 b_3 NI_3 NS_395 0 -1.1195898937057986e-04
GC_3_396 b_3 NI_3 NS_396 0 -8.4306666865705156e-04
GC_3_397 b_3 NI_3 NS_397 0 7.7280265843750603e-03
GC_3_398 b_3 NI_3 NS_398 0 9.0202204730654059e-06
GC_3_399 b_3 NI_3 NS_399 0 -9.6634488202820357e-05
GC_3_400 b_3 NI_3 NS_400 0 2.9651571857704782e-04
GC_3_401 b_3 NI_3 NS_401 0 -3.3163443963254882e-04
GC_3_402 b_3 NI_3 NS_402 0 -3.2884471614393968e-04
GC_3_403 b_3 NI_3 NS_403 0 -4.0412104358328299e-04
GC_3_404 b_3 NI_3 NS_404 0 8.6763312991390736e-05
GC_3_405 b_3 NI_3 NS_405 0 2.9350207524444187e-04
GC_3_406 b_3 NI_3 NS_406 0 -4.4776193796994859e-04
GC_3_407 b_3 NI_3 NS_407 0 6.2516853924282363e-04
GC_3_408 b_3 NI_3 NS_408 0 -1.8960918626385014e-05
GC_3_409 b_3 NI_3 NS_409 0 1.3539220472624360e-04
GC_3_410 b_3 NI_3 NS_410 0 9.4950342091591590e-05
GC_3_411 b_3 NI_3 NS_411 0 3.4862200786376843e-05
GC_3_412 b_3 NI_3 NS_412 0 1.4119830710080466e-03
GC_3_413 b_3 NI_3 NS_413 0 -1.8260134412977780e-04
GC_3_414 b_3 NI_3 NS_414 0 7.9695822135999986e-05
GC_3_415 b_3 NI_3 NS_415 0 -7.0512394795017332e-04
GC_3_416 b_3 NI_3 NS_416 0 -2.9672200172269162e-04
GC_3_417 b_3 NI_3 NS_417 0 -2.4767152799482856e-05
GC_3_418 b_3 NI_3 NS_418 0 -3.0036082031317054e-05
GC_3_419 b_3 NI_3 NS_419 0 -4.4857128750504088e-05
GC_3_420 b_3 NI_3 NS_420 0 -1.6601802972874874e-04
GC_3_421 b_3 NI_3 NS_421 0 -2.0894933548908116e-05
GC_3_422 b_3 NI_3 NS_422 0 1.3600740242838033e-04
GC_3_423 b_3 NI_3 NS_423 0 1.4084978598245678e-03
GC_3_424 b_3 NI_3 NS_424 0 1.2981759270782880e-03
GC_3_425 b_3 NI_3 NS_425 0 -3.2343135050883818e-05
GC_3_426 b_3 NI_3 NS_426 0 -1.4843822911442105e-05
GC_3_427 b_3 NI_3 NS_427 0 -5.0841242194314446e-04
GC_3_428 b_3 NI_3 NS_428 0 -9.3666150316099224e-04
GC_3_429 b_3 NI_3 NS_429 0 7.7396634298119641e-07
GC_3_430 b_3 NI_3 NS_430 0 -8.2858693472348655e-07
GC_3_431 b_3 NI_3 NS_431 0 -2.6889382336137911e-04
GC_3_432 b_3 NI_3 NS_432 0 -2.7151585645640331e-04
GC_3_433 b_3 NI_3 NS_433 0 -9.4411536699408078e-06
GC_3_434 b_3 NI_3 NS_434 0 -8.5978046102982603e-06
GC_3_435 b_3 NI_3 NS_435 0 -8.1906673591319125e-07
GC_3_436 b_3 NI_3 NS_436 0 6.8055887976788983e-08
GC_3_437 b_3 NI_3 NS_437 0 6.1738909043795916e-07
GC_3_438 b_3 NI_3 NS_438 0 -1.9212070179232509e-06
GC_3_439 b_3 NI_3 NS_439 0 -3.1984535111501502e-04
GC_3_440 b_3 NI_3 NS_440 0 -8.6008306224280180e-05
GC_3_441 b_3 NI_3 NS_441 0 -5.9553613149984001e-04
GC_3_442 b_3 NI_3 NS_442 0 9.6315189351087356e-05
GC_3_443 b_3 NI_3 NS_443 0 7.4891764804713287e-04
GC_3_444 b_3 NI_3 NS_444 0 -7.6481436722697577e-04
GC_3_445 b_3 NI_3 NS_445 0 3.9570991689186788e-04
GC_3_446 b_3 NI_3 NS_446 0 5.4605098010070770e-04
GC_3_447 b_3 NI_3 NS_447 0 -5.0914917056236054e-04
GC_3_448 b_3 NI_3 NS_448 0 -9.6590883434148774e-05
GC_3_449 b_3 NI_3 NS_449 0 1.0850139269768405e-03
GC_3_450 b_3 NI_3 NS_450 0 7.1873997539444168e-04
GC_3_451 b_3 NI_3 NS_451 0 -3.8689747566383677e-03
GC_3_452 b_3 NI_3 NS_452 0 -5.7242459464367274e-06
GC_3_453 b_3 NI_3 NS_453 0 5.7749955123705848e-04
GC_3_454 b_3 NI_3 NS_454 0 -4.5812355667677516e-04
GC_3_455 b_3 NI_3 NS_455 0 4.9505562911093788e-03
GC_3_456 b_3 NI_3 NS_456 0 -1.9110899413094711e-03
GC_3_457 b_3 NI_3 NS_457 0 2.4907722048131750e-04
GC_3_458 b_3 NI_3 NS_458 0 2.8215532031872399e-04
GC_3_459 b_3 NI_3 NS_459 0 -1.8134564186740934e-04
GC_3_460 b_3 NI_3 NS_460 0 1.2555367702898302e-03
GC_3_461 b_3 NI_3 NS_461 0 1.4635577727976294e-04
GC_3_462 b_3 NI_3 NS_462 0 -7.9921116496408328e-05
GC_3_463 b_3 NI_3 NS_463 0 1.5231733203812699e-04
GC_3_464 b_3 NI_3 NS_464 0 -6.5484773340644992e-05
GC_3_465 b_3 NI_3 NS_465 0 2.4317120255093729e-05
GC_3_466 b_3 NI_3 NS_466 0 8.2980927795174301e-05
GC_3_467 b_3 NI_3 NS_467 0 -3.1341482874231710e-03
GC_3_468 b_3 NI_3 NS_468 0 5.9087530955422383e-03
GC_3_469 b_3 NI_3 NS_469 0 2.1126459932355389e-06
GC_3_470 b_3 NI_3 NS_470 0 -1.1515540422381241e-05
GC_3_471 b_3 NI_3 NS_471 0 1.2415481697417110e-03
GC_3_472 b_3 NI_3 NS_472 0 -1.3121289262191785e-03
GC_3_473 b_3 NI_3 NS_473 0 -2.6295683726552061e-06
GC_3_474 b_3 NI_3 NS_474 0 7.2501522577720853e-07
GC_3_475 b_3 NI_3 NS_475 0 -9.4527347476437297e-05
GC_3_476 b_3 NI_3 NS_476 0 -1.5390036697602515e-03
GC_3_477 b_3 NI_3 NS_477 0 -1.0624980100645438e-05
GC_3_478 b_3 NI_3 NS_478 0 2.3213582454223141e-06
GC_3_479 b_3 NI_3 NS_479 0 -2.2320696335517259e-08
GC_3_480 b_3 NI_3 NS_480 0 4.5396607488890537e-07
GC_3_481 b_3 NI_3 NS_481 0 -2.7172503004980594e-07
GC_3_482 b_3 NI_3 NS_482 0 1.9128169239052082e-06
GC_3_483 b_3 NI_3 NS_483 0 -9.2710721307573524e-05
GC_3_484 b_3 NI_3 NS_484 0 -4.7248540664724493e-04
GC_3_485 b_3 NI_3 NS_485 0 1.2860599102839690e-02
GC_3_486 b_3 NI_3 NS_486 0 -4.7108784671294158e-05
GC_3_487 b_3 NI_3 NS_487 0 -6.3757923383382512e-04
GC_3_488 b_3 NI_3 NS_488 0 6.3611841265055183e-04
GC_3_489 b_3 NI_3 NS_489 0 -2.5329589470801694e-04
GC_3_490 b_3 NI_3 NS_490 0 -8.0152231835417011e-04
GC_3_491 b_3 NI_3 NS_491 0 -3.2284861037629073e-04
GC_3_492 b_3 NI_3 NS_492 0 -5.4335058909925536e-05
GC_3_493 b_3 NI_3 NS_493 0 5.6866688777839009e-04
GC_3_494 b_3 NI_3 NS_494 0 -1.0194718258469170e-04
GC_3_495 b_3 NI_3 NS_495 0 -4.5872329693319371e-04
GC_3_496 b_3 NI_3 NS_496 0 3.4302166777774954e-04
GC_3_497 b_3 NI_3 NS_497 0 9.8835247173617225e-05
GC_3_498 b_3 NI_3 NS_498 0 7.1405683557043716e-05
GC_3_499 b_3 NI_3 NS_499 0 -1.6623360729887987e-05
GC_3_500 b_3 NI_3 NS_500 0 8.1597706230803315e-04
GC_3_501 b_3 NI_3 NS_501 0 -1.0675188823741287e-04
GC_3_502 b_3 NI_3 NS_502 0 2.9085327367988502e-05
GC_3_503 b_3 NI_3 NS_503 0 -3.9627565687383318e-04
GC_3_504 b_3 NI_3 NS_504 0 -3.6658052500531917e-05
GC_3_505 b_3 NI_3 NS_505 0 2.4797360072531910e-05
GC_3_506 b_3 NI_3 NS_506 0 -4.9863110543331874e-05
GC_3_507 b_3 NI_3 NS_507 0 -2.5438337743798785e-05
GC_3_508 b_3 NI_3 NS_508 0 -9.6386968114607193e-05
GC_3_509 b_3 NI_3 NS_509 0 -1.7547397692856301e-05
GC_3_510 b_3 NI_3 NS_510 0 7.7928789906384812e-05
GC_3_511 b_3 NI_3 NS_511 0 2.6795502965724113e-04
GC_3_512 b_3 NI_3 NS_512 0 -3.3132577595083949e-04
GC_3_513 b_3 NI_3 NS_513 0 -1.8047884761594767e-05
GC_3_514 b_3 NI_3 NS_514 0 -3.7519022938333955e-06
GC_3_515 b_3 NI_3 NS_515 0 -4.4529983056114175e-04
GC_3_516 b_3 NI_3 NS_516 0 -1.1352623896118837e-04
GC_3_517 b_3 NI_3 NS_517 0 7.6780461513979569e-07
GC_3_518 b_3 NI_3 NS_518 0 6.1923071483191369e-07
GC_3_519 b_3 NI_3 NS_519 0 3.8876469458972182e-06
GC_3_520 b_3 NI_3 NS_520 0 -1.5897523647155986e-04
GC_3_521 b_3 NI_3 NS_521 0 -5.3256301119531560e-06
GC_3_522 b_3 NI_3 NS_522 0 -3.9141387157100451e-06
GC_3_523 b_3 NI_3 NS_523 0 -1.1739995720442399e-07
GC_3_524 b_3 NI_3 NS_524 0 4.5921977452371521e-07
GC_3_525 b_3 NI_3 NS_525 0 1.4615445195250366e-07
GC_3_526 b_3 NI_3 NS_526 0 -1.2343398222469982e-06
GC_3_527 b_3 NI_3 NS_527 0 -1.2461339215070303e-04
GC_3_528 b_3 NI_3 NS_528 0 -3.7127215250916990e-05
GD_3_1 b_3 NI_3 NA_1 0 1.4295396545135259e-03
GD_3_2 b_3 NI_3 NA_2 0 -6.4005299132180574e-02
GD_3_3 b_3 NI_3 NA_3 0 -1.3992074896311074e-01
GD_3_4 b_3 NI_3 NA_4 0 -4.1208491348131655e-02
GD_3_5 b_3 NI_3 NA_5 0 -2.4863362120756275e-03
GD_3_6 b_3 NI_3 NA_6 0 -8.5081740125845309e-02
GD_3_7 b_3 NI_3 NA_7 0 -3.3528076124901697e-02
GD_3_8 b_3 NI_3 NA_8 0 -3.8026279499973878e-02
GD_3_9 b_3 NI_3 NA_9 0 -1.4148907501163139e-02
GD_3_10 b_3 NI_3 NA_10 0 -8.7399610071584553e-03
GD_3_11 b_3 NI_3 NA_11 0 -3.1623102731393551e-03
GD_3_12 b_3 NI_3 NA_12 0 -1.2056772305497425e-02
*
* Port 4
VI_4 a_4 NI_4 0
RI_4 NI_4 b_4 5.0000000000000000e+01
GC_4_1 b_4 NI_4 NS_1 0 5.8037900911619769e-02
GC_4_2 b_4 NI_4 NS_2 0 -4.5391613580359413e-05
GC_4_3 b_4 NI_4 NS_3 0 -6.3536055289762170e-03
GC_4_4 b_4 NI_4 NS_4 0 -2.8143303559288670e-03
GC_4_5 b_4 NI_4 NS_5 0 4.5439174097504920e-03
GC_4_6 b_4 NI_4 NS_6 0 2.6349731677999659e-03
GC_4_7 b_4 NI_4 NS_7 0 -4.5415303820585143e-05
GC_4_8 b_4 NI_4 NS_8 0 -1.7645941483163141e-04
GC_4_9 b_4 NI_4 NS_9 0 1.4094138610975505e-03
GC_4_10 b_4 NI_4 NS_10 0 1.6567426437178192e-03
GC_4_11 b_4 NI_4 NS_11 0 -3.2810119542654834e-04
GC_4_12 b_4 NI_4 NS_12 0 -6.3409302560670368e-04
GC_4_13 b_4 NI_4 NS_13 0 -7.6751549017047466e-05
GC_4_14 b_4 NI_4 NS_14 0 6.6003546609637881e-05
GC_4_15 b_4 NI_4 NS_15 0 -3.9096021782227507e-03
GC_4_16 b_4 NI_4 NS_16 0 7.7685266678578617e-04
GC_4_17 b_4 NI_4 NS_17 0 -4.9588475792091185e-05
GC_4_18 b_4 NI_4 NS_18 0 -6.0471268029322489e-05
GC_4_19 b_4 NI_4 NS_19 0 -1.7887581848090588e-04
GC_4_20 b_4 NI_4 NS_20 0 8.0545532416792498e-04
GC_4_21 b_4 NI_4 NS_21 0 3.3912111282138945e-04
GC_4_22 b_4 NI_4 NS_22 0 1.0742553058750490e-04
GC_4_23 b_4 NI_4 NS_23 0 -2.2963037690875347e-05
GC_4_24 b_4 NI_4 NS_24 0 -2.3066274525423433e-05
GC_4_25 b_4 NI_4 NS_25 0 -4.0039232497656551e-05
GC_4_26 b_4 NI_4 NS_26 0 5.7029416437652149e-05
GC_4_27 b_4 NI_4 NS_27 0 -2.9145374640092737e-03
GC_4_28 b_4 NI_4 NS_28 0 -3.6207520601354471e-03
GC_4_29 b_4 NI_4 NS_29 0 1.3068746776432973e-05
GC_4_30 b_4 NI_4 NS_30 0 3.1587675471214885e-05
GC_4_31 b_4 NI_4 NS_31 0 -4.5771698929789810e-04
GC_4_32 b_4 NI_4 NS_32 0 1.9610214200766517e-03
GC_4_33 b_4 NI_4 NS_33 0 -2.2807159051902862e-07
GC_4_34 b_4 NI_4 NS_34 0 6.2996816397536069e-06
GC_4_35 b_4 NI_4 NS_35 0 8.8143137241771918e-04
GC_4_36 b_4 NI_4 NS_36 0 -3.5786971016317601e-04
GC_4_37 b_4 NI_4 NS_37 0 -7.6419218491463737e-06
GC_4_38 b_4 NI_4 NS_38 0 -7.5620559149404928e-06
GC_4_39 b_4 NI_4 NS_39 0 1.6426148499720869e-06
GC_4_40 b_4 NI_4 NS_40 0 -1.8962551873051357e-07
GC_4_41 b_4 NI_4 NS_41 0 1.4166606030741220e-06
GC_4_42 b_4 NI_4 NS_42 0 2.3011833054199314e-06
GC_4_43 b_4 NI_4 NS_43 0 1.4619905521803795e-04
GC_4_44 b_4 NI_4 NS_44 0 -9.6902802575447400e-05
GC_4_45 b_4 NI_4 NS_45 0 8.7751625081479660e-03
GC_4_46 b_4 NI_4 NS_46 0 -8.8798500395057954e-04
GC_4_47 b_4 NI_4 NS_47 0 4.0914945985556350e-03
GC_4_48 b_4 NI_4 NS_48 0 1.6307259180191370e-03
GC_4_49 b_4 NI_4 NS_49 0 -5.3014703536143270e-03
GC_4_50 b_4 NI_4 NS_50 0 -2.1301209066617232e-03
GC_4_51 b_4 NI_4 NS_51 0 2.8460769614407807e-04
GC_4_52 b_4 NI_4 NS_52 0 -2.7857758597359442e-04
GC_4_53 b_4 NI_4 NS_53 0 1.2238021831951732e-03
GC_4_54 b_4 NI_4 NS_54 0 1.5352189569616329e-04
GC_4_55 b_4 NI_4 NS_55 0 -1.1202117097799771e-04
GC_4_56 b_4 NI_4 NS_56 0 -5.2488576617233077e-04
GC_4_57 b_4 NI_4 NS_57 0 -1.8818100184081488e-05
GC_4_58 b_4 NI_4 NS_58 0 -3.7427298974799188e-05
GC_4_59 b_4 NI_4 NS_59 0 -1.1719674758648394e-03
GC_4_60 b_4 NI_4 NS_60 0 7.9808056970974873e-04
GC_4_61 b_4 NI_4 NS_61 0 2.2581156953555204e-05
GC_4_62 b_4 NI_4 NS_62 0 -1.1119962756800013e-05
GC_4_63 b_4 NI_4 NS_63 0 -3.3838560922205585e-05
GC_4_64 b_4 NI_4 NS_64 0 -6.9917908694758126e-05
GC_4_65 b_4 NI_4 NS_65 0 3.5064736479516689e-04
GC_4_66 b_4 NI_4 NS_66 0 -1.1489355437373060e-04
GC_4_67 b_4 NI_4 NS_67 0 -9.7941340620369299e-06
GC_4_68 b_4 NI_4 NS_68 0 -2.4824519236806852e-05
GC_4_69 b_4 NI_4 NS_69 0 -4.2367230508540880e-05
GC_4_70 b_4 NI_4 NS_70 0 -7.9066594814710458e-05
GC_4_71 b_4 NI_4 NS_71 0 9.9007343262649166e-04
GC_4_72 b_4 NI_4 NS_72 0 -9.7965342279545688e-04
GC_4_73 b_4 NI_4 NS_73 0 -3.3535994703154117e-05
GC_4_74 b_4 NI_4 NS_74 0 -3.7480040638335247e-05
GC_4_75 b_4 NI_4 NS_75 0 2.8908942376098124e-04
GC_4_76 b_4 NI_4 NS_76 0 -1.1664426933413635e-04
GC_4_77 b_4 NI_4 NS_77 0 -1.0500935035024947e-05
GC_4_78 b_4 NI_4 NS_78 0 1.2001480743325358e-05
GC_4_79 b_4 NI_4 NS_79 0 4.3994234631950278e-04
GC_4_80 b_4 NI_4 NS_80 0 6.7489704781433996e-05
GC_4_81 b_4 NI_4 NS_81 0 -1.8378090856609828e-07
GC_4_82 b_4 NI_4 NS_82 0 -9.7233119619739009e-06
GC_4_83 b_4 NI_4 NS_83 0 1.9425684176809202e-05
GC_4_84 b_4 NI_4 NS_84 0 2.9634541787841915e-07
GC_4_85 b_4 NI_4 NS_85 0 2.7196986588519131e-05
GC_4_86 b_4 NI_4 NS_86 0 -8.8295382142346779e-06
GC_4_87 b_4 NI_4 NS_87 0 -1.4646195798440965e-04
GC_4_88 b_4 NI_4 NS_88 0 8.9473388638158549e-05
GC_4_89 b_4 NI_4 NS_89 0 3.5592756509576370e-02
GC_4_90 b_4 NI_4 NS_90 0 1.0566342780244884e-02
GC_4_91 b_4 NI_4 NS_91 0 -1.0030245334559490e-02
GC_4_92 b_4 NI_4 NS_92 0 -3.9402786524045446e-03
GC_4_93 b_4 NI_4 NS_93 0 -9.6876630078036180e-03
GC_4_94 b_4 NI_4 NS_94 0 -1.5121362881058648e-03
GC_4_95 b_4 NI_4 NS_95 0 1.0311872886692329e-04
GC_4_96 b_4 NI_4 NS_96 0 1.2871602580839339e-04
GC_4_97 b_4 NI_4 NS_97 0 3.1272239929089115e-03
GC_4_98 b_4 NI_4 NS_98 0 2.8101416702448218e-03
GC_4_99 b_4 NI_4 NS_99 0 -2.3553740587581715e-05
GC_4_100 b_4 NI_4 NS_100 0 -1.3694868956482204e-03
GC_4_101 b_4 NI_4 NS_101 0 -3.0695226880895396e-06
GC_4_102 b_4 NI_4 NS_102 0 2.1713712327575308e-04
GC_4_103 b_4 NI_4 NS_103 0 3.8553268785384096e-03
GC_4_104 b_4 NI_4 NS_104 0 -6.7826699393733246e-04
GC_4_105 b_4 NI_4 NS_105 0 -2.0010021958702011e-05
GC_4_106 b_4 NI_4 NS_106 0 -3.8245690504303865e-05
GC_4_107 b_4 NI_4 NS_107 0 9.2898787845845001e-04
GC_4_108 b_4 NI_4 NS_108 0 8.1451531254779583e-04
GC_4_109 b_4 NI_4 NS_109 0 1.0575758980543072e-04
GC_4_110 b_4 NI_4 NS_110 0 -3.4831406172675306e-04
GC_4_111 b_4 NI_4 NS_111 0 1.9680245448349469e-05
GC_4_112 b_4 NI_4 NS_112 0 -1.2167884875337538e-05
GC_4_113 b_4 NI_4 NS_113 0 -3.1699702536433388e-05
GC_4_114 b_4 NI_4 NS_114 0 6.2682040378137229e-05
GC_4_115 b_4 NI_4 NS_115 0 -3.7150273361114656e-03
GC_4_116 b_4 NI_4 NS_116 0 -8.4011823567153616e-04
GC_4_117 b_4 NI_4 NS_117 0 1.2136870855344402e-05
GC_4_118 b_4 NI_4 NS_118 0 3.1614162054389282e-05
GC_4_119 b_4 NI_4 NS_119 0 3.2005309971982207e-04
GC_4_120 b_4 NI_4 NS_120 0 1.4242989306020137e-03
GC_4_121 b_4 NI_4 NS_121 0 7.8628303252876169e-06
GC_4_122 b_4 NI_4 NS_122 0 1.1551604683026880e-06
GC_4_123 b_4 NI_4 NS_123 0 4.2314727284380467e-06
GC_4_124 b_4 NI_4 NS_124 0 -9.4246059404437066e-04
GC_4_125 b_4 NI_4 NS_125 0 -7.4444313980296953e-06
GC_4_126 b_4 NI_4 NS_126 0 8.3986347636447364e-06
GC_4_127 b_4 NI_4 NS_127 0 -6.2998892143283251e-07
GC_4_128 b_4 NI_4 NS_128 0 -1.1435436815393905e-06
GC_4_129 b_4 NI_4 NS_129 0 2.3364262781518730e-06
GC_4_130 b_4 NI_4 NS_130 0 -4.2027290091253618e-06
GC_4_131 b_4 NI_4 NS_131 0 1.4553375233739318e-05
GC_4_132 b_4 NI_4 NS_132 0 -2.0877287906439742e-04
GC_4_133 b_4 NI_4 NS_133 0 -1.9911304066966054e-01
GC_4_134 b_4 NI_4 NS_134 0 8.5662066364841621e-03
GC_4_135 b_4 NI_4 NS_135 0 6.9162321737312113e-03
GC_4_136 b_4 NI_4 NS_136 0 3.9901198413718302e-03
GC_4_137 b_4 NI_4 NS_137 0 6.4587737558107327e-03
GC_4_138 b_4 NI_4 NS_138 0 1.8604385695946918e-03
GC_4_139 b_4 NI_4 NS_139 0 6.3282541713731780e-04
GC_4_140 b_4 NI_4 NS_140 0 6.4517715295479166e-04
GC_4_141 b_4 NI_4 NS_141 0 9.6060350324212937e-04
GC_4_142 b_4 NI_4 NS_142 0 1.8662185525905402e-03
GC_4_143 b_4 NI_4 NS_143 0 4.3552638832494292e-03
GC_4_144 b_4 NI_4 NS_144 0 3.1931408672211232e-03
GC_4_145 b_4 NI_4 NS_145 0 -2.2521520770938080e-04
GC_4_146 b_4 NI_4 NS_146 0 2.9221524527560421e-04
GC_4_147 b_4 NI_4 NS_147 0 2.1813909604553455e-03
GC_4_148 b_4 NI_4 NS_148 0 8.7749386607433918e-03
GC_4_149 b_4 NI_4 NS_149 0 -7.9100653538227724e-05
GC_4_150 b_4 NI_4 NS_150 0 1.0626401667861065e-04
GC_4_151 b_4 NI_4 NS_151 0 -4.9572244403585993e-04
GC_4_152 b_4 NI_4 NS_152 0 4.0024403045172980e-03
GC_4_153 b_4 NI_4 NS_153 0 8.1571632375715712e-04
GC_4_154 b_4 NI_4 NS_154 0 -3.3724250619521055e-04
GC_4_155 b_4 NI_4 NS_155 0 -1.3711494681792132e-04
GC_4_156 b_4 NI_4 NS_156 0 1.6679374831575291e-04
GC_4_157 b_4 NI_4 NS_157 0 2.1234104135687060e-05
GC_4_158 b_4 NI_4 NS_158 0 4.3308996291672127e-05
GC_4_159 b_4 NI_4 NS_159 0 -2.2428406684761908e-02
GC_4_160 b_4 NI_4 NS_160 0 -1.6108321009257549e-03
GC_4_161 b_4 NI_4 NS_161 0 2.2604084785632039e-05
GC_4_162 b_4 NI_4 NS_162 0 -4.6000439468082354e-05
GC_4_163 b_4 NI_4 NS_163 0 5.3358270807663697e-03
GC_4_164 b_4 NI_4 NS_164 0 6.0985148250481038e-03
GC_4_165 b_4 NI_4 NS_165 0 -3.9695378545560011e-06
GC_4_166 b_4 NI_4 NS_166 0 5.2088411556272047e-05
GC_4_167 b_4 NI_4 NS_167 0 2.0488419979492298e-03
GC_4_168 b_4 NI_4 NS_168 0 -3.3078624751465540e-03
GC_4_169 b_4 NI_4 NS_169 0 -6.5276422698008245e-05
GC_4_170 b_4 NI_4 NS_170 0 -2.5803750617077114e-05
GC_4_171 b_4 NI_4 NS_171 0 2.2030831849274082e-05
GC_4_172 b_4 NI_4 NS_172 0 -1.7377810350978173e-05
GC_4_173 b_4 NI_4 NS_173 0 5.4216390200527370e-05
GC_4_174 b_4 NI_4 NS_174 0 2.2217428770580030e-06
GC_4_175 b_4 NI_4 NS_175 0 4.3856471262557071e-04
GC_4_176 b_4 NI_4 NS_176 0 -6.4382068731820379e-04
GC_4_177 b_4 NI_4 NS_177 0 7.9090541096631467e-02
GC_4_178 b_4 NI_4 NS_178 0 -1.8753891934570854e-04
GC_4_179 b_4 NI_4 NS_179 0 -7.9628952946777555e-03
GC_4_180 b_4 NI_4 NS_180 0 -1.3312361042146998e-03
GC_4_181 b_4 NI_4 NS_181 0 4.0624094848743823e-03
GC_4_182 b_4 NI_4 NS_182 0 8.9025948188663033e-04
GC_4_183 b_4 NI_4 NS_183 0 -1.7175446058969300e-04
GC_4_184 b_4 NI_4 NS_184 0 -2.0552608254835279e-04
GC_4_185 b_4 NI_4 NS_185 0 2.2730308381595688e-03
GC_4_186 b_4 NI_4 NS_186 0 2.1453855438277629e-03
GC_4_187 b_4 NI_4 NS_187 0 -3.6129542573779469e-03
GC_4_188 b_4 NI_4 NS_188 0 8.2927294684756564e-05
GC_4_189 b_4 NI_4 NS_189 0 -6.0375578867270731e-05
GC_4_190 b_4 NI_4 NS_190 0 6.4655742863406338e-05
GC_4_191 b_4 NI_4 NS_191 0 -3.5049542933613866e-03
GC_4_192 b_4 NI_4 NS_192 0 -1.0708422061933320e-03
GC_4_193 b_4 NI_4 NS_193 0 -6.0243098770760409e-05
GC_4_194 b_4 NI_4 NS_194 0 -7.4937641499728776e-05
GC_4_195 b_4 NI_4 NS_195 0 1.2896796859445579e-04
GC_4_196 b_4 NI_4 NS_196 0 7.9264486089296044e-04
GC_4_197 b_4 NI_4 NS_197 0 3.3003245123156981e-04
GC_4_198 b_4 NI_4 NS_198 0 8.6816748827042072e-05
GC_4_199 b_4 NI_4 NS_199 0 -1.1460558929759584e-05
GC_4_200 b_4 NI_4 NS_200 0 -4.5242522304721139e-05
GC_4_201 b_4 NI_4 NS_201 0 -4.5094621905489968e-05
GC_4_202 b_4 NI_4 NS_202 0 7.2170011057056348e-05
GC_4_203 b_4 NI_4 NS_203 0 -2.2447327803743066e-03
GC_4_204 b_4 NI_4 NS_204 0 -4.1020458340130812e-03
GC_4_205 b_4 NI_4 NS_205 0 1.3778971009546602e-05
GC_4_206 b_4 NI_4 NS_206 0 3.8512360168277608e-05
GC_4_207 b_4 NI_4 NS_207 0 -7.4799408551703321e-04
GC_4_208 b_4 NI_4 NS_208 0 1.9582910052945075e-03
GC_4_209 b_4 NI_4 NS_209 0 -2.2456765653522471e-06
GC_4_210 b_4 NI_4 NS_210 0 6.3878129954961257e-06
GC_4_211 b_4 NI_4 NS_211 0 8.2569554700073831e-04
GC_4_212 b_4 NI_4 NS_212 0 -3.1208623877638326e-04
GC_4_213 b_4 NI_4 NS_213 0 -5.7576625426037623e-06
GC_4_214 b_4 NI_4 NS_214 0 -5.9278064276702181e-06
GC_4_215 b_4 NI_4 NS_215 0 1.8096092615440938e-06
GC_4_216 b_4 NI_4 NS_216 0 9.6200693197132668e-07
GC_4_217 b_4 NI_4 NS_217 0 2.2428087883872576e-06
GC_4_218 b_4 NI_4 NS_218 0 2.0329091765041225e-06
GC_4_219 b_4 NI_4 NS_219 0 1.0634100977949442e-04
GC_4_220 b_4 NI_4 NS_220 0 -1.0811605671790378e-04
GC_4_221 b_4 NI_4 NS_221 0 1.4868737222541860e-02
GC_4_222 b_4 NI_4 NS_222 0 -9.0521683786481684e-04
GC_4_223 b_4 NI_4 NS_223 0 5.1923134121618962e-03
GC_4_224 b_4 NI_4 NS_224 0 1.8804578989254039e-04
GC_4_225 b_4 NI_4 NS_225 0 -4.6846850537262067e-03
GC_4_226 b_4 NI_4 NS_226 0 -4.6334876488245873e-04
GC_4_227 b_4 NI_4 NS_227 0 -4.6875297228628213e-05
GC_4_228 b_4 NI_4 NS_228 0 3.5920032392449753e-04
GC_4_229 b_4 NI_4 NS_229 0 1.7419991386670951e-03
GC_4_230 b_4 NI_4 NS_230 0 4.6910729612522853e-04
GC_4_231 b_4 NI_4 NS_231 0 -5.9872156804480767e-04
GC_4_232 b_4 NI_4 NS_232 0 7.8370106575934484e-04
GC_4_233 b_4 NI_4 NS_233 0 -4.4853720882010063e-05
GC_4_234 b_4 NI_4 NS_234 0 -2.7051728432734727e-05
GC_4_235 b_4 NI_4 NS_235 0 -1.0481874245215784e-03
GC_4_236 b_4 NI_4 NS_236 0 7.5893148791403428e-04
GC_4_237 b_4 NI_4 NS_237 0 2.8066215579745036e-05
GC_4_238 b_4 NI_4 NS_238 0 -1.0508975046585542e-05
GC_4_239 b_4 NI_4 NS_239 0 4.0160463333257308e-05
GC_4_240 b_4 NI_4 NS_240 0 1.8963418054608085e-04
GC_4_241 b_4 NI_4 NS_241 0 5.9498363649804187e-04
GC_4_242 b_4 NI_4 NS_242 0 -3.3226303060296321e-04
GC_4_243 b_4 NI_4 NS_243 0 -2.1053218625905960e-05
GC_4_244 b_4 NI_4 NS_244 0 -2.2314748170464161e-05
GC_4_245 b_4 NI_4 NS_245 0 -6.1132345278409105e-05
GC_4_246 b_4 NI_4 NS_246 0 -1.1441393125639912e-04
GC_4_247 b_4 NI_4 NS_247 0 -1.0164192156973033e-03
GC_4_248 b_4 NI_4 NS_248 0 -9.4331324048784794e-04
GC_4_249 b_4 NI_4 NS_249 0 -4.4329838527798224e-05
GC_4_250 b_4 NI_4 NS_250 0 -5.1218545215283094e-05
GC_4_251 b_4 NI_4 NS_251 0 1.2063597043096915e-03
GC_4_252 b_4 NI_4 NS_252 0 1.2515559086610949e-04
GC_4_253 b_4 NI_4 NS_253 0 -9.0752223114982749e-06
GC_4_254 b_4 NI_4 NS_254 0 2.2441912694612616e-05
GC_4_255 b_4 NI_4 NS_255 0 7.0128225280765709e-04
GC_4_256 b_4 NI_4 NS_256 0 -4.7774977714722301e-04
GC_4_257 b_4 NI_4 NS_257 0 -8.6518861578120274e-06
GC_4_258 b_4 NI_4 NS_258 0 -1.1605988730708756e-05
GC_4_259 b_4 NI_4 NS_259 0 3.0259247740664876e-05
GC_4_260 b_4 NI_4 NS_260 0 -3.0790805676235554e-06
GC_4_261 b_4 NI_4 NS_261 0 3.8686884749681343e-05
GC_4_262 b_4 NI_4 NS_262 0 -1.5074008812057827e-05
GC_4_263 b_4 NI_4 NS_263 0 -1.4550123728449205e-04
GC_4_264 b_4 NI_4 NS_264 0 8.3127541615878319e-05
GC_4_265 b_4 NI_4 NS_265 0 3.3788776489855760e-02
GC_4_266 b_4 NI_4 NS_266 0 -2.0388118517120833e-04
GC_4_267 b_4 NI_4 NS_267 0 -5.5026168440841603e-03
GC_4_268 b_4 NI_4 NS_268 0 5.0652734122618175e-04
GC_4_269 b_4 NI_4 NS_269 0 2.6909309198925794e-03
GC_4_270 b_4 NI_4 NS_270 0 -2.3867910102454669e-03
GC_4_271 b_4 NI_4 NS_271 0 -1.5748424508111585e-04
GC_4_272 b_4 NI_4 NS_272 0 2.3007682555106667e-04
GC_4_273 b_4 NI_4 NS_273 0 2.1605684616711534e-03
GC_4_274 b_4 NI_4 NS_274 0 1.4832932339809953e-03
GC_4_275 b_4 NI_4 NS_275 0 -3.5966326719687049e-03
GC_4_276 b_4 NI_4 NS_276 0 -4.5070157856038490e-04
GC_4_277 b_4 NI_4 NS_277 0 2.6407191397333634e-05
GC_4_278 b_4 NI_4 NS_278 0 4.2459118046818802e-05
GC_4_279 b_4 NI_4 NS_279 0 -9.5021268675752018e-04
GC_4_280 b_4 NI_4 NS_280 0 7.3529008092300478e-05
GC_4_281 b_4 NI_4 NS_281 0 -3.1930639160069537e-05
GC_4_282 b_4 NI_4 NS_282 0 -4.3847887821133365e-05
GC_4_283 b_4 NI_4 NS_283 0 2.5669071476667847e-04
GC_4_284 b_4 NI_4 NS_284 0 1.8080885874418112e-04
GC_4_285 b_4 NI_4 NS_285 0 1.2241948718681259e-04
GC_4_286 b_4 NI_4 NS_286 0 6.7511183617961613e-05
GC_4_287 b_4 NI_4 NS_287 0 6.9805692799856073e-06
GC_4_288 b_4 NI_4 NS_288 0 -5.0247317021756518e-05
GC_4_289 b_4 NI_4 NS_289 0 -3.9996725251244851e-05
GC_4_290 b_4 NI_4 NS_290 0 4.8484425348060069e-05
GC_4_291 b_4 NI_4 NS_291 0 5.4138962736918685e-04
GC_4_292 b_4 NI_4 NS_292 0 -2.5242648813851684e-03
GC_4_293 b_4 NI_4 NS_293 0 -1.6793893837338612e-06
GC_4_294 b_4 NI_4 NS_294 0 2.4071648612027942e-05
GC_4_295 b_4 NI_4 NS_295 0 -8.6339595635934023e-04
GC_4_296 b_4 NI_4 NS_296 0 6.5339803165767249e-04
GC_4_297 b_4 NI_4 NS_297 0 -2.6633411344177252e-06
GC_4_298 b_4 NI_4 NS_298 0 3.2874311567234784e-06
GC_4_299 b_4 NI_4 NS_299 0 4.5084976437783741e-04
GC_4_300 b_4 NI_4 NS_300 0 1.3105409694284416e-04
GC_4_301 b_4 NI_4 NS_301 0 -3.7032606381164901e-07
GC_4_302 b_4 NI_4 NS_302 0 -5.3490604080725260e-06
GC_4_303 b_4 NI_4 NS_303 0 1.4168052287537736e-06
GC_4_304 b_4 NI_4 NS_304 0 5.8378197436501823e-07
GC_4_305 b_4 NI_4 NS_305 0 -4.2206705602281307e-07
GC_4_306 b_4 NI_4 NS_306 0 -9.7422833236169196e-07
GC_4_307 b_4 NI_4 NS_307 0 1.5117049942330119e-05
GC_4_308 b_4 NI_4 NS_308 0 -1.3826360892256054e-05
GC_4_309 b_4 NI_4 NS_309 0 1.4346644168074832e-02
GC_4_310 b_4 NI_4 NS_310 0 -3.2571209576701197e-04
GC_4_311 b_4 NI_4 NS_311 0 3.8560164645098090e-03
GC_4_312 b_4 NI_4 NS_312 0 -1.3456190142717662e-03
GC_4_313 b_4 NI_4 NS_313 0 -2.0590715975493095e-03
GC_4_314 b_4 NI_4 NS_314 0 2.4721393991260559e-03
GC_4_315 b_4 NI_4 NS_315 0 -4.7762474195825607e-04
GC_4_316 b_4 NI_4 NS_316 0 3.2548320151441599e-04
GC_4_317 b_4 NI_4 NS_317 0 9.9959767323699812e-04
GC_4_318 b_4 NI_4 NS_318 0 4.1630294474335501e-04
GC_4_319 b_4 NI_4 NS_319 0 -8.6285491435552752e-04
GC_4_320 b_4 NI_4 NS_320 0 1.3420833491334481e-03
GC_4_321 b_4 NI_4 NS_321 0 -6.3972814612053069e-05
GC_4_322 b_4 NI_4 NS_322 0 -3.3676946877136676e-05
GC_4_323 b_4 NI_4 NS_323 0 -7.0937095949161037e-04
GC_4_324 b_4 NI_4 NS_324 0 1.2971988293449437e-03
GC_4_325 b_4 NI_4 NS_325 0 2.2513531540496999e-06
GC_4_326 b_4 NI_4 NS_326 0 -1.5088578185054530e-05
GC_4_327 b_4 NI_4 NS_327 0 -3.1945186313053992e-04
GC_4_328 b_4 NI_4 NS_328 0 1.6807809343323259e-04
GC_4_329 b_4 NI_4 NS_329 0 3.6929719377991403e-04
GC_4_330 b_4 NI_4 NS_330 0 -1.5814388121801348e-04
GC_4_331 b_4 NI_4 NS_331 0 -3.4003789822325312e-05
GC_4_332 b_4 NI_4 NS_332 0 -1.8098843256076628e-05
GC_4_333 b_4 NI_4 NS_333 0 -4.3632733360996033e-05
GC_4_334 b_4 NI_4 NS_334 0 -7.0613142644086928e-05
GC_4_335 b_4 NI_4 NS_335 0 -2.4385716411181972e-03
GC_4_336 b_4 NI_4 NS_336 0 -1.9933288806851111e-03
GC_4_337 b_4 NI_4 NS_337 0 -1.8744992907818436e-05
GC_4_338 b_4 NI_4 NS_338 0 -2.2263668901252286e-05
GC_4_339 b_4 NI_4 NS_339 0 8.0829228780665563e-04
GC_4_340 b_4 NI_4 NS_340 0 6.8884903194073440e-04
GC_4_341 b_4 NI_4 NS_341 0 -2.1565200804590415e-06
GC_4_342 b_4 NI_4 NS_342 0 1.5281424704567723e-05
GC_4_343 b_4 NI_4 NS_343 0 6.3224990822832023e-04
GC_4_344 b_4 NI_4 NS_344 0 -4.6727514220131264e-04
GC_4_345 b_4 NI_4 NS_345 0 -7.4456206726498038e-06
GC_4_346 b_4 NI_4 NS_346 0 -7.5910541543065306e-06
GC_4_347 b_4 NI_4 NS_347 0 2.0564702572194485e-05
GC_4_348 b_4 NI_4 NS_348 0 -6.1114226788233746e-07
GC_4_349 b_4 NI_4 NS_349 0 1.9470775408923073e-05
GC_4_350 b_4 NI_4 NS_350 0 -2.5895216178275397e-06
GC_4_351 b_4 NI_4 NS_351 0 4.8596091408822928e-05
GC_4_352 b_4 NI_4 NS_352 0 3.8883970351115865e-05
GC_4_353 b_4 NI_4 NS_353 0 8.5315067134810550e-03
GC_4_354 b_4 NI_4 NS_354 0 1.0772723634224599e-05
GC_4_355 b_4 NI_4 NS_355 0 -8.2028579500118744e-05
GC_4_356 b_4 NI_4 NS_356 0 2.8470289855928466e-04
GC_4_357 b_4 NI_4 NS_357 0 -3.1093127014794180e-04
GC_4_358 b_4 NI_4 NS_358 0 -3.0657286207580670e-04
GC_4_359 b_4 NI_4 NS_359 0 -3.3410662522855673e-04
GC_4_360 b_4 NI_4 NS_360 0 1.0880594076358764e-04
GC_4_361 b_4 NI_4 NS_361 0 3.0336050826959056e-04
GC_4_362 b_4 NI_4 NS_362 0 -4.1443568323169539e-04
GC_4_363 b_4 NI_4 NS_363 0 7.1085970422315136e-04
GC_4_364 b_4 NI_4 NS_364 0 -1.4210419406766896e-05
GC_4_365 b_4 NI_4 NS_365 0 1.1796089934075293e-04
GC_4_366 b_4 NI_4 NS_366 0 1.2662332072705223e-04
GC_4_367 b_4 NI_4 NS_367 0 -1.8339202834724628e-05
GC_4_368 b_4 NI_4 NS_368 0 1.4343089140541603e-03
GC_4_369 b_4 NI_4 NS_369 0 -1.4176996572940750e-04
GC_4_370 b_4 NI_4 NS_370 0 6.8389848460749899e-05
GC_4_371 b_4 NI_4 NS_371 0 -6.2914179993684533e-04
GC_4_372 b_4 NI_4 NS_372 0 -1.4961658144516842e-04
GC_4_373 b_4 NI_4 NS_373 0 -1.2871117250182717e-05
GC_4_374 b_4 NI_4 NS_374 0 -4.7807577996485917e-05
GC_4_375 b_4 NI_4 NS_375 0 -3.0255667205900539e-05
GC_4_376 b_4 NI_4 NS_376 0 -1.2353373532765711e-04
GC_4_377 b_4 NI_4 NS_377 0 -3.2600878552422430e-06
GC_4_378 b_4 NI_4 NS_378 0 9.9802305100462545e-05
GC_4_379 b_4 NI_4 NS_379 0 6.6929850062252285e-04
GC_4_380 b_4 NI_4 NS_380 0 3.5611076640541784e-04
GC_4_381 b_4 NI_4 NS_381 0 -2.6654133857971154e-05
GC_4_382 b_4 NI_4 NS_382 0 -1.1439792006128005e-05
GC_4_383 b_4 NI_4 NS_383 0 -3.8522597243801379e-04
GC_4_384 b_4 NI_4 NS_384 0 -3.6760188218926528e-04
GC_4_385 b_4 NI_4 NS_385 0 3.9498711479028995e-09
GC_4_386 b_4 NI_4 NS_386 0 1.6529104081972102e-06
GC_4_387 b_4 NI_4 NS_387 0 -1.3698592798363203e-04
GC_4_388 b_4 NI_4 NS_388 0 -1.4723215144275324e-04
GC_4_389 b_4 NI_4 NS_389 0 -8.5640418505645242e-06
GC_4_390 b_4 NI_4 NS_390 0 -1.4077661444204956e-05
GC_4_391 b_4 NI_4 NS_391 0 -1.9766256340575659e-07
GC_4_392 b_4 NI_4 NS_392 0 1.2404380989621838e-06
GC_4_393 b_4 NI_4 NS_393 0 -8.8913539346097190e-07
GC_4_394 b_4 NI_4 NS_394 0 -1.4725025388982397e-06
GC_4_395 b_4 NI_4 NS_395 0 -2.1057908720284772e-04
GC_4_396 b_4 NI_4 NS_396 0 -2.6955568110038412e-05
GC_4_397 b_4 NI_4 NS_397 0 1.5261941981014114e-03
GC_4_398 b_4 NI_4 NS_398 0 -1.5319598367235623e-05
GC_4_399 b_4 NI_4 NS_399 0 -9.5775329198149084e-05
GC_4_400 b_4 NI_4 NS_400 0 -3.4024140403347722e-04
GC_4_401 b_4 NI_4 NS_401 0 3.2583761548974206e-04
GC_4_402 b_4 NI_4 NS_402 0 -7.3639757147470064e-05
GC_4_403 b_4 NI_4 NS_403 0 -3.9906035404597880e-04
GC_4_404 b_4 NI_4 NS_404 0 3.9982820502898220e-05
GC_4_405 b_4 NI_4 NS_405 0 1.5255884742074513e-04
GC_4_406 b_4 NI_4 NS_406 0 -2.6852099193982917e-04
GC_4_407 b_4 NI_4 NS_407 0 4.6393368014827291e-04
GC_4_408 b_4 NI_4 NS_408 0 -3.6411470907070148e-04
GC_4_409 b_4 NI_4 NS_409 0 1.3626390401286451e-05
GC_4_410 b_4 NI_4 NS_410 0 4.0018141947369151e-05
GC_4_411 b_4 NI_4 NS_411 0 6.6803819396953643e-04
GC_4_412 b_4 NI_4 NS_412 0 -4.2046827255124694e-04
GC_4_413 b_4 NI_4 NS_413 0 1.6906141686149965e-05
GC_4_414 b_4 NI_4 NS_414 0 -5.1056777976067540e-05
GC_4_415 b_4 NI_4 NS_415 0 8.5696231056375566e-04
GC_4_416 b_4 NI_4 NS_416 0 -3.7368037799428793e-04
GC_4_417 b_4 NI_4 NS_417 0 -2.2643100637513984e-04
GC_4_418 b_4 NI_4 NS_418 0 -3.2059432883560832e-04
GC_4_419 b_4 NI_4 NS_419 0 1.3707448885870150e-05
GC_4_420 b_4 NI_4 NS_420 0 -2.5539863199586436e-05
GC_4_421 b_4 NI_4 NS_421 0 -4.4913202416834814e-05
GC_4_422 b_4 NI_4 NS_422 0 -1.7837500363400956e-04
GC_4_423 b_4 NI_4 NS_423 0 -4.5214064158074730e-03
GC_4_424 b_4 NI_4 NS_424 0 5.5192320494758485e-03
GC_4_425 b_4 NI_4 NS_425 0 1.9681308042940423e-05
GC_4_426 b_4 NI_4 NS_426 0 1.8399778805462555e-05
GC_4_427 b_4 NI_4 NS_427 0 3.9278727568875333e-03
GC_4_428 b_4 NI_4 NS_428 0 -1.6403554226381224e-03
GC_4_429 b_4 NI_4 NS_429 0 1.8963351723398959e-05
GC_4_430 b_4 NI_4 NS_430 0 3.1967088306355990e-06
GC_4_431 b_4 NI_4 NS_431 0 -3.6724315351813224e-04
GC_4_432 b_4 NI_4 NS_432 0 -4.8547844066548459e-04
GC_4_433 b_4 NI_4 NS_433 0 -4.9843697472442049e-05
GC_4_434 b_4 NI_4 NS_434 0 1.1155930632506564e-05
GC_4_435 b_4 NI_4 NS_435 0 3.1539029017405053e-05
GC_4_436 b_4 NI_4 NS_436 0 -5.5713807446134231e-06
GC_4_437 b_4 NI_4 NS_437 0 -2.3464566286285402e-05
GC_4_438 b_4 NI_4 NS_438 0 1.3832772270725422e-05
GC_4_439 b_4 NI_4 NS_439 0 4.1989882755443387e-04
GC_4_440 b_4 NI_4 NS_440 0 1.2945206282210316e-04
GC_4_441 b_4 NI_4 NS_441 0 1.2175543499857654e-02
GC_4_442 b_4 NI_4 NS_442 0 -4.6083429603035999e-05
GC_4_443 b_4 NI_4 NS_443 0 -6.2453566370276154e-04
GC_4_444 b_4 NI_4 NS_444 0 6.3789086988907940e-04
GC_4_445 b_4 NI_4 NS_445 0 -2.7049982030935126e-04
GC_4_446 b_4 NI_4 NS_446 0 -7.8978524657718899e-04
GC_4_447 b_4 NI_4 NS_447 0 -2.7800657453891766e-04
GC_4_448 b_4 NI_4 NS_448 0 -7.8678014192119398e-05
GC_4_449 b_4 NI_4 NS_449 0 5.5570752696025647e-04
GC_4_450 b_4 NI_4 NS_450 0 -1.0487176986931883e-04
GC_4_451 b_4 NI_4 NS_451 0 -4.1408773513617448e-04
GC_4_452 b_4 NI_4 NS_452 0 3.4470204585731275e-04
GC_4_453 b_4 NI_4 NS_453 0 8.5057662413234910e-05
GC_4_454 b_4 NI_4 NS_454 0 7.9836957021941755e-05
GC_4_455 b_4 NI_4 NS_455 0 -5.9875960166428691e-05
GC_4_456 b_4 NI_4 NS_456 0 8.3159683833063515e-04
GC_4_457 b_4 NI_4 NS_457 0 -1.0066004163796856e-04
GC_4_458 b_4 NI_4 NS_458 0 3.0280993752121507e-05
GC_4_459 b_4 NI_4 NS_459 0 -4.4908456592590118e-04
GC_4_460 b_4 NI_4 NS_460 0 -2.6213334942869309e-05
GC_4_461 b_4 NI_4 NS_461 0 2.3536341430201514e-05
GC_4_462 b_4 NI_4 NS_462 0 -4.8881025380654421e-05
GC_4_463 b_4 NI_4 NS_463 0 -2.3920214847479896e-05
GC_4_464 b_4 NI_4 NS_464 0 -9.2012627954446321e-05
GC_4_465 b_4 NI_4 NS_465 0 -2.0726269113696521e-05
GC_4_466 b_4 NI_4 NS_466 0 7.3624203123458359e-05
GC_4_467 b_4 NI_4 NS_467 0 2.1980646442512459e-04
GC_4_468 b_4 NI_4 NS_468 0 -5.5910333391851613e-04
GC_4_469 b_4 NI_4 NS_469 0 -1.4806914977658869e-05
GC_4_470 b_4 NI_4 NS_470 0 -5.3585934609099017e-06
GC_4_471 b_4 NI_4 NS_471 0 -4.5281730698559775e-04
GC_4_472 b_4 NI_4 NS_472 0 -6.8227078627393410e-05
GC_4_473 b_4 NI_4 NS_473 0 -7.1565924338040763e-07
GC_4_474 b_4 NI_4 NS_474 0 -4.9648836493726108e-07
GC_4_475 b_4 NI_4 NS_475 0 6.2426543885756136e-05
GC_4_476 b_4 NI_4 NS_476 0 -1.0001616018765932e-04
GC_4_477 b_4 NI_4 NS_477 0 -4.6421494786171610e-06
GC_4_478 b_4 NI_4 NS_478 0 -8.6256922947363364e-06
GC_4_479 b_4 NI_4 NS_479 0 7.1916189844323931e-07
GC_4_480 b_4 NI_4 NS_480 0 1.2656688479656689e-08
GC_4_481 b_4 NI_4 NS_481 0 -9.5193072747027250e-07
GC_4_482 b_4 NI_4 NS_482 0 -6.3026953824664039e-08
GC_4_483 b_4 NI_4 NS_483 0 -1.0272740019320222e-04
GC_4_484 b_4 NI_4 NS_484 0 -2.6090958640876207e-05
GC_4_485 b_4 NI_4 NS_485 0 7.2567150194420831e-04
GC_4_486 b_4 NI_4 NS_486 0 -8.0781696509598381e-06
GC_4_487 b_4 NI_4 NS_487 0 3.3662973581674458e-04
GC_4_488 b_4 NI_4 NS_488 0 -6.9380013119351325e-04
GC_4_489 b_4 NI_4 NS_489 0 3.8925063164818298e-04
GC_4_490 b_4 NI_4 NS_490 0 4.9571224155920226e-04
GC_4_491 b_4 NI_4 NS_491 0 -3.5207873969822295e-04
GC_4_492 b_4 NI_4 NS_492 0 3.5471582840414126e-04
GC_4_493 b_4 NI_4 NS_493 0 2.9819382406724937e-04
GC_4_494 b_4 NI_4 NS_494 0 -8.7688023949028271e-05
GC_4_495 b_4 NI_4 NS_495 0 1.7845249464237185e-04
GC_4_496 b_4 NI_4 NS_496 0 2.3242787143991554e-04
GC_4_497 b_4 NI_4 NS_497 0 -7.9353728475845016e-06
GC_4_498 b_4 NI_4 NS_498 0 1.6355173208022105e-05
GC_4_499 b_4 NI_4 NS_499 0 3.3755574083596567e-04
GC_4_500 b_4 NI_4 NS_500 0 -1.5646858022025112e-04
GC_4_501 b_4 NI_4 NS_501 0 1.0475827515741910e-05
GC_4_502 b_4 NI_4 NS_502 0 -3.0044320080782736e-05
GC_4_503 b_4 NI_4 NS_503 0 4.1675432117365638e-04
GC_4_504 b_4 NI_4 NS_504 0 -1.9135953763998011e-04
GC_4_505 b_4 NI_4 NS_505 0 -5.3924880208338861e-05
GC_4_506 b_4 NI_4 NS_506 0 -1.8196864574411708e-04
GC_4_507 b_4 NI_4 NS_507 0 3.1612224022943859e-06
GC_4_508 b_4 NI_4 NS_508 0 -1.6726211032061179e-05
GC_4_509 b_4 NI_4 NS_509 0 -3.0790345365712247e-05
GC_4_510 b_4 NI_4 NS_510 0 -1.1130855547968180e-04
GC_4_511 b_4 NI_4 NS_511 0 -2.6624618418490081e-03
GC_4_512 b_4 NI_4 NS_512 0 2.8868612301620037e-03
GC_4_513 b_4 NI_4 NS_513 0 4.8420947191782850e-06
GC_4_514 b_4 NI_4 NS_514 0 5.8948043903717390e-06
GC_4_515 b_4 NI_4 NS_515 0 2.2756129492902421e-03
GC_4_516 b_4 NI_4 NS_516 0 -8.7878950774536425e-04
GC_4_517 b_4 NI_4 NS_517 0 6.5909470395028978e-06
GC_4_518 b_4 NI_4 NS_518 0 2.6244148314341721e-06
GC_4_519 b_4 NI_4 NS_519 0 -1.2637915667291526e-04
GC_4_520 b_4 NI_4 NS_520 0 -2.8418512985914173e-04
GC_4_521 b_4 NI_4 NS_521 0 -1.9337984037377680e-05
GC_4_522 b_4 NI_4 NS_522 0 4.2957374779766990e-06
GC_4_523 b_4 NI_4 NS_523 0 2.0232738660558289e-05
GC_4_524 b_4 NI_4 NS_524 0 -1.2019293960926881e-06
GC_4_525 b_4 NI_4 NS_525 0 -9.1170649436953674e-06
GC_4_526 b_4 NI_4 NS_526 0 4.5475276396473840e-06
GC_4_527 b_4 NI_4 NS_527 0 2.1200327349106256e-04
GC_4_528 b_4 NI_4 NS_528 0 5.1564113869493095e-05
GD_4_1 b_4 NI_4 NA_1 0 -6.1519775667100637e-02
GD_4_2 b_4 NI_4 NA_2 0 -1.5790005140183538e-02
GD_4_3 b_4 NI_4 NA_3 0 -4.1208491348117569e-02
GD_4_4 b_4 NI_4 NA_4 0 2.4887730874937283e-01
GD_4_5 b_4 NI_4 NA_5 0 -8.1131772018087647e-02
GD_4_6 b_4 NI_4 NA_6 0 -2.6996141370235122e-02
GD_4_7 b_4 NI_4 NA_7 0 -3.3792607450469921e-02
GD_4_8 b_4 NI_4 NA_8 0 -1.8322305683349256e-02
GD_4_9 b_4 NI_4 NA_9 0 -9.6793188063716371e-03
GD_4_10 b_4 NI_4 NA_10 0 -4.2863540065094866e-03
GD_4_11 b_4 NI_4 NA_11 0 -1.1170994029428290e-02
GD_4_12 b_4 NI_4 NA_12 0 -3.3553895468527795e-03
*
* Port 5
VI_5 a_5 NI_5 0
RI_5 NI_5 b_5 5.0000000000000000e+01
GC_5_1 b_5 NI_5 NS_1 0 3.2244365380994539e-02
GC_5_2 b_5 NI_5 NS_2 0 9.9828524791980861e-05
GC_5_3 b_5 NI_5 NS_3 0 6.0074318997957012e-03
GC_5_4 b_5 NI_5 NS_4 0 1.1808748036606631e-03
GC_5_5 b_5 NI_5 NS_5 0 -4.3858387871842028e-03
GC_5_6 b_5 NI_5 NS_6 0 2.6167250205370129e-03
GC_5_7 b_5 NI_5 NS_7 0 -1.9520787432520902e-04
GC_5_8 b_5 NI_5 NS_8 0 -9.2904559744207084e-04
GC_5_9 b_5 NI_5 NS_9 0 1.2072633119826243e-03
GC_5_10 b_5 NI_5 NS_10 0 6.0278955275615050e-03
GC_5_11 b_5 NI_5 NS_11 0 -1.0133194922039136e-02
GC_5_12 b_5 NI_5 NS_12 0 -1.2931473172359100e-03
GC_5_13 b_5 NI_5 NS_13 0 8.6808542155119716e-04
GC_5_14 b_5 NI_5 NS_14 0 2.4012285397789830e-04
GC_5_15 b_5 NI_5 NS_15 0 -2.6165023295145937e-03
GC_5_16 b_5 NI_5 NS_16 0 3.6605151016874459e-04
GC_5_17 b_5 NI_5 NS_17 0 -7.6933221236069439e-05
GC_5_18 b_5 NI_5 NS_18 0 1.2695582224028410e-04
GC_5_19 b_5 NI_5 NS_19 0 -1.9995731938827342e-03
GC_5_20 b_5 NI_5 NS_20 0 -3.7551143656506273e-03
GC_5_21 b_5 NI_5 NS_21 0 -9.6756900546674646e-05
GC_5_22 b_5 NI_5 NS_22 0 6.2460712246393321e-04
GC_5_23 b_5 NI_5 NS_23 0 1.5201611793014941e-04
GC_5_24 b_5 NI_5 NS_24 0 -7.2212052149075117e-05
GC_5_25 b_5 NI_5 NS_25 0 -4.6513391124261637e-06
GC_5_26 b_5 NI_5 NS_26 0 -1.0029132993935659e-04
GC_5_27 b_5 NI_5 NS_27 0 3.3711763004527916e-03
GC_5_28 b_5 NI_5 NS_28 0 -2.1823934854050841e-03
GC_5_29 b_5 NI_5 NS_29 0 -1.4940585946732025e-05
GC_5_30 b_5 NI_5 NS_30 0 -2.1910509337651751e-06
GC_5_31 b_5 NI_5 NS_31 0 -4.3001084132156074e-04
GC_5_32 b_5 NI_5 NS_32 0 -2.5085607216320193e-03
GC_5_33 b_5 NI_5 NS_33 0 -4.7110668016106179e-07
GC_5_34 b_5 NI_5 NS_34 0 -6.5528040246407808e-06
GC_5_35 b_5 NI_5 NS_35 0 1.4780811371675727e-03
GC_5_36 b_5 NI_5 NS_36 0 8.3287926240604179e-04
GC_5_37 b_5 NI_5 NS_37 0 8.6742405906214917e-06
GC_5_38 b_5 NI_5 NS_38 0 2.8103872220601476e-06
GC_5_39 b_5 NI_5 NS_39 0 1.7339333174647046e-06
GC_5_40 b_5 NI_5 NS_40 0 3.7347143987416175e-06
GC_5_41 b_5 NI_5 NS_41 0 3.9892378273707868e-07
GC_5_42 b_5 NI_5 NS_42 0 9.7631192443308858e-08
GC_5_43 b_5 NI_5 NS_43 0 1.6077375852876219e-04
GC_5_44 b_5 NI_5 NS_44 0 1.1337143098119208e-04
GC_5_45 b_5 NI_5 NS_45 0 3.9622292483443407e-02
GC_5_46 b_5 NI_5 NS_46 0 -2.3691614670306646e-04
GC_5_47 b_5 NI_5 NS_47 0 -5.6773487281087855e-03
GC_5_48 b_5 NI_5 NS_48 0 6.9768052855822757e-04
GC_5_49 b_5 NI_5 NS_49 0 2.5618358951827350e-03
GC_5_50 b_5 NI_5 NS_50 0 -2.4925754830134716e-03
GC_5_51 b_5 NI_5 NS_51 0 -9.2175038618915226e-05
GC_5_52 b_5 NI_5 NS_52 0 -2.7688128220226916e-05
GC_5_53 b_5 NI_5 NS_53 0 2.2172444865354219e-03
GC_5_54 b_5 NI_5 NS_54 0 1.5253139973632149e-03
GC_5_55 b_5 NI_5 NS_55 0 -3.9397653556183876e-03
GC_5_56 b_5 NI_5 NS_56 0 -2.6243794845758479e-04
GC_5_57 b_5 NI_5 NS_57 0 3.7947450825701729e-05
GC_5_58 b_5 NI_5 NS_58 0 2.6486134502783982e-05
GC_5_59 b_5 NI_5 NS_59 0 -5.9147239083467886e-04
GC_5_60 b_5 NI_5 NS_60 0 -3.0435858907722088e-05
GC_5_61 b_5 NI_5 NS_61 0 -3.5906261591624696e-05
GC_5_62 b_5 NI_5 NS_62 0 -6.8523126878389666e-05
GC_5_63 b_5 NI_5 NS_63 0 3.9647464963470173e-04
GC_5_64 b_5 NI_5 NS_64 0 5.8710706303311759e-04
GC_5_65 b_5 NI_5 NS_65 0 2.6985515067974402e-04
GC_5_66 b_5 NI_5 NS_66 0 9.9496333024439999e-05
GC_5_67 b_5 NI_5 NS_67 0 1.6862576875474535e-06
GC_5_68 b_5 NI_5 NS_68 0 -3.9011134413238240e-05
GC_5_69 b_5 NI_5 NS_69 0 -4.0921664144303365e-05
GC_5_70 b_5 NI_5 NS_70 0 5.9107831720709437e-05
GC_5_71 b_5 NI_5 NS_71 0 -1.1821912786363956e-03
GC_5_72 b_5 NI_5 NS_72 0 -3.6957213808795223e-03
GC_5_73 b_5 NI_5 NS_73 0 1.2454417973241905e-05
GC_5_74 b_5 NI_5 NS_74 0 3.5707535556061523e-05
GC_5_75 b_5 NI_5 NS_75 0 -7.7345298234279066e-04
GC_5_76 b_5 NI_5 NS_76 0 1.6500640224275996e-03
GC_5_77 b_5 NI_5 NS_77 0 -3.2939445416139824e-06
GC_5_78 b_5 NI_5 NS_78 0 6.0222030229246202e-06
GC_5_79 b_5 NI_5 NS_79 0 7.5502075950925108e-04
GC_5_80 b_5 NI_5 NS_80 0 -1.1755906200740002e-04
GC_5_81 b_5 NI_5 NS_81 0 -3.7668355127365563e-06
GC_5_82 b_5 NI_5 NS_82 0 -5.7648358657243210e-06
GC_5_83 b_5 NI_5 NS_83 0 1.8659211074008522e-06
GC_5_84 b_5 NI_5 NS_84 0 1.1002313748249628e-06
GC_5_85 b_5 NI_5 NS_85 0 1.6261228556296335e-06
GC_5_86 b_5 NI_5 NS_86 0 9.8172636404989763e-07
GC_5_87 b_5 NI_5 NS_87 0 7.5333039511060661e-05
GC_5_88 b_5 NI_5 NS_88 0 -9.8976170955782471e-05
GC_5_89 b_5 NI_5 NS_89 0 2.6042158903321374e-03
GC_5_90 b_5 NI_5 NS_90 0 8.9383988555531482e-05
GC_5_91 b_5 NI_5 NS_91 0 7.3168842305765154e-03
GC_5_92 b_5 NI_5 NS_92 0 3.7799779023196737e-03
GC_5_93 b_5 NI_5 NS_93 0 -5.6738793867510077e-03
GC_5_94 b_5 NI_5 NS_94 0 -2.2607660269688239e-03
GC_5_95 b_5 NI_5 NS_95 0 -5.6491116057188535e-06
GC_5_96 b_5 NI_5 NS_96 0 3.1195551134693885e-04
GC_5_97 b_5 NI_5 NS_97 0 2.1334644263685128e-03
GC_5_98 b_5 NI_5 NS_98 0 8.2163653387986747e-03
GC_5_99 b_5 NI_5 NS_99 0 -1.0559431133077907e-02
GC_5_100 b_5 NI_5 NS_100 0 -1.3285589993704975e-03
GC_5_101 b_5 NI_5 NS_101 0 1.2038340771693167e-03
GC_5_102 b_5 NI_5 NS_102 0 3.3587979404634146e-04
GC_5_103 b_5 NI_5 NS_103 0 -3.1080656922313037e-03
GC_5_104 b_5 NI_5 NS_104 0 -3.7438129827452606e-03
GC_5_105 b_5 NI_5 NS_105 0 -1.0879779738672750e-04
GC_5_106 b_5 NI_5 NS_106 0 1.6956704233102846e-04
GC_5_107 b_5 NI_5 NS_107 0 -2.8483499052597773e-03
GC_5_108 b_5 NI_5 NS_108 0 -4.7724640016430404e-03
GC_5_109 b_5 NI_5 NS_109 0 -2.0528968079450597e-04
GC_5_110 b_5 NI_5 NS_110 0 1.3525004221160498e-03
GC_5_111 b_5 NI_5 NS_111 0 2.3453680792220473e-04
GC_5_112 b_5 NI_5 NS_112 0 -1.0747945072540712e-04
GC_5_113 b_5 NI_5 NS_113 0 3.5790555353218140e-06
GC_5_114 b_5 NI_5 NS_114 0 -1.3549743494172637e-04
GC_5_115 b_5 NI_5 NS_115 0 9.4726475671575317e-03
GC_5_116 b_5 NI_5 NS_116 0 -4.0329155800449559e-04
GC_5_117 b_5 NI_5 NS_117 0 -1.8693687614478894e-05
GC_5_118 b_5 NI_5 NS_118 0 -7.4224207540062189e-06
GC_5_119 b_5 NI_5 NS_119 0 -2.5277859512197768e-04
GC_5_120 b_5 NI_5 NS_120 0 -4.4868851113488029e-03
GC_5_121 b_5 NI_5 NS_121 0 -9.9295665704392690e-06
GC_5_122 b_5 NI_5 NS_122 0 -1.0716933609920537e-05
GC_5_123 b_5 NI_5 NS_123 0 2.0753773612370210e-03
GC_5_124 b_5 NI_5 NS_124 0 2.4612096179740645e-03
GC_5_125 b_5 NI_5 NS_125 0 2.4869002600459783e-05
GC_5_126 b_5 NI_5 NS_126 0 -4.5088540019455849e-06
GC_5_127 b_5 NI_5 NS_127 0 4.0935831701061889e-06
GC_5_128 b_5 NI_5 NS_128 0 6.6436021457809100e-06
GC_5_129 b_5 NI_5 NS_129 0 -4.0065427047022509e-06
GC_5_130 b_5 NI_5 NS_130 0 1.5010664236060760e-06
GC_5_131 b_5 NI_5 NS_131 0 1.6970189876096246e-04
GC_5_132 b_5 NI_5 NS_132 0 2.9856672128604787e-04
GC_5_133 b_5 NI_5 NS_133 0 7.9090541093941188e-02
GC_5_134 b_5 NI_5 NS_134 0 -1.8753891928554770e-04
GC_5_135 b_5 NI_5 NS_135 0 -7.9628952946147122e-03
GC_5_136 b_5 NI_5 NS_136 0 -1.3312361044795426e-03
GC_5_137 b_5 NI_5 NS_137 0 4.0624094852024263e-03
GC_5_138 b_5 NI_5 NS_138 0 8.9025948184945564e-04
GC_5_139 b_5 NI_5 NS_139 0 -1.7175446087046436e-04
GC_5_140 b_5 NI_5 NS_140 0 -2.0552608256950035e-04
GC_5_141 b_5 NI_5 NS_141 0 2.2730308383067757e-03
GC_5_142 b_5 NI_5 NS_142 0 2.1453855437625455e-03
GC_5_143 b_5 NI_5 NS_143 0 -3.6129542572109208e-03
GC_5_144 b_5 NI_5 NS_144 0 8.2927294187206958e-05
GC_5_145 b_5 NI_5 NS_145 0 -6.0375578826631384e-05
GC_5_146 b_5 NI_5 NS_146 0 6.4655742876646357e-05
GC_5_147 b_5 NI_5 NS_147 0 -3.5049542923732903e-03
GC_5_148 b_5 NI_5 NS_148 0 -1.0708422063766192e-03
GC_5_149 b_5 NI_5 NS_149 0 -6.0243098756034484e-05
GC_5_150 b_5 NI_5 NS_150 0 -7.4937641487169988e-05
GC_5_151 b_5 NI_5 NS_151 0 1.2896796906850739e-04
GC_5_152 b_5 NI_5 NS_152 0 7.9264486096659490e-04
GC_5_153 b_5 NI_5 NS_153 0 3.3003245117004150e-04
GC_5_154 b_5 NI_5 NS_154 0 8.6816748608083851e-05
GC_5_155 b_5 NI_5 NS_155 0 -1.1460558907618658e-05
GC_5_156 b_5 NI_5 NS_156 0 -4.5242522289853583e-05
GC_5_157 b_5 NI_5 NS_157 0 -4.5094621889510604e-05
GC_5_158 b_5 NI_5 NS_158 0 7.2170011048356899e-05
GC_5_159 b_5 NI_5 NS_159 0 -2.2447327809589179e-03
GC_5_160 b_5 NI_5 NS_160 0 -4.1020458309214474e-03
GC_5_161 b_5 NI_5 NS_161 0 1.3778971008727520e-05
GC_5_162 b_5 NI_5 NS_162 0 3.8512360160793143e-05
GC_5_163 b_5 NI_5 NS_163 0 -7.4799408466917898e-04
GC_5_164 b_5 NI_5 NS_164 0 1.9582910047306816e-03
GC_5_165 b_5 NI_5 NS_165 0 -2.2456765588594575e-06
GC_5_166 b_5 NI_5 NS_166 0 6.3878129911746356e-06
GC_5_167 b_5 NI_5 NS_167 0 8.2569554634636863e-04
GC_5_168 b_5 NI_5 NS_168 0 -3.1208623911656254e-04
GC_5_169 b_5 NI_5 NS_169 0 -5.7576625422102723e-06
GC_5_170 b_5 NI_5 NS_170 0 -5.9278064158143056e-06
GC_5_171 b_5 NI_5 NS_171 0 1.8096092591377094e-06
GC_5_172 b_5 NI_5 NS_172 0 9.6200693185800489e-07
GC_5_173 b_5 NI_5 NS_173 0 2.2428087891106241e-06
GC_5_174 b_5 NI_5 NS_174 0 2.0329091730257411e-06
GC_5_175 b_5 NI_5 NS_175 0 1.0634100967364962e-04
GC_5_176 b_5 NI_5 NS_176 0 -1.0811605679546574e-04
GC_5_177 b_5 NI_5 NS_177 0 -3.8456946131811096e-02
GC_5_178 b_5 NI_5 NS_178 0 9.5814061555555326e-03
GC_5_179 b_5 NI_5 NS_179 0 7.6493799906160826e-03
GC_5_180 b_5 NI_5 NS_180 0 5.7441793810456190e-03
GC_5_181 b_5 NI_5 NS_181 0 8.6076412255488375e-03
GC_5_182 b_5 NI_5 NS_182 0 2.0686378237644199e-03
GC_5_183 b_5 NI_5 NS_183 0 8.1262644050416233e-04
GC_5_184 b_5 NI_5 NS_184 0 9.1524606724773449e-05
GC_5_185 b_5 NI_5 NS_185 0 1.1544344553108769e-03
GC_5_186 b_5 NI_5 NS_186 0 7.5721126809619498e-03
GC_5_187 b_5 NI_5 NS_187 0 -6.2626971072388482e-03
GC_5_188 b_5 NI_5 NS_188 0 1.4916061621861802e-03
GC_5_189 b_5 NI_5 NS_189 0 1.1402995878527294e-03
GC_5_190 b_5 NI_5 NS_190 0 4.0641770352262710e-04
GC_5_191 b_5 NI_5 NS_191 0 4.2534801013027661e-03
GC_5_192 b_5 NI_5 NS_192 0 2.0414646548285492e-03
GC_5_193 b_5 NI_5 NS_193 0 -5.3511805251271584e-05
GC_5_194 b_5 NI_5 NS_194 0 2.4218123028149456e-04
GC_5_195 b_5 NI_5 NS_195 0 -2.0724382817808472e-03
GC_5_196 b_5 NI_5 NS_196 0 -4.2349254427752041e-03
GC_5_197 b_5 NI_5 NS_197 0 -1.3638375758782562e-03
GC_5_198 b_5 NI_5 NS_198 0 8.0900049121767920e-04
GC_5_199 b_5 NI_5 NS_199 0 2.8889689461934352e-04
GC_5_200 b_5 NI_5 NS_200 0 -5.9706420541582305e-05
GC_5_201 b_5 NI_5 NS_201 0 3.9971421635026441e-05
GC_5_202 b_5 NI_5 NS_202 0 -1.5267061231940220e-04
GC_5_203 b_5 NI_5 NS_203 0 6.1987670116489943e-03
GC_5_204 b_5 NI_5 NS_204 0 1.1384055215491375e-02
GC_5_205 b_5 NI_5 NS_205 0 -2.7515882295402370e-05
GC_5_206 b_5 NI_5 NS_206 0 -2.4625761116562264e-05
GC_5_207 b_5 NI_5 NS_207 0 2.3977683675418600e-03
GC_5_208 b_5 NI_5 NS_208 0 -6.2227746184028779e-03
GC_5_209 b_5 NI_5 NS_209 0 1.2155119281200910e-06
GC_5_210 b_5 NI_5 NS_210 0 -3.1204934996252658e-05
GC_5_211 b_5 NI_5 NS_211 0 -1.3636263788745426e-03
GC_5_212 b_5 NI_5 NS_212 0 1.7061070517221176e-03
GC_5_213 b_5 NI_5 NS_213 0 3.1150972876651945e-05
GC_5_214 b_5 NI_5 NS_214 0 3.7839870360888018e-05
GC_5_215 b_5 NI_5 NS_215 0 -5.9125806847308774e-06
GC_5_216 b_5 NI_5 NS_216 0 9.2500869601109815e-06
GC_5_217 b_5 NI_5 NS_217 0 -1.7599511465735342e-06
GC_5_218 b_5 NI_5 NS_218 0 -1.3455033273787848e-05
GC_5_219 b_5 NI_5 NS_219 0 -2.9750635249231925e-04
GC_5_220 b_5 NI_5 NS_220 0 1.9931009069805385e-05
GC_5_221 b_5 NI_5 NS_221 0 3.9962027184811059e-02
GC_5_222 b_5 NI_5 NS_222 0 1.0588732470610698e-02
GC_5_223 b_5 NI_5 NS_223 0 -1.0193347271424392e-02
GC_5_224 b_5 NI_5 NS_224 0 -3.7206493005082350e-03
GC_5_225 b_5 NI_5 NS_225 0 -1.0020644056533502e-02
GC_5_226 b_5 NI_5 NS_226 0 -1.5713931515428489e-03
GC_5_227 b_5 NI_5 NS_227 0 2.4732141494451663e-04
GC_5_228 b_5 NI_5 NS_228 0 3.2125410344377810e-04
GC_5_229 b_5 NI_5 NS_229 0 3.2798571436146967e-03
GC_5_230 b_5 NI_5 NS_230 0 2.6161575250410705e-03
GC_5_231 b_5 NI_5 NS_231 0 -3.1327026533056377e-06
GC_5_232 b_5 NI_5 NS_232 0 -1.2102463877062630e-03
GC_5_233 b_5 NI_5 NS_233 0 5.6871261011407120e-05
GC_5_234 b_5 NI_5 NS_234 0 2.1753016652257322e-04
GC_5_235 b_5 NI_5 NS_235 0 3.9969428161820116e-03
GC_5_236 b_5 NI_5 NS_236 0 -7.3260214595799911e-04
GC_5_237 b_5 NI_5 NS_237 0 -6.2359911000013630e-05
GC_5_238 b_5 NI_5 NS_238 0 -5.0868083898728312e-05
GC_5_239 b_5 NI_5 NS_239 0 9.3493465713459327e-04
GC_5_240 b_5 NI_5 NS_240 0 1.0875839353701006e-03
GC_5_241 b_5 NI_5 NS_241 0 3.4693368860064228e-04
GC_5_242 b_5 NI_5 NS_242 0 -2.2630614490516665e-04
GC_5_243 b_5 NI_5 NS_243 0 1.2003658655397281e-05
GC_5_244 b_5 NI_5 NS_244 0 -3.7882926845192460e-05
GC_5_245 b_5 NI_5 NS_245 0 -3.9285558208603948e-05
GC_5_246 b_5 NI_5 NS_246 0 9.8860389115961104e-05
GC_5_247 b_5 NI_5 NS_247 0 -4.8820830484010746e-03
GC_5_248 b_5 NI_5 NS_248 0 -2.4003111667969456e-03
GC_5_249 b_5 NI_5 NS_249 0 2.1363378247568702e-05
GC_5_250 b_5 NI_5 NS_250 0 4.2602964476681926e-05
GC_5_251 b_5 NI_5 NS_251 0 1.6006805688787397e-04
GC_5_252 b_5 NI_5 NS_252 0 2.4980899428617624e-03
GC_5_253 b_5 NI_5 NS_253 0 2.4803343258633376e-06
GC_5_254 b_5 NI_5 NS_254 0 6.1212001869943332e-06
GC_5_255 b_5 NI_5 NS_255 0 5.2104534243277228e-04
GC_5_256 b_5 NI_5 NS_256 0 -1.0729617440540626e-03
GC_5_257 b_5 NI_5 NS_257 0 -1.1700289029475927e-05
GC_5_258 b_5 NI_5 NS_258 0 1.0227773336499386e-06
GC_5_259 b_5 NI_5 NS_259 0 4.1362991622832609e-07
GC_5_260 b_5 NI_5 NS_260 0 -2.5091994015230544e-07
GC_5_261 b_5 NI_5 NS_261 0 5.7644240421736841e-06
GC_5_262 b_5 NI_5 NS_262 0 -1.2770521809109405e-06
GC_5_263 b_5 NI_5 NS_263 0 3.8396977536416129e-05
GC_5_264 b_5 NI_5 NS_264 0 -3.1083180658733964e-04
GC_5_265 b_5 NI_5 NS_265 0 -2.3102765050035754e-03
GC_5_266 b_5 NI_5 NS_266 0 -5.6302554834059085e-05
GC_5_267 b_5 NI_5 NS_267 0 4.8917621372247515e-03
GC_5_268 b_5 NI_5 NS_268 0 4.5898850358825427e-03
GC_5_269 b_5 NI_5 NS_269 0 -5.2257083881593709e-03
GC_5_270 b_5 NI_5 NS_270 0 -4.9630806880663165e-03
GC_5_271 b_5 NI_5 NS_271 0 -3.1758750408598992e-05
GC_5_272 b_5 NI_5 NS_272 0 4.0982304422402822e-04
GC_5_273 b_5 NI_5 NS_273 0 1.6246603458520156e-03
GC_5_274 b_5 NI_5 NS_274 0 5.2287885909755357e-03
GC_5_275 b_5 NI_5 NS_275 0 -3.1142704505184539e-03
GC_5_276 b_5 NI_5 NS_276 0 -1.0630667122860460e-03
GC_5_277 b_5 NI_5 NS_277 0 9.4725716780622515e-04
GC_5_278 b_5 NI_5 NS_278 0 1.7721185240836477e-04
GC_5_279 b_5 NI_5 NS_279 0 -4.1398836436283828e-03
GC_5_280 b_5 NI_5 NS_280 0 -2.5394954768048314e-03
GC_5_281 b_5 NI_5 NS_281 0 -1.9713332435797364e-05
GC_5_282 b_5 NI_5 NS_282 0 1.5941970475496516e-04
GC_5_283 b_5 NI_5 NS_283 0 -2.1284931935887739e-03
GC_5_284 b_5 NI_5 NS_284 0 -2.4351069177410089e-03
GC_5_285 b_5 NI_5 NS_285 0 -1.0461556113211233e-04
GC_5_286 b_5 NI_5 NS_286 0 4.9700616758197264e-04
GC_5_287 b_5 NI_5 NS_287 0 1.8903158518676137e-04
GC_5_288 b_5 NI_5 NS_288 0 -7.4294459641910068e-05
GC_5_289 b_5 NI_5 NS_289 0 1.0810013983289087e-05
GC_5_290 b_5 NI_5 NS_290 0 -7.5591724716502943e-05
GC_5_291 b_5 NI_5 NS_291 0 6.3545869409599885e-03
GC_5_292 b_5 NI_5 NS_292 0 1.7233810253697288e-03
GC_5_293 b_5 NI_5 NS_293 0 -1.2260279587495150e-05
GC_5_294 b_5 NI_5 NS_294 0 -9.0304455070883921e-06
GC_5_295 b_5 NI_5 NS_295 0 5.8006672565003568e-04
GC_5_296 b_5 NI_5 NS_296 0 -3.3175830065427054e-03
GC_5_297 b_5 NI_5 NS_297 0 -4.5370061403508940e-07
GC_5_298 b_5 NI_5 NS_298 0 -8.1119313026556810e-06
GC_5_299 b_5 NI_5 NS_299 0 1.1037567384525532e-03
GC_5_300 b_5 NI_5 NS_300 0 8.2773916724776357e-04
GC_5_301 b_5 NI_5 NS_301 0 1.0500685485364173e-05
GC_5_302 b_5 NI_5 NS_302 0 6.2650302569019120e-06
GC_5_303 b_5 NI_5 NS_303 0 6.7421289916027836e-07
GC_5_304 b_5 NI_5 NS_304 0 4.8437550747881798e-06
GC_5_305 b_5 NI_5 NS_305 0 -1.2318448452316107e-06
GC_5_306 b_5 NI_5 NS_306 0 -1.3055735652838377e-06
GC_5_307 b_5 NI_5 NS_307 0 3.2270008807814667e-05
GC_5_308 b_5 NI_5 NS_308 0 6.8860284938117319e-05
GC_5_309 b_5 NI_5 NS_309 0 6.0421197831496125e-02
GC_5_310 b_5 NI_5 NS_310 0 -3.6827372954720063e-05
GC_5_311 b_5 NI_5 NS_311 0 -6.2389308912164324e-03
GC_5_312 b_5 NI_5 NS_312 0 -2.7366714951562571e-03
GC_5_313 b_5 NI_5 NS_313 0 4.3480874691867316e-03
GC_5_314 b_5 NI_5 NS_314 0 2.6774408416624525e-03
GC_5_315 b_5 NI_5 NS_315 0 1.1678547753811451e-05
GC_5_316 b_5 NI_5 NS_316 0 -1.7177681619933382e-04
GC_5_317 b_5 NI_5 NS_317 0 1.4030047731868240e-03
GC_5_318 b_5 NI_5 NS_318 0 1.5327719107916663e-03
GC_5_319 b_5 NI_5 NS_319 0 -1.6524998007451012e-04
GC_5_320 b_5 NI_5 NS_320 0 -5.5449878908086646e-04
GC_5_321 b_5 NI_5 NS_321 0 -4.4222879919293256e-05
GC_5_322 b_5 NI_5 NS_322 0 8.2932074075072327e-05
GC_5_323 b_5 NI_5 NS_323 0 -3.9348491179489655e-03
GC_5_324 b_5 NI_5 NS_324 0 9.0024826912425899e-04
GC_5_325 b_5 NI_5 NS_325 0 -7.6706357745706587e-05
GC_5_326 b_5 NI_5 NS_326 0 -4.7530693257353095e-05
GC_5_327 b_5 NI_5 NS_327 0 -2.6253121756213946e-04
GC_5_328 b_5 NI_5 NS_328 0 7.8548584460573522e-04
GC_5_329 b_5 NI_5 NS_329 0 3.7693847907946647e-04
GC_5_330 b_5 NI_5 NS_330 0 7.5655003878155995e-05
GC_5_331 b_5 NI_5 NS_331 0 -2.9752808522482495e-05
GC_5_332 b_5 NI_5 NS_332 0 -4.3987289641949176e-05
GC_5_333 b_5 NI_5 NS_333 0 -3.6114408051746811e-05
GC_5_334 b_5 NI_5 NS_334 0 7.8741547466039323e-05
GC_5_335 b_5 NI_5 NS_335 0 -2.9776567213243206e-03
GC_5_336 b_5 NI_5 NS_336 0 -3.4609542512370420e-03
GC_5_337 b_5 NI_5 NS_337 0 9.4828012768645293e-06
GC_5_338 b_5 NI_5 NS_338 0 2.7662340654252481e-05
GC_5_339 b_5 NI_5 NS_339 0 -5.0479588627622639e-04
GC_5_340 b_5 NI_5 NS_340 0 1.9356741741823646e-03
GC_5_341 b_5 NI_5 NS_341 0 -2.3893783596952559e-07
GC_5_342 b_5 NI_5 NS_342 0 8.3496619147057847e-06
GC_5_343 b_5 NI_5 NS_343 0 8.4947825682599306e-04
GC_5_344 b_5 NI_5 NS_344 0 -4.7265474842607868e-04
GC_5_345 b_5 NI_5 NS_345 0 -1.0503840231802794e-05
GC_5_346 b_5 NI_5 NS_346 0 -8.1324124595990232e-06
GC_5_347 b_5 NI_5 NS_347 0 1.6478068579582161e-06
GC_5_348 b_5 NI_5 NS_348 0 -1.8081853757228395e-07
GC_5_349 b_5 NI_5 NS_349 0 2.8189705286376191e-06
GC_5_350 b_5 NI_5 NS_350 0 2.2727648657738798e-06
GC_5_351 b_5 NI_5 NS_351 0 9.6821179203479760e-05
GC_5_352 b_5 NI_5 NS_352 0 -1.1669203142000675e-04
GC_5_353 b_5 NI_5 NS_353 0 2.4139312687904996e-03
GC_5_354 b_5 NI_5 NS_354 0 9.6680950481903852e-05
GC_5_355 b_5 NI_5 NS_355 0 3.1994561853517070e-04
GC_5_356 b_5 NI_5 NS_356 0 -8.7100380895429371e-04
GC_5_357 b_5 NI_5 NS_357 0 7.1087236294905621e-04
GC_5_358 b_5 NI_5 NS_358 0 1.4391781267747540e-05
GC_5_359 b_5 NI_5 NS_359 0 -7.3534902539577776e-04
GC_5_360 b_5 NI_5 NS_360 0 -1.4673971988368988e-04
GC_5_361 b_5 NI_5 NS_361 0 1.0990118954384896e-03
GC_5_362 b_5 NI_5 NS_362 0 -3.1185214881388860e-05
GC_5_363 b_5 NI_5 NS_363 0 -2.7438275141884118e-03
GC_5_364 b_5 NI_5 NS_364 0 -1.1079316845945687e-03
GC_5_365 b_5 NI_5 NS_365 0 5.9680753538581476e-04
GC_5_366 b_5 NI_5 NS_366 0 -6.5920999095061487e-04
GC_5_367 b_5 NI_5 NS_367 0 8.5310220433374457e-03
GC_5_368 b_5 NI_5 NS_368 0 -1.5952180219669157e-03
GC_5_369 b_5 NI_5 NS_369 0 4.2746865750881093e-04
GC_5_370 b_5 NI_5 NS_370 0 3.7746972261496961e-04
GC_5_371 b_5 NI_5 NS_371 0 2.6330902542843191e-04
GC_5_372 b_5 NI_5 NS_372 0 3.6143004478172967e-03
GC_5_373 b_5 NI_5 NS_373 0 6.5053959467030258e-04
GC_5_374 b_5 NI_5 NS_374 0 -2.3888047970593203e-04
GC_5_375 b_5 NI_5 NS_375 0 2.1942958590474748e-04
GC_5_376 b_5 NI_5 NS_376 0 -3.3735988990458384e-05
GC_5_377 b_5 NI_5 NS_377 0 3.3614712092204545e-05
GC_5_378 b_5 NI_5 NS_378 0 1.2776920490727245e-04
GC_5_379 b_5 NI_5 NS_379 0 -8.7398808234879066e-03
GC_5_380 b_5 NI_5 NS_380 0 8.3619022200427055e-03
GC_5_381 b_5 NI_5 NS_381 0 1.8693432768392749e-05
GC_5_382 b_5 NI_5 NS_382 0 -2.0149242822077061e-05
GC_5_383 b_5 NI_5 NS_383 0 2.5892110784207518e-03
GC_5_384 b_5 NI_5 NS_384 0 -6.9767556815147284e-04
GC_5_385 b_5 NI_5 NS_385 0 -3.4587537048955583e-07
GC_5_386 b_5 NI_5 NS_386 0 8.7176429314881436e-06
GC_5_387 b_5 NI_5 NS_387 0 -1.3654485375687043e-04
GC_5_388 b_5 NI_5 NS_388 0 -2.7337224861056567e-03
GC_5_389 b_5 NI_5 NS_389 0 -2.0591606493928745e-05
GC_5_390 b_5 NI_5 NS_390 0 -1.6458114477610213e-06
GC_5_391 b_5 NI_5 NS_391 0 2.4308058031548395e-07
GC_5_392 b_5 NI_5 NS_392 0 -2.1701123792235827e-06
GC_5_393 b_5 NI_5 NS_393 0 3.0566742261178208e-06
GC_5_394 b_5 NI_5 NS_394 0 3.7661484469844031e-06
GC_5_395 b_5 NI_5 NS_395 0 -5.1317205501389211e-05
GC_5_396 b_5 NI_5 NS_396 0 -9.0248529435821637e-04
GC_5_397 b_5 NI_5 NS_397 0 -7.1088849105676287e-04
GC_5_398 b_5 NI_5 NS_398 0 -1.0290584205003197e-05
GC_5_399 b_5 NI_5 NS_399 0 -4.1250910329876584e-04
GC_5_400 b_5 NI_5 NS_400 0 4.7815803778606113e-04
GC_5_401 b_5 NI_5 NS_401 0 -3.9399575878955941e-04
GC_5_402 b_5 NI_5 NS_402 0 -7.2278800105064094e-04
GC_5_403 b_5 NI_5 NS_403 0 1.7080006446896256e-04
GC_5_404 b_5 NI_5 NS_404 0 9.8664442876759343e-05
GC_5_405 b_5 NI_5 NS_405 0 3.6260541168672931e-04
GC_5_406 b_5 NI_5 NS_406 0 -4.4679531492165271e-04
GC_5_407 b_5 NI_5 NS_407 0 -1.3702939240224171e-04
GC_5_408 b_5 NI_5 NS_408 0 -3.3659294258125516e-04
GC_5_409 b_5 NI_5 NS_409 0 1.4010813851232366e-04
GC_5_410 b_5 NI_5 NS_410 0 9.8537587419989924e-05
GC_5_411 b_5 NI_5 NS_411 0 6.2326444065433832e-04
GC_5_412 b_5 NI_5 NS_412 0 7.9136181573167381e-04
GC_5_413 b_5 NI_5 NS_413 0 -1.7591874792000900e-04
GC_5_414 b_5 NI_5 NS_414 0 8.9003469355352776e-05
GC_5_415 b_5 NI_5 NS_415 0 -6.3010392097129339e-04
GC_5_416 b_5 NI_5 NS_416 0 -2.6044385106976562e-04
GC_5_417 b_5 NI_5 NS_417 0 1.0028196392698200e-05
GC_5_418 b_5 NI_5 NS_418 0 -5.0794922494728464e-06
GC_5_419 b_5 NI_5 NS_419 0 -3.2384806390931528e-05
GC_5_420 b_5 NI_5 NS_420 0 -1.6288168404798959e-04
GC_5_421 b_5 NI_5 NS_421 0 -2.7079363306113395e-06
GC_5_422 b_5 NI_5 NS_422 0 1.3740897235138739e-04
GC_5_423 b_5 NI_5 NS_423 0 1.7623174796124856e-03
GC_5_424 b_5 NI_5 NS_424 0 5.1534815168764530e-04
GC_5_425 b_5 NI_5 NS_425 0 -3.4570806902412952e-05
GC_5_426 b_5 NI_5 NS_426 0 -1.2429379872401744e-05
GC_5_427 b_5 NI_5 NS_427 0 -6.0693986847044717e-04
GC_5_428 b_5 NI_5 NS_428 0 -6.4955916960114527e-04
GC_5_429 b_5 NI_5 NS_429 0 -3.0075113568137578e-07
GC_5_430 b_5 NI_5 NS_430 0 2.8853001137391853e-06
GC_5_431 b_5 NI_5 NS_431 0 -1.6611803705107836e-04
GC_5_432 b_5 NI_5 NS_432 0 -1.9127878199285504e-04
GC_5_433 b_5 NI_5 NS_433 0 -1.5211829052331083e-05
GC_5_434 b_5 NI_5 NS_434 0 -2.1541416894135329e-05
GC_5_435 b_5 NI_5 NS_435 0 -1.1816764535421973e-07
GC_5_436 b_5 NI_5 NS_436 0 2.7174551912528279e-06
GC_5_437 b_5 NI_5 NS_437 0 -1.9245062661824920e-06
GC_5_438 b_5 NI_5 NS_438 0 -2.3028589209896225e-06
GC_5_439 b_5 NI_5 NS_439 0 -3.4362024833763745e-04
GC_5_440 b_5 NI_5 NS_440 0 -2.5267490539171112e-05
GC_5_441 b_5 NI_5 NS_441 0 4.8740243414620308e-03
GC_5_442 b_5 NI_5 NS_442 0 8.2133775933265985e-05
GC_5_443 b_5 NI_5 NS_443 0 1.2174357505631422e-03
GC_5_444 b_5 NI_5 NS_444 0 -2.8692723051254566e-04
GC_5_445 b_5 NI_5 NS_445 0 -6.2843474003004157e-04
GC_5_446 b_5 NI_5 NS_446 0 4.4929006328386570e-04
GC_5_447 b_5 NI_5 NS_447 0 -3.4540408631566049e-05
GC_5_448 b_5 NI_5 NS_448 0 -3.2219075221820540e-04
GC_5_449 b_5 NI_5 NS_449 0 8.3501548966014353e-04
GC_5_450 b_5 NI_5 NS_450 0 6.1005908877900176e-04
GC_5_451 b_5 NI_5 NS_451 0 -2.5776192570601854e-03
GC_5_452 b_5 NI_5 NS_452 0 -1.6176696481261608e-03
GC_5_453 b_5 NI_5 NS_453 0 5.6361992128378940e-04
GC_5_454 b_5 NI_5 NS_454 0 -4.2454792676631397e-04
GC_5_455 b_5 NI_5 NS_455 0 4.8135801902980807e-03
GC_5_456 b_5 NI_5 NS_456 0 2.5417996989340636e-04
GC_5_457 b_5 NI_5 NS_457 0 2.6020828746912647e-04
GC_5_458 b_5 NI_5 NS_458 0 2.9165246152071085e-04
GC_5_459 b_5 NI_5 NS_459 0 -2.1076434916729737e-04
GC_5_460 b_5 NI_5 NS_460 0 2.0647333764686492e-03
GC_5_461 b_5 NI_5 NS_461 0 3.3049505127314327e-04
GC_5_462 b_5 NI_5 NS_462 0 -2.8507368560661781e-04
GC_5_463 b_5 NI_5 NS_463 0 1.6354465160810084e-04
GC_5_464 b_5 NI_5 NS_464 0 -3.4625689173347250e-05
GC_5_465 b_5 NI_5 NS_465 0 2.3300170921264969e-05
GC_5_466 b_5 NI_5 NS_466 0 8.0327766767791410e-05
GC_5_467 b_5 NI_5 NS_467 0 -5.3876956411268925e-03
GC_5_468 b_5 NI_5 NS_468 0 4.4054534284285757e-03
GC_5_469 b_5 NI_5 NS_469 0 7.3753179782482502e-06
GC_5_470 b_5 NI_5 NS_470 0 -8.5812508503662017e-06
GC_5_471 b_5 NI_5 NS_471 0 1.5140669367755156e-03
GC_5_472 b_5 NI_5 NS_472 0 -6.7750671415452775e-04
GC_5_473 b_5 NI_5 NS_473 0 -1.6866880359158633e-07
GC_5_474 b_5 NI_5 NS_474 0 2.8600671414401324e-06
GC_5_475 b_5 NI_5 NS_475 0 -9.7868658616219280e-05
GC_5_476 b_5 NI_5 NS_476 0 -1.8748906601346552e-03
GC_5_477 b_5 NI_5 NS_477 0 -1.3227272428234349e-05
GC_5_478 b_5 NI_5 NS_478 0 2.6824782585082586e-06
GC_5_479 b_5 NI_5 NS_479 0 4.9111115756478873e-07
GC_5_480 b_5 NI_5 NS_480 0 -4.2338703000707321e-07
GC_5_481 b_5 NI_5 NS_481 0 1.0530280974965416e-06
GC_5_482 b_5 NI_5 NS_482 0 2.3016437855836697e-06
GC_5_483 b_5 NI_5 NS_483 0 -2.0012229930578792e-05
GC_5_484 b_5 NI_5 NS_484 0 -5.5318162044055974e-04
GC_5_485 b_5 NI_5 NS_485 0 -5.7455593048132856e-03
GC_5_486 b_5 NI_5 NS_486 0 -1.3716215621579276e-05
GC_5_487 b_5 NI_5 NS_487 0 -1.2902669175307905e-03
GC_5_488 b_5 NI_5 NS_488 0 1.8771742178124549e-04
GC_5_489 b_5 NI_5 NS_489 0 6.4514523678001602e-04
GC_5_490 b_5 NI_5 NS_490 0 -1.2038987595191445e-03
GC_5_491 b_5 NI_5 NS_491 0 2.1272691424110206e-04
GC_5_492 b_5 NI_5 NS_492 0 3.4674124185271040e-04
GC_5_493 b_5 NI_5 NS_493 0 6.6254640754180691e-04
GC_5_494 b_5 NI_5 NS_494 0 -1.1137056874215373e-04
GC_5_495 b_5 NI_5 NS_495 0 -2.1909421257070876e-04
GC_5_496 b_5 NI_5 NS_496 0 -1.0971104498881318e-03
GC_5_497 b_5 NI_5 NS_497 0 1.1271902698829315e-04
GC_5_498 b_5 NI_5 NS_498 0 1.0158079417607240e-04
GC_5_499 b_5 NI_5 NS_499 0 7.7218349984786543e-04
GC_5_500 b_5 NI_5 NS_500 0 1.1535193279813092e-03
GC_5_501 b_5 NI_5 NS_501 0 -1.0184549197056253e-04
GC_5_502 b_5 NI_5 NS_502 0 4.1168523306404628e-05
GC_5_503 b_5 NI_5 NS_503 0 -2.2789404980754876e-04
GC_5_504 b_5 NI_5 NS_504 0 -5.7001304019747188e-05
GC_5_505 b_5 NI_5 NS_505 0 4.3656688892071348e-05
GC_5_506 b_5 NI_5 NS_506 0 7.3423703404103225e-05
GC_5_507 b_5 NI_5 NS_507 0 -1.5631560600456247e-05
GC_5_508 b_5 NI_5 NS_508 0 -8.6266448429855549e-05
GC_5_509 b_5 NI_5 NS_509 0 -5.6545615455229681e-06
GC_5_510 b_5 NI_5 NS_510 0 8.0449816916865400e-05
GC_5_511 b_5 NI_5 NS_511 0 1.2320690702655051e-03
GC_5_512 b_5 NI_5 NS_512 0 -1.1378689725304187e-04
GC_5_513 b_5 NI_5 NS_513 0 -1.8359328859453610e-05
GC_5_514 b_5 NI_5 NS_514 0 -1.7125560047858077e-06
GC_5_515 b_5 NI_5 NS_515 0 -4.6257679591309072e-04
GC_5_516 b_5 NI_5 NS_516 0 -2.2343191874938216e-04
GC_5_517 b_5 NI_5 NS_517 0 -9.6214933178157316e-07
GC_5_518 b_5 NI_5 NS_518 0 1.7060879724194057e-06
GC_5_519 b_5 NI_5 NS_519 0 5.5096224065722935e-05
GC_5_520 b_5 NI_5 NS_520 0 7.9463084773843410e-06
GC_5_521 b_5 NI_5 NS_521 0 -5.7752551925015270e-06
GC_5_522 b_5 NI_5 NS_522 0 -1.0983567741154812e-05
GC_5_523 b_5 NI_5 NS_523 0 -8.6041549642901027e-08
GC_5_524 b_5 NI_5 NS_524 0 1.4999175527637077e-06
GC_5_525 b_5 NI_5 NS_525 0 -7.6507448085130989e-07
GC_5_526 b_5 NI_5 NS_526 0 -8.2473616905741955e-07
GC_5_527 b_5 NI_5 NS_527 0 -1.4442635117720728e-04
GC_5_528 b_5 NI_5 NS_528 0 -7.1193339673344635e-06
GD_5_1 b_5 NI_5 NA_1 0 -2.7144956678917524e-02
GD_5_2 b_5 NI_5 NA_2 0 -3.8919846984815723e-02
GD_5_3 b_5 NI_5 NA_3 0 -2.4863362120855904e-03
GD_5_4 b_5 NI_5 NA_4 0 -8.1131772018049497e-02
GD_5_5 b_5 NI_5 NA_5 0 -1.2762615838889130e-01
GD_5_6 b_5 NI_5 NA_6 0 -4.5682579115351507e-02
GD_5_7 b_5 NI_5 NA_7 0 3.1661145472940107e-03
GD_5_8 b_5 NI_5 NA_8 0 -6.4533380289607173e-02
GD_5_9 b_5 NI_5 NA_9 0 -1.0163011055352394e-02
GD_5_10 b_5 NI_5 NA_10 0 2.3233316772011231e-04
GD_5_11 b_5 NI_5 NA_11 0 -8.5027406839015690e-03
GD_5_12 b_5 NI_5 NA_12 0 3.8252618377322013e-03
*
* Port 6
VI_6 a_6 NI_6 0
RI_6 NI_6 b_6 5.0000000000000000e+01
GC_6_1 b_6 NI_6 NS_1 0 3.9830603410147818e-02
GC_6_2 b_6 NI_6 NS_2 0 -2.4322542854890260e-04
GC_6_3 b_6 NI_6 NS_3 0 -5.7110893755099364e-03
GC_6_4 b_6 NI_6 NS_4 0 7.2542276901784418e-04
GC_6_5 b_6 NI_6 NS_5 0 2.5474744467541845e-03
GC_6_6 b_6 NI_6 NS_6 0 -2.5373687858914425e-03
GC_6_7 b_6 NI_6 NS_7 0 -1.4254927959627729e-04
GC_6_8 b_6 NI_6 NS_8 0 -9.8480190854557357e-05
GC_6_9 b_6 NI_6 NS_9 0 2.2444319478208282e-03
GC_6_10 b_6 NI_6 NS_10 0 1.5038716765943100e-03
GC_6_11 b_6 NI_6 NS_11 0 -3.9323770329617860e-03
GC_6_12 b_6 NI_6 NS_12 0 -2.6470139855919552e-04
GC_6_13 b_6 NI_6 NS_13 0 4.0227174862792031e-05
GC_6_14 b_6 NI_6 NS_14 0 4.4920581904286438e-05
GC_6_15 b_6 NI_6 NS_15 0 -5.2289784528911922e-04
GC_6_16 b_6 NI_6 NS_16 0 4.9940666470567543e-05
GC_6_17 b_6 NI_6 NS_17 0 -3.9921698099398038e-05
GC_6_18 b_6 NI_6 NS_18 0 -6.7229226927963443e-05
GC_6_19 b_6 NI_6 NS_19 0 3.7977461246309130e-04
GC_6_20 b_6 NI_6 NS_20 0 6.0672558278264594e-04
GC_6_21 b_6 NI_6 NS_21 0 2.6790942005904233e-04
GC_6_22 b_6 NI_6 NS_22 0 9.6544193171171593e-05
GC_6_23 b_6 NI_6 NS_23 0 6.6752439891905742e-06
GC_6_24 b_6 NI_6 NS_24 0 -4.0602730927540927e-05
GC_6_25 b_6 NI_6 NS_25 0 -4.8598436737337434e-05
GC_6_26 b_6 NI_6 NS_26 0 6.2512102454711423e-05
GC_6_27 b_6 NI_6 NS_27 0 -1.3971105484155055e-03
GC_6_28 b_6 NI_6 NS_28 0 -3.7813793880914167e-03
GC_6_29 b_6 NI_6 NS_29 0 1.2454946635133655e-05
GC_6_30 b_6 NI_6 NS_30 0 3.7793609041316060e-05
GC_6_31 b_6 NI_6 NS_31 0 -7.5664292325571252e-04
GC_6_32 b_6 NI_6 NS_32 0 1.7285494982454852e-03
GC_6_33 b_6 NI_6 NS_33 0 -2.0679609820440022e-06
GC_6_34 b_6 NI_6 NS_34 0 4.9619035873791856e-06
GC_6_35 b_6 NI_6 NS_35 0 8.0168064245103262e-04
GC_6_36 b_6 NI_6 NS_36 0 -1.1023020662863690e-04
GC_6_37 b_6 NI_6 NS_37 0 -3.9683682353189376e-06
GC_6_38 b_6 NI_6 NS_38 0 -7.6300296415848966e-06
GC_6_39 b_6 NI_6 NS_39 0 1.5154235559745067e-06
GC_6_40 b_6 NI_6 NS_40 0 1.3076496074384342e-06
GC_6_41 b_6 NI_6 NS_41 0 3.0137216617609802e-07
GC_6_42 b_6 NI_6 NS_42 0 4.8592073733667445e-07
GC_6_43 b_6 NI_6 NS_43 0 8.3304624315719009e-05
GC_6_44 b_6 NI_6 NS_44 0 -1.1370974194841250e-04
GC_6_45 b_6 NI_6 NS_45 0 1.0174600218954685e-02
GC_6_46 b_6 NI_6 NS_46 0 -2.8650416274633413e-04
GC_6_47 b_6 NI_6 NS_47 0 3.9837980473669907e-03
GC_6_48 b_6 NI_6 NS_48 0 -1.4862491485228783e-03
GC_6_49 b_6 NI_6 NS_49 0 -1.9750021259970557e-03
GC_6_50 b_6 NI_6 NS_50 0 2.5692173911406116e-03
GC_6_51 b_6 NI_6 NS_51 0 -4.0285519048554409e-04
GC_6_52 b_6 NI_6 NS_52 0 5.4624486755165582e-04
GC_6_53 b_6 NI_6 NS_53 0 1.0533751763619975e-03
GC_6_54 b_6 NI_6 NS_54 0 3.9215571415958302e-04
GC_6_55 b_6 NI_6 NS_55 0 -8.0041842152921031e-04
GC_6_56 b_6 NI_6 NS_56 0 1.5810096051209783e-03
GC_6_57 b_6 NI_6 NS_57 0 -7.2381194506060466e-05
GC_6_58 b_6 NI_6 NS_58 0 -1.1174353923413688e-05
GC_6_59 b_6 NI_6 NS_59 0 -8.1638383083086142e-04
GC_6_60 b_6 NI_6 NS_60 0 1.6523830354099010e-03
GC_6_61 b_6 NI_6 NS_61 0 5.3324304212695666e-06
GC_6_62 b_6 NI_6 NS_62 0 -9.9047558826837007e-06
GC_6_63 b_6 NI_6 NS_63 0 -5.7076756896376067e-04
GC_6_64 b_6 NI_6 NS_64 0 3.5892225165992783e-04
GC_6_65 b_6 NI_6 NS_65 0 8.0492513267018480e-04
GC_6_66 b_6 NI_6 NS_66 0 -2.5425679866022830e-04
GC_6_67 b_6 NI_6 NS_67 0 -5.0150945571990952e-05
GC_6_68 b_6 NI_6 NS_68 0 -2.0214685123216745e-05
GC_6_69 b_6 NI_6 NS_69 0 -6.4779125500343988e-05
GC_6_70 b_6 NI_6 NS_70 0 -8.3375408565885056e-05
GC_6_71 b_6 NI_6 NS_71 0 -1.9983725866581110e-03
GC_6_72 b_6 NI_6 NS_72 0 -4.0871062302356110e-03
GC_6_73 b_6 NI_6 NS_73 0 -3.7151760291355864e-05
GC_6_74 b_6 NI_6 NS_74 0 -4.0640124263546837e-05
GC_6_75 b_6 NI_6 NS_75 0 4.6431047556514673e-04
GC_6_76 b_6 NI_6 NS_76 0 1.1400822470250963e-03
GC_6_77 b_6 NI_6 NS_77 0 -1.1854253224864280e-05
GC_6_78 b_6 NI_6 NS_78 0 2.8311009771546935e-05
GC_6_79 b_6 NI_6 NS_79 0 1.3271215909218361e-03
GC_6_80 b_6 NI_6 NS_80 0 -5.6138040441624495e-04
GC_6_81 b_6 NI_6 NS_81 0 -1.6263062673830376e-05
GC_6_82 b_6 NI_6 NS_82 0 -2.1206591784042912e-05
GC_6_83 b_6 NI_6 NS_83 0 2.8840060827294480e-05
GC_6_84 b_6 NI_6 NS_84 0 -5.1580401547823156e-06
GC_6_85 b_6 NI_6 NS_85 0 3.6899101272443611e-05
GC_6_86 b_6 NI_6 NS_86 0 -1.3010675946513801e-05
GC_6_87 b_6 NI_6 NS_87 0 -2.4542530501047832e-05
GC_6_88 b_6 NI_6 NS_88 0 1.0909947822692387e-04
GC_6_89 b_6 NI_6 NS_89 0 8.1634989487190543e-02
GC_6_90 b_6 NI_6 NS_90 0 -1.7855520848885707e-04
GC_6_91 b_6 NI_6 NS_91 0 -8.1217039938947574e-03
GC_6_92 b_6 NI_6 NS_92 0 -1.4130427046941366e-03
GC_6_93 b_6 NI_6 NS_93 0 4.3646354929183636e-03
GC_6_94 b_6 NI_6 NS_94 0 7.2119099458071458e-04
GC_6_95 b_6 NI_6 NS_95 0 -1.8113522918444773e-04
GC_6_96 b_6 NI_6 NS_96 0 -1.6145934090534071e-04
GC_6_97 b_6 NI_6 NS_97 0 2.5751373575947124e-03
GC_6_98 b_6 NI_6 NS_98 0 2.0530627791015142e-03
GC_6_99 b_6 NI_6 NS_99 0 -3.6491066352041883e-03
GC_6_100 b_6 NI_6 NS_100 0 7.0375491691996610e-05
GC_6_101 b_6 NI_6 NS_101 0 2.6301012340195487e-06
GC_6_102 b_6 NI_6 NS_102 0 8.5417228931749777e-05
GC_6_103 b_6 NI_6 NS_103 0 -2.8536830694483981e-03
GC_6_104 b_6 NI_6 NS_104 0 -4.3976365300399655e-04
GC_6_105 b_6 NI_6 NS_105 0 -7.1372657804810426e-05
GC_6_106 b_6 NI_6 NS_106 0 -9.3882816993163273e-05
GC_6_107 b_6 NI_6 NS_107 0 3.2933766697634917e-04
GC_6_108 b_6 NI_6 NS_108 0 1.1937540401921708e-03
GC_6_109 b_6 NI_6 NS_109 0 2.9779979134300410e-04
GC_6_110 b_6 NI_6 NS_110 0 6.9897393737391878e-05
GC_6_111 b_6 NI_6 NS_111 0 -1.0138278225086331e-05
GC_6_112 b_6 NI_6 NS_112 0 -5.8810761896895306e-05
GC_6_113 b_6 NI_6 NS_113 0 -7.3616762325398453e-05
GC_6_114 b_6 NI_6 NS_114 0 9.6077852787415318e-05
GC_6_115 b_6 NI_6 NS_115 0 -3.5047392211565729e-03
GC_6_116 b_6 NI_6 NS_116 0 -4.6442490854770938e-03
GC_6_117 b_6 NI_6 NS_117 0 1.5227540021690968e-05
GC_6_118 b_6 NI_6 NS_118 0 5.2820572140949044e-05
GC_6_119 b_6 NI_6 NS_119 0 -6.9522072569494020e-04
GC_6_120 b_6 NI_6 NS_120 0 2.6562085571492249e-03
GC_6_121 b_6 NI_6 NS_121 0 1.6594180217862189e-06
GC_6_122 b_6 NI_6 NS_122 0 1.0312508174849725e-05
GC_6_123 b_6 NI_6 NS_123 0 9.8502296552702476e-04
GC_6_124 b_6 NI_6 NS_124 0 -5.1952539190437750e-04
GC_6_125 b_6 NI_6 NS_125 0 -1.1041367157635248e-05
GC_6_126 b_6 NI_6 NS_126 0 -6.1479352927901222e-06
GC_6_127 b_6 NI_6 NS_127 0 2.4642040308282564e-06
GC_6_128 b_6 NI_6 NS_128 0 -1.0710691384717275e-06
GC_6_129 b_6 NI_6 NS_129 0 1.5538657259898591e-06
GC_6_130 b_6 NI_6 NS_130 0 -1.9821850099313737e-06
GC_6_131 b_6 NI_6 NS_131 0 1.2731390756076059e-04
GC_6_132 b_6 NI_6 NS_132 0 -1.9349184096370106e-04
GC_6_133 b_6 NI_6 NS_133 0 1.4868737219190844e-02
GC_6_134 b_6 NI_6 NS_134 0 -9.0521683784051509e-04
GC_6_135 b_6 NI_6 NS_135 0 5.1923134121647334e-03
GC_6_136 b_6 NI_6 NS_136 0 1.8804578979169832e-04
GC_6_137 b_6 NI_6 NS_137 0 -4.6846850536250758e-03
GC_6_138 b_6 NI_6 NS_138 0 -4.6334876493114185e-04
GC_6_139 b_6 NI_6 NS_139 0 -4.6875297217060257e-05
GC_6_140 b_6 NI_6 NS_140 0 3.5920032473963666e-04
GC_6_141 b_6 NI_6 NS_141 0 1.7419991386864232e-03
GC_6_142 b_6 NI_6 NS_142 0 4.6910729608585686e-04
GC_6_143 b_6 NI_6 NS_143 0 -5.9872156819448634e-04
GC_6_144 b_6 NI_6 NS_144 0 7.8370106566356501e-04
GC_6_145 b_6 NI_6 NS_145 0 -4.4853720878413514e-05
GC_6_146 b_6 NI_6 NS_146 0 -2.7051728445257702e-05
GC_6_147 b_6 NI_6 NS_147 0 -1.0481874246076844e-03
GC_6_148 b_6 NI_6 NS_148 0 7.5893148745671780e-04
GC_6_149 b_6 NI_6 NS_149 0 2.8066215583145067e-05
GC_6_150 b_6 NI_6 NS_150 0 -1.0508975054603258e-05
GC_6_151 b_6 NI_6 NS_151 0 4.0160463309880764e-05
GC_6_152 b_6 NI_6 NS_152 0 1.8963418027127465e-04
GC_6_153 b_6 NI_6 NS_153 0 5.9498363634590706e-04
GC_6_154 b_6 NI_6 NS_154 0 -3.3226303041736943e-04
GC_6_155 b_6 NI_6 NS_155 0 -2.1053218621853619e-05
GC_6_156 b_6 NI_6 NS_156 0 -2.2314748186781000e-05
GC_6_157 b_6 NI_6 NS_157 0 -6.1132345286946642e-05
GC_6_158 b_6 NI_6 NS_158 0 -1.1441393126431592e-04
GC_6_159 b_6 NI_6 NS_159 0 -1.0164192132145632e-03
GC_6_160 b_6 NI_6 NS_160 0 -9.4331324072360542e-04
GC_6_161 b_6 NI_6 NS_161 0 -4.4329838532056313e-05
GC_6_162 b_6 NI_6 NS_162 0 -5.1218545212960035e-05
GC_6_163 b_6 NI_6 NS_163 0 1.2063597037327480e-03
GC_6_164 b_6 NI_6 NS_164 0 1.2515559041430873e-04
GC_6_165 b_6 NI_6 NS_165 0 -9.0752223173963567e-06
GC_6_166 b_6 NI_6 NS_166 0 2.2441912691963291e-05
GC_6_167 b_6 NI_6 NS_167 0 7.0128225278336934e-04
GC_6_168 b_6 NI_6 NS_168 0 -4.7774977648062440e-04
GC_6_169 b_6 NI_6 NS_169 0 -8.6518861492922990e-06
GC_6_170 b_6 NI_6 NS_170 0 -1.1605988735471779e-05
GC_6_171 b_6 NI_6 NS_171 0 3.0259247741440890e-05
GC_6_172 b_6 NI_6 NS_172 0 -3.0790805659628177e-06
GC_6_173 b_6 NI_6 NS_173 0 3.8686884746829200e-05
GC_6_174 b_6 NI_6 NS_174 0 -1.5074008811312458e-05
GC_6_175 b_6 NI_6 NS_175 0 -1.4550123730524067e-04
GC_6_176 b_6 NI_6 NS_176 0 8.3127541719150270e-05
GC_6_177 b_6 NI_6 NS_177 0 3.9962027181927824e-02
GC_6_178 b_6 NI_6 NS_178 0 1.0588732470662204e-02
GC_6_179 b_6 NI_6 NS_179 0 -1.0193347271344862e-02
GC_6_180 b_6 NI_6 NS_180 0 -3.7206493006669743e-03
GC_6_181 b_6 NI_6 NS_181 0 -1.0020644056348359e-02
GC_6_182 b_6 NI_6 NS_182 0 -1.5713931515257721e-03
GC_6_183 b_6 NI_6 NS_183 0 2.4732141498164952e-04
GC_6_184 b_6 NI_6 NS_184 0 3.2125410369983012e-04
GC_6_185 b_6 NI_6 NS_185 0 3.2798571436834186e-03
GC_6_186 b_6 NI_6 NS_186 0 2.6161575250191718e-03
GC_6_187 b_6 NI_6 NS_187 0 -3.1327026197680793e-06
GC_6_188 b_6 NI_6 NS_188 0 -1.2102463879049125e-03
GC_6_189 b_6 NI_6 NS_189 0 5.6871261025697176e-05
GC_6_190 b_6 NI_6 NS_190 0 2.1753016652436286e-04
GC_6_191 b_6 NI_6 NS_191 0 3.9969428165071760e-03
GC_6_192 b_6 NI_6 NS_192 0 -7.3260214614694421e-04
GC_6_193 b_6 NI_6 NS_193 0 -6.2359910994036613e-05
GC_6_194 b_6 NI_6 NS_194 0 -5.0868083896777622e-05
GC_6_195 b_6 NI_6 NS_195 0 9.3493465729481179e-04
GC_6_196 b_6 NI_6 NS_196 0 1.0875839353178427e-03
GC_6_197 b_6 NI_6 NS_197 0 3.4693368855255775e-04
GC_6_198 b_6 NI_6 NS_198 0 -2.2630614492804953e-04
GC_6_199 b_6 NI_6 NS_199 0 1.2003658664690462e-05
GC_6_200 b_6 NI_6 NS_200 0 -3.7882926843930740e-05
GC_6_201 b_6 NI_6 NS_201 0 -3.9285558205074666e-05
GC_6_202 b_6 NI_6 NS_202 0 9.8860389111435305e-05
GC_6_203 b_6 NI_6 NS_203 0 -4.8820830478935500e-03
GC_6_204 b_6 NI_6 NS_204 0 -2.4003111658503357e-03
GC_6_205 b_6 NI_6 NS_205 0 2.1363378246382507e-05
GC_6_206 b_6 NI_6 NS_206 0 4.2602964474998445e-05
GC_6_207 b_6 NI_6 NS_207 0 1.6006805700589932e-04
GC_6_208 b_6 NI_6 NS_208 0 2.4980899425545576e-03
GC_6_209 b_6 NI_6 NS_209 0 2.4803343266547476e-06
GC_6_210 b_6 NI_6 NS_210 0 6.1212001849789140e-06
GC_6_211 b_6 NI_6 NS_211 0 5.2104534221729620e-04
GC_6_212 b_6 NI_6 NS_212 0 -1.0729617439953767e-03
GC_6_213 b_6 NI_6 NS_213 0 -1.1700289027278051e-05
GC_6_214 b_6 NI_6 NS_214 0 1.0227773365315870e-06
GC_6_215 b_6 NI_6 NS_215 0 4.1362991567403323e-07
GC_6_216 b_6 NI_6 NS_216 0 -2.5091993960977189e-07
GC_6_217 b_6 NI_6 NS_217 0 5.7644240416330535e-06
GC_6_218 b_6 NI_6 NS_218 0 -1.2770521820352859e-06
GC_6_219 b_6 NI_6 NS_219 0 3.8396977493448139e-05
GC_6_220 b_6 NI_6 NS_220 0 -3.1083180658393584e-04
GC_6_221 b_6 NI_6 NS_221 0 -2.1916729752687131e-01
GC_6_222 b_6 NI_6 NS_222 0 8.8019172797176599e-03
GC_6_223 b_6 NI_6 NS_223 0 7.0519108771433915e-03
GC_6_224 b_6 NI_6 NS_224 0 3.4545754907558072e-03
GC_6_225 b_6 NI_6 NS_225 0 7.1607832722372800e-03
GC_6_226 b_6 NI_6 NS_226 0 1.4578431379371069e-03
GC_6_227 b_6 NI_6 NS_227 0 1.1804171169549483e-03
GC_6_228 b_6 NI_6 NS_228 0 1.0386009368080627e-03
GC_6_229 b_6 NI_6 NS_229 0 1.2144100099967413e-03
GC_6_230 b_6 NI_6 NS_230 0 1.5788920679182547e-03
GC_6_231 b_6 NI_6 NS_231 0 4.5630578186509011e-03
GC_6_232 b_6 NI_6 NS_232 0 2.5390110653844529e-03
GC_6_233 b_6 NI_6 NS_233 0 -1.8111055768406251e-04
GC_6_234 b_6 NI_6 NS_234 0 3.0919646243102790e-04
GC_6_235 b_6 NI_6 NS_235 0 3.0893147003397798e-03
GC_6_236 b_6 NI_6 NS_236 0 7.9359172882505977e-03
GC_6_237 b_6 NI_6 NS_237 0 -4.0915269204910056e-05
GC_6_238 b_6 NI_6 NS_238 0 9.1472366830577532e-05
GC_6_239 b_6 NI_6 NS_239 0 1.6472460704121405e-05
GC_6_240 b_6 NI_6 NS_240 0 3.5421431018332222e-03
GC_6_241 b_6 NI_6 NS_241 0 1.0622569443642996e-03
GC_6_242 b_6 NI_6 NS_242 0 -6.8296720483817109e-04
GC_6_243 b_6 NI_6 NS_243 0 -1.0930764459769772e-04
GC_6_244 b_6 NI_6 NS_244 0 1.2954531047062299e-04
GC_6_245 b_6 NI_6 NS_245 0 -2.4238715312639600e-05
GC_6_246 b_6 NI_6 NS_246 0 -6.2752423449305810e-05
GC_6_247 b_6 NI_6 NS_247 0 -1.7997447536087154e-02
GC_6_248 b_6 NI_6 NS_248 0 1.9517406458543507e-03
GC_6_249 b_6 NI_6 NS_249 0 -1.8159402171433099e-05
GC_6_250 b_6 NI_6 NS_250 0 -7.2519743057649036e-05
GC_6_251 b_6 NI_6 NS_251 0 5.9759781521052571e-03
GC_6_252 b_6 NI_6 NS_252 0 3.9996779207515489e-03
GC_6_253 b_6 NI_6 NS_253 0 -7.1397312165802025e-06
GC_6_254 b_6 NI_6 NS_254 0 5.9657260318116979e-05
GC_6_255 b_6 NI_6 NS_255 0 1.6480597010149899e-03
GC_6_256 b_6 NI_6 NS_256 0 -2.9127911423027248e-03
GC_6_257 b_6 NI_6 NS_257 0 -6.6257646500060273e-05
GC_6_258 b_6 NI_6 NS_258 0 -2.5827409180625481e-05
GC_6_259 b_6 NI_6 NS_259 0 4.1008145540848061e-05
GC_6_260 b_6 NI_6 NS_260 0 -2.1742914390407809e-05
GC_6_261 b_6 NI_6 NS_261 0 6.5751443806159169e-05
GC_6_262 b_6 NI_6 NS_262 0 -2.1094771611080387e-05
GC_6_263 b_6 NI_6 NS_263 0 1.5161659985092951e-04
GC_6_264 b_6 NI_6 NS_264 0 -3.6616603539102471e-04
GC_6_265 b_6 NI_6 NS_265 0 5.9277590838375097e-02
GC_6_266 b_6 NI_6 NS_266 0 -2.7475158416143431e-05
GC_6_267 b_6 NI_6 NS_267 0 -6.3572684074957421e-03
GC_6_268 b_6 NI_6 NS_268 0 -2.7885077927858959e-03
GC_6_269 b_6 NI_6 NS_269 0 4.5424974237903227e-03
GC_6_270 b_6 NI_6 NS_270 0 2.5253523132831744e-03
GC_6_271 b_6 NI_6 NS_271 0 -9.3193455285250066e-05
GC_6_272 b_6 NI_6 NS_272 0 -9.3032552141541048e-06
GC_6_273 b_6 NI_6 NS_273 0 1.5993141753560831e-03
GC_6_274 b_6 NI_6 NS_274 0 1.4580953562381125e-03
GC_6_275 b_6 NI_6 NS_275 0 -2.8701040068948065e-04
GC_6_276 b_6 NI_6 NS_276 0 -6.3420842027111916e-04
GC_6_277 b_6 NI_6 NS_277 0 -1.1034372346330829e-05
GC_6_278 b_6 NI_6 NS_278 0 8.4701987232064558e-05
GC_6_279 b_6 NI_6 NS_279 0 -3.5420564190410961e-03
GC_6_280 b_6 NI_6 NS_280 0 1.1662922820359428e-03
GC_6_281 b_6 NI_6 NS_281 0 -8.5346020860497458e-05
GC_6_282 b_6 NI_6 NS_282 0 -5.6139264978598483e-05
GC_6_283 b_6 NI_6 NS_283 0 -1.6726118345553390e-04
GC_6_284 b_6 NI_6 NS_284 0 9.3040813197838685e-04
GC_6_285 b_6 NI_6 NS_285 0 3.2255186671266146e-04
GC_6_286 b_6 NI_6 NS_286 0 7.3322217666168618e-05
GC_6_287 b_6 NI_6 NS_287 0 -2.6835730194517945e-05
GC_6_288 b_6 NI_6 NS_288 0 -5.6552671435283881e-05
GC_6_289 b_6 NI_6 NS_289 0 -5.6342788325116567e-05
GC_6_290 b_6 NI_6 NS_290 0 9.0721114310191061e-05
GC_6_291 b_6 NI_6 NS_291 0 -3.0380232212207587e-03
GC_6_292 b_6 NI_6 NS_292 0 -3.5983006084404946e-03
GC_6_293 b_6 NI_6 NS_293 0 6.1954298309832121e-06
GC_6_294 b_6 NI_6 NS_294 0 3.5318192628800297e-05
GC_6_295 b_6 NI_6 NS_295 0 -5.3321561707320435e-04
GC_6_296 b_6 NI_6 NS_296 0 2.1117743705272181e-03
GC_6_297 b_6 NI_6 NS_297 0 -1.1845645591959225e-06
GC_6_298 b_6 NI_6 NS_298 0 9.0485614613806269e-06
GC_6_299 b_6 NI_6 NS_299 0 8.9383790627042673e-04
GC_6_300 b_6 NI_6 NS_300 0 -4.6641889262250111e-04
GC_6_301 b_6 NI_6 NS_301 0 -1.0904722203280007e-05
GC_6_302 b_6 NI_6 NS_302 0 -8.7298638010968662e-06
GC_6_303 b_6 NI_6 NS_303 0 2.4742799153883301e-06
GC_6_304 b_6 NI_6 NS_304 0 -1.9522346992084102e-06
GC_6_305 b_6 NI_6 NS_305 0 2.5702271722069605e-06
GC_6_306 b_6 NI_6 NS_306 0 -5.3615507651314731e-07
GC_6_307 b_6 NI_6 NS_307 0 9.3122811888528758e-05
GC_6_308 b_6 NI_6 NS_308 0 -1.4546258529250070e-04
GC_6_309 b_6 NI_6 NS_309 0 5.1376735144672177e-03
GC_6_310 b_6 NI_6 NS_310 0 -8.5693344052372193e-04
GC_6_311 b_6 NI_6 NS_311 0 4.0087013484621957e-03
GC_6_312 b_6 NI_6 NS_312 0 1.4684993441549845e-03
GC_6_313 b_6 NI_6 NS_313 0 -5.0365459478129903e-03
GC_6_314 b_6 NI_6 NS_314 0 -2.2501676135626672e-03
GC_6_315 b_6 NI_6 NS_315 0 8.8585647777355078e-05
GC_6_316 b_6 NI_6 NS_316 0 -4.7111936328809839e-05
GC_6_317 b_6 NI_6 NS_317 0 1.2781738230755234e-03
GC_6_318 b_6 NI_6 NS_318 0 7.9183488293869874e-05
GC_6_319 b_6 NI_6 NS_319 0 -6.1023622501290825e-05
GC_6_320 b_6 NI_6 NS_320 0 -6.7361576683503852e-04
GC_6_321 b_6 NI_6 NS_321 0 -1.5335861991374395e-05
GC_6_322 b_6 NI_6 NS_322 0 -3.8568167418822492e-05
GC_6_323 b_6 NI_6 NS_323 0 -9.7886818352386552e-04
GC_6_324 b_6 NI_6 NS_324 0 2.9189571122630498e-04
GC_6_325 b_6 NI_6 NS_325 0 3.3318511217508879e-05
GC_6_326 b_6 NI_6 NS_326 0 -2.7505581611665406e-05
GC_6_327 b_6 NI_6 NS_327 0 2.7376445228166060e-04
GC_6_328 b_6 NI_6 NS_328 0 -3.4607185237523966e-04
GC_6_329 b_6 NI_6 NS_329 0 2.5238630268626365e-04
GC_6_330 b_6 NI_6 NS_330 0 -1.6497682043695270e-04
GC_6_331 b_6 NI_6 NS_331 0 4.9667981131509945e-06
GC_6_332 b_6 NI_6 NS_332 0 -4.0538677631279679e-05
GC_6_333 b_6 NI_6 NS_333 0 -5.4313372911997898e-05
GC_6_334 b_6 NI_6 NS_334 0 -1.2916412901304612e-04
GC_6_335 b_6 NI_6 NS_335 0 1.4019882907441330e-03
GC_6_336 b_6 NI_6 NS_336 0 1.0625811330597654e-03
GC_6_337 b_6 NI_6 NS_337 0 -3.6553139039786101e-05
GC_6_338 b_6 NI_6 NS_338 0 -3.5152318726458940e-05
GC_6_339 b_6 NI_6 NS_339 0 1.1014908675308710e-03
GC_6_340 b_6 NI_6 NS_340 0 -1.0003693782859890e-03
GC_6_341 b_6 NI_6 NS_341 0 -4.7847417900245465e-06
GC_6_342 b_6 NI_6 NS_342 0 1.2027907655571776e-05
GC_6_343 b_6 NI_6 NS_343 0 1.7371194810321554e-04
GC_6_344 b_6 NI_6 NS_344 0 1.6458802072935713e-04
GC_6_345 b_6 NI_6 NS_345 0 -3.6207438456807786e-06
GC_6_346 b_6 NI_6 NS_346 0 -6.1269579384187236e-06
GC_6_347 b_6 NI_6 NS_347 0 2.6885551537093056e-05
GC_6_348 b_6 NI_6 NS_348 0 -1.7410672224629665e-07
GC_6_349 b_6 NI_6 NS_349 0 2.0594390266189919e-05
GC_6_350 b_6 NI_6 NS_350 0 -1.0279336532064359e-05
GC_6_351 b_6 NI_6 NS_351 0 -1.2397257946063613e-04
GC_6_352 b_6 NI_6 NS_352 0 1.7605344121446033e-04
GC_6_353 b_6 NI_6 NS_353 0 1.4261314013675171e-03
GC_6_354 b_6 NI_6 NS_354 0 -6.7033253027303681e-06
GC_6_355 b_6 NI_6 NS_355 0 -4.0969191184713394e-04
GC_6_356 b_6 NI_6 NS_356 0 4.6129996941727354e-04
GC_6_357 b_6 NI_6 NS_357 0 -3.7193509193635506e-04
GC_6_358 b_6 NI_6 NS_358 0 -7.2968885137358322e-04
GC_6_359 b_6 NI_6 NS_359 0 -3.0997807845427585e-05
GC_6_360 b_6 NI_6 NS_360 0 2.8271282081989351e-04
GC_6_361 b_6 NI_6 NS_361 0 3.7364201469673784e-04
GC_6_362 b_6 NI_6 NS_362 0 -4.5726431904445945e-04
GC_6_363 b_6 NI_6 NS_363 0 -1.3928557292169861e-04
GC_6_364 b_6 NI_6 NS_364 0 -4.0307293929535653e-04
GC_6_365 b_6 NI_6 NS_365 0 1.4612912619455299e-04
GC_6_366 b_6 NI_6 NS_366 0 9.8407616569496707e-05
GC_6_367 b_6 NI_6 NS_367 0 7.3128165221715276e-04
GC_6_368 b_6 NI_6 NS_368 0 7.1015589117140714e-04
GC_6_369 b_6 NI_6 NS_369 0 -1.7533806806157838e-04
GC_6_370 b_6 NI_6 NS_370 0 8.7703986869635880e-05
GC_6_371 b_6 NI_6 NS_371 0 -5.5700440717348562e-04
GC_6_372 b_6 NI_6 NS_372 0 -3.1092007879362973e-04
GC_6_373 b_6 NI_6 NS_373 0 -4.0364246139326242e-05
GC_6_374 b_6 NI_6 NS_374 0 -5.7661532819735310e-07
GC_6_375 b_6 NI_6 NS_375 0 -2.6374630329792578e-05
GC_6_376 b_6 NI_6 NS_376 0 -1.6347356146472261e-04
GC_6_377 b_6 NI_6 NS_377 0 -7.2801185811186911e-07
GC_6_378 b_6 NI_6 NS_378 0 1.3419482376214964e-04
GC_6_379 b_6 NI_6 NS_379 0 2.0646318574329314e-03
GC_6_380 b_6 NI_6 NS_380 0 1.0799052118371075e-03
GC_6_381 b_6 NI_6 NS_381 0 -3.5532406587675479e-05
GC_6_382 b_6 NI_6 NS_382 0 -1.4195518965399246e-05
GC_6_383 b_6 NI_6 NS_383 0 -5.4147212509371033e-04
GC_6_384 b_6 NI_6 NS_384 0 -8.3310959628123777e-04
GC_6_385 b_6 NI_6 NS_385 0 -6.7268862332531227e-07
GC_6_386 b_6 NI_6 NS_386 0 2.0299725601371080e-06
GC_6_387 b_6 NI_6 NS_387 0 -2.8595469569032251e-04
GC_6_388 b_6 NI_6 NS_388 0 -1.3148419610101373e-04
GC_6_389 b_6 NI_6 NS_389 0 -1.3820329669696083e-05
GC_6_390 b_6 NI_6 NS_390 0 -2.1115572382647261e-05
GC_6_391 b_6 NI_6 NS_391 0 -4.4101161008105011e-07
GC_6_392 b_6 NI_6 NS_392 0 3.2097387335878071e-06
GC_6_393 b_6 NI_6 NS_393 0 -2.0199105055665310e-06
GC_6_394 b_6 NI_6 NS_394 0 -3.4269797520103543e-06
GC_6_395 b_6 NI_6 NS_395 0 -3.7162045615700179e-04
GC_6_396 b_6 NI_6 NS_396 0 -2.5400512145005682e-05
GC_6_397 b_6 NI_6 NS_397 0 -1.6129938179184479e-03
GC_6_398 b_6 NI_6 NS_398 0 -1.1216280374692098e-06
GC_6_399 b_6 NI_6 NS_399 0 8.6298601442825359e-05
GC_6_400 b_6 NI_6 NS_400 0 -6.0149869369217305e-04
GC_6_401 b_6 NI_6 NS_401 0 4.6217613371854678e-04
GC_6_402 b_6 NI_6 NS_402 0 1.7239974561086789e-04
GC_6_403 b_6 NI_6 NS_403 0 -6.4557502754674604e-04
GC_6_404 b_6 NI_6 NS_404 0 1.3454361190154656e-05
GC_6_405 b_6 NI_6 NS_405 0 1.9087915044525069e-04
GC_6_406 b_6 NI_6 NS_406 0 -2.3417011386435606e-04
GC_6_407 b_6 NI_6 NS_407 0 1.7009027506395113e-04
GC_6_408 b_6 NI_6 NS_408 0 -3.9750363413545579e-04
GC_6_409 b_6 NI_6 NS_409 0 2.5851660907411725e-05
GC_6_410 b_6 NI_6 NS_410 0 4.2872190148582236e-05
GC_6_411 b_6 NI_6 NS_411 0 1.0420958346208508e-03
GC_6_412 b_6 NI_6 NS_412 0 -8.8542226357826086e-04
GC_6_413 b_6 NI_6 NS_413 0 2.3399744822301506e-05
GC_6_414 b_6 NI_6 NS_414 0 -6.5819520446056234e-05
GC_6_415 b_6 NI_6 NS_415 0 1.1041828901481555e-03
GC_6_416 b_6 NI_6 NS_416 0 -4.9338505119980085e-04
GC_6_417 b_6 NI_6 NS_417 0 -3.7362382505429795e-04
GC_6_418 b_6 NI_6 NS_418 0 -5.0906320589109077e-04
GC_6_419 b_6 NI_6 NS_419 0 1.4981476835176925e-05
GC_6_420 b_6 NI_6 NS_420 0 -3.7130324349898189e-05
GC_6_421 b_6 NI_6 NS_421 0 -7.2096742130301340e-05
GC_6_422 b_6 NI_6 NS_422 0 -2.3775088355210662e-04
GC_6_423 b_6 NI_6 NS_423 0 -5.3620413423775852e-03
GC_6_424 b_6 NI_6 NS_424 0 7.4549018751145970e-03
GC_6_425 b_6 NI_6 NS_425 0 2.3383017597085474e-05
GC_6_426 b_6 NI_6 NS_426 0 2.3332420278995572e-05
GC_6_427 b_6 NI_6 NS_427 0 5.0524938007056180e-03
GC_6_428 b_6 NI_6 NS_428 0 -2.4214348915860729e-03
GC_6_429 b_6 NI_6 NS_429 0 3.4032351581274262e-05
GC_6_430 b_6 NI_6 NS_430 0 4.7094825644498306e-06
GC_6_431 b_6 NI_6 NS_431 0 -6.0307805619445865e-04
GC_6_432 b_6 NI_6 NS_432 0 -5.4086150589779838e-04
GC_6_433 b_6 NI_6 NS_433 0 -7.7108763443060039e-05
GC_6_434 b_6 NI_6 NS_434 0 2.0771886408506818e-05
GC_6_435 b_6 NI_6 NS_435 0 4.4023055567359980e-05
GC_6_436 b_6 NI_6 NS_436 0 -1.2450719914009934e-05
GC_6_437 b_6 NI_6 NS_437 0 -2.6682140053410156e-05
GC_6_438 b_6 NI_6 NS_438 0 2.4203943022263110e-05
GC_6_439 b_6 NI_6 NS_439 0 5.9698486964600837e-04
GC_6_440 b_6 NI_6 NS_440 0 2.0364815574433964e-04
GC_6_441 b_6 NI_6 NS_441 0 -4.2622168612487391e-03
GC_6_442 b_6 NI_6 NS_442 0 -1.8702595842776447e-05
GC_6_443 b_6 NI_6 NS_443 0 -1.2972508191197523e-03
GC_6_444 b_6 NI_6 NS_444 0 2.2387696940233379e-04
GC_6_445 b_6 NI_6 NS_445 0 6.0737820138401374e-04
GC_6_446 b_6 NI_6 NS_446 0 -1.2187294176997398e-03
GC_6_447 b_6 NI_6 NS_447 0 -2.8443767277755778e-05
GC_6_448 b_6 NI_6 NS_448 0 1.5685281224036603e-04
GC_6_449 b_6 NI_6 NS_449 0 6.8039264115879515e-04
GC_6_450 b_6 NI_6 NS_450 0 -1.4008572729733829e-04
GC_6_451 b_6 NI_6 NS_451 0 -2.4018327499072918e-04
GC_6_452 b_6 NI_6 NS_452 0 -1.0944691643645350e-03
GC_6_453 b_6 NI_6 NS_453 0 1.2252475684124435e-04
GC_6_454 b_6 NI_6 NS_454 0 9.3166855023312076e-05
GC_6_455 b_6 NI_6 NS_455 0 9.6116463624006142e-04
GC_6_456 b_6 NI_6 NS_456 0 1.2705264054194243e-03
GC_6_457 b_6 NI_6 NS_457 0 -1.2482948934993546e-04
GC_6_458 b_6 NI_6 NS_458 0 4.8405549862692550e-05
GC_6_459 b_6 NI_6 NS_459 0 -2.5231909942981088e-04
GC_6_460 b_6 NI_6 NS_460 0 -5.5638004726569957e-05
GC_6_461 b_6 NI_6 NS_461 0 -1.2047343992583138e-05
GC_6_462 b_6 NI_6 NS_462 0 4.2813796517522313e-05
GC_6_463 b_6 NI_6 NS_463 0 -1.9209038448738522e-05
GC_6_464 b_6 NI_6 NS_464 0 -1.0859384247396916e-04
GC_6_465 b_6 NI_6 NS_465 0 -2.1956983040740757e-05
GC_6_466 b_6 NI_6 NS_466 0 1.0095892929448008e-04
GC_6_467 b_6 NI_6 NS_467 0 1.0425907919263090e-03
GC_6_468 b_6 NI_6 NS_468 0 7.4111169177215337e-04
GC_6_469 b_6 NI_6 NS_469 0 -1.8694169599223877e-05
GC_6_470 b_6 NI_6 NS_470 0 -6.7359230752824077e-06
GC_6_471 b_6 NI_6 NS_471 0 -3.0562213693831255e-04
GC_6_472 b_6 NI_6 NS_472 0 -5.2287179528384426e-04
GC_6_473 b_6 NI_6 NS_473 0 -1.7539255782784296e-06
GC_6_474 b_6 NI_6 NS_474 0 -1.4693677281763799e-06
GC_6_475 b_6 NI_6 NS_475 0 -3.9879059939977138e-05
GC_6_476 b_6 NI_6 NS_476 0 -1.4014732454265826e-04
GC_6_477 b_6 NI_6 NS_477 0 -8.1771730056874770e-06
GC_6_478 b_6 NI_6 NS_478 0 -1.1988129325785360e-05
GC_6_479 b_6 NI_6 NS_479 0 1.6414955000622858e-07
GC_6_480 b_6 NI_6 NS_480 0 -5.1072690272563863e-07
GC_6_481 b_6 NI_6 NS_481 0 -4.9584215512914680e-07
GC_6_482 b_6 NI_6 NS_482 0 -9.0816035651892502e-07
GC_6_483 b_6 NI_6 NS_483 0 -1.9937568316974561e-04
GC_6_484 b_6 NI_6 NS_484 0 -7.4310487947240215e-05
GC_6_485 b_6 NI_6 NS_485 0 1.2540202005088580e-03
GC_6_486 b_6 NI_6 NS_486 0 -3.2026248879287399e-05
GC_6_487 b_6 NI_6 NS_487 0 8.1546736481515904e-04
GC_6_488 b_6 NI_6 NS_488 0 -5.7894156629346484e-04
GC_6_489 b_6 NI_6 NS_489 0 -2.7239275217817238e-04
GC_6_490 b_6 NI_6 NS_490 0 7.7376690267265012e-04
GC_6_491 b_6 NI_6 NS_491 0 -6.0919698983267221e-04
GC_6_492 b_6 NI_6 NS_492 0 1.2902447373881986e-04
GC_6_493 b_6 NI_6 NS_493 0 1.7009403279741848e-04
GC_6_494 b_6 NI_6 NS_494 0 -1.4359737392369837e-04
GC_6_495 b_6 NI_6 NS_495 0 -1.4322674764686403e-04
GC_6_496 b_6 NI_6 NS_496 0 -1.9327103583475759e-04
GC_6_497 b_6 NI_6 NS_497 0 -7.5152624414637542e-06
GC_6_498 b_6 NI_6 NS_498 0 1.8486941659858916e-05
GC_6_499 b_6 NI_6 NS_499 0 5.1042155090203118e-04
GC_6_500 b_6 NI_6 NS_500 0 -7.9716883458515634e-05
GC_6_501 b_6 NI_6 NS_501 0 1.4250158379019971e-05
GC_6_502 b_6 NI_6 NS_502 0 -4.2994163224837802e-05
GC_6_503 b_6 NI_6 NS_503 0 4.8058563417986802e-04
GC_6_504 b_6 NI_6 NS_504 0 -3.1871655519444389e-04
GC_6_505 b_6 NI_6 NS_505 0 -8.9583996024427120e-05
GC_6_506 b_6 NI_6 NS_506 0 -2.2334874757592725e-04
GC_6_507 b_6 NI_6 NS_507 0 1.6604558158687174e-06
GC_6_508 b_6 NI_6 NS_508 0 -2.8920547493064642e-05
GC_6_509 b_6 NI_6 NS_509 0 -4.7202523302081558e-05
GC_6_510 b_6 NI_6 NS_510 0 -1.4992322040080472e-04
GC_6_511 b_6 NI_6 NS_511 0 -3.0985337913214130e-03
GC_6_512 b_6 NI_6 NS_512 0 3.2699874763168057e-03
GC_6_513 b_6 NI_6 NS_513 0 6.7883969185989973e-06
GC_6_514 b_6 NI_6 NS_514 0 5.2403618437626842e-06
GC_6_515 b_6 NI_6 NS_515 0 2.8197714176916478e-03
GC_6_516 b_6 NI_6 NS_516 0 -1.1144627610881123e-03
GC_6_517 b_6 NI_6 NS_517 0 1.1482132041537219e-05
GC_6_518 b_6 NI_6 NS_518 0 5.4142568331144456e-06
GC_6_519 b_6 NI_6 NS_519 0 -4.5566564097796303e-05
GC_6_520 b_6 NI_6 NS_520 0 -2.6279788251409115e-04
GC_6_521 b_6 NI_6 NS_521 0 -3.3524201685262749e-05
GC_6_522 b_6 NI_6 NS_522 0 3.0850583765467052e-06
GC_6_523 b_6 NI_6 NS_523 0 2.8178598698449791e-05
GC_6_524 b_6 NI_6 NS_524 0 -3.9493520627439564e-06
GC_6_525 b_6 NI_6 NS_525 0 -1.1068944764827016e-05
GC_6_526 b_6 NI_6 NS_526 0 8.6936063233646166e-06
GC_6_527 b_6 NI_6 NS_527 0 2.9997972068650610e-04
GC_6_528 b_6 NI_6 NS_528 0 1.2609752803919799e-04
GD_6_1 b_6 NI_6 NA_1 0 -3.8611709331058917e-02
GD_6_2 b_6 NI_6 NA_2 0 -1.9402984504318918e-02
GD_6_3 b_6 NI_6 NA_3 0 -8.5081740125850264e-02
GD_6_4 b_6 NI_6 NA_4 0 -2.6996141370273997e-02
GD_6_5 b_6 NI_6 NA_5 0 -4.5682579115256035e-02
GD_6_6 b_6 NI_6 NA_6 0 2.4591321146872933e-01
GD_6_7 b_6 NI_6 NA_7 0 -6.3855611028977077e-02
GD_6_8 b_6 NI_6 NA_8 0 -1.5472297387371610e-02
GD_6_9 b_6 NI_6 NA_9 0 -2.9442930721125258e-03
GD_6_10 b_6 NI_6 NA_10 0 -1.1283511704917291e-03
GD_6_11 b_6 NI_6 NA_11 0 3.3959406975204456e-03
GD_6_12 b_6 NI_6 NA_12 0 -3.3694698103710597e-03
*
* Port 7
VI_7 a_7 NI_7 0
RI_7 NI_7 b_7 5.0000000000000000e+01
GC_7_1 b_7 NI_7 NS_1 0 5.9439141061517322e-03
GC_7_2 b_7 NI_7 NS_2 0 2.1847207596614084e-04
GC_7_3 b_7 NI_7 NS_3 0 3.9291690159699456e-03
GC_7_4 b_7 NI_7 NS_4 0 -1.0764521587849746e-03
GC_7_5 b_7 NI_7 NS_5 0 -1.1873467966992629e-03
GC_7_6 b_7 NI_7 NS_6 0 3.8898348436914956e-03
GC_7_7 b_7 NI_7 NS_7 0 -5.8511401949246080e-05
GC_7_8 b_7 NI_7 NS_8 0 9.3949177831428461e-05
GC_7_9 b_7 NI_7 NS_9 0 1.0192425276705573e-03
GC_7_10 b_7 NI_7 NS_10 0 4.4797091585656104e-03
GC_7_11 b_7 NI_7 NS_11 0 -1.1924405994122813e-02
GC_7_12 b_7 NI_7 NS_12 0 -9.9346967053355931e-04
GC_7_13 b_7 NI_7 NS_13 0 6.9198140465335470e-04
GC_7_14 b_7 NI_7 NS_14 0 8.6915782290582076e-05
GC_7_15 b_7 NI_7 NS_15 0 2.5020735856144056e-03
GC_7_16 b_7 NI_7 NS_16 0 -2.0610917873215909e-03
GC_7_17 b_7 NI_7 NS_17 0 -1.3573399581325375e-05
GC_7_18 b_7 NI_7 NS_18 0 9.8333464695988309e-05
GC_7_19 b_7 NI_7 NS_19 0 -1.0167624825276774e-03
GC_7_20 b_7 NI_7 NS_20 0 -3.1477886592925553e-03
GC_7_21 b_7 NI_7 NS_21 0 -1.5179162231568179e-04
GC_7_22 b_7 NI_7 NS_22 0 1.1321621591393962e-03
GC_7_23 b_7 NI_7 NS_23 0 1.3200640895982799e-04
GC_7_24 b_7 NI_7 NS_24 0 -8.2116949279960354e-05
GC_7_25 b_7 NI_7 NS_25 0 -1.0844656258320520e-05
GC_7_26 b_7 NI_7 NS_26 0 -6.6003135295787633e-05
GC_7_27 b_7 NI_7 NS_27 0 4.3543271238076628e-03
GC_7_28 b_7 NI_7 NS_28 0 -1.1807794079106522e-03
GC_7_29 b_7 NI_7 NS_29 0 -1.2831524223698284e-05
GC_7_30 b_7 NI_7 NS_30 0 1.3708259124627471e-06
GC_7_31 b_7 NI_7 NS_31 0 -9.4374339341009208e-04
GC_7_32 b_7 NI_7 NS_32 0 -2.1709858009766815e-03
GC_7_33 b_7 NI_7 NS_33 0 -8.8601880379515323e-06
GC_7_34 b_7 NI_7 NS_34 0 -3.6726130169973089e-06
GC_7_35 b_7 NI_7 NS_35 0 1.2863760193210600e-03
GC_7_36 b_7 NI_7 NS_36 0 1.6432059901724844e-03
GC_7_37 b_7 NI_7 NS_37 0 1.4652244937660880e-05
GC_7_38 b_7 NI_7 NS_38 0 -6.3341415228459764e-06
GC_7_39 b_7 NI_7 NS_39 0 2.6462469595512812e-06
GC_7_40 b_7 NI_7 NS_40 0 5.0865518996177130e-06
GC_7_41 b_7 NI_7 NS_41 0 -4.2435176395824786e-06
GC_7_42 b_7 NI_7 NS_42 0 1.4705365648533031e-06
GC_7_43 b_7 NI_7 NS_43 0 6.4674498431806243e-05
GC_7_44 b_7 NI_7 NS_44 0 2.0173185713240373e-04
GC_7_45 b_7 NI_7 NS_45 0 2.3421754060697925e-02
GC_7_46 b_7 NI_7 NS_46 0 -2.5744160039516806e-04
GC_7_47 b_7 NI_7 NS_47 0 -3.1492332532555701e-03
GC_7_48 b_7 NI_7 NS_48 0 2.0868689764298809e-03
GC_7_49 b_7 NI_7 NS_49 0 -4.7099148723427878e-05
GC_7_50 b_7 NI_7 NS_50 0 -3.0612636009240135e-03
GC_7_51 b_7 NI_7 NS_51 0 1.8864770714304853e-04
GC_7_52 b_7 NI_7 NS_52 0 6.7951159702872319e-05
GC_7_53 b_7 NI_7 NS_53 0 1.5603791899529099e-03
GC_7_54 b_7 NI_7 NS_54 0 8.3668656893529656e-04
GC_7_55 b_7 NI_7 NS_55 0 -5.1453057171495144e-03
GC_7_56 b_7 NI_7 NS_56 0 8.9095471934515160e-04
GC_7_57 b_7 NI_7 NS_57 0 5.5190051680566597e-05
GC_7_58 b_7 NI_7 NS_58 0 -1.6637660310999658e-05
GC_7_59 b_7 NI_7 NS_59 0 4.4096880992025117e-04
GC_7_60 b_7 NI_7 NS_60 0 -2.0968202351476567e-03
GC_7_61 b_7 NI_7 NS_61 0 -1.8612084072054220e-05
GC_7_62 b_7 NI_7 NS_62 0 -4.8223265364785141e-05
GC_7_63 b_7 NI_7 NS_63 0 4.1823346922071752e-04
GC_7_64 b_7 NI_7 NS_64 0 9.3471779186359996e-06
GC_7_65 b_7 NI_7 NS_65 0 2.4959788655034171e-05
GC_7_66 b_7 NI_7 NS_66 0 4.9544013231237725e-05
GC_7_67 b_7 NI_7 NS_67 0 1.4606028207415028e-05
GC_7_68 b_7 NI_7 NS_68 0 -5.2036211392318819e-05
GC_7_69 b_7 NI_7 NS_69 0 -4.0054349091419820e-05
GC_7_70 b_7 NI_7 NS_70 0 3.5301421246226519e-05
GC_7_71 b_7 NI_7 NS_71 0 1.2943919321089614e-03
GC_7_72 b_7 NI_7 NS_72 0 -2.6457135426925455e-03
GC_7_73 b_7 NI_7 NS_73 0 -3.0503865609536689e-06
GC_7_74 b_7 NI_7 NS_74 0 2.3441240390873434e-05
GC_7_75 b_7 NI_7 NS_75 0 -9.6046850693487366e-04
GC_7_76 b_7 NI_7 NS_76 0 4.3628075591360297e-04
GC_7_77 b_7 NI_7 NS_77 0 -3.6554029447310160e-06
GC_7_78 b_7 NI_7 NS_78 0 2.1266828979296259e-06
GC_7_79 b_7 NI_7 NS_79 0 3.3213154638935119e-04
GC_7_80 b_7 NI_7 NS_80 0 2.8075420759839223e-04
GC_7_81 b_7 NI_7 NS_81 0 1.7568629403513460e-06
GC_7_82 b_7 NI_7 NS_82 0 -4.7935201506672608e-06
GC_7_83 b_7 NI_7 NS_83 0 1.4472919115040033e-06
GC_7_84 b_7 NI_7 NS_84 0 9.2826859798322778e-07
GC_7_85 b_7 NI_7 NS_85 0 -1.2266856706023291e-06
GC_7_86 b_7 NI_7 NS_86 0 -1.4451505818684560e-06
GC_7_87 b_7 NI_7 NS_87 0 -2.2064618631452007e-06
GC_7_88 b_7 NI_7 NS_88 0 -1.2790581488882601e-06
GC_7_89 b_7 NI_7 NS_89 0 3.6231626107672693e-02
GC_7_90 b_7 NI_7 NS_90 0 1.5138667923208845e-04
GC_7_91 b_7 NI_7 NS_91 0 5.9839007046610000e-03
GC_7_92 b_7 NI_7 NS_92 0 1.2391252333414017e-03
GC_7_93 b_7 NI_7 NS_93 0 -4.2692852410159887e-03
GC_7_94 b_7 NI_7 NS_94 0 2.4099803366335448e-03
GC_7_95 b_7 NI_7 NS_95 0 -1.8580069002251427e-04
GC_7_96 b_7 NI_7 NS_96 0 -8.7100542170489301e-04
GC_7_97 b_7 NI_7 NS_97 0 1.3876197649330881e-03
GC_7_98 b_7 NI_7 NS_98 0 6.0150671935242364e-03
GC_7_99 b_7 NI_7 NS_99 0 -1.0172212263051676e-02
GC_7_100 b_7 NI_7 NS_100 0 -1.3505052452387617e-03
GC_7_101 b_7 NI_7 NS_101 0 9.3708588828123453e-04
GC_7_102 b_7 NI_7 NS_102 0 1.5662942157510323e-04
GC_7_103 b_7 NI_7 NS_103 0 -1.4485518766621257e-03
GC_7_104 b_7 NI_7 NS_104 0 3.5854117452970794e-04
GC_7_105 b_7 NI_7 NS_105 0 -4.7419853035915228e-05
GC_7_106 b_7 NI_7 NS_106 0 1.3954276661689845e-04
GC_7_107 b_7 NI_7 NS_107 0 -1.9605622258680503e-03
GC_7_108 b_7 NI_7 NS_108 0 -3.0129734996269257e-03
GC_7_109 b_7 NI_7 NS_109 0 -9.1329852567328319e-05
GC_7_110 b_7 NI_7 NS_110 0 5.5448636407292391e-04
GC_7_111 b_7 NI_7 NS_111 0 1.5028063213180337e-04
GC_7_112 b_7 NI_7 NS_112 0 -9.0394723584491941e-05
GC_7_113 b_7 NI_7 NS_113 0 -6.3512238769862386e-06
GC_7_114 b_7 NI_7 NS_114 0 -5.3563262495730585e-05
GC_7_115 b_7 NI_7 NS_115 0 1.5528939188632351e-03
GC_7_116 b_7 NI_7 NS_116 0 -1.7847901804522387e-03
GC_7_117 b_7 NI_7 NS_117 0 -5.4102261688958868e-06
GC_7_118 b_7 NI_7 NS_118 0 1.0647019392077615e-07
GC_7_119 b_7 NI_7 NS_119 0 9.8253138992989640e-05
GC_7_120 b_7 NI_7 NS_120 0 -1.9582777913004818e-03
GC_7_121 b_7 NI_7 NS_121 0 3.9378267394752841e-07
GC_7_122 b_7 NI_7 NS_122 0 -4.4113111950412442e-06
GC_7_123 b_7 NI_7 NS_123 0 1.5333070809383119e-03
GC_7_124 b_7 NI_7 NS_124 0 3.4475709693679042e-04
GC_7_125 b_7 NI_7 NS_125 0 2.5739790537335242e-06
GC_7_126 b_7 NI_7 NS_126 0 2.1758756797359121e-06
GC_7_127 b_7 NI_7 NS_127 0 1.8069203400319066e-06
GC_7_128 b_7 NI_7 NS_128 0 2.7659732112035587e-06
GC_7_129 b_7 NI_7 NS_129 0 1.1298204587340375e-06
GC_7_130 b_7 NI_7 NS_130 0 9.3955426964680420e-07
GC_7_131 b_7 NI_7 NS_131 0 1.4884658142473619e-04
GC_7_132 b_7 NI_7 NS_132 0 1.9234487314637752e-05
GC_7_133 b_7 NI_7 NS_133 0 3.3788776492737121e-02
GC_7_134 b_7 NI_7 NS_134 0 -2.0388118518869242e-04
GC_7_135 b_7 NI_7 NS_135 0 -5.5026168440733408e-03
GC_7_136 b_7 NI_7 NS_136 0 5.0652734130573161e-04
GC_7_137 b_7 NI_7 NS_137 0 2.6909309198139696e-03
GC_7_138 b_7 NI_7 NS_138 0 -2.3867910101861437e-03
GC_7_139 b_7 NI_7 NS_139 0 -1.5748424516710995e-04
GC_7_140 b_7 NI_7 NS_140 0 2.3007682487844228e-04
GC_7_141 b_7 NI_7 NS_141 0 2.1605684616547312e-03
GC_7_142 b_7 NI_7 NS_142 0 1.4832932340275234e-03
GC_7_143 b_7 NI_7 NS_143 0 -3.5966326718437263e-03
GC_7_144 b_7 NI_7 NS_144 0 -4.5070157842589021e-04
GC_7_145 b_7 NI_7 NS_145 0 2.6407191388053029e-05
GC_7_146 b_7 NI_7 NS_146 0 4.2459118057071248e-05
GC_7_147 b_7 NI_7 NS_147 0 -9.5021268680580871e-04
GC_7_148 b_7 NI_7 NS_148 0 7.3529008469964320e-05
GC_7_149 b_7 NI_7 NS_149 0 -3.1930639164977246e-05
GC_7_150 b_7 NI_7 NS_150 0 -4.3847887817200422e-05
GC_7_151 b_7 NI_7 NS_151 0 2.5669071472464428e-04
GC_7_152 b_7 NI_7 NS_152 0 1.8080885891674225e-04
GC_7_153 b_7 NI_7 NS_153 0 1.2241948725387865e-04
GC_7_154 b_7 NI_7 NS_154 0 6.7511183462780149e-05
GC_7_155 b_7 NI_7 NS_155 0 6.9805692748253691e-06
GC_7_156 b_7 NI_7 NS_156 0 -5.0247317014538246e-05
GC_7_157 b_7 NI_7 NS_157 0 -3.9996725247957170e-05
GC_7_158 b_7 NI_7 NS_158 0 4.8484425352641372e-05
GC_7_159 b_7 NI_7 NS_159 0 5.4138962585919268e-04
GC_7_160 b_7 NI_7 NS_160 0 -2.5242648812577773e-03
GC_7_161 b_7 NI_7 NS_161 0 -1.6793893815166864e-06
GC_7_162 b_7 NI_7 NS_162 0 2.4071648611053088e-05
GC_7_163 b_7 NI_7 NS_163 0 -8.6339595605048323e-04
GC_7_164 b_7 NI_7 NS_164 0 6.5339803193640190e-04
GC_7_165 b_7 NI_7 NS_165 0 -2.6633411307241567e-06
GC_7_166 b_7 NI_7 NS_166 0 3.2874311568619628e-06
GC_7_167 b_7 NI_7 NS_167 0 4.5084976431734018e-04
GC_7_168 b_7 NI_7 NS_168 0 1.3105409654359907e-04
GC_7_169 b_7 NI_7 NS_169 0 -3.7032606737620257e-07
GC_7_170 b_7 NI_7 NS_170 0 -5.3490604046251028e-06
GC_7_171 b_7 NI_7 NS_171 0 1.4168052283244437e-06
GC_7_172 b_7 NI_7 NS_172 0 5.8378197348837311e-07
GC_7_173 b_7 NI_7 NS_173 0 -4.2206705466282581e-07
GC_7_174 b_7 NI_7 NS_174 0 -9.7422833278502886e-07
GC_7_175 b_7 NI_7 NS_175 0 1.5117049950528037e-05
GC_7_176 b_7 NI_7 NS_176 0 -1.3826360948128436e-05
GC_7_177 b_7 NI_7 NS_177 0 -2.3102765054898600e-03
GC_7_178 b_7 NI_7 NS_178 0 -5.6302554827866204e-05
GC_7_179 b_7 NI_7 NS_179 0 4.8917621372270865e-03
GC_7_180 b_7 NI_7 NS_180 0 4.5898850358533820e-03
GC_7_181 b_7 NI_7 NS_181 0 -5.2257083881258977e-03
GC_7_182 b_7 NI_7 NS_182 0 -4.9630806880778082e-03
GC_7_183 b_7 NI_7 NS_183 0 -3.1758750525029789e-05
GC_7_184 b_7 NI_7 NS_184 0 4.0982304428894845e-04
GC_7_185 b_7 NI_7 NS_185 0 1.6246603458643760e-03
GC_7_186 b_7 NI_7 NS_186 0 5.2287885909636407e-03
GC_7_187 b_7 NI_7 NS_187 0 -3.1142704505303692e-03
GC_7_188 b_7 NI_7 NS_188 0 -1.0630667123437936e-03
GC_7_189 b_7 NI_7 NS_189 0 9.4725716781049365e-04
GC_7_190 b_7 NI_7 NS_190 0 1.7721185240702870e-04
GC_7_191 b_7 NI_7 NS_191 0 -4.1398836435463876e-03
GC_7_192 b_7 NI_7 NS_192 0 -2.5394954768980520e-03
GC_7_193 b_7 NI_7 NS_193 0 -1.9713332433680704e-05
GC_7_194 b_7 NI_7 NS_194 0 1.5941970475476767e-04
GC_7_195 b_7 NI_7 NS_195 0 -2.1284931935396088e-03
GC_7_196 b_7 NI_7 NS_196 0 -2.4351069177824371e-03
GC_7_197 b_7 NI_7 NS_197 0 -1.0461556118051425e-04
GC_7_198 b_7 NI_7 NS_198 0 4.9700616757469699e-04
GC_7_199 b_7 NI_7 NS_199 0 1.8903158519031538e-04
GC_7_200 b_7 NI_7 NS_200 0 -7.4294459643291450e-05
GC_7_201 b_7 NI_7 NS_201 0 1.0810013983657165e-05
GC_7_202 b_7 NI_7 NS_202 0 -7.5591724719156758e-05
GC_7_203 b_7 NI_7 NS_203 0 6.3545869413145079e-03
GC_7_204 b_7 NI_7 NS_204 0 1.7233810257730841e-03
GC_7_205 b_7 NI_7 NS_205 0 -1.2260279588459924e-05
GC_7_206 b_7 NI_7 NS_206 0 -9.0304455076240320e-06
GC_7_207 b_7 NI_7 NS_207 0 5.8006672565822704e-04
GC_7_208 b_7 NI_7 NS_208 0 -3.3175830067033035e-03
GC_7_209 b_7 NI_7 NS_209 0 -4.5370061416517539e-07
GC_7_210 b_7 NI_7 NS_210 0 -8.1119313040742241e-06
GC_7_211 b_7 NI_7 NS_211 0 1.1037567383314750e-03
GC_7_212 b_7 NI_7 NS_212 0 8.2773916732083804e-04
GC_7_213 b_7 NI_7 NS_213 0 1.0500685487296867e-05
GC_7_214 b_7 NI_7 NS_214 0 6.2650302579076899e-06
GC_7_215 b_7 NI_7 NS_215 0 6.7421289897777093e-07
GC_7_216 b_7 NI_7 NS_216 0 4.8437550751310926e-06
GC_7_217 b_7 NI_7 NS_217 0 -1.2318448457263625e-06
GC_7_218 b_7 NI_7 NS_218 0 -1.3055735657052743e-06
GC_7_219 b_7 NI_7 NS_219 0 3.2270008786896775e-05
GC_7_220 b_7 NI_7 NS_220 0 6.8860284947307586e-05
GC_7_221 b_7 NI_7 NS_221 0 5.9277590836364580e-02
GC_7_222 b_7 NI_7 NS_222 0 -2.7475158407972991e-05
GC_7_223 b_7 NI_7 NS_223 0 -6.3572684075049032e-03
GC_7_224 b_7 NI_7 NS_224 0 -2.7885077928212036e-03
GC_7_225 b_7 NI_7 NS_225 0 4.5424974238212320e-03
GC_7_226 b_7 NI_7 NS_226 0 2.5253523132497853e-03
GC_7_227 b_7 NI_7 NS_227 0 -9.3193455074473222e-05
GC_7_228 b_7 NI_7 NS_228 0 -9.3032547894338991e-06
GC_7_229 b_7 NI_7 NS_229 0 1.5993141753580054e-03
GC_7_230 b_7 NI_7 NS_230 0 1.4580953562150609e-03
GC_7_231 b_7 NI_7 NS_231 0 -2.8701040077193309e-04
GC_7_232 b_7 NI_7 NS_232 0 -6.3420842031165271e-04
GC_7_233 b_7 NI_7 NS_233 0 -1.1034372344341867e-05
GC_7_234 b_7 NI_7 NS_234 0 8.4701987225579783e-05
GC_7_235 b_7 NI_7 NS_235 0 -3.5420564190981048e-03
GC_7_236 b_7 NI_7 NS_236 0 1.1662922818368056e-03
GC_7_237 b_7 NI_7 NS_237 0 -8.5346020859039572e-05
GC_7_238 b_7 NI_7 NS_238 0 -5.6139264981744174e-05
GC_7_239 b_7 NI_7 NS_239 0 -1.6726118347777994e-04
GC_7_240 b_7 NI_7 NS_240 0 9.3040813187772280e-04
GC_7_241 b_7 NI_7 NS_241 0 3.2255186671226882e-04
GC_7_242 b_7 NI_7 NS_242 0 7.3322217775050340e-05
GC_7_243 b_7 NI_7 NS_243 0 -2.6835730194153883e-05
GC_7_244 b_7 NI_7 NS_244 0 -5.6552671440687646e-05
GC_7_245 b_7 NI_7 NS_245 0 -5.6342788328570036e-05
GC_7_246 b_7 NI_7 NS_246 0 9.0721114308469971e-05
GC_7_247 b_7 NI_7 NS_247 0 -3.0380232203784355e-03
GC_7_248 b_7 NI_7 NS_248 0 -3.5983006088756569e-03
GC_7_249 b_7 NI_7 NS_249 0 6.1954298298330490e-06
GC_7_250 b_7 NI_7 NS_250 0 3.5318192629975518e-05
GC_7_251 b_7 NI_7 NS_251 0 -5.3321561732109514e-04
GC_7_252 b_7 NI_7 NS_252 0 2.1117743704417236e-03
GC_7_253 b_7 NI_7 NS_253 0 -1.1845645614010351e-06
GC_7_254 b_7 NI_7 NS_254 0 9.0485614621172880e-06
GC_7_255 b_7 NI_7 NS_255 0 8.9383790640334472e-04
GC_7_256 b_7 NI_7 NS_256 0 -4.6641889240103194e-04
GC_7_257 b_7 NI_7 NS_257 0 -1.0904722201934424e-05
GC_7_258 b_7 NI_7 NS_258 0 -8.7298638041021899e-06
GC_7_259 b_7 NI_7 NS_259 0 2.4742799158168492e-06
GC_7_260 b_7 NI_7 NS_260 0 -1.9522346988261633e-06
GC_7_261 b_7 NI_7 NS_261 0 2.5702271715648011e-06
GC_7_262 b_7 NI_7 NS_262 0 -5.3615507586756008e-07
GC_7_263 b_7 NI_7 NS_263 0 9.3122811898031194e-05
GC_7_264 b_7 NI_7 NS_264 0 -1.4546258525853303e-04
GC_7_265 b_7 NI_7 NS_265 0 -6.6494762477659369e-02
GC_7_266 b_7 NI_7 NS_266 0 9.5222185336713665e-03
GC_7_267 b_7 NI_7 NS_267 0 3.3251563225004002e-03
GC_7_268 b_7 NI_7 NS_268 0 6.1666298301850169e-03
GC_7_269 b_7 NI_7 NS_269 0 1.1107800458305147e-02
GC_7_270 b_7 NI_7 NS_270 0 -2.0149036987123408e-03
GC_7_271 b_7 NI_7 NS_271 0 1.3498531998863538e-03
GC_7_272 b_7 NI_7 NS_272 0 2.9521017623217774e-04
GC_7_273 b_7 NI_7 NS_273 0 4.8846429154445880e-04
GC_7_274 b_7 NI_7 NS_274 0 3.2727632371526479e-03
GC_7_275 b_7 NI_7 NS_275 0 2.8251501620791264e-03
GC_7_276 b_7 NI_7 NS_276 0 1.8041991044350596e-03
GC_7_277 b_7 NI_7 NS_277 0 5.9160532635601311e-04
GC_7_278 b_7 NI_7 NS_278 0 2.4409710067768174e-04
GC_7_279 b_7 NI_7 NS_279 0 6.8785585268744493e-03
GC_7_280 b_7 NI_7 NS_280 0 1.7164826902234382e-03
GC_7_281 b_7 NI_7 NS_281 0 9.9251747402730264e-06
GC_7_282 b_7 NI_7 NS_282 0 1.8677444277298373e-04
GC_7_283 b_7 NI_7 NS_283 0 -2.9258037410407196e-04
GC_7_284 b_7 NI_7 NS_284 0 -1.7103636201394644e-04
GC_7_285 b_7 NI_7 NS_285 0 -8.4508225671216014e-04
GC_7_286 b_7 NI_7 NS_286 0 -4.8324404273654612e-05
GC_7_287 b_7 NI_7 NS_287 0 1.7314882799633410e-04
GC_7_288 b_7 NI_7 NS_288 0 1.9594268058376846e-05
GC_7_289 b_7 NI_7 NS_289 0 5.7380937927632977e-05
GC_7_290 b_7 NI_7 NS_290 0 -3.5219650554357396e-05
GC_7_291 b_7 NI_7 NS_291 0 1.8926565137964351e-04
GC_7_292 b_7 NI_7 NS_292 0 1.3528903667732005e-02
GC_7_293 b_7 NI_7 NS_293 0 -2.6458324386558524e-06
GC_7_294 b_7 NI_7 NS_294 0 -2.3999964122856930e-05
GC_7_295 b_7 NI_7 NS_295 0 3.7524971306963036e-03
GC_7_296 b_7 NI_7 NS_296 0 -3.5266096927151942e-03
GC_7_297 b_7 NI_7 NS_297 0 7.7463329619347689e-06
GC_7_298 b_7 NI_7 NS_298 0 -2.3390922074122061e-05
GC_7_299 b_7 NI_7 NS_299 0 -2.4081133114190034e-03
GC_7_300 b_7 NI_7 NS_300 0 2.3176199539476339e-04
GC_7_301 b_7 NI_7 NS_301 0 1.6776462230667103e-05
GC_7_302 b_7 NI_7 NS_302 0 3.7607295901718968e-05
GC_7_303 b_7 NI_7 NS_303 0 -7.0258918117164391e-06
GC_7_304 b_7 NI_7 NS_304 0 3.9133226425838692e-06
GC_7_305 b_7 NI_7 NS_305 0 -1.5806428880474016e-07
GC_7_306 b_7 NI_7 NS_306 0 -1.2355249164985502e-05
GC_7_307 b_7 NI_7 NS_307 0 -3.8022028875125231e-04
GC_7_308 b_7 NI_7 NS_308 0 -2.0923481084399824e-04
GC_7_309 b_7 NI_7 NS_309 0 -4.5821523658044283e-03
GC_7_310 b_7 NI_7 NS_310 0 1.0788925958565686e-02
GC_7_311 b_7 NI_7 NS_311 0 -6.5333831447196766e-03
GC_7_312 b_7 NI_7 NS_312 0 -5.4371970102081116e-03
GC_7_313 b_7 NI_7 NS_313 0 -1.0914481872779833e-02
GC_7_314 b_7 NI_7 NS_314 0 1.2736385743768552e-03
GC_7_315 b_7 NI_7 NS_315 0 -9.4819069836860580e-05
GC_7_316 b_7 NI_7 NS_316 0 3.9069242484353627e-04
GC_7_317 b_7 NI_7 NS_317 0 1.4774361920882365e-03
GC_7_318 b_7 NI_7 NS_318 0 1.4368899447882041e-03
GC_7_319 b_7 NI_7 NS_319 0 3.6435127131149783e-03
GC_7_320 b_7 NI_7 NS_320 0 -1.8516237880199630e-03
GC_7_321 b_7 NI_7 NS_321 0 2.6133282809248685e-05
GC_7_322 b_7 NI_7 NS_322 0 2.1621467225545540e-04
GC_7_323 b_7 NI_7 NS_323 0 3.9921421230628210e-03
GC_7_324 b_7 NI_7 NS_324 0 -7.4621132918073767e-04
GC_7_325 b_7 NI_7 NS_325 0 -3.0089941978086058e-05
GC_7_326 b_7 NI_7 NS_326 0 6.8046501633328924e-06
GC_7_327 b_7 NI_7 NS_327 0 5.6442616583170571e-04
GC_7_328 b_7 NI_7 NS_328 0 4.3238635481732303e-04
GC_7_329 b_7 NI_7 NS_329 0 -1.2482521398954970e-04
GC_7_330 b_7 NI_7 NS_330 0 -1.7680257590173658e-04
GC_7_331 b_7 NI_7 NS_331 0 1.1211226811617114e-05
GC_7_332 b_7 NI_7 NS_332 0 -1.6761100512086912e-05
GC_7_333 b_7 NI_7 NS_333 0 -1.2439218072072848e-05
GC_7_334 b_7 NI_7 NS_334 0 4.9587571208924681e-05
GC_7_335 b_7 NI_7 NS_335 0 -1.6187039380390774e-03
GC_7_336 b_7 NI_7 NS_336 0 1.4493921262166637e-03
GC_7_337 b_7 NI_7 NS_337 0 1.2389723295603609e-07
GC_7_338 b_7 NI_7 NS_338 0 9.2817258227532540e-06
GC_7_339 b_7 NI_7 NS_339 0 4.2359656730646487e-04
GC_7_340 b_7 NI_7 NS_340 0 3.4854987842622469e-04
GC_7_341 b_7 NI_7 NS_341 0 3.0184122581906815e-06
GC_7_342 b_7 NI_7 NS_342 0 -3.0791218879052865e-06
GC_7_343 b_7 NI_7 NS_343 0 -4.3096361546171157e-04
GC_7_344 b_7 NI_7 NS_344 0 -4.5112539915902937e-04
GC_7_345 b_7 NI_7 NS_345 0 -1.1581514634486947e-06
GC_7_346 b_7 NI_7 NS_346 0 6.1494073705939346e-06
GC_7_347 b_7 NI_7 NS_347 0 -1.0684323054328656e-06
GC_7_348 b_7 NI_7 NS_348 0 -4.0127851117258884e-07
GC_7_349 b_7 NI_7 NS_349 0 1.0169324583284768e-06
GC_7_350 b_7 NI_7 NS_350 0 -3.7111724868456058e-06
GC_7_351 b_7 NI_7 NS_351 0 -8.8087432341110068e-05
GC_7_352 b_7 NI_7 NS_352 0 -1.2028649345859139e-04
GC_7_353 b_7 NI_7 NS_353 0 3.5834678521060532e-03
GC_7_354 b_7 NI_7 NS_354 0 8.0313721368173964e-05
GC_7_355 b_7 NI_7 NS_355 0 1.2125857014403337e-03
GC_7_356 b_7 NI_7 NS_356 0 -2.7628360310693044e-04
GC_7_357 b_7 NI_7 NS_357 0 -6.4692423473338291e-04
GC_7_358 b_7 NI_7 NS_358 0 4.4659637773701133e-04
GC_7_359 b_7 NI_7 NS_359 0 2.1428901980793000e-04
GC_7_360 b_7 NI_7 NS_360 0 -2.5603165591254746e-04
GC_7_361 b_7 NI_7 NS_361 0 8.2635413568237686e-04
GC_7_362 b_7 NI_7 NS_362 0 6.1218140992108986e-04
GC_7_363 b_7 NI_7 NS_363 0 -2.6080396907017965e-03
GC_7_364 b_7 NI_7 NS_364 0 -1.5666489054060174e-03
GC_7_365 b_7 NI_7 NS_365 0 5.5976536102705584e-04
GC_7_366 b_7 NI_7 NS_366 0 -4.2694680618673021e-04
GC_7_367 b_7 NI_7 NS_367 0 4.7026602460860873e-03
GC_7_368 b_7 NI_7 NS_368 0 2.6472777831841566e-04
GC_7_369 b_7 NI_7 NS_369 0 2.5844773429801603e-04
GC_7_370 b_7 NI_7 NS_370 0 2.9271130743307983e-04
GC_7_371 b_7 NI_7 NS_371 0 -2.8765856144508735e-04
GC_7_372 b_7 NI_7 NS_372 0 2.0760526355505476e-03
GC_7_373 b_7 NI_7 NS_373 0 3.8090031711596195e-04
GC_7_374 b_7 NI_7 NS_374 0 -2.4005240876429377e-04
GC_7_375 b_7 NI_7 NS_375 0 1.5716287449247428e-04
GC_7_376 b_7 NI_7 NS_376 0 -3.5218565516665886e-05
GC_7_377 b_7 NI_7 NS_377 0 2.0202027053944267e-05
GC_7_378 b_7 NI_7 NS_378 0 8.2366507970074157e-05
GC_7_379 b_7 NI_7 NS_379 0 -5.3580682666611833e-03
GC_7_380 b_7 NI_7 NS_380 0 3.7167113723961969e-03
GC_7_381 b_7 NI_7 NS_381 0 7.9503335385362543e-06
GC_7_382 b_7 NI_7 NS_382 0 -7.0044734454111343e-06
GC_7_383 b_7 NI_7 NS_383 0 1.3621321753052209e-03
GC_7_384 b_7 NI_7 NS_384 0 -5.3201538374183924e-04
GC_7_385 b_7 NI_7 NS_385 0 -9.0546419352635080e-07
GC_7_386 b_7 NI_7 NS_386 0 4.3015069194720401e-06
GC_7_387 b_7 NI_7 NS_387 0 7.7188888909667154e-05
GC_7_388 b_7 NI_7 NS_388 0 -1.8474386960385981e-03
GC_7_389 b_7 NI_7 NS_389 0 -1.4193057448472648e-05
GC_7_390 b_7 NI_7 NS_390 0 4.7812196329167757e-07
GC_7_391 b_7 NI_7 NS_391 0 9.7442154904529834e-07
GC_7_392 b_7 NI_7 NS_392 0 -5.4921797321363542e-07
GC_7_393 b_7 NI_7 NS_393 0 1.0258930376172071e-06
GC_7_394 b_7 NI_7 NS_394 0 3.0913345035619029e-06
GC_7_395 b_7 NI_7 NS_395 0 6.4165385829198158e-06
GC_7_396 b_7 NI_7 NS_396 0 -5.4179235905194001e-04
GC_7_397 b_7 NI_7 NS_397 0 -6.2322634912590378e-03
GC_7_398 b_7 NI_7 NS_398 0 -1.2416071891481447e-05
GC_7_399 b_7 NI_7 NS_399 0 -1.3035774726316519e-03
GC_7_400 b_7 NI_7 NS_400 0 1.9884360932651425e-04
GC_7_401 b_7 NI_7 NS_401 0 6.2664041871043550e-04
GC_7_402 b_7 NI_7 NS_402 0 -1.2431051798743077e-03
GC_7_403 b_7 NI_7 NS_403 0 1.7210278963165896e-04
GC_7_404 b_7 NI_7 NS_404 0 4.2920511801935069e-04
GC_7_405 b_7 NI_7 NS_405 0 6.8009317943040553e-04
GC_7_406 b_7 NI_7 NS_406 0 -1.5853185863710567e-04
GC_7_407 b_7 NI_7 NS_407 0 -3.0814038139756966e-04
GC_7_408 b_7 NI_7 NS_408 0 -1.1173399442914852e-03
GC_7_409 b_7 NI_7 NS_409 0 1.2333963613156033e-04
GC_7_410 b_7 NI_7 NS_410 0 8.7534403680851556e-05
GC_7_411 b_7 NI_7 NS_411 0 9.0830992530396783e-04
GC_7_412 b_7 NI_7 NS_412 0 1.1149235050858196e-03
GC_7_413 b_7 NI_7 NS_413 0 -1.2352304983248894e-04
GC_7_414 b_7 NI_7 NS_414 0 4.6413235105364170e-05
GC_7_415 b_7 NI_7 NS_415 0 -2.7408836361522470e-04
GC_7_416 b_7 NI_7 NS_416 0 -1.3257425720715135e-04
GC_7_417 b_7 NI_7 NS_417 0 -8.6050522862137377e-06
GC_7_418 b_7 NI_7 NS_418 0 1.0950272477430510e-04
GC_7_419 b_7 NI_7 NS_419 0 -1.8675625068203713e-05
GC_7_420 b_7 NI_7 NS_420 0 -1.1250038395602193e-04
GC_7_421 b_7 NI_7 NS_421 0 -2.4144023940579036e-05
GC_7_422 b_7 NI_7 NS_422 0 1.0005723471235129e-04
GC_7_423 b_7 NI_7 NS_423 0 1.6840836981850476e-03
GC_7_424 b_7 NI_7 NS_424 0 4.0776072417039369e-04
GC_7_425 b_7 NI_7 NS_425 0 -1.9460197963427897e-05
GC_7_426 b_7 NI_7 NS_426 0 -5.2366315431364974e-06
GC_7_427 b_7 NI_7 NS_427 0 -5.0767072267578434e-04
GC_7_428 b_7 NI_7 NS_428 0 -5.8499862185243910e-04
GC_7_429 b_7 NI_7 NS_429 0 -2.9905042436320838e-06
GC_7_430 b_7 NI_7 NS_430 0 -1.1786801177474877e-06
GC_7_431 b_7 NI_7 NS_431 0 4.1730246312260866e-05
GC_7_432 b_7 NI_7 NS_432 0 1.3928214582228655e-05
GC_7_433 b_7 NI_7 NS_433 0 -7.3520328696277384e-06
GC_7_434 b_7 NI_7 NS_434 0 -1.3797200575740811e-05
GC_7_435 b_7 NI_7 NS_435 0 2.5650292630520437e-07
GC_7_436 b_7 NI_7 NS_436 0 -2.1526931200278170e-07
GC_7_437 b_7 NI_7 NS_437 0 -7.7261866481780742e-07
GC_7_438 b_7 NI_7 NS_438 0 -4.5527832812121016e-07
GC_7_439 b_7 NI_7 NS_439 0 -1.9540881946221276e-04
GC_7_440 b_7 NI_7 NS_440 0 -4.7659893093569407e-05
GC_7_441 b_7 NI_7 NS_441 0 -2.1746756486062023e-02
GC_7_442 b_7 NI_7 NS_442 0 5.8937899901301319e-05
GC_7_443 b_7 NI_7 NS_443 0 1.0843242476638178e-03
GC_7_444 b_7 NI_7 NS_444 0 9.6537558233263359e-04
GC_7_445 b_7 NI_7 NS_445 0 -1.0198865006342684e-03
GC_7_446 b_7 NI_7 NS_446 0 -2.3849025650808779e-03
GC_7_447 b_7 NI_7 NS_447 0 1.4595521117558656e-04
GC_7_448 b_7 NI_7 NS_448 0 2.5884633111860689e-04
GC_7_449 b_7 NI_7 NS_449 0 8.4426091525658352e-04
GC_7_450 b_7 NI_7 NS_450 0 6.7751307326670545e-04
GC_7_451 b_7 NI_7 NS_451 0 -2.4390665898987263e-04
GC_7_452 b_7 NI_7 NS_452 0 -2.0975094874955847e-03
GC_7_453 b_7 NI_7 NS_453 0 4.5037889464466090e-04
GC_7_454 b_7 NI_7 NS_454 0 -1.9869603242855737e-04
GC_7_455 b_7 NI_7 NS_455 0 3.5419877997764169e-03
GC_7_456 b_7 NI_7 NS_456 0 -1.3881278338688673e-03
GC_7_457 b_7 NI_7 NS_457 0 1.5488187442919073e-04
GC_7_458 b_7 NI_7 NS_458 0 2.3487517886527007e-04
GC_7_459 b_7 NI_7 NS_459 0 6.6774674880512343e-06
GC_7_460 b_7 NI_7 NS_460 0 1.7467335404571670e-03
GC_7_461 b_7 NI_7 NS_461 0 4.4000232228377664e-04
GC_7_462 b_7 NI_7 NS_462 0 -9.5748361107440545e-05
GC_7_463 b_7 NI_7 NS_463 0 1.3346714377526913e-04
GC_7_464 b_7 NI_7 NS_464 0 -8.4655146310459243e-06
GC_7_465 b_7 NI_7 NS_465 0 2.9929389938409207e-05
GC_7_466 b_7 NI_7 NS_466 0 4.9975086173554425e-05
GC_7_467 b_7 NI_7 NS_467 0 -1.4185634012040078e-03
GC_7_468 b_7 NI_7 NS_468 0 4.3874626584350859e-03
GC_7_469 b_7 NI_7 NS_469 0 2.7557404677616182e-06
GC_7_470 b_7 NI_7 NS_470 0 -1.0689923345248595e-05
GC_7_471 b_7 NI_7 NS_471 0 1.2492459767292031e-03
GC_7_472 b_7 NI_7 NS_472 0 -1.2779703733938749e-03
GC_7_473 b_7 NI_7 NS_473 0 -2.2594999772547222e-06
GC_7_474 b_7 NI_7 NS_474 0 6.3091793563155254e-07
GC_7_475 b_7 NI_7 NS_475 0 -2.3206754678886394e-04
GC_7_476 b_7 NI_7 NS_476 0 -6.1637128587119173e-04
GC_7_477 b_7 NI_7 NS_477 0 -4.3786769071513617e-06
GC_7_478 b_7 NI_7 NS_478 0 2.9645673122955204e-06
GC_7_479 b_7 NI_7 NS_479 0 -4.9355590017084711e-07
GC_7_480 b_7 NI_7 NS_480 0 9.8927474165977298e-07
GC_7_481 b_7 NI_7 NS_481 0 -6.7785015205748306e-07
GC_7_482 b_7 NI_7 NS_482 0 2.1152219998159034e-07
GC_7_483 b_7 NI_7 NS_483 0 -8.3278584173612029e-05
GC_7_484 b_7 NI_7 NS_484 0 -3.2379209763017992e-04
GC_7_485 b_7 NI_7 NS_485 0 2.7416821051744677e-03
GC_7_486 b_7 NI_7 NS_486 0 4.1168496060369298e-05
GC_7_487 b_7 NI_7 NS_487 0 -1.7998031526982130e-03
GC_7_488 b_7 NI_7 NS_488 0 -1.0956975879269052e-03
GC_7_489 b_7 NI_7 NS_489 0 1.4061287677669702e-03
GC_7_490 b_7 NI_7 NS_490 0 7.0213036244794430e-04
GC_7_491 b_7 NI_7 NS_491 0 4.4494701196522576e-05
GC_7_492 b_7 NI_7 NS_492 0 6.0761409587553249e-05
GC_7_493 b_7 NI_7 NS_493 0 4.0868527090343640e-04
GC_7_494 b_7 NI_7 NS_494 0 2.8035047528832149e-05
GC_7_495 b_7 NI_7 NS_495 0 6.1039431010325243e-04
GC_7_496 b_7 NI_7 NS_496 0 -1.3317933062690285e-03
GC_7_497 b_7 NI_7 NS_497 0 4.2358957621109143e-05
GC_7_498 b_7 NI_7 NS_498 0 1.2273835103457644e-04
GC_7_499 b_7 NI_7 NS_499 0 9.7907625504608243e-06
GC_7_500 b_7 NI_7 NS_500 0 7.0033702328739012e-04
GC_7_501 b_7 NI_7 NS_501 0 -8.1819293742038611e-05
GC_7_502 b_7 NI_7 NS_502 0 2.7092583159589771e-05
GC_7_503 b_7 NI_7 NS_503 0 -2.0444835460940776e-04
GC_7_504 b_7 NI_7 NS_504 0 2.8030879045222912e-04
GC_7_505 b_7 NI_7 NS_505 0 -4.0192522846451143e-05
GC_7_506 b_7 NI_7 NS_506 0 1.2817891199304503e-04
GC_7_507 b_7 NI_7 NS_507 0 -1.8759764288480388e-05
GC_7_508 b_7 NI_7 NS_508 0 -5.5203906826557110e-05
GC_7_509 b_7 NI_7 NS_509 0 -1.2490526482841677e-05
GC_7_510 b_7 NI_7 NS_510 0 6.3122935733742955e-05
GC_7_511 b_7 NI_7 NS_511 0 1.9078896463457667e-04
GC_7_512 b_7 NI_7 NS_512 0 4.4062811585763624e-04
GC_7_513 b_7 NI_7 NS_513 0 -9.5864328014227382e-06
GC_7_514 b_7 NI_7 NS_514 0 -2.3338414428524787e-06
GC_7_515 b_7 NI_7 NS_515 0 -9.9191687010027974e-05
GC_7_516 b_7 NI_7 NS_516 0 -3.7418946817470170e-05
GC_7_517 b_7 NI_7 NS_517 0 -1.0967008857644201e-06
GC_7_518 b_7 NI_7 NS_518 0 -6.6645484055876929e-07
GC_7_519 b_7 NI_7 NS_519 0 -4.7273373326054193e-05
GC_7_520 b_7 NI_7 NS_520 0 -8.4486612936809791e-05
GC_7_521 b_7 NI_7 NS_521 0 -3.2869429489985182e-06
GC_7_522 b_7 NI_7 NS_522 0 -5.2571843707229419e-06
GC_7_523 b_7 NI_7 NS_523 0 2.8977119062965852e-08
GC_7_524 b_7 NI_7 NS_524 0 -1.8341953377811822e-07
GC_7_525 b_7 NI_7 NS_525 0 -1.9804352512996423e-07
GC_7_526 b_7 NI_7 NS_526 0 -6.8285135728515926e-07
GC_7_527 b_7 NI_7 NS_527 0 -8.7484558678843332e-05
GC_7_528 b_7 NI_7 NS_528 0 -3.9080144657133506e-05
GD_7_1 b_7 NI_7 NA_1 0 -7.3137574930142359e-03
GD_7_2 b_7 NI_7 NA_2 0 -1.9300869900852460e-02
GD_7_3 b_7 NI_7 NA_3 0 -3.3528076124910648e-02
GD_7_4 b_7 NI_7 NA_4 0 -3.3792607450468061e-02
GD_7_5 b_7 NI_7 NA_5 0 3.1661145475003721e-03
GD_7_6 b_7 NI_7 NA_6 0 -6.3855611028907952e-02
GD_7_7 b_7 NI_7 NA_7 0 -1.0515167052926983e-01
GD_7_8 b_7 NI_7 NA_8 0 2.2066460413501855e-03
GD_7_9 b_7 NI_7 NA_9 0 -7.4851737810537637e-03
GD_7_10 b_7 NI_7 NA_10 0 4.0000538907056550e-03
GD_7_11 b_7 NI_7 NA_11 0 1.5477922166694339e-02
GD_7_12 b_7 NI_7 NA_12 0 -4.8329132536223162e-03
*
* Port 8
VI_8 a_8 NI_8 0
RI_8 NI_8 b_8 5.0000000000000000e+01
GC_8_1 b_8 NI_8 NS_1 0 2.4593395635663318e-02
GC_8_2 b_8 NI_8 NS_2 0 -2.7114935219866605e-04
GC_8_3 b_8 NI_8 NS_3 0 -3.1075014061171932e-03
GC_8_4 b_8 NI_8 NS_4 0 2.1556221558027121e-03
GC_8_5 b_8 NI_8 NS_5 0 -1.6908285272954388e-04
GC_8_6 b_8 NI_8 NS_6 0 -2.9744396168026625e-03
GC_8_7 b_8 NI_8 NS_7 0 7.5991706571492936e-05
GC_8_8 b_8 NI_8 NS_8 0 -2.4659598439688205e-04
GC_8_9 b_8 NI_8 NS_9 0 1.4466916131144097e-03
GC_8_10 b_8 NI_8 NS_10 0 9.0058273375874726e-04
GC_8_11 b_8 NI_8 NS_11 0 -5.0460613125547097e-03
GC_8_12 b_8 NI_8 NS_12 0 8.7682714812494303e-04
GC_8_13 b_8 NI_8 NS_13 0 3.0130002312446856e-05
GC_8_14 b_8 NI_8 NS_14 0 4.0039850070300280e-07
GC_8_15 b_8 NI_8 NS_15 0 1.8645445617464980e-04
GC_8_16 b_8 NI_8 NS_16 0 -1.9818018239608063e-03
GC_8_17 b_8 NI_8 NS_17 0 -2.0176917698719751e-05
GC_8_18 b_8 NI_8 NS_18 0 -3.9507402810761220e-05
GC_8_19 b_8 NI_8 NS_19 0 2.8860100237410876e-04
GC_8_20 b_8 NI_8 NS_20 0 -4.9452534621776642e-06
GC_8_21 b_8 NI_8 NS_21 0 7.1942322661314954e-05
GC_8_22 b_8 NI_8 NS_22 0 3.7908807969966141e-06
GC_8_23 b_8 NI_8 NS_23 0 1.1194651049055135e-05
GC_8_24 b_8 NI_8 NS_24 0 -4.4453585838356961e-05
GC_8_25 b_8 NI_8 NS_25 0 -3.1554967380579020e-05
GC_8_26 b_8 NI_8 NS_26 0 3.3040657505303318e-05
GC_8_27 b_8 NI_8 NS_27 0 9.3944094738243654e-04
GC_8_28 b_8 NI_8 NS_28 0 -2.6364004916283475e-03
GC_8_29 b_8 NI_8 NS_29 0 -1.2270495974473855e-07
GC_8_30 b_8 NI_8 NS_30 0 1.9316389583385848e-05
GC_8_31 b_8 NI_8 NS_31 0 -8.6168010273659362e-04
GC_8_32 b_8 NI_8 NS_32 0 4.2423950693609139e-04
GC_8_33 b_8 NI_8 NS_33 0 -1.8533796811325924e-06
GC_8_34 b_8 NI_8 NS_34 0 6.8712208291206232e-07
GC_8_35 b_8 NI_8 NS_35 0 3.4391126449299930e-04
GC_8_36 b_8 NI_8 NS_36 0 1.6790993967036010e-04
GC_8_37 b_8 NI_8 NS_37 0 8.0359013757229361e-07
GC_8_38 b_8 NI_8 NS_38 0 -5.0402799774972350e-06
GC_8_39 b_8 NI_8 NS_39 0 5.9990434497557396e-07
GC_8_40 b_8 NI_8 NS_40 0 1.8242004973731380e-06
GC_8_41 b_8 NI_8 NS_41 0 -1.2684532558888763e-06
GC_8_42 b_8 NI_8 NS_42 0 3.3700600991404728e-07
GC_8_43 b_8 NI_8 NS_43 0 1.1952390334586036e-05
GC_8_44 b_8 NI_8 NS_44 0 -4.1352774876995469e-06
GC_8_45 b_8 NI_8 NS_45 0 8.6673466856446914e-03
GC_8_46 b_8 NI_8 NS_46 0 -2.9984941057195073e-05
GC_8_47 b_8 NI_8 NS_47 0 2.1816743945560772e-03
GC_8_48 b_8 NI_8 NS_48 0 -2.1543335272455554e-03
GC_8_49 b_8 NI_8 NS_49 0 4.7628283025565185e-04
GC_8_50 b_8 NI_8 NS_50 0 2.8951595500022100e-03
GC_8_51 b_8 NI_8 NS_51 0 -6.1397029163312415e-04
GC_8_52 b_8 NI_8 NS_52 0 1.0765340969343003e-03
GC_8_53 b_8 NI_8 NS_53 0 8.2212247297831526e-04
GC_8_54 b_8 NI_8 NS_54 0 5.1234698847225349e-04
GC_8_55 b_8 NI_8 NS_55 0 -7.4259407369527358e-04
GC_8_56 b_8 NI_8 NS_56 0 2.1129567376339635e-03
GC_8_57 b_8 NI_8 NS_57 0 -6.1191759673204988e-05
GC_8_58 b_8 NI_8 NS_58 0 1.4744946937292393e-05
GC_8_59 b_8 NI_8 NS_59 0 -2.2804571893777318e-04
GC_8_60 b_8 NI_8 NS_60 0 6.5316934905777183e-04
GC_8_61 b_8 NI_8 NS_61 0 -1.5995759626839670e-06
GC_8_62 b_8 NI_8 NS_62 0 -1.2931702807115667e-06
GC_8_63 b_8 NI_8 NS_63 0 -2.8228159302209118e-04
GC_8_64 b_8 NI_8 NS_64 0 4.2644225259329011e-04
GC_8_65 b_8 NI_8 NS_65 0 3.8310011445206115e-04
GC_8_66 b_8 NI_8 NS_66 0 -1.1535321348205964e-04
GC_8_67 b_8 NI_8 NS_67 0 -3.4956354091090015e-05
GC_8_68 b_8 NI_8 NS_68 0 1.4524549544787352e-08
GC_8_69 b_8 NI_8 NS_69 0 -3.1199052874975391e-05
GC_8_70 b_8 NI_8 NS_70 0 -5.2999155684376183e-05
GC_8_71 b_8 NI_8 NS_71 0 -3.2585180293578713e-03
GC_8_72 b_8 NI_8 NS_72 0 -2.4625876749988567e-03
GC_8_73 b_8 NI_8 NS_73 0 -1.2474920979436765e-05
GC_8_74 b_8 NI_8 NS_74 0 -2.2356700288140441e-05
GC_8_75 b_8 NI_8 NS_75 0 8.9320177560216381e-04
GC_8_76 b_8 NI_8 NS_76 0 1.1299644973896659e-03
GC_8_77 b_8 NI_8 NS_77 0 -6.0030462613161338e-06
GC_8_78 b_8 NI_8 NS_78 0 1.6306029807388328e-05
GC_8_79 b_8 NI_8 NS_79 0 8.9863476524265542e-04
GC_8_80 b_8 NI_8 NS_80 0 -5.2531439816253282e-04
GC_8_81 b_8 NI_8 NS_81 0 -1.6778739700989552e-05
GC_8_82 b_8 NI_8 NS_82 0 -1.4778186090356306e-05
GC_8_83 b_8 NI_8 NS_83 0 1.8946097026276836e-05
GC_8_84 b_8 NI_8 NS_84 0 -2.7209500099856703e-06
GC_8_85 b_8 NI_8 NS_85 0 1.9862635423631519e-05
GC_8_86 b_8 NI_8 NS_86 0 -1.9588298801400901e-06
GC_8_87 b_8 NI_8 NS_87 0 9.0585069250316013e-05
GC_8_88 b_8 NI_8 NS_88 0 7.8226261893442641e-06
GC_8_89 b_8 NI_8 NS_89 0 3.9278846319616319e-02
GC_8_90 b_8 NI_8 NS_90 0 -2.3265152077309051e-04
GC_8_91 b_8 NI_8 NS_91 0 -5.5253451610276366e-03
GC_8_92 b_8 NI_8 NS_92 0 6.2104283207451024e-04
GC_8_93 b_8 NI_8 NS_93 0 2.5852580646764265e-03
GC_8_94 b_8 NI_8 NS_94 0 -2.3322111819087297e-03
GC_8_95 b_8 NI_8 NS_95 0 -1.2110043366567674e-04
GC_8_96 b_8 NI_8 NS_96 0 -1.0841748016520446e-04
GC_8_97 b_8 NI_8 NS_97 0 2.1251555571973470e-03
GC_8_98 b_8 NI_8 NS_98 0 1.5334216510319613e-03
GC_8_99 b_8 NI_8 NS_99 0 -3.5719108322565776e-03
GC_8_100 b_8 NI_8 NS_100 0 -2.5194945395030921e-04
GC_8_101 b_8 NI_8 NS_101 0 2.5534493275795878e-05
GC_8_102 b_8 NI_8 NS_102 0 5.0696215903984527e-05
GC_8_103 b_8 NI_8 NS_103 0 -1.1603657122755098e-03
GC_8_104 b_8 NI_8 NS_104 0 4.3393020805183435e-04
GC_8_105 b_8 NI_8 NS_105 0 -4.0767606299660926e-05
GC_8_106 b_8 NI_8 NS_106 0 -4.9184528492342711e-05
GC_8_107 b_8 NI_8 NS_107 0 1.6115967684340282e-04
GC_8_108 b_8 NI_8 NS_108 0 3.2723857613347268e-04
GC_8_109 b_8 NI_8 NS_109 0 1.7364231065572722e-04
GC_8_110 b_8 NI_8 NS_110 0 2.0402195792500321e-05
GC_8_111 b_8 NI_8 NS_111 0 -1.9107067325678238e-06
GC_8_112 b_8 NI_8 NS_112 0 -5.3476859258656551e-05
GC_8_113 b_8 NI_8 NS_113 0 -4.4206306558365556e-05
GC_8_114 b_8 NI_8 NS_114 0 5.9070667225187056e-05
GC_8_115 b_8 NI_8 NS_115 0 -4.5025573590962652e-04
GC_8_116 b_8 NI_8 NS_116 0 -3.1591330044269603e-03
GC_8_117 b_8 NI_8 NS_117 0 1.9145429707028403e-06
GC_8_118 b_8 NI_8 NS_118 0 2.6495128071926067e-05
GC_8_119 b_8 NI_8 NS_119 0 -8.6230308353456406e-04
GC_8_120 b_8 NI_8 NS_120 0 1.0286235613800731e-03
GC_8_121 b_8 NI_8 NS_121 0 2.6847871015320964e-07
GC_8_122 b_8 NI_8 NS_122 0 5.0567698566009330e-06
GC_8_123 b_8 NI_8 NS_123 0 5.7311274975334608e-04
GC_8_124 b_8 NI_8 NS_124 0 -1.0736585803470242e-04
GC_8_125 b_8 NI_8 NS_125 0 -4.3512627396367627e-06
GC_8_126 b_8 NI_8 NS_126 0 -4.8626484643761261e-06
GC_8_127 b_8 NI_8 NS_127 0 1.4331945468825050e-06
GC_8_128 b_8 NI_8 NS_128 0 2.7487829662134382e-07
GC_8_129 b_8 NI_8 NS_129 0 -2.4890050151989451e-07
GC_8_130 b_8 NI_8 NS_130 0 -5.5507407408408238e-07
GC_8_131 b_8 NI_8 NS_131 0 4.3337950634625972e-05
GC_8_132 b_8 NI_8 NS_132 0 -4.9008439799148626e-05
GC_8_133 b_8 NI_8 NS_133 0 1.4346644166532216e-02
GC_8_134 b_8 NI_8 NS_134 0 -3.2571209575321788e-04
GC_8_135 b_8 NI_8 NS_135 0 3.8560164645142767e-03
GC_8_136 b_8 NI_8 NS_136 0 -1.3456190143291361e-03
GC_8_137 b_8 NI_8 NS_137 0 -2.0590715974895522e-03
GC_8_138 b_8 NI_8 NS_138 0 2.4721393991014276e-03
GC_8_139 b_8 NI_8 NS_139 0 -4.7762474198232493e-04
GC_8_140 b_8 NI_8 NS_140 0 3.2548320179989624e-04
GC_8_141 b_8 NI_8 NS_141 0 9.9959767325172593e-04
GC_8_142 b_8 NI_8 NS_142 0 4.1630294471912461e-04
GC_8_143 b_8 NI_8 NS_143 0 -8.6285491442327422e-04
GC_8_144 b_8 NI_8 NS_144 0 1.3420833490423521e-03
GC_8_145 b_8 NI_8 NS_145 0 -6.3972814605936325e-05
GC_8_146 b_8 NI_8 NS_146 0 -3.3676946883496105e-05
GC_8_147 b_8 NI_8 NS_147 0 -7.0937095941846478e-04
GC_8_148 b_8 NI_8 NS_148 0 1.2971988290964578e-03
GC_8_149 b_8 NI_8 NS_149 0 2.2513531581429358e-06
GC_8_150 b_8 NI_8 NS_150 0 -1.5088578187585105e-05
GC_8_151 b_8 NI_8 NS_151 0 -3.1945186306644129e-04
GC_8_152 b_8 NI_8 NS_152 0 1.6807809331141404e-04
GC_8_153 b_8 NI_8 NS_153 0 3.6929719372194293e-04
GC_8_154 b_8 NI_8 NS_154 0 -1.5814388119498530e-04
GC_8_155 b_8 NI_8 NS_155 0 -3.4003789816100142e-05
GC_8_156 b_8 NI_8 NS_156 0 -1.8098843261341727e-05
GC_8_157 b_8 NI_8 NS_157 0 -4.3632733361989075e-05
GC_8_158 b_8 NI_8 NS_158 0 -7.0613142649465993e-05
GC_8_159 b_8 NI_8 NS_159 0 -2.4385716402016383e-03
GC_8_160 b_8 NI_8 NS_160 0 -1.9933288802154473e-03
GC_8_161 b_8 NI_8 NS_161 0 -1.8744992910007925e-05
GC_8_162 b_8 NI_8 NS_162 0 -2.2263668901584967e-05
GC_8_163 b_8 NI_8 NS_163 0 8.0829228771176756e-04
GC_8_164 b_8 NI_8 NS_164 0 6.8884903163412387e-04
GC_8_165 b_8 NI_8 NS_165 0 -2.1565200809653787e-06
GC_8_166 b_8 NI_8 NS_166 0 1.5281424702645663e-05
GC_8_167 b_8 NI_8 NS_167 0 6.3224990808630904e-04
GC_8_168 b_8 NI_8 NS_168 0 -4.6727514202602979e-04
GC_8_169 b_8 NI_8 NS_169 0 -7.4456206692949951e-06
GC_8_170 b_8 NI_8 NS_170 0 -7.5910541532498553e-06
GC_8_171 b_8 NI_8 NS_171 0 2.0564702571969638e-05
GC_8_172 b_8 NI_8 NS_172 0 -6.1114226711786471e-07
GC_8_173 b_8 NI_8 NS_173 0 1.9470775407895717e-05
GC_8_174 b_8 NI_8 NS_174 0 -2.5895216184176408e-06
GC_8_175 b_8 NI_8 NS_175 0 4.8596091375417920e-05
GC_8_176 b_8 NI_8 NS_176 0 3.8883970377356919e-05
GC_8_177 b_8 NI_8 NS_177 0 6.0421197827840410e-02
GC_8_178 b_8 NI_8 NS_178 0 -3.6827372911797645e-05
GC_8_179 b_8 NI_8 NS_179 0 -6.2389308911892640e-03
GC_8_180 b_8 NI_8 NS_180 0 -2.7366714953431250e-03
GC_8_181 b_8 NI_8 NS_181 0 4.3480874694045634e-03
GC_8_182 b_8 NI_8 NS_182 0 2.6774408416081366e-03
GC_8_183 b_8 NI_8 NS_183 0 1.1678547841684981e-05
GC_8_184 b_8 NI_8 NS_184 0 -1.7177681576738694e-04
GC_8_185 b_8 NI_8 NS_185 0 1.4030047732710585e-03
GC_8_186 b_8 NI_8 NS_186 0 1.5327719107316314e-03
GC_8_187 b_8 NI_8 NS_187 0 -1.6524998006924496e-04
GC_8_188 b_8 NI_8 NS_188 0 -5.5449878940516965e-04
GC_8_189 b_8 NI_8 NS_189 0 -4.4222879893705305e-05
GC_8_190 b_8 NI_8 NS_190 0 8.2932074075282283e-05
GC_8_191 b_8 NI_8 NS_191 0 -3.9348491174446970e-03
GC_8_192 b_8 NI_8 NS_192 0 9.0024826881519968e-04
GC_8_193 b_8 NI_8 NS_193 0 -7.6706357735892891e-05
GC_8_194 b_8 NI_8 NS_194 0 -4.7530693253196230e-05
GC_8_195 b_8 NI_8 NS_195 0 -2.6253121731623449e-04
GC_8_196 b_8 NI_8 NS_196 0 7.8548584454826329e-04
GC_8_197 b_8 NI_8 NS_197 0 3.7693847905193479e-04
GC_8_198 b_8 NI_8 NS_198 0 7.5655003871510690e-05
GC_8_199 b_8 NI_8 NS_199 0 -2.9752808509463622e-05
GC_8_200 b_8 NI_8 NS_200 0 -4.3987289638661705e-05
GC_8_201 b_8 NI_8 NS_201 0 -3.6114408045871269e-05
GC_8_202 b_8 NI_8 NS_202 0 7.8741547459712543e-05
GC_8_203 b_8 NI_8 NS_203 0 -2.9776567208377883e-03
GC_8_204 b_8 NI_8 NS_204 0 -3.4609542499809743e-03
GC_8_205 b_8 NI_8 NS_205 0 9.4828012754501486e-06
GC_8_206 b_8 NI_8 NS_206 0 2.7662340651239988e-05
GC_8_207 b_8 NI_8 NS_207 0 -5.0479588604570419e-04
GC_8_208 b_8 NI_8 NS_208 0 1.9356741737958899e-03
GC_8_209 b_8 NI_8 NS_209 0 -2.3893783463969064e-07
GC_8_210 b_8 NI_8 NS_210 0 8.3496619134356910e-06
GC_8_211 b_8 NI_8 NS_211 0 8.4947825661724804e-04
GC_8_212 b_8 NI_8 NS_212 0 -4.7265474840161041e-04
GC_8_213 b_8 NI_8 NS_213 0 -1.0503840230757291e-05
GC_8_214 b_8 NI_8 NS_214 0 -8.1324124562096361e-06
GC_8_215 b_8 NI_8 NS_215 0 1.6478068570531525e-06
GC_8_216 b_8 NI_8 NS_216 0 -1.8081853728059508e-07
GC_8_217 b_8 NI_8 NS_217 0 2.8189705285236246e-06
GC_8_218 b_8 NI_8 NS_218 0 2.2727648644739650e-06
GC_8_219 b_8 NI_8 NS_219 0 9.6821179156039342e-05
GC_8_220 b_8 NI_8 NS_220 0 -1.1669203143134337e-04
GC_8_221 b_8 NI_8 NS_221 0 5.1376735148024226e-03
GC_8_222 b_8 NI_8 NS_222 0 -8.5693344052351940e-04
GC_8_223 b_8 NI_8 NS_223 0 4.0087013484640241e-03
GC_8_224 b_8 NI_8 NS_224 0 1.4684993441502275e-03
GC_8_225 b_8 NI_8 NS_225 0 -5.0365459478060558e-03
GC_8_226 b_8 NI_8 NS_226 0 -2.2501676135610483e-03
GC_8_227 b_8 NI_8 NS_227 0 8.8585647604431716e-05
GC_8_228 b_8 NI_8 NS_228 0 -4.7111936342334970e-05
GC_8_229 b_8 NI_8 NS_229 0 1.2781738230788844e-03
GC_8_230 b_8 NI_8 NS_230 0 7.9183488293519921e-05
GC_8_231 b_8 NI_8 NS_231 0 -6.1023622498442992e-05
GC_8_232 b_8 NI_8 NS_232 0 -6.7361576684991616e-04
GC_8_233 b_8 NI_8 NS_233 0 -1.5335861990188664e-05
GC_8_234 b_8 NI_8 NS_234 0 -3.8568167418970045e-05
GC_8_235 b_8 NI_8 NS_235 0 -9.7886818348638031e-04
GC_8_236 b_8 NI_8 NS_236 0 2.9189571120701399e-04
GC_8_237 b_8 NI_8 NS_237 0 3.3318511218339737e-05
GC_8_238 b_8 NI_8 NS_238 0 -2.7505581611540140e-05
GC_8_239 b_8 NI_8 NS_239 0 2.7376445230532895e-04
GC_8_240 b_8 NI_8 NS_240 0 -3.4607185238368733e-04
GC_8_241 b_8 NI_8 NS_241 0 2.5238630264112809e-04
GC_8_242 b_8 NI_8 NS_242 0 -1.6497682043412640e-04
GC_8_243 b_8 NI_8 NS_243 0 4.9667981146136705e-06
GC_8_244 b_8 NI_8 NS_244 0 -4.0538677631256138e-05
GC_8_245 b_8 NI_8 NS_245 0 -5.4313372911559373e-05
GC_8_246 b_8 NI_8 NS_246 0 -1.2916412901387993e-04
GC_8_247 b_8 NI_8 NS_247 0 1.4019882908662630e-03
GC_8_248 b_8 NI_8 NS_248 0 1.0625811332673066e-03
GC_8_249 b_8 NI_8 NS_249 0 -3.6553139040063846e-05
GC_8_250 b_8 NI_8 NS_250 0 -3.5152318726719637e-05
GC_8_251 b_8 NI_8 NS_251 0 1.1014908675481740e-03
GC_8_252 b_8 NI_8 NS_252 0 -1.0003693783473568e-03
GC_8_253 b_8 NI_8 NS_253 0 -4.7847417906557266e-06
GC_8_254 b_8 NI_8 NS_254 0 1.2027907655017784e-05
GC_8_255 b_8 NI_8 NS_255 0 1.7371194804376654e-04
GC_8_256 b_8 NI_8 NS_256 0 1.6458802078227148e-04
GC_8_257 b_8 NI_8 NS_257 0 -3.6207438447946017e-06
GC_8_258 b_8 NI_8 NS_258 0 -6.1269579384206531e-06
GC_8_259 b_8 NI_8 NS_259 0 2.6885551537030461e-05
GC_8_260 b_8 NI_8 NS_260 0 -1.7410672214440041e-07
GC_8_261 b_8 NI_8 NS_261 0 2.0594390266007675e-05
GC_8_262 b_8 NI_8 NS_262 0 -1.0279336532168936e-05
GC_8_263 b_8 NI_8 NS_263 0 -1.2397257946827225e-04
GC_8_264 b_8 NI_8 NS_264 0 1.7605344121835294e-04
GC_8_265 b_8 NI_8 NS_265 0 -4.5821523693421011e-03
GC_8_266 b_8 NI_8 NS_266 0 1.0788925958635483e-02
GC_8_267 b_8 NI_8 NS_267 0 -6.5333831445965199e-03
GC_8_268 b_8 NI_8 NS_268 0 -5.4371970104120848e-03
GC_8_269 b_8 NI_8 NS_269 0 -1.0914481872538680e-02
GC_8_270 b_8 NI_8 NS_270 0 1.2736385744278806e-03
GC_8_271 b_8 NI_8 NS_271 0 -9.4819069602320897e-05
GC_8_272 b_8 NI_8 NS_272 0 3.9069242513460319e-04
GC_8_273 b_8 NI_8 NS_273 0 1.4774361921807715e-03
GC_8_274 b_8 NI_8 NS_274 0 1.4368899447768082e-03
GC_8_275 b_8 NI_8 NS_275 0 3.6435127132210974e-03
GC_8_276 b_8 NI_8 NS_276 0 -1.8516237882379538e-03
GC_8_277 b_8 NI_8 NS_277 0 2.6133282825083650e-05
GC_8_278 b_8 NI_8 NS_278 0 2.1621467226400591e-04
GC_8_279 b_8 NI_8 NS_279 0 3.9921421234583457e-03
GC_8_280 b_8 NI_8 NS_280 0 -7.4621132924849694e-04
GC_8_281 b_8 NI_8 NS_281 0 -3.0089941973406912e-05
GC_8_282 b_8 NI_8 NS_282 0 6.8046501682177704e-06
GC_8_283 b_8 NI_8 NS_283 0 5.6442616599018192e-04
GC_8_284 b_8 NI_8 NS_284 0 4.3238635484186243e-04
GC_8_285 b_8 NI_8 NS_285 0 -1.2482521396169936e-04
GC_8_286 b_8 NI_8 NS_286 0 -1.7680257592016176e-04
GC_8_287 b_8 NI_8 NS_287 0 1.1211226818374743e-05
GC_8_288 b_8 NI_8 NS_288 0 -1.6761100506634154e-05
GC_8_289 b_8 NI_8 NS_289 0 -1.2439218067149084e-05
GC_8_290 b_8 NI_8 NS_290 0 4.9587571207105600e-05
GC_8_291 b_8 NI_8 NS_291 0 -1.6187039380756050e-03
GC_8_292 b_8 NI_8 NS_292 0 1.4493921269564329e-03
GC_8_293 b_8 NI_8 NS_293 0 1.2389723297253635e-07
GC_8_294 b_8 NI_8 NS_294 0 9.2817258208298607e-06
GC_8_295 b_8 NI_8 NS_295 0 4.2359656752067156e-04
GC_8_296 b_8 NI_8 NS_296 0 3.4854987827485142e-04
GC_8_297 b_8 NI_8 NS_297 0 3.0184122599443057e-06
GC_8_298 b_8 NI_8 NS_298 0 -3.0791218879930976e-06
GC_8_299 b_8 NI_8 NS_299 0 -4.3096361555056497e-04
GC_8_300 b_8 NI_8 NS_300 0 -4.5112539923784729e-04
GC_8_301 b_8 NI_8 NS_301 0 -1.1581514642817726e-06
GC_8_302 b_8 NI_8 NS_302 0 6.1494073731193219e-06
GC_8_303 b_8 NI_8 NS_303 0 -1.0684323060365693e-06
GC_8_304 b_8 NI_8 NS_304 0 -4.0127851121547984e-07
GC_8_305 b_8 NI_8 NS_305 0 1.0169324586937280e-06
GC_8_306 b_8 NI_8 NS_306 0 -3.7111724876794081e-06
GC_8_307 b_8 NI_8 NS_307 0 -8.8087432364060419e-05
GC_8_308 b_8 NI_8 NS_308 0 -1.2028649347907900e-04
GC_8_309 b_8 NI_8 NS_309 0 -2.1113478665757726e-01
GC_8_310 b_8 NI_8 NS_310 0 8.5660017210819200e-03
GC_8_311 b_8 NI_8 NS_311 0 4.0113681753027510e-03
GC_8_312 b_8 NI_8 NS_312 0 6.1391632821758404e-03
GC_8_313 b_8 NI_8 NS_313 0 6.6340605226096177e-03
GC_8_314 b_8 NI_8 NS_314 0 -1.4582428328252866e-03
GC_8_315 b_8 NI_8 NS_315 0 9.6516091993271525e-04
GC_8_316 b_8 NI_8 NS_316 0 -5.7822442219214152e-05
GC_8_317 b_8 NI_8 NS_317 0 1.4947863348180879e-04
GC_8_318 b_8 NI_8 NS_318 0 1.3893338081767521e-03
GC_8_319 b_8 NI_8 NS_319 0 4.9776329198209764e-03
GC_8_320 b_8 NI_8 NS_320 0 1.7638386187156436e-03
GC_8_321 b_8 NI_8 NS_321 0 -1.8932257614757327e-04
GC_8_322 b_8 NI_8 NS_322 0 2.9236482145448791e-04
GC_8_323 b_8 NI_8 NS_323 0 1.9617007500600117e-03
GC_8_324 b_8 NI_8 NS_324 0 7.3227104377111647e-03
GC_8_325 b_8 NI_8 NS_325 0 -7.3092588562402683e-05
GC_8_326 b_8 NI_8 NS_326 0 8.9723684537196575e-05
GC_8_327 b_8 NI_8 NS_327 0 -2.0782257059445868e-04
GC_8_328 b_8 NI_8 NS_328 0 3.3803981562061615e-03
GC_8_329 b_8 NI_8 NS_329 0 4.4141950030329187e-04
GC_8_330 b_8 NI_8 NS_330 0 -2.1456447925159131e-04
GC_8_331 b_8 NI_8 NS_331 0 -1.0785138575826919e-04
GC_8_332 b_8 NI_8 NS_332 0 1.4691137816012748e-04
GC_8_333 b_8 NI_8 NS_333 0 2.8120152879036509e-05
GC_8_334 b_8 NI_8 NS_334 0 2.9699388309969230e-05
GC_8_335 b_8 NI_8 NS_335 0 -1.9232751362500404e-02
GC_8_336 b_8 NI_8 NS_336 0 5.9467325243440692e-04
GC_8_337 b_8 NI_8 NS_337 0 3.1217608364754775e-05
GC_8_338 b_8 NI_8 NS_338 0 -2.2994374581603267e-05
GC_8_339 b_8 NI_8 NS_339 0 5.0846771120718988e-03
GC_8_340 b_8 NI_8 NS_340 0 4.6998071121847167e-03
GC_8_341 b_8 NI_8 NS_341 0 -2.4279142284932220e-07
GC_8_342 b_8 NI_8 NS_342 0 3.7834919412460354e-05
GC_8_343 b_8 NI_8 NS_343 0 1.4188869934566883e-03
GC_8_344 b_8 NI_8 NS_344 0 -2.5314470789937586e-03
GC_8_345 b_8 NI_8 NS_345 0 -5.5946119718608327e-05
GC_8_346 b_8 NI_8 NS_346 0 -1.9037153344232468e-05
GC_8_347 b_8 NI_8 NS_347 0 1.8118124101075809e-05
GC_8_348 b_8 NI_8 NS_348 0 -1.4358066116576021e-05
GC_8_349 b_8 NI_8 NS_349 0 3.1017329145465499e-05
GC_8_350 b_8 NI_8 NS_350 0 5.8871032118776386e-06
GC_8_351 b_8 NI_8 NS_351 0 4.6828400934348884e-04
GC_8_352 b_8 NI_8 NS_352 0 -5.1619220031633454e-04
GC_8_353 b_8 NI_8 NS_353 0 -3.3596046312003814e-03
GC_8_354 b_8 NI_8 NS_354 0 -1.5357282886155885e-05
GC_8_355 b_8 NI_8 NS_355 0 -1.2853688887098922e-03
GC_8_356 b_8 NI_8 NS_356 0 1.9144836475557033e-04
GC_8_357 b_8 NI_8 NS_357 0 6.4740289862914619e-04
GC_8_358 b_8 NI_8 NS_358 0 -1.1924884174172236e-03
GC_8_359 b_8 NI_8 NS_359 0 4.2127835039369701e-05
GC_8_360 b_8 NI_8 NS_360 0 3.5526847894747928e-04
GC_8_361 b_8 NI_8 NS_361 0 6.6890344636583252e-04
GC_8_362 b_8 NI_8 NS_362 0 -1.0341192240949039e-04
GC_8_363 b_8 NI_8 NS_363 0 -1.8170804303906235e-04
GC_8_364 b_8 NI_8 NS_364 0 -1.1073483359259556e-03
GC_8_365 b_8 NI_8 NS_365 0 1.1320629413702615e-04
GC_8_366 b_8 NI_8 NS_366 0 1.0476172109529106e-04
GC_8_367 b_8 NI_8 NS_367 0 8.3200918954854243e-04
GC_8_368 b_8 NI_8 NS_368 0 1.2040721077215249e-03
GC_8_369 b_8 NI_8 NS_369 0 -1.0147887174600907e-04
GC_8_370 b_8 NI_8 NS_370 0 4.2035797425393133e-05
GC_8_371 b_8 NI_8 NS_371 0 -1.9983718934942028e-04
GC_8_372 b_8 NI_8 NS_372 0 -2.9893821264334980e-05
GC_8_373 b_8 NI_8 NS_373 0 2.2020248797864871e-05
GC_8_374 b_8 NI_8 NS_374 0 5.8965112007747697e-05
GC_8_375 b_8 NI_8 NS_375 0 -1.4937242476196734e-05
GC_8_376 b_8 NI_8 NS_376 0 -8.3901333612622454e-05
GC_8_377 b_8 NI_8 NS_377 0 -4.7296432233853782e-06
GC_8_378 b_8 NI_8 NS_378 0 8.0424174036672932e-05
GC_8_379 b_8 NI_8 NS_379 0 1.0974276174671703e-03
GC_8_380 b_8 NI_8 NS_380 0 1.4494282332578982e-04
GC_8_381 b_8 NI_8 NS_381 0 -1.8372063949728332e-05
GC_8_382 b_8 NI_8 NS_382 0 -2.6850224727397426e-06
GC_8_383 b_8 NI_8 NS_383 0 -3.8023420969606755e-04
GC_8_384 b_8 NI_8 NS_384 0 -2.4029551609091500e-04
GC_8_385 b_8 NI_8 NS_385 0 -8.9435495031103380e-07
GC_8_386 b_8 NI_8 NS_386 0 1.3958817058645732e-06
GC_8_387 b_8 NI_8 NS_387 0 -2.5819851643427248e-06
GC_8_388 b_8 NI_8 NS_388 0 -1.0925382282421013e-05
GC_8_389 b_8 NI_8 NS_389 0 -5.5669719443155555e-06
GC_8_390 b_8 NI_8 NS_390 0 -1.0627986222534553e-05
GC_8_391 b_8 NI_8 NS_391 0 -2.3114210635278910e-07
GC_8_392 b_8 NI_8 NS_392 0 1.5466960949473566e-06
GC_8_393 b_8 NI_8 NS_393 0 -6.4514413684816150e-07
GC_8_394 b_8 NI_8 NS_394 0 -1.2572882377336663e-06
GC_8_395 b_8 NI_8 NS_395 0 -1.5171645924969059e-04
GC_8_396 b_8 NI_8 NS_396 0 -1.4717975322435192e-05
GC_8_397 b_8 NI_8 NS_397 0 -2.3345115047256014e-04
GC_8_398 b_8 NI_8 NS_398 0 -3.2970542038658449e-05
GC_8_399 b_8 NI_8 NS_399 0 8.1136508213380733e-04
GC_8_400 b_8 NI_8 NS_400 0 -5.7431833983557514e-04
GC_8_401 b_8 NI_8 NS_401 0 -2.7931887907723627e-04
GC_8_402 b_8 NI_8 NS_402 0 7.6862165704357649e-04
GC_8_403 b_8 NI_8 NS_403 0 -5.3118289761842582e-04
GC_8_404 b_8 NI_8 NS_404 0 7.8733510748291404e-05
GC_8_405 b_8 NI_8 NS_405 0 1.6731011812601642e-04
GC_8_406 b_8 NI_8 NS_406 0 -1.4298139967554229e-04
GC_8_407 b_8 NI_8 NS_407 0 -1.4733629587225717e-04
GC_8_408 b_8 NI_8 NS_408 0 -1.7551594527536414e-04
GC_8_409 b_8 NI_8 NS_409 0 -9.1393439145907078e-06
GC_8_410 b_8 NI_8 NS_410 0 1.8521895863060328e-05
GC_8_411 b_8 NI_8 NS_411 0 4.6414426212986007e-04
GC_8_412 b_8 NI_8 NS_412 0 -5.5381479116483633e-05
GC_8_413 b_8 NI_8 NS_413 0 1.3031382761236514e-05
GC_8_414 b_8 NI_8 NS_414 0 -4.2861688096145277e-05
GC_8_415 b_8 NI_8 NS_415 0 4.4991053652783695e-04
GC_8_416 b_8 NI_8 NS_416 0 -3.0860129067544111e-04
GC_8_417 b_8 NI_8 NS_417 0 -6.4627580253418735e-05
GC_8_418 b_8 NI_8 NS_418 0 -2.0303595032190226e-04
GC_8_419 b_8 NI_8 NS_419 0 -1.3024353460578898e-07
GC_8_420 b_8 NI_8 NS_420 0 -2.9082176289912082e-05
GC_8_421 b_8 NI_8 NS_421 0 -4.7331757059329788e-05
GC_8_422 b_8 NI_8 NS_422 0 -1.4943585407730322e-04
GC_8_423 b_8 NI_8 NS_423 0 -3.2088715493229884e-03
GC_8_424 b_8 NI_8 NS_424 0 2.9751852937223151e-03
GC_8_425 b_8 NI_8 NS_425 0 6.9811125761412180e-06
GC_8_426 b_8 NI_8 NS_426 0 5.8153286823260506e-06
GC_8_427 b_8 NI_8 NS_427 0 2.7935002120222708e-03
GC_8_428 b_8 NI_8 NS_428 0 -1.0271068467940247e-03
GC_8_429 b_8 NI_8 NS_429 0 1.1192633568573385e-05
GC_8_430 b_8 NI_8 NS_430 0 6.5893740730623478e-06
GC_8_431 b_8 NI_8 NS_431 0 4.5241610782323802e-05
GC_8_432 b_8 NI_8 NS_432 0 -2.7697856887010634e-04
GC_8_433 b_8 NI_8 NS_433 0 -3.4507818243987188e-05
GC_8_434 b_8 NI_8 NS_434 0 1.8608654449272834e-06
GC_8_435 b_8 NI_8 NS_435 0 2.8555673918546639e-05
GC_8_436 b_8 NI_8 NS_436 0 -3.8266426293290861e-06
GC_8_437 b_8 NI_8 NS_437 0 -1.0952885268107529e-05
GC_8_438 b_8 NI_8 NS_438 0 8.9524069303394480e-06
GC_8_439 b_8 NI_8 NS_439 0 3.1196288951872381e-04
GC_8_440 b_8 NI_8 NS_440 0 1.2630031373859661e-04
GC_8_441 b_8 NI_8 NS_441 0 3.6983307980224993e-03
GC_8_442 b_8 NI_8 NS_442 0 3.9376601155199612e-05
GC_8_443 b_8 NI_8 NS_443 0 -1.7988795077153827e-03
GC_8_444 b_8 NI_8 NS_444 0 -1.0939128926076905e-03
GC_8_445 b_8 NI_8 NS_445 0 1.4015306841865822e-03
GC_8_446 b_8 NI_8 NS_446 0 7.0587049622438422e-04
GC_8_447 b_8 NI_8 NS_447 0 -2.2953689107977449e-05
GC_8_448 b_8 NI_8 NS_448 0 1.1614350863459133e-04
GC_8_449 b_8 NI_8 NS_449 0 4.0637789565206074e-04
GC_8_450 b_8 NI_8 NS_450 0 3.1642458149146990e-05
GC_8_451 b_8 NI_8 NS_451 0 6.1325648672609114e-04
GC_8_452 b_8 NI_8 NS_452 0 -1.3287104761042813e-03
GC_8_453 b_8 NI_8 NS_453 0 4.1404832731776599e-05
GC_8_454 b_8 NI_8 NS_454 0 1.2227939958522836e-04
GC_8_455 b_8 NI_8 NS_455 0 5.0954432078513106e-06
GC_8_456 b_8 NI_8 NS_456 0 6.8254233759740095e-04
GC_8_457 b_8 NI_8 NS_457 0 -8.0991991923683664e-05
GC_8_458 b_8 NI_8 NS_458 0 2.6628114778313386e-05
GC_8_459 b_8 NI_8 NS_459 0 -1.9810162686942367e-04
GC_8_460 b_8 NI_8 NS_460 0 2.6959461393542383e-04
GC_8_461 b_8 NI_8 NS_461 0 -5.4364225168979975e-05
GC_8_462 b_8 NI_8 NS_462 0 1.3713015731147633e-04
GC_8_463 b_8 NI_8 NS_463 0 -1.8322208204072464e-05
GC_8_464 b_8 NI_8 NS_464 0 -5.5537144300232469e-05
GC_8_465 b_8 NI_8 NS_465 0 -1.3234449291264797e-05
GC_8_466 b_8 NI_8 NS_466 0 6.2432784437886461e-05
GC_8_467 b_8 NI_8 NS_467 0 2.7168476450573862e-04
GC_8_468 b_8 NI_8 NS_468 0 5.1435504235666622e-04
GC_8_469 b_8 NI_8 NS_469 0 -9.9147809345207669e-06
GC_8_470 b_8 NI_8 NS_470 0 -2.7125789585324150e-06
GC_8_471 b_8 NI_8 NS_471 0 -9.8472937326628601e-05
GC_8_472 b_8 NI_8 NS_472 0 -7.1571949366725041e-05
GC_8_473 b_8 NI_8 NS_473 0 -1.3734911853709993e-06
GC_8_474 b_8 NI_8 NS_474 0 -8.0815576004514630e-07
GC_8_475 b_8 NI_8 NS_475 0 -6.0327746652318092e-05
GC_8_476 b_8 NI_8 NS_476 0 -5.7714251284654566e-05
GC_8_477 b_8 NI_8 NS_477 0 -2.8623358256090717e-06
GC_8_478 b_8 NI_8 NS_478 0 -5.3798795692023060e-06
GC_8_479 b_8 NI_8 NS_479 0 1.3944909274021752e-07
GC_8_480 b_8 NI_8 NS_480 0 -5.4613466000379097e-08
GC_8_481 b_8 NI_8 NS_481 0 -3.7581453636501627e-07
GC_8_482 b_8 NI_8 NS_482 0 -8.1654791595564893e-07
GC_8_483 b_8 NI_8 NS_483 0 -9.0194584966714971e-05
GC_8_484 b_8 NI_8 NS_484 0 -3.6865693235548075e-05
GC_8_485 b_8 NI_8 NS_485 0 -2.0376969200563708e-03
GC_8_486 b_8 NI_8 NS_486 0 -2.6979148551402511e-04
GC_8_487 b_8 NI_8 NS_487 0 9.8746942026919460e-04
GC_8_488 b_8 NI_8 NS_488 0 6.2089334501431526e-04
GC_8_489 b_8 NI_8 NS_489 0 -1.6023503573559992e-03
GC_8_490 b_8 NI_8 NS_490 0 -1.0182016742790909e-03
GC_8_491 b_8 NI_8 NS_491 0 -1.5221769095373708e-04
GC_8_492 b_8 NI_8 NS_492 0 -3.5021747076024247e-04
GC_8_493 b_8 NI_8 NS_493 0 2.7047197216827139e-04
GC_8_494 b_8 NI_8 NS_494 0 -1.3273472072047545e-04
GC_8_495 b_8 NI_8 NS_495 0 1.8394262142209721e-05
GC_8_496 b_8 NI_8 NS_496 0 -7.8835916884693435e-04
GC_8_497 b_8 NI_8 NS_497 0 1.1315950061779080e-06
GC_8_498 b_8 NI_8 NS_498 0 2.5322931789875400e-05
GC_8_499 b_8 NI_8 NS_499 0 1.9640154350910604e-04
GC_8_500 b_8 NI_8 NS_500 0 -3.7604674859442137e-04
GC_8_501 b_8 NI_8 NS_501 0 1.6413426707313411e-05
GC_8_502 b_8 NI_8 NS_502 0 -2.2490592157640993e-05
GC_8_503 b_8 NI_8 NS_503 0 4.6980028007335723e-04
GC_8_504 b_8 NI_8 NS_504 0 -2.8035645500171127e-04
GC_8_505 b_8 NI_8 NS_505 0 -5.2532684295386703e-05
GC_8_506 b_8 NI_8 NS_506 0 -1.2391619075578417e-04
GC_8_507 b_8 NI_8 NS_507 0 1.1188319459244365e-05
GC_8_508 b_8 NI_8 NS_508 0 -1.7939387655076858e-05
GC_8_509 b_8 NI_8 NS_509 0 -2.4806303415376573e-05
GC_8_510 b_8 NI_8 NS_510 0 -1.0140405251345679e-04
GC_8_511 b_8 NI_8 NS_511 0 -1.0091146191824774e-03
GC_8_512 b_8 NI_8 NS_512 0 2.6860199448676572e-03
GC_8_513 b_8 NI_8 NS_513 0 -1.3367844719751132e-06
GC_8_514 b_8 NI_8 NS_514 0 -8.5138660201484172e-07
GC_8_515 b_8 NI_8 NS_515 0 1.7787760505881885e-03
GC_8_516 b_8 NI_8 NS_516 0 -1.0063314776989545e-03
GC_8_517 b_8 NI_8 NS_517 0 3.9880543844080053e-06
GC_8_518 b_8 NI_8 NS_518 0 2.0130104600302771e-06
GC_8_519 b_8 NI_8 NS_519 0 -1.2995156884474643e-04
GC_8_520 b_8 NI_8 NS_520 0 -3.9594108524536858e-06
GC_8_521 b_8 NI_8 NS_521 0 -9.3783845154687570e-06
GC_8_522 b_8 NI_8 NS_522 0 3.0116554135362462e-06
GC_8_523 b_8 NI_8 NS_523 0 1.7798938505784383e-05
GC_8_524 b_8 NI_8 NS_524 0 2.4251323766619211e-07
GC_8_525 b_8 NI_8 NS_525 0 -4.5695707038171263e-06
GC_8_526 b_8 NI_8 NS_526 0 2.4362469575008091e-06
GC_8_527 b_8 NI_8 NS_527 0 1.2410760116051358e-04
GC_8_528 b_8 NI_8 NS_528 0 6.9885891927635820e-05
GD_8_1 b_8 NI_8 NA_1 0 -1.8618147620898955e-02
GD_8_2 b_8 NI_8 NA_2 0 -1.1805446344122346e-02
GD_8_3 b_8 NI_8 NA_3 0 -3.8026279499986590e-02
GD_8_4 b_8 NI_8 NA_4 0 -1.8322305683301718e-02
GD_8_5 b_8 NI_8 NA_5 0 -6.4533380289556311e-02
GD_8_6 b_8 NI_8 NA_6 0 -1.5472297387311994e-02
GD_8_7 b_8 NI_8 NA_7 0 2.2066460413552795e-03
GD_8_8 b_8 NI_8 NA_8 0 2.6570761232874396e-01
GD_8_9 b_8 NI_8 NA_9 0 1.3218788982330152e-03
GD_8_10 b_8 NI_8 NA_10 0 -1.3222267236412642e-03
GD_8_11 b_8 NI_8 NA_11 0 -5.9634419064444862e-03
GD_8_12 b_8 NI_8 NA_12 0 -2.1945666339029030e-04
*
* Port 9
VI_9 a_9 NI_9 0
RI_9 NI_9 b_9 5.0000000000000000e+01
GC_9_1 b_9 NI_9 NS_1 0 1.2161754773099645e-02
GC_9_2 b_9 NI_9 NS_2 0 2.9743901560926960e-05
GC_9_3 b_9 NI_9 NS_3 0 -8.0268601604319568e-05
GC_9_4 b_9 NI_9 NS_4 0 -3.8275723532876533e-04
GC_9_5 b_9 NI_9 NS_5 0 5.0603859991743365e-04
GC_9_6 b_9 NI_9 NS_6 0 -3.1256005231946346e-04
GC_9_7 b_9 NI_9 NS_7 0 -6.7844626111423654e-04
GC_9_8 b_9 NI_9 NS_8 0 -7.6615536918423510e-05
GC_9_9 b_9 NI_9 NS_9 0 8.2391435272929816e-04
GC_9_10 b_9 NI_9 NS_10 0 -3.4301927393391425e-04
GC_9_11 b_9 NI_9 NS_11 0 -3.8630160293515279e-04
GC_9_12 b_9 NI_9 NS_12 0 7.9971579167091968e-05
GC_9_13 b_9 NI_9 NS_13 0 4.1339530172817575e-04
GC_9_14 b_9 NI_9 NS_14 0 -5.0204318453922708e-04
GC_9_15 b_9 NI_9 NS_15 0 4.5638961827993924e-03
GC_9_16 b_9 NI_9 NS_16 0 -3.0340001920336302e-04
GC_9_17 b_9 NI_9 NS_17 0 3.0315089964349032e-04
GC_9_18 b_9 NI_9 NS_18 0 2.6717916448729719e-04
GC_9_19 b_9 NI_9 NS_19 0 -1.1764918185559171e-04
GC_9_20 b_9 NI_9 NS_20 0 2.6577146494903233e-03
GC_9_21 b_9 NI_9 NS_21 0 3.7125976346548932e-04
GC_9_22 b_9 NI_9 NS_22 0 -3.2361049428798077e-04
GC_9_23 b_9 NI_9 NS_23 0 1.2111192952132933e-04
GC_9_24 b_9 NI_9 NS_24 0 -2.2611626583080682e-05
GC_9_25 b_9 NI_9 NS_25 0 2.2635844585305873e-05
GC_9_26 b_9 NI_9 NS_26 0 1.1332281423392591e-04
GC_9_27 b_9 NI_9 NS_27 0 -6.9718390859677386e-03
GC_9_28 b_9 NI_9 NS_28 0 5.8338761726857884e-03
GC_9_29 b_9 NI_9 NS_29 0 1.3223443970424284e-05
GC_9_30 b_9 NI_9 NS_30 0 -1.0943210253097955e-05
GC_9_31 b_9 NI_9 NS_31 0 1.9431588743285713e-03
GC_9_32 b_9 NI_9 NS_32 0 -1.5744097609214557e-04
GC_9_33 b_9 NI_9 NS_33 0 4.6981066944375941e-06
GC_9_34 b_9 NI_9 NS_34 0 8.4502206082711448e-06
GC_9_35 b_9 NI_9 NS_35 0 -3.6496771295242529e-05
GC_9_36 b_9 NI_9 NS_36 0 -2.6828697374069862e-03
GC_9_37 b_9 NI_9 NS_37 0 -2.5651202033223720e-05
GC_9_38 b_9 NI_9 NS_38 0 5.1753396868897984e-06
GC_9_39 b_9 NI_9 NS_39 0 -1.6607257807269245e-06
GC_9_40 b_9 NI_9 NS_40 0 -2.6004079990906647e-06
GC_9_41 b_9 NI_9 NS_41 0 4.4174125239708836e-06
GC_9_42 b_9 NI_9 NS_42 0 1.8743929862647062e-06
GC_9_43 b_9 NI_9 NS_43 0 -5.3721009391869094e-05
GC_9_44 b_9 NI_9 NS_44 0 -6.8479971901771368e-04
GC_9_45 b_9 NI_9 NS_45 0 1.0870601564304205e-02
GC_9_46 b_9 NI_9 NS_46 0 1.2683920773059339e-05
GC_9_47 b_9 NI_9 NS_47 0 5.2885786629354156e-05
GC_9_48 b_9 NI_9 NS_48 0 1.1568908029124325e-04
GC_9_49 b_9 NI_9 NS_49 0 -1.5750037883566239e-04
GC_9_50 b_9 NI_9 NS_50 0 -4.0872092959585028e-05
GC_9_51 b_9 NI_9 NS_51 0 -4.8227685786262660e-04
GC_9_52 b_9 NI_9 NS_52 0 4.6562153026052393e-05
GC_9_53 b_9 NI_9 NS_53 0 1.8156450060677554e-04
GC_9_54 b_9 NI_9 NS_54 0 -2.7879076984154328e-04
GC_9_55 b_9 NI_9 NS_55 0 9.2224055984269960e-04
GC_9_56 b_9 NI_9 NS_56 0 8.0881795329622636e-05
GC_9_57 b_9 NI_9 NS_57 0 8.6181904775834841e-05
GC_9_58 b_9 NI_9 NS_58 0 6.4647132230620245e-05
GC_9_59 b_9 NI_9 NS_59 0 -2.1132938265746600e-04
GC_9_60 b_9 NI_9 NS_60 0 1.6262901390715449e-03
GC_9_61 b_9 NI_9 NS_61 0 -1.3064987932563931e-04
GC_9_62 b_9 NI_9 NS_62 0 6.0058879276137848e-05
GC_9_63 b_9 NI_9 NS_63 0 -5.6746966409917683e-04
GC_9_64 b_9 NI_9 NS_64 0 -1.3590971363418842e-04
GC_9_65 b_9 NI_9 NS_65 0 4.7008698275640580e-06
GC_9_66 b_9 NI_9 NS_66 0 -9.8943493853762034e-05
GC_9_67 b_9 NI_9 NS_67 0 -3.1885075063585268e-05
GC_9_68 b_9 NI_9 NS_68 0 -1.0495393743851835e-04
GC_9_69 b_9 NI_9 NS_69 0 -3.1288021028945983e-06
GC_9_70 b_9 NI_9 NS_70 0 9.4842169187206167e-05
GC_9_71 b_9 NI_9 NS_71 0 6.0029511585859054e-05
GC_9_72 b_9 NI_9 NS_72 0 3.8375889912076969e-04
GC_9_73 b_9 NI_9 NS_73 0 -2.2343874718566364e-05
GC_9_74 b_9 NI_9 NS_74 0 -1.1997769890853945e-05
GC_9_75 b_9 NI_9 NS_75 0 -2.2102137077803388e-04
GC_9_76 b_9 NI_9 NS_76 0 -1.8404117038051118e-04
GC_9_77 b_9 NI_9 NS_77 0 4.5603143395521223e-07
GC_9_78 b_9 NI_9 NS_78 0 2.4999756906066381e-06
GC_9_79 b_9 NI_9 NS_79 0 -6.2589325193952814e-05
GC_9_80 b_9 NI_9 NS_80 0 -2.4324721605504322e-04
GC_9_81 b_9 NI_9 NS_81 0 -1.0946832818994846e-05
GC_9_82 b_9 NI_9 NS_82 0 -1.6208402770865455e-05
GC_9_83 b_9 NI_9 NS_83 0 -2.3535191915758593e-07
GC_9_84 b_9 NI_9 NS_84 0 1.2084763953168231e-06
GC_9_85 b_9 NI_9 NS_85 0 -4.9809921916408984e-07
GC_9_86 b_9 NI_9 NS_86 0 -1.3863858263100164e-06
GC_9_87 b_9 NI_9 NS_87 0 -2.1116633731439128e-04
GC_9_88 b_9 NI_9 NS_88 0 -4.4890192160091162e-05
GC_9_89 b_9 NI_9 NS_89 0 6.6558836823774614e-03
GC_9_90 b_9 NI_9 NS_90 0 7.2037377053766778e-05
GC_9_91 b_9 NI_9 NS_91 0 7.7325136216140475e-06
GC_9_92 b_9 NI_9 NS_92 0 -7.3280918763234289e-04
GC_9_93 b_9 NI_9 NS_93 0 7.9624033450338314e-04
GC_9_94 b_9 NI_9 NS_94 0 -3.2506063197561269e-04
GC_9_95 b_9 NI_9 NS_95 0 -1.1197732187520468e-03
GC_9_96 b_9 NI_9 NS_96 0 1.8635816200616716e-04
GC_9_97 b_9 NI_9 NS_97 0 1.1683215654314540e-03
GC_9_98 b_9 NI_9 NS_98 0 -3.2146532527721093e-04
GC_9_99 b_9 NI_9 NS_99 0 -1.7507408033464406e-03
GC_9_100 b_9 NI_9 NS_100 0 -2.5742536920201546e-04
GC_9_101 b_9 NI_9 NS_101 0 5.7845458146642975e-04
GC_9_102 b_9 NI_9 NS_102 0 -6.8230827729747531e-04
GC_9_103 b_9 NI_9 NS_103 0 7.2709872965402858e-03
GC_9_104 b_9 NI_9 NS_104 0 -1.6936100436079401e-03
GC_9_105 b_9 NI_9 NS_105 0 4.0505317000387079e-04
GC_9_106 b_9 NI_9 NS_106 0 3.9573834929403833e-04
GC_9_107 b_9 NI_9 NS_107 0 -1.6840727706978641e-05
GC_9_108 b_9 NI_9 NS_108 0 3.4144445070573982e-03
GC_9_109 b_9 NI_9 NS_109 0 4.6607954031386900e-04
GC_9_110 b_9 NI_9 NS_110 0 -3.4889675089399695e-04
GC_9_111 b_9 NI_9 NS_111 0 2.0083092384290518e-04
GC_9_112 b_9 NI_9 NS_112 0 -7.4041779309955765e-05
GC_9_113 b_9 NI_9 NS_113 0 3.7699005103411359e-05
GC_9_114 b_9 NI_9 NS_114 0 1.3194479967360527e-04
GC_9_115 b_9 NI_9 NS_115 0 -7.2294081533616538e-03
GC_9_116 b_9 NI_9 NS_116 0 8.8351753128317716e-03
GC_9_117 b_9 NI_9 NS_117 0 9.4168030262795573e-06
GC_9_118 b_9 NI_9 NS_118 0 -1.8238204868149572e-05
GC_9_119 b_9 NI_9 NS_119 0 2.3124639190924426e-03
GC_9_120 b_9 NI_9 NS_120 0 -1.0858815281433766e-03
GC_9_121 b_9 NI_9 NS_121 0 -2.2710860775659603e-06
GC_9_122 b_9 NI_9 NS_122 0 6.2393270376437589e-06
GC_9_123 b_9 NI_9 NS_123 0 -2.9346244144622325e-04
GC_9_124 b_9 NI_9 NS_124 0 -2.7375782709969823e-03
GC_9_125 b_9 NI_9 NS_125 0 -2.3823606196989841e-05
GC_9_126 b_9 NI_9 NS_126 0 7.0564506394605772e-07
GC_9_127 b_9 NI_9 NS_127 0 -4.5845482435394924e-07
GC_9_128 b_9 NI_9 NS_128 0 -2.3108276892485427e-06
GC_9_129 b_9 NI_9 NS_129 0 2.5409493165338796e-06
GC_9_130 b_9 NI_9 NS_130 0 3.3613287519374331e-06
GC_9_131 b_9 NI_9 NS_131 0 -1.1195898938226832e-04
GC_9_132 b_9 NI_9 NS_132 0 -8.4306666866020648e-04
GC_9_133 b_9 NI_9 NS_133 0 8.5315067141513087e-03
GC_9_134 b_9 NI_9 NS_134 0 1.0772723631049934e-05
GC_9_135 b_9 NI_9 NS_135 0 -8.2028579496581453e-05
GC_9_136 b_9 NI_9 NS_136 0 2.8470289857292973e-04
GC_9_137 b_9 NI_9 NS_137 0 -3.1093127015946248e-04
GC_9_138 b_9 NI_9 NS_138 0 -3.0657286206216012e-04
GC_9_139 b_9 NI_9 NS_139 0 -3.3410662526607256e-04
GC_9_140 b_9 NI_9 NS_140 0 1.0880594062745147e-04
GC_9_141 b_9 NI_9 NS_141 0 3.0336050826921320e-04
GC_9_142 b_9 NI_9 NS_142 0 -4.1443568322086123e-04
GC_9_143 b_9 NI_9 NS_143 0 7.1085970425959974e-04
GC_9_144 b_9 NI_9 NS_144 0 -1.4210419379702384e-05
GC_9_145 b_9 NI_9 NS_145 0 1.1796089933875008e-04
GC_9_146 b_9 NI_9 NS_146 0 1.2662332073008390e-04
GC_9_147 b_9 NI_9 NS_147 0 -1.8339202834380932e-05
GC_9_148 b_9 NI_9 NS_148 0 1.4343089141500964e-03
GC_9_149 b_9 NI_9 NS_149 0 -1.4176996573033525e-04
GC_9_150 b_9 NI_9 NS_150 0 6.8389848462040222e-05
GC_9_151 b_9 NI_9 NS_151 0 -6.2914179994444386e-04
GC_9_152 b_9 NI_9 NS_152 0 -1.4961658139380450e-04
GC_9_153 b_9 NI_9 NS_153 0 -1.2871117239019329e-05
GC_9_154 b_9 NI_9 NS_154 0 -4.7807578019794360e-05
GC_9_155 b_9 NI_9 NS_155 0 -3.0255667207690058e-05
GC_9_156 b_9 NI_9 NS_156 0 -1.2353373532478953e-04
GC_9_157 b_9 NI_9 NS_157 0 -3.2600878545211723e-06
GC_9_158 b_9 NI_9 NS_158 0 9.9802305102526689e-05
GC_9_159 b_9 NI_9 NS_159 0 6.6929850026039358e-04
GC_9_160 b_9 NI_9 NS_160 0 3.5611076636833232e-04
GC_9_161 b_9 NI_9 NS_161 0 -2.6654133857284736e-05
GC_9_162 b_9 NI_9 NS_162 0 -1.1439792006077319e-05
GC_9_163 b_9 NI_9 NS_163 0 -3.8522597237421890e-04
GC_9_164 b_9 NI_9 NS_164 0 -3.6760188209892028e-04
GC_9_165 b_9 NI_9 NS_165 0 3.9498715625751564e-09
GC_9_166 b_9 NI_9 NS_166 0 1.6529104084264056e-06
GC_9_167 b_9 NI_9 NS_167 0 -1.3698592797299191e-04
GC_9_168 b_9 NI_9 NS_168 0 -1.4723215151569771e-04
GC_9_169 b_9 NI_9 NS_169 0 -8.5640418514025532e-06
GC_9_170 b_9 NI_9 NS_170 0 -1.4077661444153333e-05
GC_9_171 b_9 NI_9 NS_171 0 -1.9766256345940988e-07
GC_9_172 b_9 NI_9 NS_172 0 1.2404380986910700e-06
GC_9_173 b_9 NI_9 NS_173 0 -8.8913539306545071e-07
GC_9_174 b_9 NI_9 NS_174 0 -1.4725025387726742e-06
GC_9_175 b_9 NI_9 NS_175 0 -2.1057908719550008e-04
GC_9_176 b_9 NI_9 NS_176 0 -2.6955568122266091e-05
GC_9_177 b_9 NI_9 NS_177 0 2.4139312681306412e-03
GC_9_178 b_9 NI_9 NS_178 0 9.6680950485263713e-05
GC_9_179 b_9 NI_9 NS_179 0 3.1994561853024327e-04
GC_9_180 b_9 NI_9 NS_180 0 -8.7100380896955657e-04
GC_9_181 b_9 NI_9 NS_181 0 7.1087236296235579e-04
GC_9_182 b_9 NI_9 NS_182 0 1.4391781251235134e-05
GC_9_183 b_9 NI_9 NS_183 0 -7.3534902540049382e-04
GC_9_184 b_9 NI_9 NS_184 0 -1.4673971971647986e-04
GC_9_185 b_9 NI_9 NS_185 0 1.0990118954392388e-03
GC_9_186 b_9 NI_9 NS_186 0 -3.1185214893761647e-05
GC_9_187 b_9 NI_9 NS_187 0 -2.7438275142306731e-03
GC_9_188 b_9 NI_9 NS_188 0 -1.1079316846233091e-03
GC_9_189 b_9 NI_9 NS_189 0 5.9680753538759145e-04
GC_9_190 b_9 NI_9 NS_190 0 -6.5920999095400842e-04
GC_9_191 b_9 NI_9 NS_191 0 8.5310220433288137e-03
GC_9_192 b_9 NI_9 NS_192 0 -1.5952180220836934e-03
GC_9_193 b_9 NI_9 NS_193 0 4.2746865751006530e-04
GC_9_194 b_9 NI_9 NS_194 0 3.7746972261309936e-04
GC_9_195 b_9 NI_9 NS_195 0 2.6330902543408679e-04
GC_9_196 b_9 NI_9 NS_196 0 3.6143004477540994e-03
GC_9_197 b_9 NI_9 NS_197 0 6.5053959463734837e-04
GC_9_198 b_9 NI_9 NS_198 0 -2.3888047967161709e-04
GC_9_199 b_9 NI_9 NS_199 0 2.1942958590614024e-04
GC_9_200 b_9 NI_9 NS_200 0 -3.3735988993723581e-05
GC_9_201 b_9 NI_9 NS_201 0 3.3614712090549626e-05
GC_9_202 b_9 NI_9 NS_202 0 1.2776920490539963e-04
GC_9_203 b_9 NI_9 NS_203 0 -8.7398808229486279e-03
GC_9_204 b_9 NI_9 NS_204 0 8.3619022200682996e-03
GC_9_205 b_9 NI_9 NS_205 0 1.8693432767334181e-05
GC_9_206 b_9 NI_9 NS_206 0 -2.0149242821608713e-05
GC_9_207 b_9 NI_9 NS_207 0 2.5892110783086735e-03
GC_9_208 b_9 NI_9 NS_208 0 -6.9767556827055055e-04
GC_9_209 b_9 NI_9 NS_209 0 -3.4587537152880438e-07
GC_9_210 b_9 NI_9 NS_210 0 8.7176429309332658e-06
GC_9_211 b_9 NI_9 NS_211 0 -1.3654485377959314e-04
GC_9_212 b_9 NI_9 NS_212 0 -2.7337224859746889e-03
GC_9_213 b_9 NI_9 NS_213 0 -2.0591606492199513e-05
GC_9_214 b_9 NI_9 NS_214 0 -1.6458114482527407e-06
GC_9_215 b_9 NI_9 NS_215 0 2.4308058035740027e-07
GC_9_216 b_9 NI_9 NS_216 0 -2.1701123788410292e-06
GC_9_217 b_9 NI_9 NS_217 0 3.0566742254987261e-06
GC_9_218 b_9 NI_9 NS_218 0 3.7661484470120329e-06
GC_9_219 b_9 NI_9 NS_219 0 -5.1317205510064739e-05
GC_9_220 b_9 NI_9 NS_220 0 -9.0248529433808046e-04
GC_9_221 b_9 NI_9 NS_221 0 1.4261314005657637e-03
GC_9_222 b_9 NI_9 NS_222 0 -6.7033252988336709e-06
GC_9_223 b_9 NI_9 NS_223 0 -4.0969191185085427e-04
GC_9_224 b_9 NI_9 NS_224 0 4.6129996940063174e-04
GC_9_225 b_9 NI_9 NS_225 0 -3.7193509192184974e-04
GC_9_226 b_9 NI_9 NS_226 0 -7.2968885138887188e-04
GC_9_227 b_9 NI_9 NS_227 0 -3.0997807785260422e-05
GC_9_228 b_9 NI_9 NS_228 0 2.8271282100559176e-04
GC_9_229 b_9 NI_9 NS_229 0 3.7364201469781581e-04
GC_9_230 b_9 NI_9 NS_230 0 -4.5726431905588624e-04
GC_9_231 b_9 NI_9 NS_231 0 -1.3928557296147105e-04
GC_9_232 b_9 NI_9 NS_232 0 -4.0307293931965968e-04
GC_9_233 b_9 NI_9 NS_233 0 1.4612912619615845e-04
GC_9_234 b_9 NI_9 NS_234 0 9.8407616566267614e-05
GC_9_235 b_9 NI_9 NS_235 0 7.3128165219896548e-04
GC_9_236 b_9 NI_9 NS_236 0 7.1015589107148230e-04
GC_9_237 b_9 NI_9 NS_237 0 -1.7533806806115589e-04
GC_9_238 b_9 NI_9 NS_238 0 8.7703986868127226e-05
GC_9_239 b_9 NI_9 NS_239 0 -5.5700440718160359e-04
GC_9_240 b_9 NI_9 NS_240 0 -3.1092007885116048e-04
GC_9_241 b_9 NI_9 NS_241 0 -4.0364246150819856e-05
GC_9_242 b_9 NI_9 NS_242 0 -5.7661528876527086e-07
GC_9_243 b_9 NI_9 NS_243 0 -2.6374630329052356e-05
GC_9_244 b_9 NI_9 NS_244 0 -1.6347356146842316e-04
GC_9_245 b_9 NI_9 NS_245 0 -7.2801185992670951e-07
GC_9_246 b_9 NI_9 NS_246 0 1.3419482376026169e-04
GC_9_247 b_9 NI_9 NS_247 0 2.0646318579023953e-03
GC_9_248 b_9 NI_9 NS_248 0 1.0799052117643399e-03
GC_9_249 b_9 NI_9 NS_249 0 -3.5532406588555106e-05
GC_9_250 b_9 NI_9 NS_250 0 -1.4195518965058892e-05
GC_9_251 b_9 NI_9 NS_251 0 -5.4147212520699558e-04
GC_9_252 b_9 NI_9 NS_252 0 -8.3310959636911962e-04
GC_9_253 b_9 NI_9 NS_253 0 -6.7268862415105981e-07
GC_9_254 b_9 NI_9 NS_254 0 2.0299725600112224e-06
GC_9_255 b_9 NI_9 NS_255 0 -2.8595469567507760e-04
GC_9_256 b_9 NI_9 NS_256 0 -1.3148419599512718e-04
GC_9_257 b_9 NI_9 NS_257 0 -1.3820329668716023e-05
GC_9_258 b_9 NI_9 NS_258 0 -2.1115572383413484e-05
GC_9_259 b_9 NI_9 NS_259 0 -4.4101160994088077e-07
GC_9_260 b_9 NI_9 NS_260 0 3.2097387339354278e-06
GC_9_261 b_9 NI_9 NS_261 0 -2.0199105060333220e-06
GC_9_262 b_9 NI_9 NS_262 0 -3.4269797520560149e-06
GC_9_263 b_9 NI_9 NS_263 0 -3.7162045616204620e-04
GC_9_264 b_9 NI_9 NS_264 0 -2.5400512127395654e-05
GC_9_265 b_9 NI_9 NS_265 0 3.5834678516367372e-03
GC_9_266 b_9 NI_9 NS_266 0 8.0313721371873357e-05
GC_9_267 b_9 NI_9 NS_267 0 1.2125857014380378e-03
GC_9_268 b_9 NI_9 NS_268 0 -2.7628360312396554e-04
GC_9_269 b_9 NI_9 NS_269 0 -6.4692423471594406e-04
GC_9_270 b_9 NI_9 NS_270 0 4.4659637772397688e-04
GC_9_271 b_9 NI_9 NS_271 0 2.1428901978077971e-04
GC_9_272 b_9 NI_9 NS_272 0 -2.5603165580087784e-04
GC_9_273 b_9 NI_9 NS_273 0 8.2635413568686762e-04
GC_9_274 b_9 NI_9 NS_274 0 6.1218140991048376e-04
GC_9_275 b_9 NI_9 NS_275 0 -2.6080396907278850e-03
GC_9_276 b_9 NI_9 NS_276 0 -1.5666489054400733e-03
GC_9_277 b_9 NI_9 NS_277 0 5.5976536102930394e-04
GC_9_278 b_9 NI_9 NS_278 0 -4.2694680618903983e-04
GC_9_279 b_9 NI_9 NS_279 0 4.7026602461107559e-03
GC_9_280 b_9 NI_9 NS_280 0 2.6472777822684785e-04
GC_9_281 b_9 NI_9 NS_281 0 2.5844773429946322e-04
GC_9_282 b_9 NI_9 NS_282 0 2.9271130743222434e-04
GC_9_283 b_9 NI_9 NS_283 0 -2.8765856142495740e-04
GC_9_284 b_9 NI_9 NS_284 0 2.0760526355052978e-03
GC_9_285 b_9 NI_9 NS_285 0 3.8090031708854210e-04
GC_9_286 b_9 NI_9 NS_286 0 -2.4005240874845643e-04
GC_9_287 b_9 NI_9 NS_287 0 1.5716287449452776e-04
GC_9_288 b_9 NI_9 NS_288 0 -3.5218565518884665e-05
GC_9_289 b_9 NI_9 NS_289 0 2.0202027053361928e-05
GC_9_290 b_9 NI_9 NS_290 0 8.2366507968036290e-05
GC_9_291 b_9 NI_9 NS_291 0 -5.3580682663034633e-03
GC_9_292 b_9 NI_9 NS_292 0 3.7167113725431245e-03
GC_9_293 b_9 NI_9 NS_293 0 7.9503335376660228e-06
GC_9_294 b_9 NI_9 NS_294 0 -7.0044734455260419e-06
GC_9_295 b_9 NI_9 NS_295 0 1.3621321752628681e-03
GC_9_296 b_9 NI_9 NS_296 0 -5.3201538385273274e-04
GC_9_297 b_9 NI_9 NS_297 0 -9.0546419405520450e-07
GC_9_298 b_9 NI_9 NS_298 0 4.3015069188338549e-06
GC_9_299 b_9 NI_9 NS_299 0 7.7188888867490361e-05
GC_9_300 b_9 NI_9 NS_300 0 -1.8474386959577984e-03
GC_9_301 b_9 NI_9 NS_301 0 -1.4193057447242855e-05
GC_9_302 b_9 NI_9 NS_302 0 4.7812196325175680e-07
GC_9_303 b_9 NI_9 NS_303 0 9.7442154900942755e-07
GC_9_304 b_9 NI_9 NS_304 0 -5.4921797296610507e-07
GC_9_305 b_9 NI_9 NS_305 0 1.0258930372469946e-06
GC_9_306 b_9 NI_9 NS_306 0 3.0913345034165156e-06
GC_9_307 b_9 NI_9 NS_307 0 6.4165385727105785e-06
GC_9_308 b_9 NI_9 NS_308 0 -5.4179235904114743e-04
GC_9_309 b_9 NI_9 NS_309 0 -3.3596046330365754e-03
GC_9_310 b_9 NI_9 NS_310 0 -1.5357282876484801e-05
GC_9_311 b_9 NI_9 NS_311 0 -1.2853688887160793e-03
GC_9_312 b_9 NI_9 NS_312 0 1.9144836471412502e-04
GC_9_313 b_9 NI_9 NS_313 0 6.4740289866826561e-04
GC_9_314 b_9 NI_9 NS_314 0 -1.1924884174498852e-03
GC_9_315 b_9 NI_9 NS_315 0 4.2127835191561179e-05
GC_9_316 b_9 NI_9 NS_316 0 3.5526847929452209e-04
GC_9_317 b_9 NI_9 NS_317 0 6.6890344637202158e-04
GC_9_318 b_9 NI_9 NS_318 0 -1.0341192243477801e-04
GC_9_319 b_9 NI_9 NS_319 0 -1.8170804311608320e-04
GC_9_320 b_9 NI_9 NS_320 0 -1.1073483359935017e-03
GC_9_321 b_9 NI_9 NS_321 0 1.1320629414164313e-04
GC_9_322 b_9 NI_9 NS_322 0 1.0476172108883145e-04
GC_9_323 b_9 NI_9 NS_323 0 8.3200918956199672e-04
GC_9_324 b_9 NI_9 NS_324 0 1.2040721075074949e-03
GC_9_325 b_9 NI_9 NS_325 0 -1.0147887174316338e-04
GC_9_326 b_9 NI_9 NS_326 0 4.2035797423002684e-05
GC_9_327 b_9 NI_9 NS_327 0 -1.9983718932669025e-04
GC_9_328 b_9 NI_9 NS_328 0 -2.9893821359294221e-05
GC_9_329 b_9 NI_9 NS_329 0 2.2020248785983658e-05
GC_9_330 b_9 NI_9 NS_330 0 5.8965112076539864e-05
GC_9_331 b_9 NI_9 NS_331 0 -1.4937242473338253e-05
GC_9_332 b_9 NI_9 NS_332 0 -8.3901333616260250e-05
GC_9_333 b_9 NI_9 NS_333 0 -4.7296432253495857e-06
GC_9_334 b_9 NI_9 NS_334 0 8.0424174034312583e-05
GC_9_335 b_9 NI_9 NS_335 0 1.0974276182127919e-03
GC_9_336 b_9 NI_9 NS_336 0 1.4494282324601916e-04
GC_9_337 b_9 NI_9 NS_337 0 -1.8372063950990509e-05
GC_9_338 b_9 NI_9 NS_338 0 -2.6850224722801285e-06
GC_9_339 b_9 NI_9 NS_339 0 -3.8023420985216361e-04
GC_9_340 b_9 NI_9 NS_340 0 -2.4029551623610011e-04
GC_9_341 b_9 NI_9 NS_341 0 -8.9435495160535128e-07
GC_9_342 b_9 NI_9 NS_342 0 1.3958817058058782e-06
GC_9_343 b_9 NI_9 NS_343 0 -2.5819851275692963e-06
GC_9_344 b_9 NI_9 NS_344 0 -1.0925382112013293e-05
GC_9_345 b_9 NI_9 NS_345 0 -5.5669719427201816e-06
GC_9_346 b_9 NI_9 NS_346 0 -1.0627986223883534e-05
GC_9_347 b_9 NI_9 NS_347 0 -2.3114210621941944e-07
GC_9_348 b_9 NI_9 NS_348 0 1.5466960953935360e-06
GC_9_349 b_9 NI_9 NS_349 0 -6.4514413740663690e-07
GC_9_350 b_9 NI_9 NS_350 0 -1.2572882375781853e-06
GC_9_351 b_9 NI_9 NS_351 0 -1.5171645925483252e-04
GC_9_352 b_9 NI_9 NS_352 0 -1.4717975297335839e-05
GC_9_353 b_9 NI_9 NS_353 0 -5.0986361188087970e-02
GC_9_354 b_9 NI_9 NS_354 0 9.8082259587425960e-03
GC_9_355 b_9 NI_9 NS_355 0 7.9168814016099230e-03
GC_9_356 b_9 NI_9 NS_356 0 5.0389555984185165e-03
GC_9_357 b_9 NI_9 NS_357 0 9.4829047764393194e-03
GC_9_358 b_9 NI_9 NS_358 0 1.9785524727485479e-03
GC_9_359 b_9 NI_9 NS_359 0 -6.0007190672912861e-04
GC_9_360 b_9 NI_9 NS_360 0 7.8263633744156641e-04
GC_9_361 b_9 NI_9 NS_361 0 1.5437764904947030e-03
GC_9_362 b_9 NI_9 NS_362 0 7.4012733849043739e-03
GC_9_363 b_9 NI_9 NS_363 0 -6.0620505266434834e-03
GC_9_364 b_9 NI_9 NS_364 0 2.6382358250863377e-04
GC_9_365 b_9 NI_9 NS_365 0 1.2329501210911844e-03
GC_9_366 b_9 NI_9 NS_366 0 4.2810565178545500e-04
GC_9_367 b_9 NI_9 NS_367 0 6.3440656110471116e-03
GC_9_368 b_9 NI_9 NS_368 0 9.4522862418090683e-04
GC_9_369 b_9 NI_9 NS_369 0 -1.7350750785645542e-05
GC_9_370 b_9 NI_9 NS_370 0 2.5749619088246230e-04
GC_9_371 b_9 NI_9 NS_371 0 -1.0055108721650804e-03
GC_9_372 b_9 NI_9 NS_372 0 -4.5230088600222412e-03
GC_9_373 b_9 NI_9 NS_373 0 -2.0191780150629729e-03
GC_9_374 b_9 NI_9 NS_374 0 5.9249302140784808e-04
GC_9_375 b_9 NI_9 NS_375 0 3.4441612341796270e-04
GC_9_376 b_9 NI_9 NS_376 0 -4.9308068080902694e-05
GC_9_377 b_9 NI_9 NS_377 0 6.1177253401625150e-05
GC_9_378 b_9 NI_9 NS_378 0 -1.8446806183367872e-04
GC_9_379 b_9 NI_9 NS_379 0 9.3450561577715623e-03
GC_9_380 b_9 NI_9 NS_380 0 1.8620811597075820e-02
GC_9_381 b_9 NI_9 NS_381 0 -3.7034328142528691e-05
GC_9_382 b_9 NI_9 NS_382 0 -3.5656298377191646e-05
GC_9_383 b_9 NI_9 NS_383 0 3.3466507888062643e-03
GC_9_384 b_9 NI_9 NS_384 0 -8.3994019331495081e-03
GC_9_385 b_9 NI_9 NS_385 0 8.8505617125210881e-07
GC_9_386 b_9 NI_9 NS_386 0 -4.7891736177095839e-05
GC_9_387 b_9 NI_9 NS_387 0 -3.1578015545850905e-03
GC_9_388 b_9 NI_9 NS_388 0 2.2820894111749796e-03
GC_9_389 b_9 NI_9 NS_389 0 4.8782950964600653e-05
GC_9_390 b_9 NI_9 NS_390 0 5.5323618325058681e-05
GC_9_391 b_9 NI_9 NS_391 0 -1.0339004954193335e-05
GC_9_392 b_9 NI_9 NS_392 0 1.2644204611104499e-05
GC_9_393 b_9 NI_9 NS_393 0 -5.2829366108426465e-06
GC_9_394 b_9 NI_9 NS_394 0 -2.0865007676213934e-05
GC_9_395 b_9 NI_9 NS_395 0 -6.0270757932994335e-04
GC_9_396 b_9 NI_9 NS_396 0 3.6077027959281097e-05
GC_9_397 b_9 NI_9 NS_397 0 5.5079885173182068e-02
GC_9_398 b_9 NI_9 NS_398 0 1.0249097508341872e-02
GC_9_399 b_9 NI_9 NS_399 0 -1.0900785196341170e-02
GC_9_400 b_9 NI_9 NS_400 0 -2.8075048843151404e-03
GC_9_401 b_9 NI_9 NS_401 0 -1.1111934901381208e-02
GC_9_402 b_9 NI_9 NS_402 0 -2.0162350986878000e-03
GC_9_403 b_9 NI_9 NS_403 0 3.4216451652439227e-04
GC_9_404 b_9 NI_9 NS_404 0 1.7538471465930900e-04
GC_9_405 b_9 NI_9 NS_405 0 2.8570119427276529e-03
GC_9_406 b_9 NI_9 NS_406 0 2.5669763841477569e-03
GC_9_407 b_9 NI_9 NS_407 0 -7.1641143582970481e-04
GC_9_408 b_9 NI_9 NS_408 0 -3.7785910780989320e-04
GC_9_409 b_9 NI_9 NS_409 0 -3.2407103709410412e-06
GC_9_410 b_9 NI_9 NS_410 0 1.6235831739973056e-04
GC_9_411 b_9 NI_9 NS_411 0 2.1652453145106689e-03
GC_9_412 b_9 NI_9 NS_412 0 -9.3477382890688537e-04
GC_9_413 b_9 NI_9 NS_413 0 -7.9759638715941404e-05
GC_9_414 b_9 NI_9 NS_414 0 -7.8221968491712252e-05
GC_9_415 b_9 NI_9 NS_415 0 2.2662088453650472e-04
GC_9_416 b_9 NI_9 NS_416 0 7.5012201212576663e-04
GC_9_417 b_9 NI_9 NS_417 0 4.5585921897400036e-04
GC_9_418 b_9 NI_9 NS_418 0 9.5807685428941926e-06
GC_9_419 b_9 NI_9 NS_419 0 -1.1372072976730736e-05
GC_9_420 b_9 NI_9 NS_420 0 -7.2075787769774316e-05
GC_9_421 b_9 NI_9 NS_421 0 -6.4692380210474659e-05
GC_9_422 b_9 NI_9 NS_422 0 1.0151464244118120e-04
GC_9_423 b_9 NI_9 NS_423 0 -3.7213129836945898e-03
GC_9_424 b_9 NI_9 NS_424 0 -6.3818399000517730e-03
GC_9_425 b_9 NI_9 NS_425 0 1.9441165279835976e-05
GC_9_426 b_9 NI_9 NS_426 0 5.0541321237142331e-05
GC_9_427 b_9 NI_9 NS_427 0 -1.0614296185994989e-03
GC_9_428 b_9 NI_9 NS_428 0 2.9857789214100105e-03
GC_9_429 b_9 NI_9 NS_429 0 -3.5376691686443600e-06
GC_9_430 b_9 NI_9 NS_430 0 1.0088123398121202e-05
GC_9_431 b_9 NI_9 NS_431 0 1.2771011861475445e-03
GC_9_432 b_9 NI_9 NS_432 0 -6.9238023682800592e-04
GC_9_433 b_9 NI_9 NS_433 0 -1.0835274676604775e-05
GC_9_434 b_9 NI_9 NS_434 0 -1.1871256966619453e-05
GC_9_435 b_9 NI_9 NS_435 0 3.1750992784676096e-06
GC_9_436 b_9 NI_9 NS_436 0 1.5686657785292131e-07
GC_9_437 b_9 NI_9 NS_437 0 4.0891112544934762e-06
GC_9_438 b_9 NI_9 NS_438 0 2.5456789688210091e-06
GC_9_439 b_9 NI_9 NS_439 0 1.5524175379744170e-04
GC_9_440 b_9 NI_9 NS_440 0 -2.0845533502672991e-04
GC_9_441 b_9 NI_9 NS_441 0 -7.1368608610331060e-03
GC_9_442 b_9 NI_9 NS_442 0 1.6911409837844351e-05
GC_9_443 b_9 NI_9 NS_443 0 4.9589846136580112e-03
GC_9_444 b_9 NI_9 NS_444 0 4.3009851005016272e-03
GC_9_445 b_9 NI_9 NS_445 0 -4.8726242306803480e-03
GC_9_446 b_9 NI_9 NS_446 0 -5.0308499535408986e-03
GC_9_447 b_9 NI_9 NS_447 0 -6.8510161916888481e-04
GC_9_448 b_9 NI_9 NS_448 0 6.7883526952786197e-04
GC_9_449 b_9 NI_9 NS_449 0 1.7789404043728079e-03
GC_9_450 b_9 NI_9 NS_450 0 5.1569106671690021e-03
GC_9_451 b_9 NI_9 NS_451 0 -3.0496667159804021e-03
GC_9_452 b_9 NI_9 NS_452 0 -1.5564734572627950e-03
GC_9_453 b_9 NI_9 NS_453 0 9.8324904594770512e-04
GC_9_454 b_9 NI_9 NS_454 0 1.8005064269863152e-04
GC_9_455 b_9 NI_9 NS_455 0 -3.3298236192449006e-03
GC_9_456 b_9 NI_9 NS_456 0 -3.0004590503739416e-03
GC_9_457 b_9 NI_9 NS_457 0 -4.5982348547055682e-06
GC_9_458 b_9 NI_9 NS_458 0 1.6643701797551590e-04
GC_9_459 b_9 NI_9 NS_459 0 -1.7248145320885046e-03
GC_9_460 b_9 NI_9 NS_460 0 -2.5695238669702879e-03
GC_9_461 b_9 NI_9 NS_461 0 -4.3288848925954925e-04
GC_9_462 b_9 NI_9 NS_462 0 4.1891790230309903e-04
GC_9_463 b_9 NI_9 NS_463 0 2.1078437320663220e-04
GC_9_464 b_9 NI_9 NS_464 0 -7.3375779825501057e-05
GC_9_465 b_9 NI_9 NS_465 0 1.7773460080877991e-05
GC_9_466 b_9 NI_9 NS_466 0 -8.9595572023375145e-05
GC_9_467 b_9 NI_9 NS_467 0 7.9792399367571657e-03
GC_9_468 b_9 NI_9 NS_468 0 4.4950600667203943e-03
GC_9_469 b_9 NI_9 NS_469 0 -1.6110559709327304e-05
GC_9_470 b_9 NI_9 NS_470 0 -1.3105727796451883e-05
GC_9_471 b_9 NI_9 NS_471 0 8.6073305163032363e-04
GC_9_472 b_9 NI_9 NS_472 0 -4.2071176952506026e-03
GC_9_473 b_9 NI_9 NS_473 0 -2.3354229611255937e-06
GC_9_474 b_9 NI_9 NS_474 0 -1.6822606718590027e-05
GC_9_475 b_9 NI_9 NS_475 0 3.4135262751364755e-04
GC_9_476 b_9 NI_9 NS_476 0 1.2274243237997235e-03
GC_9_477 b_9 NI_9 NS_477 0 2.1127925244962802e-05
GC_9_478 b_9 NI_9 NS_478 0 1.1437367675874946e-05
GC_9_479 b_9 NI_9 NS_479 0 -5.2955422678998639e-07
GC_9_480 b_9 NI_9 NS_480 0 6.3789583716281013e-06
GC_9_481 b_9 NI_9 NS_481 0 -3.5556222103933835e-06
GC_9_482 b_9 NI_9 NS_482 0 -3.5517433913476649e-06
GC_9_483 b_9 NI_9 NS_483 0 -8.3306625096499890e-05
GC_9_484 b_9 NI_9 NS_484 0 1.0471443468128497e-04
GC_9_485 b_9 NI_9 NS_485 0 6.2350542204722373e-02
GC_9_486 b_9 NI_9 NS_486 0 -7.6655238724899512e-05
GC_9_487 b_9 NI_9 NS_487 0 -6.3061911194348145e-03
GC_9_488 b_9 NI_9 NS_488 0 -2.5760123202549176e-03
GC_9_489 b_9 NI_9 NS_489 0 4.1561119706079765e-03
GC_9_490 b_9 NI_9 NS_490 0 2.6622431684155934e-03
GC_9_491 b_9 NI_9 NS_491 0 1.8528782169450468e-05
GC_9_492 b_9 NI_9 NS_492 0 1.7264093034512670e-05
GC_9_493 b_9 NI_9 NS_493 0 1.3250795596053181e-03
GC_9_494 b_9 NI_9 NS_494 0 1.5410622118971747e-03
GC_9_495 b_9 NI_9 NS_495 0 -3.0663438042944605e-04
GC_9_496 b_9 NI_9 NS_496 0 -3.0277794366041707e-04
GC_9_497 b_9 NI_9 NS_497 0 -6.5925268971414209e-05
GC_9_498 b_9 NI_9 NS_498 0 7.1505999992965509e-05
GC_9_499 b_9 NI_9 NS_499 0 -4.4716097058221001e-03
GC_9_500 b_9 NI_9 NS_500 0 9.1005488819941179e-04
GC_9_501 b_9 NI_9 NS_501 0 -8.4331119162080027e-05
GC_9_502 b_9 NI_9 NS_502 0 -5.7373344947339092e-05
GC_9_503 b_9 NI_9 NS_503 0 -5.0364603611441437e-04
GC_9_504 b_9 NI_9 NS_504 0 6.7167669742950148e-04
GC_9_505 b_9 NI_9 NS_505 0 3.8218817592004198e-04
GC_9_506 b_9 NI_9 NS_506 0 2.1974337081503590e-04
GC_9_507 b_9 NI_9 NS_507 0 -3.8368825835013048e-05
GC_9_508 b_9 NI_9 NS_508 0 -5.5206536580870244e-05
GC_9_509 b_9 NI_9 NS_509 0 -4.5984203314077033e-05
GC_9_510 b_9 NI_9 NS_510 0 8.1003859134061334e-05
GC_9_511 b_9 NI_9 NS_511 0 -2.2101035513941484e-03
GC_9_512 b_9 NI_9 NS_512 0 -4.9286261330822529e-03
GC_9_513 b_9 NI_9 NS_513 0 8.8201569380158888e-06
GC_9_514 b_9 NI_9 NS_514 0 3.1308145197649062e-05
GC_9_515 b_9 NI_9 NS_515 0 -1.0172721444234585e-03
GC_9_516 b_9 NI_9 NS_516 0 2.0857168390285268e-03
GC_9_517 b_9 NI_9 NS_517 0 -3.9419795722248717e-06
GC_9_518 b_9 NI_9 NS_518 0 9.8955693875705696e-06
GC_9_519 b_9 NI_9 NS_519 0 1.1473988216288279e-03
GC_9_520 b_9 NI_9 NS_520 0 -1.9937430991743757e-04
GC_9_521 b_9 NI_9 NS_521 0 -9.1484455364567383e-06
GC_9_522 b_9 NI_9 NS_522 0 -1.4434541503985502e-05
GC_9_523 b_9 NI_9 NS_523 0 2.8249065377721478e-06
GC_9_524 b_9 NI_9 NS_524 0 2.5727351529563681e-07
GC_9_525 b_9 NI_9 NS_525 0 1.9039410044481964e-06
GC_9_526 b_9 NI_9 NS_526 0 3.8167548274189859e-06
GC_9_527 b_9 NI_9 NS_527 0 1.3994629961598518e-04
GC_9_528 b_9 NI_9 NS_528 0 -6.3155412284953425e-05
GD_9_1 b_9 NI_9 NA_1 0 -1.6578067018801879e-02
GD_9_2 b_9 NI_9 NA_2 0 -1.1751497739157821e-02
GD_9_3 b_9 NI_9 NA_3 0 -1.4148907501164348e-02
GD_9_4 b_9 NI_9 NA_4 0 -9.6793188063905126e-03
GD_9_5 b_9 NI_9 NA_5 0 -1.0163011055385002e-02
GD_9_6 b_9 NI_9 NA_6 0 -2.9442930721581295e-03
GD_9_7 b_9 NI_9 NA_7 0 -7.4851737810938505e-03
GD_9_8 b_9 NI_9 NA_8 0 1.3218788982517673e-03
GD_9_9 b_9 NI_9 NA_9 0 -1.2318079883968620e-01
GD_9_10 b_9 NI_9 NA_10 0 -5.2577009914565022e-02
GD_9_11 b_9 NI_9 NA_11 0 4.8325391675808210e-03
GD_9_12 b_9 NI_9 NA_12 0 -6.4891693247782961e-02
*
* Port 10
VI_10 a_10 NI_10 0
RI_10 NI_10 b_10 5.0000000000000000e+01
GC_10_1 b_10 NI_10 NS_1 0 1.0445798345885047e-02
GC_10_2 b_10 NI_10 NS_2 0 1.1156105786918765e-05
GC_10_3 b_10 NI_10 NS_3 0 5.2714340756841015e-05
GC_10_4 b_10 NI_10 NS_4 0 1.2181908853733979e-04
GC_10_5 b_10 NI_10 NS_5 0 -1.6323517218127628e-04
GC_10_6 b_10 NI_10 NS_6 0 -3.8764789145001790e-05
GC_10_7 b_10 NI_10 NS_7 0 -5.0431481608412753e-04
GC_10_8 b_10 NI_10 NS_8 0 -1.4340181294824101e-04
GC_10_9 b_10 NI_10 NS_9 0 1.8245941052621038e-04
GC_10_10 b_10 NI_10 NS_10 0 -2.8130670805904222e-04
GC_10_11 b_10 NI_10 NS_11 0 9.4346780596813839e-04
GC_10_12 b_10 NI_10 NS_12 0 6.3595592624551825e-05
GC_10_13 b_10 NI_10 NS_13 0 9.3702367669087441e-05
GC_10_14 b_10 NI_10 NS_14 0 6.1330313913874181e-05
GC_10_15 b_10 NI_10 NS_15 0 -1.2731414047712891e-04
GC_10_16 b_10 NI_10 NS_16 0 1.7312365815903888e-03
GC_10_17 b_10 NI_10 NS_17 0 -1.3386865054446114e-04
GC_10_18 b_10 NI_10 NS_18 0 6.5364885657529919e-05
GC_10_19 b_10 NI_10 NS_19 0 -5.9194929116525373e-04
GC_10_20 b_10 NI_10 NS_20 0 -7.9692111299013471e-05
GC_10_21 b_10 NI_10 NS_21 0 2.6351458292519991e-05
GC_10_22 b_10 NI_10 NS_22 0 -1.3989659762863761e-04
GC_10_23 b_10 NI_10 NS_23 0 -3.3709172044034054e-05
GC_10_24 b_10 NI_10 NS_24 0 -1.0934840339557836e-04
GC_10_25 b_10 NI_10 NS_25 0 -5.2985295736003403e-06
GC_10_26 b_10 NI_10 NS_26 0 1.0607258538668135e-04
GC_10_27 b_10 NI_10 NS_27 0 -2.3076863559121937e-04
GC_10_28 b_10 NI_10 NS_28 0 5.7415774002555966e-04
GC_10_29 b_10 NI_10 NS_29 0 -2.2802594025743819e-05
GC_10_30 b_10 NI_10 NS_30 0 -1.2185415448913340e-05
GC_10_31 b_10 NI_10 NS_31 0 -1.6734881734211727e-04
GC_10_32 b_10 NI_10 NS_32 0 -1.8254091192345772e-04
GC_10_33 b_10 NI_10 NS_33 0 1.4834463485302082e-06
GC_10_34 b_10 NI_10 NS_34 0 1.1010844430736774e-06
GC_10_35 b_10 NI_10 NS_35 0 -1.1480178822815268e-04
GC_10_36 b_10 NI_10 NS_36 0 -3.8368668690194835e-04
GC_10_37 b_10 NI_10 NS_37 0 -9.8078584142739244e-06
GC_10_38 b_10 NI_10 NS_38 0 -8.7495988509323613e-06
GC_10_39 b_10 NI_10 NS_39 0 -1.0728586460362626e-06
GC_10_40 b_10 NI_10 NS_40 0 1.2891761204566895e-06
GC_10_41 b_10 NI_10 NS_41 0 2.1697494960998458e-06
GC_10_42 b_10 NI_10 NS_42 0 -2.0403189741341821e-06
GC_10_43 b_10 NI_10 NS_43 0 -2.2730625127488280e-04
GC_10_44 b_10 NI_10 NS_44 0 -7.0817492633489228e-05
GC_10_45 b_10 NI_10 NS_45 0 3.1392042270284317e-03
GC_10_46 b_10 NI_10 NS_46 0 -1.4727048154197602e-05
GC_10_47 b_10 NI_10 NS_47 0 -1.1665231639379699e-04
GC_10_48 b_10 NI_10 NS_48 0 -1.2814012631827943e-04
GC_10_49 b_10 NI_10 NS_49 0 1.4448570206008728e-04
GC_10_50 b_10 NI_10 NS_50 0 -1.4445975474569381e-04
GC_10_51 b_10 NI_10 NS_51 0 -3.9538377913743417e-04
GC_10_52 b_10 NI_10 NS_52 0 -2.4173288850168250e-04
GC_10_53 b_10 NI_10 NS_53 0 7.3811167200999765e-05
GC_10_54 b_10 NI_10 NS_54 0 -2.2448948768730056e-04
GC_10_55 b_10 NI_10 NS_55 0 4.2540236478463589e-04
GC_10_56 b_10 NI_10 NS_56 0 -3.9300490848977469e-04
GC_10_57 b_10 NI_10 NS_57 0 1.4198989478178900e-05
GC_10_58 b_10 NI_10 NS_58 0 1.9463010674277963e-05
GC_10_59 b_10 NI_10 NS_59 0 5.4659502947086128e-04
GC_10_60 b_10 NI_10 NS_60 0 -1.8602978418755950e-04
GC_10_61 b_10 NI_10 NS_61 0 1.3269887275813519e-05
GC_10_62 b_10 NI_10 NS_62 0 -4.7731187553466309e-05
GC_10_63 b_10 NI_10 NS_63 0 6.8516055778491643e-04
GC_10_64 b_10 NI_10 NS_64 0 -2.9954464366731157e-04
GC_10_65 b_10 NI_10 NS_65 0 -2.9310255717654470e-04
GC_10_66 b_10 NI_10 NS_66 0 -3.4750843296683888e-04
GC_10_67 b_10 NI_10 NS_67 0 9.3111115450081387e-06
GC_10_68 b_10 NI_10 NS_68 0 -2.3233505324903272e-05
GC_10_69 b_10 NI_10 NS_69 0 -4.3855666996701468e-05
GC_10_70 b_10 NI_10 NS_70 0 -1.5810115206241866e-04
GC_10_71 b_10 NI_10 NS_71 0 -3.9515666254281564e-03
GC_10_72 b_10 NI_10 NS_72 0 4.6472531506407504e-03
GC_10_73 b_10 NI_10 NS_73 0 2.0019926849919699e-05
GC_10_74 b_10 NI_10 NS_74 0 2.0213601388854061e-05
GC_10_75 b_10 NI_10 NS_75 0 3.3768989065141469e-03
GC_10_76 b_10 NI_10 NS_76 0 -1.3815276327511930e-03
GC_10_77 b_10 NI_10 NS_77 0 2.2583083982312909e-05
GC_10_78 b_10 NI_10 NS_78 0 9.3600499611548355e-07
GC_10_79 b_10 NI_10 NS_79 0 -4.3990879312169086e-04
GC_10_80 b_10 NI_10 NS_80 0 -3.0573733414790823e-04
GC_10_81 b_10 NI_10 NS_81 0 -5.3083223840708894e-05
GC_10_82 b_10 NI_10 NS_82 0 1.0412448028611301e-05
GC_10_83 b_10 NI_10 NS_83 0 2.8754363054863343e-05
GC_10_84 b_10 NI_10 NS_84 0 -6.5451805268049171e-06
GC_10_85 b_10 NI_10 NS_85 0 -2.2397670208755304e-05
GC_10_86 b_10 NI_10 NS_86 0 1.6570121379749851e-05
GC_10_87 b_10 NI_10 NS_87 0 4.1369151991113123e-04
GC_10_88 b_10 NI_10 NS_88 0 1.6392327746066551e-04
GC_10_89 b_10 NI_10 NS_89 0 7.7280265844021107e-03
GC_10_90 b_10 NI_10 NS_90 0 9.0202204725899222e-06
GC_10_91 b_10 NI_10 NS_91 0 -9.6634488202786178e-05
GC_10_92 b_10 NI_10 NS_92 0 2.9651571857918001e-04
GC_10_93 b_10 NI_10 NS_93 0 -3.3163443963492615e-04
GC_10_94 b_10 NI_10 NS_94 0 -3.2884471614253862e-04
GC_10_95 b_10 NI_10 NS_95 0 -4.0412104358282687e-04
GC_10_96 b_10 NI_10 NS_96 0 8.6763312997064393e-05
GC_10_97 b_10 NI_10 NS_97 0 2.9350207524351423e-04
GC_10_98 b_10 NI_10 NS_98 0 -4.4776193796840246e-04
GC_10_99 b_10 NI_10 NS_99 0 6.2516853924440418e-04
GC_10_100 b_10 NI_10 NS_100 0 -1.8960918618451483e-05
GC_10_101 b_10 NI_10 NS_101 0 1.3539220472553418e-04
GC_10_102 b_10 NI_10 NS_102 0 9.4950342091780864e-05
GC_10_103 b_10 NI_10 NS_103 0 3.4862200771518415e-05
GC_10_104 b_10 NI_10 NS_104 0 1.4119830710187695e-03
GC_10_105 b_10 NI_10 NS_105 0 -1.8260134413015220e-04
GC_10_106 b_10 NI_10 NS_106 0 7.9695822135996991e-05
GC_10_107 b_10 NI_10 NS_107 0 -7.0512394796178469e-04
GC_10_108 b_10 NI_10 NS_108 0 -2.9672200171936512e-04
GC_10_109 b_10 NI_10 NS_109 0 -2.4767152800182374e-05
GC_10_110 b_10 NI_10 NS_110 0 -3.0036082024539753e-05
GC_10_111 b_10 NI_10 NS_111 0 -4.4857128751441353e-05
GC_10_112 b_10 NI_10 NS_112 0 -1.6601802972889676e-04
GC_10_113 b_10 NI_10 NS_113 0 -2.0894933549451156e-05
GC_10_114 b_10 NI_10 NS_114 0 1.3600740242876888e-04
GC_10_115 b_10 NI_10 NS_115 0 1.4084978598438199e-03
GC_10_116 b_10 NI_10 NS_116 0 1.2981759269940078e-03
GC_10_117 b_10 NI_10 NS_117 0 -3.2343135050856313e-05
GC_10_118 b_10 NI_10 NS_118 0 -1.4843822911213776e-05
GC_10_119 b_10 NI_10 NS_119 0 -5.0841242196674439e-04
GC_10_120 b_10 NI_10 NS_120 0 -9.3666150314275281e-04
GC_10_121 b_10 NI_10 NS_121 0 7.7396634277976096e-07
GC_10_122 b_10 NI_10 NS_122 0 -8.2858693465808597e-07
GC_10_123 b_10 NI_10 NS_123 0 -2.6889382334608199e-04
GC_10_124 b_10 NI_10 NS_124 0 -2.7151585644144397e-04
GC_10_125 b_10 NI_10 NS_125 0 -9.4411536697898700e-06
GC_10_126 b_10 NI_10 NS_126 0 -8.5978046106090909e-06
GC_10_127 b_10 NI_10 NS_127 0 -8.1906673581318271e-07
GC_10_128 b_10 NI_10 NS_128 0 6.8055887963105734e-08
GC_10_129 b_10 NI_10 NS_129 0 6.1738909035151140e-07
GC_10_130 b_10 NI_10 NS_130 0 -1.9212070177800825e-06
GC_10_131 b_10 NI_10 NS_131 0 -3.1984535111148773e-04
GC_10_132 b_10 NI_10 NS_132 0 -8.6008306220954701e-05
GC_10_133 b_10 NI_10 NS_133 0 1.5261941977131553e-03
GC_10_134 b_10 NI_10 NS_134 0 -1.5319598366534696e-05
GC_10_135 b_10 NI_10 NS_135 0 -9.5775329199510612e-05
GC_10_136 b_10 NI_10 NS_136 0 -3.4024140403571707e-04
GC_10_137 b_10 NI_10 NS_137 0 3.2583761549048046e-04
GC_10_138 b_10 NI_10 NS_138 0 -7.3639757150750223e-05
GC_10_139 b_10 NI_10 NS_139 0 -3.9906035393941404e-04
GC_10_140 b_10 NI_10 NS_140 0 3.9982820593259139e-05
GC_10_141 b_10 NI_10 NS_141 0 1.5255884741934594e-04
GC_10_142 b_10 NI_10 NS_142 0 -2.6852099194122156e-04
GC_10_143 b_10 NI_10 NS_143 0 4.6393368013922281e-04
GC_10_144 b_10 NI_10 NS_144 0 -3.6411470906455150e-04
GC_10_145 b_10 NI_10 NS_145 0 1.3626390400658627e-05
GC_10_146 b_10 NI_10 NS_146 0 4.0018141946860694e-05
GC_10_147 b_10 NI_10 NS_147 0 6.6803819393916315e-04
GC_10_148 b_10 NI_10 NS_148 0 -4.2046827255571813e-04
GC_10_149 b_10 NI_10 NS_149 0 1.6906141685769878e-05
GC_10_150 b_10 NI_10 NS_150 0 -5.1056777976307996e-05
GC_10_151 b_10 NI_10 NS_151 0 8.5696231054348834e-04
GC_10_152 b_10 NI_10 NS_152 0 -3.7368037799422792e-04
GC_10_153 b_10 NI_10 NS_153 0 -2.2643100634554131e-04
GC_10_154 b_10 NI_10 NS_154 0 -3.2059432880596791e-04
GC_10_155 b_10 NI_10 NS_155 0 1.3707448884581506e-05
GC_10_156 b_10 NI_10 NS_156 0 -2.5539863199719088e-05
GC_10_157 b_10 NI_10 NS_157 0 -4.4913202417474277e-05
GC_10_158 b_10 NI_10 NS_158 0 -1.7837500363309590e-04
GC_10_159 b_10 NI_10 NS_159 0 -4.5214064157944392e-03
GC_10_160 b_10 NI_10 NS_160 0 5.5192320492071295e-03
GC_10_161 b_10 NI_10 NS_161 0 1.9681308043240201e-05
GC_10_162 b_10 NI_10 NS_162 0 1.8399778805863191e-05
GC_10_163 b_10 NI_10 NS_163 0 3.9278727568378569e-03
GC_10_164 b_10 NI_10 NS_164 0 -1.6403554225812066e-03
GC_10_165 b_10 NI_10 NS_165 0 1.8963351723394253e-05
GC_10_166 b_10 NI_10 NS_166 0 3.1967088314425952e-06
GC_10_167 b_10 NI_10 NS_167 0 -3.6724315343308596e-04
GC_10_168 b_10 NI_10 NS_168 0 -4.8547844065716968e-04
GC_10_169 b_10 NI_10 NS_169 0 -4.9843697472967616e-05
GC_10_170 b_10 NI_10 NS_170 0 1.1155930631541816e-05
GC_10_171 b_10 NI_10 NS_171 0 3.1539029017627301e-05
GC_10_172 b_10 NI_10 NS_172 0 -5.5713807446737285e-06
GC_10_173 b_10 NI_10 NS_173 0 -2.3464566286205734e-05
GC_10_174 b_10 NI_10 NS_174 0 1.3832772271025872e-05
GC_10_175 b_10 NI_10 NS_175 0 4.1989882756594907e-04
GC_10_176 b_10 NI_10 NS_176 0 1.2945206282543610e-04
GC_10_177 b_10 NI_10 NS_177 0 -7.1088849107401480e-04
GC_10_178 b_10 NI_10 NS_178 0 -1.0290584205598624e-05
GC_10_179 b_10 NI_10 NS_179 0 -4.1250910329951329e-04
GC_10_180 b_10 NI_10 NS_180 0 4.7815803778895129e-04
GC_10_181 b_10 NI_10 NS_181 0 -3.9399575879368008e-04
GC_10_182 b_10 NI_10 NS_182 0 -7.2278800105011619e-04
GC_10_183 b_10 NI_10 NS_183 0 1.7080006447711593e-04
GC_10_184 b_10 NI_10 NS_184 0 9.8664442907403017e-05
GC_10_185 b_10 NI_10 NS_185 0 3.6260541168386587e-04
GC_10_186 b_10 NI_10 NS_186 0 -4.4679531492043949e-04
GC_10_187 b_10 NI_10 NS_187 0 -1.3702939240883738e-04
GC_10_188 b_10 NI_10 NS_188 0 -3.3659294257144801e-04
GC_10_189 b_10 NI_10 NS_189 0 1.4010813851147782e-04
GC_10_190 b_10 NI_10 NS_190 0 9.8537587419488115e-05
GC_10_191 b_10 NI_10 NS_191 0 6.2326444062824667e-04
GC_10_192 b_10 NI_10 NS_192 0 7.9136181572986763e-04
GC_10_193 b_10 NI_10 NS_193 0 -1.7591874792036079e-04
GC_10_194 b_10 NI_10 NS_194 0 8.9003469355087702e-05
GC_10_195 b_10 NI_10 NS_195 0 -6.3010392098775396e-04
GC_10_196 b_10 NI_10 NS_196 0 -2.6044385107369564e-04
GC_10_197 b_10 NI_10 NS_197 0 1.0028196390046543e-05
GC_10_198 b_10 NI_10 NS_198 0 -5.0794922346877499e-06
GC_10_199 b_10 NI_10 NS_199 0 -3.2384806391991925e-05
GC_10_200 b_10 NI_10 NS_200 0 -1.6288168404863772e-04
GC_10_201 b_10 NI_10 NS_201 0 -2.7079363314778665e-06
GC_10_202 b_10 NI_10 NS_202 0 1.3740897235171512e-04
GC_10_203 b_10 NI_10 NS_203 0 1.7623174796984188e-03
GC_10_204 b_10 NI_10 NS_204 0 5.1534815155813637e-04
GC_10_205 b_10 NI_10 NS_205 0 -3.4570806902445220e-05
GC_10_206 b_10 NI_10 NS_206 0 -1.2429379872037578e-05
GC_10_207 b_10 NI_10 NS_207 0 -6.0693986851777324e-04
GC_10_208 b_10 NI_10 NS_208 0 -6.4955916958582636e-04
GC_10_209 b_10 NI_10 NS_209 0 -3.0075113612795246e-07
GC_10_210 b_10 NI_10 NS_210 0 2.8853001138273780e-06
GC_10_211 b_10 NI_10 NS_211 0 -1.6611803702613163e-04
GC_10_212 b_10 NI_10 NS_212 0 -1.9127878195845293e-04
GC_10_213 b_10 NI_10 NS_213 0 -1.5211829052091201e-05
GC_10_214 b_10 NI_10 NS_214 0 -2.1541416894725795e-05
GC_10_215 b_10 NI_10 NS_215 0 -1.1816764519110102e-07
GC_10_216 b_10 NI_10 NS_216 0 2.7174551912918689e-06
GC_10_217 b_10 NI_10 NS_217 0 -1.9245062663532437e-06
GC_10_218 b_10 NI_10 NS_218 0 -2.3028589208291682e-06
GC_10_219 b_10 NI_10 NS_219 0 -3.4362024833352106e-04
GC_10_220 b_10 NI_10 NS_220 0 -2.5267490532350786e-05
GC_10_221 b_10 NI_10 NS_221 0 -1.6129938180432196e-03
GC_10_222 b_10 NI_10 NS_222 0 -1.1216280371254019e-06
GC_10_223 b_10 NI_10 NS_223 0 8.6298601442430276e-05
GC_10_224 b_10 NI_10 NS_224 0 -6.0149869369356332e-04
GC_10_225 b_10 NI_10 NS_225 0 4.6217613371958761e-04
GC_10_226 b_10 NI_10 NS_226 0 1.7239974560952228e-04
GC_10_227 b_10 NI_10 NS_227 0 -6.4557502753025521e-04
GC_10_228 b_10 NI_10 NS_228 0 1.3454361216322893e-05
GC_10_229 b_10 NI_10 NS_229 0 1.9087915044508892e-04
GC_10_230 b_10 NI_10 NS_230 0 -2.3417011386519667e-04
GC_10_231 b_10 NI_10 NS_231 0 1.7009027506019261e-04
GC_10_232 b_10 NI_10 NS_232 0 -3.9750363413603855e-04
GC_10_233 b_10 NI_10 NS_233 0 2.5851660907433988e-05
GC_10_234 b_10 NI_10 NS_234 0 4.2872190148310921e-05
GC_10_235 b_10 NI_10 NS_235 0 1.0420958346157112e-03
GC_10_236 b_10 NI_10 NS_236 0 -8.8542226358457297e-04
GC_10_237 b_10 NI_10 NS_237 0 2.3399744822299513e-05
GC_10_238 b_10 NI_10 NS_238 0 -6.5819520446154802e-05
GC_10_239 b_10 NI_10 NS_239 0 1.1041828901449985e-03
GC_10_240 b_10 NI_10 NS_240 0 -4.9338505120226090e-04
GC_10_241 b_10 NI_10 NS_241 0 -3.7362382505032722e-04
GC_10_242 b_10 NI_10 NS_242 0 -5.0906320588126074e-04
GC_10_243 b_10 NI_10 NS_243 0 1.4981476835019626e-05
GC_10_244 b_10 NI_10 NS_244 0 -3.7130324350036486e-05
GC_10_245 b_10 NI_10 NS_245 0 -7.2096742130449469e-05
GC_10_246 b_10 NI_10 NS_246 0 -2.3775088355202371e-04
GC_10_247 b_10 NI_10 NS_247 0 -5.3620413423565473e-03
GC_10_248 b_10 NI_10 NS_248 0 7.4549018750605109e-03
GC_10_249 b_10 NI_10 NS_249 0 2.3383017597113849e-05
GC_10_250 b_10 NI_10 NS_250 0 2.3332420279071107e-05
GC_10_251 b_10 NI_10 NS_251 0 5.0524938006929199e-03
GC_10_252 b_10 NI_10 NS_252 0 -2.4214348915788482e-03
GC_10_253 b_10 NI_10 NS_253 0 3.4032351581172340e-05
GC_10_254 b_10 NI_10 NS_254 0 4.7094825646912173e-06
GC_10_255 b_10 NI_10 NS_255 0 -6.0307805617413257e-04
GC_10_256 b_10 NI_10 NS_256 0 -5.4086150588994713e-04
GC_10_257 b_10 NI_10 NS_257 0 -7.7108763443179762e-05
GC_10_258 b_10 NI_10 NS_258 0 2.0771886408219758e-05
GC_10_259 b_10 NI_10 NS_259 0 4.4023055567395630e-05
GC_10_260 b_10 NI_10 NS_260 0 -1.2450719914018006e-05
GC_10_261 b_10 NI_10 NS_261 0 -2.6682140053387920e-05
GC_10_262 b_10 NI_10 NS_262 0 2.4203943022340418e-05
GC_10_263 b_10 NI_10 NS_263 0 5.9698486964844131e-04
GC_10_264 b_10 NI_10 NS_264 0 2.0364815574528436e-04
GC_10_265 b_10 NI_10 NS_265 0 -6.2322634914589127e-03
GC_10_266 b_10 NI_10 NS_266 0 -1.2416071890693732e-05
GC_10_267 b_10 NI_10 NS_267 0 -1.3035774726329198e-03
GC_10_268 b_10 NI_10 NS_268 0 1.9884360932291247e-04
GC_10_269 b_10 NI_10 NS_269 0 6.2664041871335211e-04
GC_10_270 b_10 NI_10 NS_270 0 -1.2431051798781848e-03
GC_10_271 b_10 NI_10 NS_271 0 1.7210278963663753e-04
GC_10_272 b_10 NI_10 NS_272 0 4.2920511807441059e-04
GC_10_273 b_10 NI_10 NS_273 0 6.8009317943017330e-04
GC_10_274 b_10 NI_10 NS_274 0 -1.5853185863977159e-04
GC_10_275 b_10 NI_10 NS_275 0 -3.0814038140888715e-04
GC_10_276 b_10 NI_10 NS_276 0 -1.1173399442954981e-03
GC_10_277 b_10 NI_10 NS_277 0 1.2333963613170610e-04
GC_10_278 b_10 NI_10 NS_278 0 8.7534403679941680e-05
GC_10_279 b_10 NI_10 NS_279 0 9.0830992529413910e-04
GC_10_280 b_10 NI_10 NS_280 0 1.1149235050586252e-03
GC_10_281 b_10 NI_10 NS_281 0 -1.2352304983233219e-04
GC_10_282 b_10 NI_10 NS_282 0 4.6413235104859305e-05
GC_10_283 b_10 NI_10 NS_283 0 -2.7408836361905665e-04
GC_10_284 b_10 NI_10 NS_284 0 -1.3257425722241619e-04
GC_10_285 b_10 NI_10 NS_285 0 -8.6050522928789891e-06
GC_10_286 b_10 NI_10 NS_286 0 1.0950272478977466e-04
GC_10_287 b_10 NI_10 NS_287 0 -1.8675625068171725e-05
GC_10_288 b_10 NI_10 NS_288 0 -1.1250038395683270e-04
GC_10_289 b_10 NI_10 NS_289 0 -2.4144023941194704e-05
GC_10_290 b_10 NI_10 NS_290 0 1.0005723471211786e-04
GC_10_291 b_10 NI_10 NS_291 0 1.6840836983295772e-03
GC_10_292 b_10 NI_10 NS_292 0 4.0776072411999060e-04
GC_10_293 b_10 NI_10 NS_293 0 -1.9460197963634631e-05
GC_10_294 b_10 NI_10 NS_294 0 -5.2366315429151821e-06
GC_10_295 b_10 NI_10 NS_295 0 -5.0767072271653429e-04
GC_10_296 b_10 NI_10 NS_296 0 -5.8499862186993520e-04
GC_10_297 b_10 NI_10 NS_297 0 -2.9905042440611839e-06
GC_10_298 b_10 NI_10 NS_298 0 -1.1786801177763678e-06
GC_10_299 b_10 NI_10 NS_299 0 4.1730246322955097e-05
GC_10_300 b_10 NI_10 NS_300 0 1.3928214623579125e-05
GC_10_301 b_10 NI_10 NS_301 0 -7.3520328692516829e-06
GC_10_302 b_10 NI_10 NS_302 0 -1.3797200576220196e-05
GC_10_303 b_10 NI_10 NS_303 0 2.5650292637822131e-07
GC_10_304 b_10 NI_10 NS_304 0 -2.1526931190488012e-07
GC_10_305 b_10 NI_10 NS_305 0 -7.7261866494944046e-07
GC_10_306 b_10 NI_10 NS_306 0 -4.5527832805265814e-07
GC_10_307 b_10 NI_10 NS_307 0 -1.9540881946200755e-04
GC_10_308 b_10 NI_10 NS_308 0 -4.7659893087259750e-05
GC_10_309 b_10 NI_10 NS_309 0 -2.3345115037887051e-04
GC_10_310 b_10 NI_10 NS_310 0 -3.2970542042603271e-05
GC_10_311 b_10 NI_10 NS_311 0 8.1136508213154233e-04
GC_10_312 b_10 NI_10 NS_312 0 -5.7431833981704569e-04
GC_10_313 b_10 NI_10 NS_313 0 -2.7931887909861256e-04
GC_10_314 b_10 NI_10 NS_314 0 7.6862165704999670e-04
GC_10_315 b_10 NI_10 NS_315 0 -5.3118289745463757e-04
GC_10_316 b_10 NI_10 NS_316 0 7.8733510734157596e-05
GC_10_317 b_10 NI_10 NS_317 0 1.6731011811870175e-04
GC_10_318 b_10 NI_10 NS_318 0 -1.4298139966765851e-04
GC_10_319 b_10 NI_10 NS_319 0 -1.4733629585662501e-04
GC_10_320 b_10 NI_10 NS_320 0 -1.7551594523040480e-04
GC_10_321 b_10 NI_10 NS_321 0 -9.1393439180958911e-06
GC_10_322 b_10 NI_10 NS_322 0 1.8521895865082134e-05
GC_10_323 b_10 NI_10 NS_323 0 4.6414426205551449e-04
GC_10_324 b_10 NI_10 NS_324 0 -5.5381479028079292e-05
GC_10_325 b_10 NI_10 NS_325 0 1.3031382758941844e-05
GC_10_326 b_10 NI_10 NS_326 0 -4.2861688095860301e-05
GC_10_327 b_10 NI_10 NS_327 0 4.4991053647490056e-04
GC_10_328 b_10 NI_10 NS_328 0 -3.0860129063767060e-04
GC_10_329 b_10 NI_10 NS_329 0 -6.4627580193048014e-05
GC_10_330 b_10 NI_10 NS_330 0 -2.0303595030685015e-04
GC_10_331 b_10 NI_10 NS_331 0 -1.3024353841261244e-07
GC_10_332 b_10 NI_10 NS_332 0 -2.9082176289076277e-05
GC_10_333 b_10 NI_10 NS_333 0 -4.7331757060001566e-05
GC_10_334 b_10 NI_10 NS_334 0 -1.4943585407488946e-04
GC_10_335 b_10 NI_10 NS_335 0 -3.2088715496302357e-03
GC_10_336 b_10 NI_10 NS_336 0 2.9751852932857641e-03
GC_10_337 b_10 NI_10 NS_337 0 6.9811125770703691e-06
GC_10_338 b_10 NI_10 NS_338 0 5.8153286828863824e-06
GC_10_339 b_10 NI_10 NS_339 0 2.7935002119964382e-03
GC_10_340 b_10 NI_10 NS_340 0 -1.0271068466381852e-03
GC_10_341 b_10 NI_10 NS_341 0 1.1192633568933525e-05
GC_10_342 b_10 NI_10 NS_342 0 6.5893740746664054e-06
GC_10_343 b_10 NI_10 NS_343 0 4.5241610918166637e-05
GC_10_344 b_10 NI_10 NS_344 0 -2.7697856894458946e-04
GC_10_345 b_10 NI_10 NS_345 0 -3.4507818246039386e-05
GC_10_346 b_10 NI_10 NS_346 0 1.8608654439488064e-06
GC_10_347 b_10 NI_10 NS_347 0 2.8555673918684445e-05
GC_10_348 b_10 NI_10 NS_348 0 -3.8266426295816841e-06
GC_10_349 b_10 NI_10 NS_349 0 -1.0952885267552230e-05
GC_10_350 b_10 NI_10 NS_350 0 8.9524069307029082e-06
GC_10_351 b_10 NI_10 NS_351 0 3.1196288953861089e-04
GC_10_352 b_10 NI_10 NS_352 0 1.2630031372981809e-04
GC_10_353 b_10 NI_10 NS_353 0 5.5079885172447919e-02
GC_10_354 b_10 NI_10 NS_354 0 1.0249097508377991e-02
GC_10_355 b_10 NI_10 NS_355 0 -1.0900785196268838e-02
GC_10_356 b_10 NI_10 NS_356 0 -2.8075048844162964e-03
GC_10_357 b_10 NI_10 NS_357 0 -1.1111934901257428e-02
GC_10_358 b_10 NI_10 NS_358 0 -2.0162350986476928e-03
GC_10_359 b_10 NI_10 NS_359 0 3.4216451632230484e-04
GC_10_360 b_10 NI_10 NS_360 0 1.7538471475903641e-04
GC_10_361 b_10 NI_10 NS_361 0 2.8570119427780362e-03
GC_10_362 b_10 NI_10 NS_362 0 2.5669763841480232e-03
GC_10_363 b_10 NI_10 NS_363 0 -7.1641143575622637e-04
GC_10_364 b_10 NI_10 NS_364 0 -3.7785910792755559e-04
GC_10_365 b_10 NI_10 NS_365 0 -3.2407103621816219e-06
GC_10_366 b_10 NI_10 NS_366 0 1.6235831740495508e-04
GC_10_367 b_10 NI_10 NS_367 0 2.1652453147647235e-03
GC_10_368 b_10 NI_10 NS_368 0 -9.3477382892972669e-04
GC_10_369 b_10 NI_10 NS_369 0 -7.9759638712865522e-05
GC_10_370 b_10 NI_10 NS_370 0 -7.8221968488663068e-05
GC_10_371 b_10 NI_10 NS_371 0 2.2662088464850874e-04
GC_10_372 b_10 NI_10 NS_372 0 7.5012201214202728e-04
GC_10_373 b_10 NI_10 NS_373 0 4.5585921892430428e-04
GC_10_374 b_10 NI_10 NS_374 0 9.5807685245857957e-06
GC_10_375 b_10 NI_10 NS_375 0 -1.1372072971644708e-05
GC_10_376 b_10 NI_10 NS_376 0 -7.2075787766220735e-05
GC_10_377 b_10 NI_10 NS_377 0 -6.4692380207092870e-05
GC_10_378 b_10 NI_10 NS_378 0 1.0151464243961415e-04
GC_10_379 b_10 NI_10 NS_379 0 -3.7213129836263484e-03
GC_10_380 b_10 NI_10 NS_380 0 -6.3818398993294931e-03
GC_10_381 b_10 NI_10 NS_381 0 1.9441165279643429e-05
GC_10_382 b_10 NI_10 NS_382 0 5.0541321235856596e-05
GC_10_383 b_10 NI_10 NS_383 0 -1.0614296184469343e-03
GC_10_384 b_10 NI_10 NS_384 0 2.9857789212590687e-03
GC_10_385 b_10 NI_10 NS_385 0 -3.5376691682339988e-06
GC_10_386 b_10 NI_10 NS_386 0 1.0088123397015968e-05
GC_10_387 b_10 NI_10 NS_387 0 1.2771011859919698e-03
GC_10_388 b_10 NI_10 NS_388 0 -6.9238023681688211e-04
GC_10_389 b_10 NI_10 NS_389 0 -1.0835274675704923e-05
GC_10_390 b_10 NI_10 NS_390 0 -1.1871256964783165e-05
GC_10_391 b_10 NI_10 NS_391 0 3.1750992780380276e-06
GC_10_392 b_10 NI_10 NS_392 0 1.5686657802304954e-07
GC_10_393 b_10 NI_10 NS_393 0 4.0891112544078022e-06
GC_10_394 b_10 NI_10 NS_394 0 2.5456789681106572e-06
GC_10_395 b_10 NI_10 NS_395 0 1.5524175377189942e-04
GC_10_396 b_10 NI_10 NS_396 0 -2.0845533503360120e-04
GC_10_397 b_10 NI_10 NS_397 0 -2.2594991372161166e-01
GC_10_398 b_10 NI_10 NS_398 0 8.6660674240525218e-03
GC_10_399 b_10 NI_10 NS_399 0 6.7697058097671327e-03
GC_10_400 b_10 NI_10 NS_400 0 3.8640470424665262e-03
GC_10_401 b_10 NI_10 NS_401 0 6.5718810672321286e-03
GC_10_402 b_10 NI_10 NS_402 0 1.3051872703833984e-03
GC_10_403 b_10 NI_10 NS_403 0 5.6335443569257096e-04
GC_10_404 b_10 NI_10 NS_404 0 4.7947529670119084e-04
GC_10_405 b_10 NI_10 NS_405 0 9.0876663309351737e-04
GC_10_406 b_10 NI_10 NS_406 0 1.5388210835884542e-03
GC_10_407 b_10 NI_10 NS_407 0 3.6633670430259928e-03
GC_10_408 b_10 NI_10 NS_408 0 3.0569328822583957e-03
GC_10_409 b_10 NI_10 NS_409 0 -2.2551832938010443e-04
GC_10_410 b_10 NI_10 NS_410 0 2.2724878003699440e-04
GC_10_411 b_10 NI_10 NS_411 0 1.6182731767061273e-03
GC_10_412 b_10 NI_10 NS_412 0 6.6640288325254459e-03
GC_10_413 b_10 NI_10 NS_413 0 -3.7817987807735173e-05
GC_10_414 b_10 NI_10 NS_414 0 4.8565874584353256e-05
GC_10_415 b_10 NI_10 NS_415 0 -3.1950958883331576e-04
GC_10_416 b_10 NI_10 NS_416 0 2.6071868680712534e-03
GC_10_417 b_10 NI_10 NS_417 0 6.0669916634225620e-04
GC_10_418 b_10 NI_10 NS_418 0 -7.5363185558610928e-04
GC_10_419 b_10 NI_10 NS_419 0 -9.8274742934651070e-05
GC_10_420 b_10 NI_10 NS_420 0 6.6838678576504177e-05
GC_10_421 b_10 NI_10 NS_421 0 -5.4808534642788891e-05
GC_10_422 b_10 NI_10 NS_422 0 -9.2846201909563096e-05
GC_10_423 b_10 NI_10 NS_423 0 -1.2172973660900621e-02
GC_10_424 b_10 NI_10 NS_424 0 2.2199131643503350e-03
GC_10_425 b_10 NI_10 NS_425 0 -3.4721488122913720e-05
GC_10_426 b_10 NI_10 NS_426 0 -6.5719987601377088e-05
GC_10_427 b_10 NI_10 NS_427 0 4.4681399320561097e-03
GC_10_428 b_10 NI_10 NS_428 0 2.5739181964929440e-03
GC_10_429 b_10 NI_10 NS_429 0 -1.1531561899430571e-05
GC_10_430 b_10 NI_10 NS_430 0 4.1333828548032238e-05
GC_10_431 b_10 NI_10 NS_431 0 7.1163705974267260e-04
GC_10_432 b_10 NI_10 NS_432 0 -1.7507861894730762e-03
GC_10_433 b_10 NI_10 NS_433 0 -3.7794415655995020e-05
GC_10_434 b_10 NI_10 NS_434 0 -2.0920320113600984e-05
GC_10_435 b_10 NI_10 NS_435 0 4.2973572794328960e-05
GC_10_436 b_10 NI_10 NS_436 0 -1.4590100852312617e-05
GC_10_437 b_10 NI_10 NS_437 0 5.6852970271972966e-05
GC_10_438 b_10 NI_10 NS_438 0 -2.3624179613460209e-05
GC_10_439 b_10 NI_10 NS_439 0 -2.8925798074105040e-05
GC_10_440 b_10 NI_10 NS_440 0 -1.0648096240312378e-04
GC_10_441 b_10 NI_10 NS_441 0 6.4982097490885571e-02
GC_10_442 b_10 NI_10 NS_442 0 -7.9954499781859006e-05
GC_10_443 b_10 NI_10 NS_443 0 -6.4095691830123418e-03
GC_10_444 b_10 NI_10 NS_444 0 -2.5862470334362519e-03
GC_10_445 b_10 NI_10 NS_445 0 4.2953376586868201e-03
GC_10_446 b_10 NI_10 NS_446 0 2.5496217089306097e-03
GC_10_447 b_10 NI_10 NS_447 0 -5.7986871121683866e-04
GC_10_448 b_10 NI_10 NS_448 0 -1.6472860858913487e-04
GC_10_449 b_10 NI_10 NS_449 0 1.5068227882712093e-03
GC_10_450 b_10 NI_10 NS_450 0 1.4953588887499098e-03
GC_10_451 b_10 NI_10 NS_451 0 -3.7977882160690073e-04
GC_10_452 b_10 NI_10 NS_452 0 -3.5978180221914532e-04
GC_10_453 b_10 NI_10 NS_453 0 -3.2659321816183206e-05
GC_10_454 b_10 NI_10 NS_454 0 7.4286695375952810e-05
GC_10_455 b_10 NI_10 NS_455 0 -4.0075330787572418e-03
GC_10_456 b_10 NI_10 NS_456 0 1.2348966679987009e-03
GC_10_457 b_10 NI_10 NS_457 0 -9.1324357043464911e-05
GC_10_458 b_10 NI_10 NS_458 0 -6.2364289763663897e-05
GC_10_459 b_10 NI_10 NS_459 0 -3.3852922119164834e-04
GC_10_460 b_10 NI_10 NS_460 0 8.5603857269848785e-04
GC_10_461 b_10 NI_10 NS_461 0 2.4651681906619346e-04
GC_10_462 b_10 NI_10 NS_462 0 1.0827517631606996e-04
GC_10_463 b_10 NI_10 NS_463 0 -3.1782974450842318e-05
GC_10_464 b_10 NI_10 NS_464 0 -6.4690402410939293e-05
GC_10_465 b_10 NI_10 NS_465 0 -6.4035102106578054e-05
GC_10_466 b_10 NI_10 NS_466 0 9.1653122159372649e-05
GC_10_467 b_10 NI_10 NS_467 0 -2.6102522623337263e-03
GC_10_468 b_10 NI_10 NS_468 0 -4.1099696298636506e-03
GC_10_469 b_10 NI_10 NS_469 0 4.9953670316701259e-06
GC_10_470 b_10 NI_10 NS_470 0 3.7688567736705239e-05
GC_10_471 b_10 NI_10 NS_471 0 -8.1465011928799830e-04
GC_10_472 b_10 NI_10 NS_472 0 2.1208816920138588e-03
GC_10_473 b_10 NI_10 NS_473 0 -3.3555708982125822e-06
GC_10_474 b_10 NI_10 NS_474 0 8.1496787466711667e-06
GC_10_475 b_10 NI_10 NS_475 0 9.0173225529161427e-04
GC_10_476 b_10 NI_10 NS_476 0 -2.9734244345509532e-04
GC_10_477 b_10 NI_10 NS_477 0 -8.8935394864351826e-06
GC_10_478 b_10 NI_10 NS_478 0 -1.0945848085526002e-05
GC_10_479 b_10 NI_10 NS_479 0 3.1108562994119338e-06
GC_10_480 b_10 NI_10 NS_480 0 -1.3430618940631939e-06
GC_10_481 b_10 NI_10 NS_481 0 1.9687573311095929e-06
GC_10_482 b_10 NI_10 NS_482 0 -4.8428928986882495e-07
GC_10_483 b_10 NI_10 NS_483 0 9.6562432086327765e-05
GC_10_484 b_10 NI_10 NS_484 0 -1.1241070115940110e-04
GC_10_485 b_10 NI_10 NS_485 0 2.4173200761658286e-03
GC_10_486 b_10 NI_10 NS_486 0 -8.9963953401236670e-04
GC_10_487 b_10 NI_10 NS_487 0 3.9215896045234093e-03
GC_10_488 b_10 NI_10 NS_488 0 1.5934910655745719e-03
GC_10_489 b_10 NI_10 NS_489 0 -5.1951684060271217e-03
GC_10_490 b_10 NI_10 NS_490 0 -2.2950835618088445e-03
GC_10_491 b_10 NI_10 NS_491 0 -1.9306587540382142e-05
GC_10_492 b_10 NI_10 NS_492 0 -3.2372028021262231e-04
GC_10_493 b_10 NI_10 NS_493 0 1.2198672017075325e-03
GC_10_494 b_10 NI_10 NS_494 0 7.2025048436841115e-05
GC_10_495 b_10 NI_10 NS_495 0 -1.1882254252938921e-04
GC_10_496 b_10 NI_10 NS_496 0 -4.9216401063620656e-04
GC_10_497 b_10 NI_10 NS_497 0 -3.0545348095281630e-05
GC_10_498 b_10 NI_10 NS_498 0 -3.9662352826719827e-05
GC_10_499 b_10 NI_10 NS_499 0 -1.4006382870501034e-03
GC_10_500 b_10 NI_10 NS_500 0 4.2432315911990589e-04
GC_10_501 b_10 NI_10 NS_501 0 2.4952484395984276e-05
GC_10_502 b_10 NI_10 NS_502 0 -3.2409263638301085e-05
GC_10_503 b_10 NI_10 NS_503 0 2.3828704999755765e-05
GC_10_504 b_10 NI_10 NS_504 0 -3.6215976704653385e-04
GC_10_505 b_10 NI_10 NS_505 0 1.8587166348127976e-04
GC_10_506 b_10 NI_10 NS_506 0 -6.1147365088913720e-05
GC_10_507 b_10 NI_10 NS_507 0 -8.6207219937669595e-06
GC_10_508 b_10 NI_10 NS_508 0 -4.8737169577157984e-05
GC_10_509 b_10 NI_10 NS_509 0 -6.4513434789059828e-05
GC_10_510 b_10 NI_10 NS_510 0 -1.2458553949252428e-04
GC_10_511 b_10 NI_10 NS_511 0 1.8961261743094657e-03
GC_10_512 b_10 NI_10 NS_512 0 -4.9493402687591224e-04
GC_10_513 b_10 NI_10 NS_513 0 -3.6844538246327047e-05
GC_10_514 b_10 NI_10 NS_514 0 -3.0272954604987923e-05
GC_10_515 b_10 NI_10 NS_515 0 6.2331791867573918e-04
GC_10_516 b_10 NI_10 NS_516 0 -7.2798220574652882e-04
GC_10_517 b_10 NI_10 NS_517 0 -1.0089473556631406e-05
GC_10_518 b_10 NI_10 NS_518 0 1.2150397114906538e-05
GC_10_519 b_10 NI_10 NS_519 0 4.2947275605289192e-04
GC_10_520 b_10 NI_10 NS_520 0 4.8341743772909829e-04
GC_10_521 b_10 NI_10 NS_521 0 -6.9441857692106417e-07
GC_10_522 b_10 NI_10 NS_522 0 -1.4088778969981107e-05
GC_10_523 b_10 NI_10 NS_523 0 2.8826109086968210e-05
GC_10_524 b_10 NI_10 NS_524 0 4.8882504842541647e-07
GC_10_525 b_10 NI_10 NS_525 0 1.9709692659308813e-05
GC_10_526 b_10 NI_10 NS_526 0 -7.9146041122049262e-06
GC_10_527 b_10 NI_10 NS_527 0 -6.7909410010081919e-05
GC_10_528 b_10 NI_10 NS_528 0 2.3598926368808900e-04
GD_10_1 b_10 NI_10 NA_1 0 -1.0469193834709857e-02
GD_10_2 b_10 NI_10 NA_2 0 -4.5743763923065135e-03
GD_10_3 b_10 NI_10 NA_3 0 -8.7399610071455108e-03
GD_10_4 b_10 NI_10 NA_4 0 -4.2863540065084527e-03
GD_10_5 b_10 NI_10 NA_5 0 2.3233316769428501e-04
GD_10_6 b_10 NI_10 NA_6 0 -1.1283511704556078e-03
GD_10_7 b_10 NI_10 NA_7 0 4.0000538907200853e-03
GD_10_8 b_10 NI_10 NA_8 0 -1.3222267237333494e-03
GD_10_9 b_10 NI_10 NA_9 0 -5.2577009914532208e-02
GD_10_10 b_10 NI_10 NA_10 0 2.6126986647181832e-01
GD_10_11 b_10 NI_10 NA_11 0 -6.6001193440252529e-02
GD_10_12 b_10 NI_10 NA_12 0 -8.6526583902597261e-03
*
* Port 11
VI_11 a_11 NI_11 0
RI_11 NI_11 b_11 5.0000000000000000e+01
GC_11_1 b_11 NI_11 NS_1 0 -4.8473916816486901e-03
GC_11_2 b_11 NI_11 NS_2 0 5.8193002899248519e-05
GC_11_3 b_11 NI_11 NS_3 0 2.5851860320959041e-04
GC_11_4 b_11 NI_11 NS_4 0 -6.1696650161226652e-04
GC_11_5 b_11 NI_11 NS_5 0 6.0893005020969874e-04
GC_11_6 b_11 NI_11 NS_6 0 2.5700322186662523e-04
GC_11_7 b_11 NI_11 NS_7 0 -1.7215809547936796e-04
GC_11_8 b_11 NI_11 NS_8 0 3.9989942727391466e-04
GC_11_9 b_11 NI_11 NS_9 0 8.3994807589277565e-04
GC_11_10 b_11 NI_11 NS_10 0 4.8884773325229877e-04
GC_11_11 b_11 NI_11 NS_11 0 -3.1212609639156880e-03
GC_11_12 b_11 NI_11 NS_12 0 9.1896700909737089e-04
GC_11_13 b_11 NI_11 NS_13 0 4.3581395274862848e-04
GC_11_14 b_11 NI_11 NS_14 0 -3.5686710409470521e-04
GC_11_15 b_11 NI_11 NS_15 0 3.0565703427418750e-03
GC_11_16 b_11 NI_11 NS_16 0 -2.4852298295363613e-03
GC_11_17 b_11 NI_11 NS_17 0 1.9537278461159393e-04
GC_11_18 b_11 NI_11 NS_18 0 1.9681133655354550e-04
GC_11_19 b_11 NI_11 NS_19 0 -2.6528209069482257e-04
GC_11_20 b_11 NI_11 NS_20 0 5.8143462088788183e-04
GC_11_21 b_11 NI_11 NS_21 0 1.9205127424194618e-04
GC_11_22 b_11 NI_11 NS_22 0 2.1095558443439777e-04
GC_11_23 b_11 NI_11 NS_23 0 1.0190831681233970e-04
GC_11_24 b_11 NI_11 NS_24 0 -5.0656230314694526e-05
GC_11_25 b_11 NI_11 NS_25 0 9.5731218469189356e-06
GC_11_26 b_11 NI_11 NS_26 0 6.0035205396192469e-05
GC_11_27 b_11 NI_11 NS_27 0 -1.7194347522501788e-03
GC_11_28 b_11 NI_11 NS_28 0 3.4195686874279527e-03
GC_11_29 b_11 NI_11 NS_29 0 2.2758905214588842e-06
GC_11_30 b_11 NI_11 NS_30 0 -4.2636900077783701e-06
GC_11_31 b_11 NI_11 NS_31 0 7.5314323528132921e-04
GC_11_32 b_11 NI_11 NS_32 0 -8.1751453311105886e-04
GC_11_33 b_11 NI_11 NS_33 0 -2.9690206859266314e-06
GC_11_34 b_11 NI_11 NS_34 0 4.5026133950992717e-06
GC_11_35 b_11 NI_11 NS_35 0 6.2327514253621955e-04
GC_11_36 b_11 NI_11 NS_36 0 -1.0591643280888055e-03
GC_11_37 b_11 NI_11 NS_37 0 -1.0813235041945276e-05
GC_11_38 b_11 NI_11 NS_38 0 -4.9049726034075299e-06
GC_11_39 b_11 NI_11 NS_39 0 1.1004026911715506e-06
GC_11_40 b_11 NI_11 NS_40 0 -1.0385899988455831e-07
GC_11_41 b_11 NI_11 NS_41 0 2.0437311014530864e-07
GC_11_42 b_11 NI_11 NS_42 0 3.5235791938011765e-06
GC_11_43 b_11 NI_11 NS_43 0 1.3478051522298464e-05
GC_11_44 b_11 NI_11 NS_44 0 -3.0832416697631430e-04
GC_11_45 b_11 NI_11 NS_45 0 1.5906152990963315e-02
GC_11_46 b_11 NI_11 NS_46 0 -4.0320958788108356e-05
GC_11_47 b_11 NI_11 NS_47 0 -1.3164639886722765e-04
GC_11_48 b_11 NI_11 NS_48 0 5.5101531541139749e-04
GC_11_49 b_11 NI_11 NS_49 0 -4.9856300340342711e-04
GC_11_50 b_11 NI_11 NS_50 0 -2.2826786249129032e-04
GC_11_51 b_11 NI_11 NS_51 0 -2.8765696173072328e-04
GC_11_52 b_11 NI_11 NS_52 0 -2.4519609645056909e-04
GC_11_53 b_11 NI_11 NS_53 0 3.1290750932331195e-04
GC_11_54 b_11 NI_11 NS_54 0 -3.7855692010178899e-05
GC_11_55 b_11 NI_11 NS_55 0 -2.9433566054198424e-04
GC_11_56 b_11 NI_11 NS_56 0 1.1003663910486448e-03
GC_11_57 b_11 NI_11 NS_57 0 6.2766487939072788e-05
GC_11_58 b_11 NI_11 NS_58 0 2.4802187766282737e-05
GC_11_59 b_11 NI_11 NS_59 0 -8.8249458763517245e-04
GC_11_60 b_11 NI_11 NS_60 0 3.7653877627055916e-04
GC_11_61 b_11 NI_11 NS_61 0 -9.2341021477939790e-05
GC_11_62 b_11 NI_11 NS_62 0 2.0573036701748738e-05
GC_11_63 b_11 NI_11 NS_63 0 -3.9481746080616856e-04
GC_11_64 b_11 NI_11 NS_64 0 -1.7241590937985623e-04
GC_11_65 b_11 NI_11 NS_65 0 2.6955932888297992e-05
GC_11_66 b_11 NI_11 NS_66 0 -7.4548020952796794e-05
GC_11_67 b_11 NI_11 NS_67 0 -2.3087067414518383e-05
GC_11_68 b_11 NI_11 NS_68 0 -8.4196444767580328e-05
GC_11_69 b_11 NI_11 NS_69 0 -2.3650398469350850e-05
GC_11_70 b_11 NI_11 NS_70 0 6.6120774689987138e-05
GC_11_71 b_11 NI_11 NS_71 0 -9.0195344052302503e-05
GC_11_72 b_11 NI_11 NS_72 0 -6.9243516545292386e-04
GC_11_73 b_11 NI_11 NS_73 0 -1.2485816604811515e-05
GC_11_74 b_11 NI_11 NS_74 0 -4.1085535300380027e-06
GC_11_75 b_11 NI_11 NS_75 0 -3.9465721502978128e-04
GC_11_76 b_11 NI_11 NS_76 0 -3.0741204990555362e-05
GC_11_77 b_11 NI_11 NS_77 0 -1.3312791490378983e-06
GC_11_78 b_11 NI_11 NS_78 0 4.3627742540086445e-07
GC_11_79 b_11 NI_11 NS_79 0 1.6509918587782237e-04
GC_11_80 b_11 NI_11 NS_80 0 -9.4789060487510918e-05
GC_11_81 b_11 NI_11 NS_81 0 -6.6463075017691510e-06
GC_11_82 b_11 NI_11 NS_82 0 -1.1071355172716636e-05
GC_11_83 b_11 NI_11 NS_83 0 7.2949670897624421e-07
GC_11_84 b_11 NI_11 NS_84 0 -8.3041486991790649e-07
GC_11_85 b_11 NI_11 NS_85 0 -2.1488601094022766e-07
GC_11_86 b_11 NI_11 NS_86 0 6.2332904511402137e-07
GC_11_87 b_11 NI_11 NS_87 0 -9.0268000838774915e-05
GC_11_88 b_11 NI_11 NS_88 0 -4.7819389251902389e-05
GC_11_89 b_11 NI_11 NS_89 0 -5.9553613092421420e-04
GC_11_90 b_11 NI_11 NS_90 0 9.6315189348237937e-05
GC_11_91 b_11 NI_11 NS_91 0 7.4891764805083889e-04
GC_11_92 b_11 NI_11 NS_92 0 -7.6481436721418652e-04
GC_11_93 b_11 NI_11 NS_93 0 3.9570991688048560e-04
GC_11_94 b_11 NI_11 NS_94 0 5.4605098011381407e-04
GC_11_95 b_11 NI_11 NS_95 0 -5.0914917058913914e-04
GC_11_96 b_11 NI_11 NS_96 0 -9.6590883566043730e-05
GC_11_97 b_11 NI_11 NS_97 0 1.0850139269758209e-03
GC_11_98 b_11 NI_11 NS_98 0 7.1873997540433253e-04
GC_11_99 b_11 NI_11 NS_99 0 -3.8689747566065641e-03
GC_11_100 b_11 NI_11 NS_100 0 -5.7242459219297451e-06
GC_11_101 b_11 NI_11 NS_101 0 5.7749955123540604e-04
GC_11_102 b_11 NI_11 NS_102 0 -4.5812355667414981e-04
GC_11_103 b_11 NI_11 NS_103 0 4.9505562911086555e-03
GC_11_104 b_11 NI_11 NS_104 0 -1.9110899412229548e-03
GC_11_105 b_11 NI_11 NS_105 0 2.4907722048023075e-04
GC_11_106 b_11 NI_11 NS_106 0 2.8215532031986571e-04
GC_11_107 b_11 NI_11 NS_107 0 -1.8134564187503868e-04
GC_11_108 b_11 NI_11 NS_108 0 1.2555367703311264e-03
GC_11_109 b_11 NI_11 NS_109 0 1.4635577729383469e-04
GC_11_110 b_11 NI_11 NS_110 0 -7.9921116520999822e-05
GC_11_111 b_11 NI_11 NS_111 0 1.5231733203705883e-04
GC_11_112 b_11 NI_11 NS_112 0 -6.5484773338806700e-05
GC_11_113 b_11 NI_11 NS_113 0 2.4317120255918722e-05
GC_11_114 b_11 NI_11 NS_114 0 8.2980927796277165e-05
GC_11_115 b_11 NI_11 NS_115 0 -3.1341482877728696e-03
GC_11_116 b_11 NI_11 NS_116 0 5.9087530955524263e-03
GC_11_117 b_11 NI_11 NS_117 0 2.1126459937742844e-06
GC_11_118 b_11 NI_11 NS_118 0 -1.1515540422665280e-05
GC_11_119 b_11 NI_11 NS_119 0 1.2415481698153619e-03
GC_11_120 b_11 NI_11 NS_120 0 -1.3121289261499606e-03
GC_11_121 b_11 NI_11 NS_121 0 -2.6295683721150993e-06
GC_11_122 b_11 NI_11 NS_122 0 7.2501522615996949e-07
GC_11_123 b_11 NI_11 NS_123 0 -9.4527347470653282e-05
GC_11_124 b_11 NI_11 NS_124 0 -1.5390036698441428e-03
GC_11_125 b_11 NI_11 NS_125 0 -1.0624980101825879e-05
GC_11_126 b_11 NI_11 NS_126 0 2.3213582458333377e-06
GC_11_127 b_11 NI_11 NS_127 0 -2.2320696414036981e-08
GC_11_128 b_11 NI_11 NS_128 0 4.5396607463796143e-07
GC_11_129 b_11 NI_11 NS_129 0 -2.7172502966045566e-07
GC_11_130 b_11 NI_11 NS_130 0 1.9128169238481216e-06
GC_11_131 b_11 NI_11 NS_131 0 -9.2710721303375886e-05
GC_11_132 b_11 NI_11 NS_132 0 -4.7248540666092702e-04
GC_11_133 b_11 NI_11 NS_133 0 1.2175543500142393e-02
GC_11_134 b_11 NI_11 NS_134 0 -4.6083429604602163e-05
GC_11_135 b_11 NI_11 NS_135 0 -6.2453566370166357e-04
GC_11_136 b_11 NI_11 NS_136 0 6.3789086989598587e-04
GC_11_137 b_11 NI_11 NS_137 0 -2.7049982031591161e-04
GC_11_138 b_11 NI_11 NS_138 0 -7.8978524657164081e-04
GC_11_139 b_11 NI_11 NS_139 0 -2.7800657455873801e-04
GC_11_140 b_11 NI_11 NS_140 0 -7.8678014251573698e-05
GC_11_141 b_11 NI_11 NS_141 0 5.5570752695911687e-04
GC_11_142 b_11 NI_11 NS_142 0 -1.0487176986489938e-04
GC_11_143 b_11 NI_11 NS_143 0 -4.1408773512406069e-04
GC_11_144 b_11 NI_11 NS_144 0 3.4470204586987263e-04
GC_11_145 b_11 NI_11 NS_145 0 8.5057662412298511e-05
GC_11_146 b_11 NI_11 NS_146 0 7.9836957022920072e-05
GC_11_147 b_11 NI_11 NS_147 0 -5.9875960170998887e-05
GC_11_148 b_11 NI_11 NS_148 0 8.3159683836512774e-04
GC_11_149 b_11 NI_11 NS_149 0 -1.0066004163839410e-04
GC_11_150 b_11 NI_11 NS_150 0 3.0280993752481032e-05
GC_11_151 b_11 NI_11 NS_151 0 -4.4908456593020454e-04
GC_11_152 b_11 NI_11 NS_152 0 -2.6213334927214514e-05
GC_11_153 b_11 NI_11 NS_153 0 2.3536341432113718e-05
GC_11_154 b_11 NI_11 NS_154 0 -4.8881025392956274e-05
GC_11_155 b_11 NI_11 NS_155 0 -2.3920214848039649e-05
GC_11_156 b_11 NI_11 NS_156 0 -9.2012627953800421e-05
GC_11_157 b_11 NI_11 NS_157 0 -2.0726269113469926e-05
GC_11_158 b_11 NI_11 NS_158 0 7.3624203123926884e-05
GC_11_159 b_11 NI_11 NS_159 0 2.1980646430524501e-04
GC_11_160 b_11 NI_11 NS_160 0 -5.5910333391176708e-04
GC_11_161 b_11 NI_11 NS_161 0 -1.4806914977460900e-05
GC_11_162 b_11 NI_11 NS_162 0 -5.3585934609506863e-06
GC_11_163 b_11 NI_11 NS_163 0 -4.5281730696261445e-04
GC_11_164 b_11 NI_11 NS_164 0 -6.8227078602587949e-05
GC_11_165 b_11 NI_11 NS_165 0 -7.1565924317990572e-07
GC_11_166 b_11 NI_11 NS_166 0 -4.9648836498395653e-07
GC_11_167 b_11 NI_11 NS_167 0 6.2426543879364331e-05
GC_11_168 b_11 NI_11 NS_168 0 -1.0001616021447374e-04
GC_11_169 b_11 NI_11 NS_169 0 -4.6421494788094875e-06
GC_11_170 b_11 NI_11 NS_170 0 -8.6256922945594454e-06
GC_11_171 b_11 NI_11 NS_171 0 7.1916189841873084e-07
GC_11_172 b_11 NI_11 NS_172 0 1.2656688409645950e-08
GC_11_173 b_11 NI_11 NS_173 0 -9.5193072737060160e-07
GC_11_174 b_11 NI_11 NS_174 0 -6.3026953828910334e-08
GC_11_175 b_11 NI_11 NS_175 0 -1.0272740019213592e-04
GC_11_176 b_11 NI_11 NS_176 0 -2.6090958644801927e-05
GC_11_177 b_11 NI_11 NS_177 0 4.8740243412646852e-03
GC_11_178 b_11 NI_11 NS_178 0 8.2133775933485549e-05
GC_11_179 b_11 NI_11 NS_179 0 1.2174357505626123e-03
GC_11_180 b_11 NI_11 NS_180 0 -2.8692723051302276e-04
GC_11_181 b_11 NI_11 NS_181 0 -6.2843474003024984e-04
GC_11_182 b_11 NI_11 NS_182 0 4.4929006328279668e-04
GC_11_183 b_11 NI_11 NS_183 0 -3.4540408579284017e-05
GC_11_184 b_11 NI_11 NS_184 0 -3.2219075219804813e-04
GC_11_185 b_11 NI_11 NS_185 0 8.3501548965939716e-04
GC_11_186 b_11 NI_11 NS_186 0 6.1005908877862500e-04
GC_11_187 b_11 NI_11 NS_187 0 -2.5776192570633101e-03
GC_11_188 b_11 NI_11 NS_188 0 -1.6176696481230424e-03
GC_11_189 b_11 NI_11 NS_189 0 5.6361992128348473e-04
GC_11_190 b_11 NI_11 NS_190 0 -4.2454792676645270e-04
GC_11_191 b_11 NI_11 NS_191 0 4.8135801902857598e-03
GC_11_192 b_11 NI_11 NS_192 0 2.5417996989332971e-04
GC_11_193 b_11 NI_11 NS_193 0 2.6020828746895760e-04
GC_11_194 b_11 NI_11 NS_194 0 2.9165246152061084e-04
GC_11_195 b_11 NI_11 NS_195 0 -2.1076434917483122e-04
GC_11_196 b_11 NI_11 NS_196 0 2.0647333764688973e-03
GC_11_197 b_11 NI_11 NS_197 0 3.3049505128633362e-04
GC_11_198 b_11 NI_11 NS_198 0 -2.8507368560049440e-04
GC_11_199 b_11 NI_11 NS_199 0 1.6354465160765803e-04
GC_11_200 b_11 NI_11 NS_200 0 -3.4625689173422467e-05
GC_11_201 b_11 NI_11 NS_201 0 2.3300170921067410e-05
GC_11_202 b_11 NI_11 NS_202 0 8.0327766768051821e-05
GC_11_203 b_11 NI_11 NS_203 0 -5.3876956411418537e-03
GC_11_204 b_11 NI_11 NS_204 0 4.4054534283433167e-03
GC_11_205 b_11 NI_11 NS_205 0 7.3753179783290724e-06
GC_11_206 b_11 NI_11 NS_206 0 -8.5812508502474934e-06
GC_11_207 b_11 NI_11 NS_207 0 1.5140669367630076e-03
GC_11_208 b_11 NI_11 NS_208 0 -6.7750671413527969e-04
GC_11_209 b_11 NI_11 NS_209 0 -1.6866880353627764e-07
GC_11_210 b_11 NI_11 NS_210 0 2.8600671417588014e-06
GC_11_211 b_11 NI_11 NS_211 0 -9.7868658587895623e-05
GC_11_212 b_11 NI_11 NS_212 0 -1.8748906601420668e-03
GC_11_213 b_11 NI_11 NS_213 0 -1.3227272428558525e-05
GC_11_214 b_11 NI_11 NS_214 0 2.6824782583262397e-06
GC_11_215 b_11 NI_11 NS_215 0 4.9111115760074644e-07
GC_11_216 b_11 NI_11 NS_216 0 -4.2338703004343962e-07
GC_11_217 b_11 NI_11 NS_217 0 1.0530280975533955e-06
GC_11_218 b_11 NI_11 NS_218 0 2.3016437856605078e-06
GC_11_219 b_11 NI_11 NS_219 0 -2.0012229927153625e-05
GC_11_220 b_11 NI_11 NS_220 0 -5.5318162044093173e-04
GC_11_221 b_11 NI_11 NS_221 0 -4.2622168612154185e-03
GC_11_222 b_11 NI_11 NS_222 0 -1.8702595843060220e-05
GC_11_223 b_11 NI_11 NS_223 0 -1.2972508191197269e-03
GC_11_224 b_11 NI_11 NS_224 0 2.2387696940363291e-04
GC_11_225 b_11 NI_11 NS_225 0 6.0737820138261295e-04
GC_11_226 b_11 NI_11 NS_226 0 -1.2187294176990034e-03
GC_11_227 b_11 NI_11 NS_227 0 -2.8443767277868362e-05
GC_11_228 b_11 NI_11 NS_228 0 1.5685281223579988e-04
GC_11_229 b_11 NI_11 NS_229 0 6.8039264115834033e-04
GC_11_230 b_11 NI_11 NS_230 0 -1.4008572729662166e-04
GC_11_231 b_11 NI_11 NS_231 0 -2.4018327499005922e-04
GC_11_232 b_11 NI_11 NS_232 0 -1.0944691643615110e-03
GC_11_233 b_11 NI_11 NS_233 0 1.2252475684100260e-04
GC_11_234 b_11 NI_11 NS_234 0 9.3166855023343179e-05
GC_11_235 b_11 NI_11 NS_235 0 9.6116463623624113e-04
GC_11_236 b_11 NI_11 NS_236 0 1.2705264054232595e-03
GC_11_237 b_11 NI_11 NS_237 0 -1.2482948935002873e-04
GC_11_238 b_11 NI_11 NS_238 0 4.8405549862681478e-05
GC_11_239 b_11 NI_11 NS_239 0 -2.5231909943176939e-04
GC_11_240 b_11 NI_11 NS_240 0 -5.5638004725413174e-05
GC_11_241 b_11 NI_11 NS_241 0 -1.2047343991792150e-05
GC_11_242 b_11 NI_11 NS_242 0 4.2813796517225872e-05
GC_11_243 b_11 NI_11 NS_243 0 -1.9209038448847786e-05
GC_11_244 b_11 NI_11 NS_244 0 -1.0859384247395714e-04
GC_11_245 b_11 NI_11 NS_245 0 -2.1956983040759900e-05
GC_11_246 b_11 NI_11 NS_246 0 1.0095892929455341e-04
GC_11_247 b_11 NI_11 NS_247 0 1.0425907919162573e-03
GC_11_248 b_11 NI_11 NS_248 0 7.4111169176200719e-04
GC_11_249 b_11 NI_11 NS_249 0 -1.8694169599199215e-05
GC_11_250 b_11 NI_11 NS_250 0 -6.7359230752629141e-06
GC_11_251 b_11 NI_11 NS_251 0 -3.0562213693880049e-04
GC_11_252 b_11 NI_11 NS_252 0 -5.2287179527942484e-04
GC_11_253 b_11 NI_11 NS_253 0 -1.7539255782719392e-06
GC_11_254 b_11 NI_11 NS_254 0 -1.4693677281556255e-06
GC_11_255 b_11 NI_11 NS_255 0 -3.9879059937983236e-05
GC_11_256 b_11 NI_11 NS_256 0 -1.4014732454458150e-04
GC_11_257 b_11 NI_11 NS_257 0 -8.1771730057211415e-06
GC_11_258 b_11 NI_11 NS_258 0 -1.1988129325798755e-05
GC_11_259 b_11 NI_11 NS_259 0 1.6414955001313328e-07
GC_11_260 b_11 NI_11 NS_260 0 -5.1072690273237900e-07
GC_11_261 b_11 NI_11 NS_261 0 -4.9584215512322265e-07
GC_11_262 b_11 NI_11 NS_262 0 -9.0816035651091780e-07
GC_11_263 b_11 NI_11 NS_263 0 -1.9937568316929214e-04
GC_11_264 b_11 NI_11 NS_264 0 -7.4310487947378369e-05
GC_11_265 b_11 NI_11 NS_265 0 -2.1746756487583244e-02
GC_11_266 b_11 NI_11 NS_266 0 5.8937899911553711e-05
GC_11_267 b_11 NI_11 NS_267 0 1.0843242476627274e-03
GC_11_268 b_11 NI_11 NS_268 0 9.6537558228928101e-04
GC_11_269 b_11 NI_11 NS_269 0 -1.0198865005901241e-03
GC_11_270 b_11 NI_11 NS_270 0 -2.3849025651063549e-03
GC_11_271 b_11 NI_11 NS_271 0 1.4595521127601979e-04
GC_11_272 b_11 NI_11 NS_272 0 2.5884633141142502e-04
GC_11_273 b_11 NI_11 NS_273 0 8.4426091526746837e-04
GC_11_274 b_11 NI_11 NS_274 0 6.7751307324535794e-04
GC_11_275 b_11 NI_11 NS_275 0 -2.4390665904233612e-04
GC_11_276 b_11 NI_11 NS_276 0 -2.0975094875629210e-03
GC_11_277 b_11 NI_11 NS_277 0 4.5037889464928931e-04
GC_11_278 b_11 NI_11 NS_278 0 -1.9869603243294646e-04
GC_11_279 b_11 NI_11 NS_279 0 3.5419877998135165e-03
GC_11_280 b_11 NI_11 NS_280 0 -1.3881278340416091e-03
GC_11_281 b_11 NI_11 NS_281 0 1.5488187443168076e-04
GC_11_282 b_11 NI_11 NS_282 0 2.3487517886360205e-04
GC_11_283 b_11 NI_11 NS_283 0 6.6774675186744129e-06
GC_11_284 b_11 NI_11 NS_284 0 1.7467335403790675e-03
GC_11_285 b_11 NI_11 NS_285 0 4.4000232227352172e-04
GC_11_286 b_11 NI_11 NS_286 0 -9.5748361049160667e-05
GC_11_287 b_11 NI_11 NS_287 0 1.3346714377869388e-04
GC_11_288 b_11 NI_11 NS_288 0 -8.4655146342736806e-06
GC_11_289 b_11 NI_11 NS_289 0 2.9929389937720576e-05
GC_11_290 b_11 NI_11 NS_290 0 4.9975086170690512e-05
GC_11_291 b_11 NI_11 NS_291 0 -1.4185634006509702e-03
GC_11_292 b_11 NI_11 NS_292 0 4.3874626584628025e-03
GC_11_293 b_11 NI_11 NS_293 0 2.7557404667068856e-06
GC_11_294 b_11 NI_11 NS_294 0 -1.0689923345412538e-05
GC_11_295 b_11 NI_11 NS_295 0 1.2492459766449387e-03
GC_11_296 b_11 NI_11 NS_296 0 -1.2779703735278562e-03
GC_11_297 b_11 NI_11 NS_297 0 -2.2594999782985963e-06
GC_11_298 b_11 NI_11 NS_298 0 6.3091793581868139e-07
GC_11_299 b_11 NI_11 NS_299 0 -2.3206754675861256e-04
GC_11_300 b_11 NI_11 NS_300 0 -6.1637128574562193e-04
GC_11_301 b_11 NI_11 NS_301 0 -4.3786769062957034e-06
GC_11_302 b_11 NI_11 NS_302 0 2.9645673111996195e-06
GC_11_303 b_11 NI_11 NS_303 0 -4.9355590015686620e-07
GC_11_304 b_11 NI_11 NS_304 0 9.8927474189929674e-07
GC_11_305 b_11 NI_11 NS_305 0 -6.7785015231702709e-07
GC_11_306 b_11 NI_11 NS_306 0 2.1152220007887991e-07
GC_11_307 b_11 NI_11 NS_307 0 -8.3278584178038664e-05
GC_11_308 b_11 NI_11 NS_308 0 -3.2379209761565790e-04
GC_11_309 b_11 NI_11 NS_309 0 3.6983307955014500e-03
GC_11_310 b_11 NI_11 NS_310 0 3.9376601175259182e-05
GC_11_311 b_11 NI_11 NS_311 0 -1.7988795077156980e-03
GC_11_312 b_11 NI_11 NS_312 0 -1.0939128926970075e-03
GC_11_313 b_11 NI_11 NS_313 0 1.4015306842828765e-03
GC_11_314 b_11 NI_11 NS_314 0 7.0587049617706855e-04
GC_11_315 b_11 NI_11 NS_315 0 -2.2953689030297298e-05
GC_11_316 b_11 NI_11 NS_316 0 1.1614350910287452e-04
GC_11_317 b_11 NI_11 NS_317 0 4.0637789568130720e-04
GC_11_318 b_11 NI_11 NS_318 0 3.1642458108544358e-05
GC_11_319 b_11 NI_11 NS_319 0 6.1325648665298013e-04
GC_11_320 b_11 NI_11 NS_320 0 -1.3287104762564226e-03
GC_11_321 b_11 NI_11 NS_321 0 4.1404832742828855e-05
GC_11_322 b_11 NI_11 NS_322 0 1.2227939957896292e-04
GC_11_323 b_11 NI_11 NS_323 0 5.0954433542250379e-06
GC_11_324 b_11 NI_11 NS_324 0 6.8254233729813274e-04
GC_11_325 b_11 NI_11 NS_325 0 -8.0991991918249629e-05
GC_11_326 b_11 NI_11 NS_326 0 2.6628114776831065e-05
GC_11_327 b_11 NI_11 NS_327 0 -1.9810162678146062e-04
GC_11_328 b_11 NI_11 NS_328 0 2.6959461381573300e-04
GC_11_329 b_11 NI_11 NS_329 0 -5.4364225212232059e-05
GC_11_330 b_11 NI_11 NS_330 0 1.3713015738887969e-04
GC_11_331 b_11 NI_11 NS_331 0 -1.8322208197344000e-05
GC_11_332 b_11 NI_11 NS_332 0 -5.5537144304284966e-05
GC_11_333 b_11 NI_11 NS_333 0 -1.3234449291475681e-05
GC_11_334 b_11 NI_11 NS_334 0 6.2432784432787526e-05
GC_11_335 b_11 NI_11 NS_335 0 2.7168476546137680e-04
GC_11_336 b_11 NI_11 NS_336 0 5.1435504266352699e-04
GC_11_337 b_11 NI_11 NS_337 0 -9.9147809363127701e-06
GC_11_338 b_11 NI_11 NS_338 0 -2.7125789590891232e-06
GC_11_339 b_11 NI_11 NS_339 0 -9.8472937423196564e-05
GC_11_340 b_11 NI_11 NS_340 0 -7.1571949641039385e-05
GC_11_341 b_11 NI_11 NS_341 0 -1.3734911868987022e-06
GC_11_342 b_11 NI_11 NS_342 0 -8.0815576055735517e-07
GC_11_343 b_11 NI_11 NS_343 0 -6.0327746684209038e-05
GC_11_344 b_11 NI_11 NS_344 0 -5.7714251067674629e-05
GC_11_345 b_11 NI_11 NS_345 0 -2.8623358233340280e-06
GC_11_346 b_11 NI_11 NS_346 0 -5.3798795699797036e-06
GC_11_347 b_11 NI_11 NS_347 0 1.3944909266611797e-07
GC_11_348 b_11 NI_11 NS_348 0 -5.4613465504597631e-08
GC_11_349 b_11 NI_11 NS_349 0 -3.7581453712602672e-07
GC_11_350 b_11 NI_11 NS_350 0 -8.1654791606260728e-07
GC_11_351 b_11 NI_11 NS_351 0 -9.0194584984776573e-05
GC_11_352 b_11 NI_11 NS_352 0 -3.6865693209927279e-05
GC_11_353 b_11 NI_11 NS_353 0 -7.1368608618871720e-03
GC_11_354 b_11 NI_11 NS_354 0 1.6911409838723812e-05
GC_11_355 b_11 NI_11 NS_355 0 4.9589846136544298e-03
GC_11_356 b_11 NI_11 NS_356 0 4.3009851005010565e-03
GC_11_357 b_11 NI_11 NS_357 0 -4.8726242306839068e-03
GC_11_358 b_11 NI_11 NS_358 0 -5.0308499535476172e-03
GC_11_359 b_11 NI_11 NS_359 0 -6.8510161897372007e-04
GC_11_360 b_11 NI_11 NS_360 0 6.7883526962910141e-04
GC_11_361 b_11 NI_11 NS_361 0 1.7789404043676528e-03
GC_11_362 b_11 NI_11 NS_362 0 5.1569106671660028e-03
GC_11_363 b_11 NI_11 NS_363 0 -3.0496667160052394e-03
GC_11_364 b_11 NI_11 NS_364 0 -1.5564734572486841e-03
GC_11_365 b_11 NI_11 NS_365 0 9.8324904594626942e-04
GC_11_366 b_11 NI_11 NS_366 0 1.8005064269697242e-04
GC_11_367 b_11 NI_11 NS_367 0 -3.3298236193101023e-03
GC_11_368 b_11 NI_11 NS_368 0 -3.0004590503988661e-03
GC_11_369 b_11 NI_11 NS_369 0 -4.5982348553156081e-06
GC_11_370 b_11 NI_11 NS_370 0 1.6643701797450461e-04
GC_11_371 b_11 NI_11 NS_371 0 -1.7248145321240554e-03
GC_11_372 b_11 NI_11 NS_372 0 -2.5695238669855686e-03
GC_11_373 b_11 NI_11 NS_373 0 -4.3288848922389819e-04
GC_11_374 b_11 NI_11 NS_374 0 4.1891790233515813e-04
GC_11_375 b_11 NI_11 NS_375 0 2.1078437320487298e-04
GC_11_376 b_11 NI_11 NS_376 0 -7.3375779826941108e-05
GC_11_377 b_11 NI_11 NS_377 0 1.7773460079401569e-05
GC_11_378 b_11 NI_11 NS_378 0 -8.9595572022739843e-05
GC_11_379 b_11 NI_11 NS_379 0 7.9792399368521193e-03
GC_11_380 b_11 NI_11 NS_380 0 4.4950600663542454e-03
GC_11_381 b_11 NI_11 NS_381 0 -1.6110559709277877e-05
GC_11_382 b_11 NI_11 NS_382 0 -1.3105727795788610e-05
GC_11_383 b_11 NI_11 NS_383 0 8.6073305154012669e-04
GC_11_384 b_11 NI_11 NS_384 0 -4.2071176951978704e-03
GC_11_385 b_11 NI_11 NS_385 0 -2.3354229614930904e-06
GC_11_386 b_11 NI_11 NS_386 0 -1.6822606717712558e-05
GC_11_387 b_11 NI_11 NS_387 0 3.4135262761920797e-04
GC_11_388 b_11 NI_11 NS_388 0 1.2274243238206970e-03
GC_11_389 b_11 NI_11 NS_389 0 2.1127925244411042e-05
GC_11_390 b_11 NI_11 NS_390 0 1.1437367674626053e-05
GC_11_391 b_11 NI_11 NS_391 0 -5.2955422656063348e-07
GC_11_392 b_11 NI_11 NS_392 0 6.3789583715842360e-06
GC_11_393 b_11 NI_11 NS_393 0 -3.5556222103709464e-06
GC_11_394 b_11 NI_11 NS_394 0 -3.5517433909585515e-06
GC_11_395 b_11 NI_11 NS_395 0 -8.3306625083272637e-05
GC_11_396 b_11 NI_11 NS_396 0 1.0471443468748322e-04
GC_11_397 b_11 NI_11 NS_397 0 6.4982097491443569e-02
GC_11_398 b_11 NI_11 NS_398 0 -7.9954499788883850e-05
GC_11_399 b_11 NI_11 NS_399 0 -6.4095691830151728e-03
GC_11_400 b_11 NI_11 NS_400 0 -2.5862470334039930e-03
GC_11_401 b_11 NI_11 NS_401 0 4.2953376586496199e-03
GC_11_402 b_11 NI_11 NS_402 0 2.5496217089425572e-03
GC_11_403 b_11 NI_11 NS_403 0 -5.7986871117690012e-04
GC_11_404 b_11 NI_11 NS_404 0 -1.6472860870375648e-04
GC_11_405 b_11 NI_11 NS_405 0 1.5068227882573957e-03
GC_11_406 b_11 NI_11 NS_406 0 1.4953588887618150e-03
GC_11_407 b_11 NI_11 NS_407 0 -3.7977882159983813e-04
GC_11_408 b_11 NI_11 NS_408 0 -3.5978180216083211e-04
GC_11_409 b_11 NI_11 NS_409 0 -3.2659321820648493e-05
GC_11_410 b_11 NI_11 NS_410 0 7.4286695376632510e-05
GC_11_411 b_11 NI_11 NS_411 0 -4.0075330788390384e-03
GC_11_412 b_11 NI_11 NS_412 0 1.2348966680736442e-03
GC_11_413 b_11 NI_11 NS_413 0 -9.1324357045341015e-05
GC_11_414 b_11 NI_11 NS_414 0 -6.2364289763961579e-05
GC_11_415 b_11 NI_11 NS_415 0 -3.3852922123323091e-04
GC_11_416 b_11 NI_11 NS_416 0 8.5603857272232350e-04
GC_11_417 b_11 NI_11 NS_417 0 2.4651681908877381e-04
GC_11_418 b_11 NI_11 NS_418 0 1.0827517630279023e-04
GC_11_419 b_11 NI_11 NS_419 0 -3.1782974453268336e-05
GC_11_420 b_11 NI_11 NS_420 0 -6.4690402410667443e-05
GC_11_421 b_11 NI_11 NS_421 0 -6.4035102107093457e-05
GC_11_422 b_11 NI_11 NS_422 0 9.1653122160889868e-05
GC_11_423 b_11 NI_11 NS_423 0 -2.6102522625645885e-03
GC_11_424 b_11 NI_11 NS_424 0 -4.1099696300817001e-03
GC_11_425 b_11 NI_11 NS_425 0 4.9953670321646839e-06
GC_11_426 b_11 NI_11 NS_426 0 3.7688567737097009e-05
GC_11_427 b_11 NI_11 NS_427 0 -8.1465011929632259e-04
GC_11_428 b_11 NI_11 NS_428 0 2.1208816921077442e-03
GC_11_429 b_11 NI_11 NS_429 0 -3.3555708979129820e-06
GC_11_430 b_11 NI_11 NS_430 0 8.1496787470558129e-06
GC_11_431 b_11 NI_11 NS_431 0 9.0173225533300109e-04
GC_11_432 b_11 NI_11 NS_432 0 -2.9734244350858660e-04
GC_11_433 b_11 NI_11 NS_433 0 -8.8935394871977257e-06
GC_11_434 b_11 NI_11 NS_434 0 -1.0945848085690160e-05
GC_11_435 b_11 NI_11 NS_435 0 3.1108562995193253e-06
GC_11_436 b_11 NI_11 NS_436 0 -1.3430618942046999e-06
GC_11_437 b_11 NI_11 NS_437 0 1.9687573313011719e-06
GC_11_438 b_11 NI_11 NS_438 0 -4.8428928971553327e-07
GC_11_439 b_11 NI_11 NS_439 0 9.6562432095580970e-05
GC_11_440 b_11 NI_11 NS_440 0 -1.1241070116390910e-04
GC_11_441 b_11 NI_11 NS_441 0 -7.2251377908674377e-02
GC_11_442 b_11 NI_11 NS_442 0 9.5756757326165842e-03
GC_11_443 b_11 NI_11 NS_443 0 3.3337563193697648e-03
GC_11_444 b_11 NI_11 NS_444 0 6.0058542265168831e-03
GC_11_445 b_11 NI_11 NS_445 0 1.1330062064927321e-02
GC_11_446 b_11 NI_11 NS_446 0 -2.0684838351827479e-03
GC_11_447 b_11 NI_11 NS_447 0 1.9754488554744954e-03
GC_11_448 b_11 NI_11 NS_448 0 1.0437980053288366e-03
GC_11_449 b_11 NI_11 NS_449 0 5.4869452473285478e-04
GC_11_450 b_11 NI_11 NS_450 0 3.2297975174149607e-03
GC_11_451 b_11 NI_11 NS_451 0 2.8064383175218930e-03
GC_11_452 b_11 NI_11 NS_452 0 1.6738031459691155e-03
GC_11_453 b_11 NI_11 NS_453 0 5.9593247742983240e-04
GC_11_454 b_11 NI_11 NS_454 0 2.4187453574720525e-04
GC_11_455 b_11 NI_11 NS_455 0 6.9390190342620188e-03
GC_11_456 b_11 NI_11 NS_456 0 1.4514386354166613e-03
GC_11_457 b_11 NI_11 NS_457 0 1.3064157357756768e-05
GC_11_458 b_11 NI_11 NS_458 0 1.8521429556360989e-04
GC_11_459 b_11 NI_11 NS_459 0 -3.1409023937183545e-04
GC_11_460 b_11 NI_11 NS_460 0 -2.7498543871318855e-04
GC_11_461 b_11 NI_11 NS_461 0 -8.3027304562673142e-04
GC_11_462 b_11 NI_11 NS_462 0 1.1721834142224093e-04
GC_11_463 b_11 NI_11 NS_463 0 1.7281715350511741e-04
GC_11_464 b_11 NI_11 NS_464 0 1.3729886454881147e-05
GC_11_465 b_11 NI_11 NS_465 0 5.2815088455860287e-05
GC_11_466 b_11 NI_11 NS_466 0 -3.6563034177065971e-05
GC_11_467 b_11 NI_11 NS_467 0 1.4385765147950356e-03
GC_11_468 b_11 NI_11 NS_468 0 1.2721758072665448e-02
GC_11_469 b_11 NI_11 NS_469 0 -3.2945308631773206e-06
GC_11_470 b_11 NI_11 NS_470 0 -2.1904043972166083e-05
GC_11_471 b_11 NI_11 NS_471 0 3.3840670438723829e-03
GC_11_472 b_11 NI_11 NS_472 0 -3.5850565357352124e-03
GC_11_473 b_11 NI_11 NS_473 0 3.7686121305685306e-06
GC_11_474 b_11 NI_11 NS_474 0 -2.2577459892852937e-05
GC_11_475 b_11 NI_11 NS_475 0 -2.1631867099908084e-03
GC_11_476 b_11 NI_11 NS_476 0 5.9560949651113666e-04
GC_11_477 b_11 NI_11 NS_477 0 1.9281288156849463e-05
GC_11_478 b_11 NI_11 NS_478 0 3.1987069010540172e-05
GC_11_479 b_11 NI_11 NS_479 0 -6.0159578382041318e-06
GC_11_480 b_11 NI_11 NS_480 0 4.3104012577967023e-06
GC_11_481 b_11 NI_11 NS_481 0 -1.3198435273751016e-06
GC_11_482 b_11 NI_11 NS_482 0 -1.0843448799993137e-05
GC_11_483 b_11 NI_11 NS_483 0 -3.5179520678514761e-04
GC_11_484 b_11 NI_11 NS_484 0 -1.5087778121561786e-04
GC_11_485 b_11 NI_11 NS_485 0 -4.2708164812436640e-04
GC_11_486 b_11 NI_11 NS_486 0 1.0643826866946010e-02
GC_11_487 b_11 NI_11 NS_487 0 -6.8704980320695294e-03
GC_11_488 b_11 NI_11 NS_488 0 -5.0120136606930732e-03
GC_11_489 b_11 NI_11 NS_489 0 -1.1447835455600174e-02
GC_11_490 b_11 NI_11 NS_490 0 1.0735562467553417e-03
GC_11_491 b_11 NI_11 NS_491 0 -7.3720616838292513e-06
GC_11_492 b_11 NI_11 NS_492 0 4.4728455451812477e-04
GC_11_493 b_11 NI_11 NS_493 0 1.2785105033416265e-03
GC_11_494 b_11 NI_11 NS_494 0 1.3899937933259741e-03
GC_11_495 b_11 NI_11 NS_495 0 3.2307851457087284e-03
GC_11_496 b_11 NI_11 NS_496 0 -1.4843900157391293e-03
GC_11_497 b_11 NI_11 NS_497 0 -1.3201530190827158e-06
GC_11_498 b_11 NI_11 NS_498 0 1.8361673199347180e-04
GC_11_499 b_11 NI_11 NS_499 0 3.0586200534853968e-03
GC_11_500 b_11 NI_11 NS_500 0 -1.0036044362863766e-03
GC_11_501 b_11 NI_11 NS_501 0 -3.6793167563891336e-05
GC_11_502 b_11 NI_11 NS_502 0 -8.9992844759134675e-06
GC_11_503 b_11 NI_11 NS_503 0 2.2235484115564079e-04
GC_11_504 b_11 NI_11 NS_504 0 2.0825856963776834e-04
GC_11_505 b_11 NI_11 NS_505 0 -9.1313663225325446e-05
GC_11_506 b_11 NI_11 NS_506 0 -1.7871925303208364e-07
GC_11_507 b_11 NI_11 NS_507 0 1.0552693715349388e-06
GC_11_508 b_11 NI_11 NS_508 0 -3.6284964868518227e-05
GC_11_509 b_11 NI_11 NS_509 0 -2.6579763599819773e-05
GC_11_510 b_11 NI_11 NS_510 0 4.9701355719157042e-05
GC_11_511 b_11 NI_11 NS_511 0 -5.4520826562979218e-04
GC_11_512 b_11 NI_11 NS_512 0 -6.7363334604601550e-04
GC_11_513 b_11 NI_11 NS_513 0 -1.5672381782841033e-06
GC_11_514 b_11 NI_11 NS_514 0 1.4085058368062036e-05
GC_11_515 b_11 NI_11 NS_515 0 -3.0121106138439286e-04
GC_11_516 b_11 NI_11 NS_516 0 5.2550430816867915e-04
GC_11_517 b_11 NI_11 NS_517 0 -1.4415676557714632e-06
GC_11_518 b_11 NI_11 NS_518 0 -7.4825902998341545e-07
GC_11_519 b_11 NI_11 NS_519 0 -5.8512334563309224e-06
GC_11_520 b_11 NI_11 NS_520 0 -1.2587912898982521e-04
GC_11_521 b_11 NI_11 NS_521 0 -7.1245039433874950e-09
GC_11_522 b_11 NI_11 NS_522 0 -1.6376168560634635e-06
GC_11_523 b_11 NI_11 NS_523 0 6.1888673428340872e-07
GC_11_524 b_11 NI_11 NS_524 0 8.9686813013682783e-08
GC_11_525 b_11 NI_11 NS_525 0 4.5856719546742315e-09
GC_11_526 b_11 NI_11 NS_526 0 -1.6803763436704656e-06
GC_11_527 b_11 NI_11 NS_527 0 -2.9751339531045461e-05
GC_11_528 b_11 NI_11 NS_528 0 -4.9532285568089859e-05
GD_11_1 b_11 NI_11 NA_1 0 1.6877265313241325e-03
GD_11_2 b_11 NI_11 NA_2 0 -1.4025804121701650e-02
GD_11_3 b_11 NI_11 NA_3 0 -3.1623102731116459e-03
GD_11_4 b_11 NI_11 NA_4 0 -1.1170994029427310e-02
GD_11_5 b_11 NI_11 NA_5 0 -8.5027406838459225e-03
GD_11_6 b_11 NI_11 NA_6 0 3.3959406975185690e-03
GD_11_7 b_11 NI_11 NA_7 0 1.5477922166692991e-02
GD_11_8 b_11 NI_11 NA_8 0 -5.9634419064440326e-03
GD_11_9 b_11 NI_11 NA_9 0 4.8325391677784234e-03
GD_11_10 b_11 NI_11 NA_10 0 -6.6001193440231920e-02
GD_11_11 b_11 NI_11 NA_11 0 -1.0471486148806908e-01
GD_11_12 b_11 NI_11 NA_12 0 2.2570012411050732e-03
*
* Port 12
VI_12 a_12 NI_12 0
RI_12 NI_12 b_12 5.0000000000000000e+01
GC_12_1 b_12 NI_12 NS_1 0 1.6296100570072559e-02
GC_12_2 b_12 NI_12 NS_2 0 -4.1214930758902265e-05
GC_12_3 b_12 NI_12 NS_3 0 -1.2942858891053103e-04
GC_12_4 b_12 NI_12 NS_4 0 5.5166694214806239e-04
GC_12_5 b_12 NI_12 NS_5 0 -4.9372937054849471e-04
GC_12_6 b_12 NI_12 NS_6 0 -2.2001000782951736e-04
GC_12_7 b_12 NI_12 NS_7 0 -2.9651335720224943e-04
GC_12_8 b_12 NI_12 NS_8 0 -2.6444772321876337e-04
GC_12_9 b_12 NI_12 NS_9 0 3.1164403721793731e-04
GC_12_10 b_12 NI_12 NS_10 0 -1.7842808434656532e-05
GC_12_11 b_12 NI_12 NS_11 0 -2.9608771829533695e-04
GC_12_12 b_12 NI_12 NS_12 0 1.0793521325067426e-03
GC_12_13 b_12 NI_12 NS_13 0 6.5206642068206693e-05
GC_12_14 b_12 NI_12 NS_14 0 3.2526449929247092e-05
GC_12_15 b_12 NI_12 NS_15 0 -8.6557103877793213e-04
GC_12_16 b_12 NI_12 NS_16 0 3.8880528827430302e-04
GC_12_17 b_12 NI_12 NS_17 0 -7.9355488105041874e-05
GC_12_18 b_12 NI_12 NS_18 0 1.9610232944851709e-05
GC_12_19 b_12 NI_12 NS_19 0 -3.6832062913798205e-04
GC_12_20 b_12 NI_12 NS_20 0 -1.0776770032875378e-04
GC_12_21 b_12 NI_12 NS_21 0 3.4176600057025599e-05
GC_12_22 b_12 NI_12 NS_22 0 -1.0181431009186025e-04
GC_12_23 b_12 NI_12 NS_23 0 -1.9440086224067240e-05
GC_12_24 b_12 NI_12 NS_24 0 -7.0944857015557361e-05
GC_12_25 b_12 NI_12 NS_25 0 -1.2758381870270887e-05
GC_12_26 b_12 NI_12 NS_26 0 5.8006996865788240e-05
GC_12_27 b_12 NI_12 NS_27 0 -2.6139701429820749e-04
GC_12_28 b_12 NI_12 NS_28 0 -8.9675752220006540e-04
GC_12_29 b_12 NI_12 NS_29 0 -1.2869092278433975e-05
GC_12_30 b_12 NI_12 NS_30 0 -1.3641917638963077e-06
GC_12_31 b_12 NI_12 NS_31 0 -3.7957515311054524e-04
GC_12_32 b_12 NI_12 NS_32 0 1.4095067300021809e-04
GC_12_33 b_12 NI_12 NS_33 0 -7.3520098428275446e-08
GC_12_34 b_12 NI_12 NS_34 0 1.2107210600389248e-06
GC_12_35 b_12 NI_12 NS_35 0 1.2449040020716455e-04
GC_12_36 b_12 NI_12 NS_36 0 -1.0300443839756642e-04
GC_12_37 b_12 NI_12 NS_37 0 -4.9067850404748891e-06
GC_12_38 b_12 NI_12 NS_38 0 -6.2409973308884862e-06
GC_12_39 b_12 NI_12 NS_39 0 -2.0865144618302342e-07
GC_12_40 b_12 NI_12 NS_40 0 4.1086273013360840e-07
GC_12_41 b_12 NI_12 NS_41 0 1.0466101575983042e-06
GC_12_42 b_12 NI_12 NS_42 0 -1.1962861370387606e-07
GC_12_43 b_12 NI_12 NS_43 0 -7.0941532996994655e-05
GC_12_44 b_12 NI_12 NS_44 0 -2.8922823969945004e-05
GC_12_45 b_12 NI_12 NS_45 0 3.5220261812522237e-04
GC_12_46 b_12 NI_12 NS_46 0 -8.7579771986352259e-07
GC_12_47 b_12 NI_12 NS_47 0 2.2948473627564558e-05
GC_12_48 b_12 NI_12 NS_48 0 -4.6155101834590204e-04
GC_12_49 b_12 NI_12 NS_49 0 4.6433028186661197e-04
GC_12_50 b_12 NI_12 NS_50 0 1.2267897827002687e-04
GC_12_51 b_12 NI_12 NS_51 0 -1.0891672106660176e-04
GC_12_52 b_12 NI_12 NS_52 0 4.1163610797680117e-04
GC_12_53 b_12 NI_12 NS_53 0 2.6657530170384698e-04
GC_12_54 b_12 NI_12 NS_54 0 -8.3139522775878879e-05
GC_12_55 b_12 NI_12 NS_55 0 3.1627686207135255e-04
GC_12_56 b_12 NI_12 NS_56 0 2.9248871819634960e-04
GC_12_57 b_12 NI_12 NS_57 0 6.4677128967219958e-06
GC_12_58 b_12 NI_12 NS_58 0 8.6588215480677794e-06
GC_12_59 b_12 NI_12 NS_59 0 7.4413225133270554e-05
GC_12_60 b_12 NI_12 NS_60 0 -2.1320762982845256e-04
GC_12_61 b_12 NI_12 NS_61 0 1.1842537556772910e-05
GC_12_62 b_12 NI_12 NS_62 0 -2.6766013677686951e-05
GC_12_63 b_12 NI_12 NS_63 0 3.7253633749675474e-04
GC_12_64 b_12 NI_12 NS_64 0 -1.5572727543174667e-04
GC_12_65 b_12 NI_12 NS_65 0 -7.4389146644681257e-05
GC_12_66 b_12 NI_12 NS_66 0 -1.3788867618173619e-04
GC_12_67 b_12 NI_12 NS_67 0 3.4360858481865310e-06
GC_12_68 b_12 NI_12 NS_68 0 -1.3216125934832868e-05
GC_12_69 b_12 NI_12 NS_69 0 -2.5993779586443113e-05
GC_12_70 b_12 NI_12 NS_70 0 -9.7663551508892377e-05
GC_12_71 b_12 NI_12 NS_71 0 -2.1904077921484446e-03
GC_12_72 b_12 NI_12 NS_72 0 2.0228372329646272e-03
GC_12_73 b_12 NI_12 NS_73 0 7.2443997939307334e-06
GC_12_74 b_12 NI_12 NS_74 0 4.9913088756208761e-06
GC_12_75 b_12 NI_12 NS_75 0 1.8971031711518321e-03
GC_12_76 b_12 NI_12 NS_76 0 -5.9841340000738735e-04
GC_12_77 b_12 NI_12 NS_77 0 7.5215563620410523e-06
GC_12_78 b_12 NI_12 NS_78 0 2.6488480223230879e-06
GC_12_79 b_12 NI_12 NS_79 0 -6.5665550032859417e-05
GC_12_80 b_12 NI_12 NS_80 0 -1.6379777749302830e-04
GC_12_81 b_12 NI_12 NS_81 0 -2.3493216194306740e-05
GC_12_82 b_12 NI_12 NS_82 0 1.7814404483826381e-07
GC_12_83 b_12 NI_12 NS_83 0 1.7964554907133169e-05
GC_12_84 b_12 NI_12 NS_84 0 -1.4685968396108438e-06
GC_12_85 b_12 NI_12 NS_85 0 -9.4303416138731226e-06
GC_12_86 b_12 NI_12 NS_86 0 5.6555931641100405e-06
GC_12_87 b_12 NI_12 NS_87 0 1.9716278086841170e-04
GC_12_88 b_12 NI_12 NS_88 0 9.8075526287332140e-05
GC_12_89 b_12 NI_12 NS_89 0 1.2860599102344000e-02
GC_12_90 b_12 NI_12 NS_90 0 -4.7108784667063974e-05
GC_12_91 b_12 NI_12 NS_91 0 -6.3757923383500766e-04
GC_12_92 b_12 NI_12 NS_92 0 6.3611841263142216e-04
GC_12_93 b_12 NI_12 NS_93 0 -2.5329589468787593e-04
GC_12_94 b_12 NI_12 NS_94 0 -8.0152231836678838e-04
GC_12_95 b_12 NI_12 NS_95 0 -3.2284861038009611e-04
GC_12_96 b_12 NI_12 NS_96 0 -5.4335058832852612e-05
GC_12_97 b_12 NI_12 NS_97 0 5.6866688778439082e-04
GC_12_98 b_12 NI_12 NS_98 0 -1.0194718259631077e-04
GC_12_99 b_12 NI_12 NS_99 0 -4.5872329695339559e-04
GC_12_100 b_12 NI_12 NS_100 0 3.4302166773113264e-04
GC_12_101 b_12 NI_12 NS_101 0 9.8835247177443618e-05
GC_12_102 b_12 NI_12 NS_102 0 7.1405683555249606e-05
GC_12_103 b_12 NI_12 NS_103 0 -1.6623360670808832e-05
GC_12_104 b_12 NI_12 NS_104 0 8.1597706222589605e-04
GC_12_105 b_12 NI_12 NS_105 0 -1.0675188823557793e-04
GC_12_106 b_12 NI_12 NS_106 0 2.9085327367720213e-05
GC_12_107 b_12 NI_12 NS_107 0 -3.9627565683372724e-04
GC_12_108 b_12 NI_12 NS_108 0 -3.6658052530096979e-05
GC_12_109 b_12 NI_12 NS_109 0 2.4797360059311451e-05
GC_12_110 b_12 NI_12 NS_110 0 -4.9863110541182036e-05
GC_12_111 b_12 NI_12 NS_111 0 -2.5438337740890820e-05
GC_12_112 b_12 NI_12 NS_112 0 -9.6386968114896960e-05
GC_12_113 b_12 NI_12 NS_113 0 -1.7547397692194710e-05
GC_12_114 b_12 NI_12 NS_114 0 7.7928789904796591e-05
GC_12_115 b_12 NI_12 NS_115 0 2.6795502983591461e-04
GC_12_116 b_12 NI_12 NS_116 0 -3.3132577572410902e-04
GC_12_117 b_12 NI_12 NS_117 0 -1.8047884762092043e-05
GC_12_118 b_12 NI_12 NS_118 0 -3.7519022942936757e-06
GC_12_119 b_12 NI_12 NS_119 0 -4.4529983054255820e-04
GC_12_120 b_12 NI_12 NS_120 0 -1.1352623905441370e-04
GC_12_121 b_12 NI_12 NS_121 0 7.6780461511745964e-07
GC_12_122 b_12 NI_12 NS_122 0 6.1923071445899240e-07
GC_12_123 b_12 NI_12 NS_123 0 3.8876469028603770e-06
GC_12_124 b_12 NI_12 NS_124 0 -1.5897523644660985e-04
GC_12_125 b_12 NI_12 NS_125 0 -5.3256301115523925e-06
GC_12_126 b_12 NI_12 NS_126 0 -3.9141387153141318e-06
GC_12_127 b_12 NI_12 NS_127 0 -1.1739995739584002e-07
GC_12_128 b_12 NI_12 NS_128 0 4.5921977467791629e-07
GC_12_129 b_12 NI_12 NS_129 0 1.4615445191271789e-07
GC_12_130 b_12 NI_12 NS_130 0 -1.2343398225296612e-06
GC_12_131 b_12 NI_12 NS_131 0 -1.2461339216163843e-04
GC_12_132 b_12 NI_12 NS_132 0 -3.7127215250479765e-05
GC_12_133 b_12 NI_12 NS_133 0 7.2567150189499442e-04
GC_12_134 b_12 NI_12 NS_134 0 -8.0781696506196679e-06
GC_12_135 b_12 NI_12 NS_135 0 3.3662973581544402e-04
GC_12_136 b_12 NI_12 NS_136 0 -6.9380013119524819e-04
GC_12_137 b_12 NI_12 NS_137 0 3.8925063164922170e-04
GC_12_138 b_12 NI_12 NS_138 0 4.9571224155613093e-04
GC_12_139 b_12 NI_12 NS_139 0 -3.5207873975382013e-04
GC_12_140 b_12 NI_12 NS_140 0 3.5471582843129044e-04
GC_12_141 b_12 NI_12 NS_141 0 2.9819382406643606e-04
GC_12_142 b_12 NI_12 NS_142 0 -8.7688023951149974e-05
GC_12_143 b_12 NI_12 NS_143 0 1.7845249462958507e-04
GC_12_144 b_12 NI_12 NS_144 0 2.3242787143737978e-04
GC_12_145 b_12 NI_12 NS_145 0 -7.9353728476505312e-06
GC_12_146 b_12 NI_12 NS_146 0 1.6355173206886091e-05
GC_12_147 b_12 NI_12 NS_147 0 3.3755574082370242e-04
GC_12_148 b_12 NI_12 NS_148 0 -1.5646858025457740e-04
GC_12_149 b_12 NI_12 NS_149 0 1.0475827515915413e-05
GC_12_150 b_12 NI_12 NS_150 0 -3.0044320081514190e-05
GC_12_151 b_12 NI_12 NS_151 0 4.1675432116952818e-04
GC_12_152 b_12 NI_12 NS_152 0 -1.9135953766420758e-04
GC_12_153 b_12 NI_12 NS_153 0 -5.3924880243516539e-05
GC_12_154 b_12 NI_12 NS_154 0 -1.8196864573496844e-04
GC_12_155 b_12 NI_12 NS_155 0 3.1612224025039707e-06
GC_12_156 b_12 NI_12 NS_156 0 -1.6726211033698121e-05
GC_12_157 b_12 NI_12 NS_157 0 -3.0790345366581852e-05
GC_12_158 b_12 NI_12 NS_158 0 -1.1130855548045588e-04
GC_12_159 b_12 NI_12 NS_159 0 -2.6624618415890498e-03
GC_12_160 b_12 NI_12 NS_160 0 2.8868612301797738e-03
GC_12_161 b_12 NI_12 NS_161 0 4.8420947188108014e-06
GC_12_162 b_12 NI_12 NS_162 0 5.8948043907289878e-06
GC_12_163 b_12 NI_12 NS_163 0 2.2756129492309970e-03
GC_12_164 b_12 NI_12 NS_164 0 -8.7878950779607813e-04
GC_12_165 b_12 NI_12 NS_165 0 6.5909470385630775e-06
GC_12_166 b_12 NI_12 NS_166 0 2.6244148307796147e-06
GC_12_167 b_12 NI_12 NS_167 0 -1.2637915670277332e-04
GC_12_168 b_12 NI_12 NS_168 0 -2.8418512977650221e-04
GC_12_169 b_12 NI_12 NS_169 0 -1.9337984036027726e-05
GC_12_170 b_12 NI_12 NS_170 0 4.2957374774286102e-06
GC_12_171 b_12 NI_12 NS_171 0 2.0232738660593380e-05
GC_12_172 b_12 NI_12 NS_172 0 -1.2019293958744443e-06
GC_12_173 b_12 NI_12 NS_173 0 -9.1170649440262913e-06
GC_12_174 b_12 NI_12 NS_174 0 4.5475276397333925e-06
GC_12_175 b_12 NI_12 NS_175 0 2.1200327348689900e-04
GC_12_176 b_12 NI_12 NS_176 0 5.1564113881334040e-05
GC_12_177 b_12 NI_12 NS_177 0 -5.7455593047236212e-03
GC_12_178 b_12 NI_12 NS_178 0 -1.3716215621066976e-05
GC_12_179 b_12 NI_12 NS_179 0 -1.2902669175292433e-03
GC_12_180 b_12 NI_12 NS_180 0 1.8771742177895430e-04
GC_12_181 b_12 NI_12 NS_181 0 6.4514523678384987e-04
GC_12_182 b_12 NI_12 NS_182 0 -1.2038987595180384e-03
GC_12_183 b_12 NI_12 NS_183 0 2.1272691423020770e-04
GC_12_184 b_12 NI_12 NS_184 0 3.4674124179603222e-04
GC_12_185 b_12 NI_12 NS_185 0 6.6254640754457466e-04
GC_12_186 b_12 NI_12 NS_186 0 -1.1137056874241261e-04
GC_12_187 b_12 NI_12 NS_187 0 -2.1909421256192588e-04
GC_12_188 b_12 NI_12 NS_188 0 -1.0971104498991428e-03
GC_12_189 b_12 NI_12 NS_189 0 1.1271902698941213e-04
GC_12_190 b_12 NI_12 NS_190 0 1.0158079417665466e-04
GC_12_191 b_12 NI_12 NS_191 0 7.7218349988356289e-04
GC_12_192 b_12 NI_12 NS_192 0 1.1535193279889227e-03
GC_12_193 b_12 NI_12 NS_193 0 -1.0184549197007561e-04
GC_12_194 b_12 NI_12 NS_194 0 4.1168523307042905e-05
GC_12_195 b_12 NI_12 NS_195 0 -2.2789404978802277e-04
GC_12_196 b_12 NI_12 NS_196 0 -5.7001304009919288e-05
GC_12_197 b_12 NI_12 NS_197 0 4.3656688895393764e-05
GC_12_198 b_12 NI_12 NS_198 0 7.3423703378600324e-05
GC_12_199 b_12 NI_12 NS_199 0 -1.5631560599607354e-05
GC_12_200 b_12 NI_12 NS_200 0 -8.6266448429086267e-05
GC_12_201 b_12 NI_12 NS_201 0 -5.6545615446022195e-06
GC_12_202 b_12 NI_12 NS_202 0 8.0449816916416215e-05
GC_12_203 b_12 NI_12 NS_203 0 1.2320690701419421e-03
GC_12_204 b_12 NI_12 NS_204 0 -1.1378689707318044e-04
GC_12_205 b_12 NI_12 NS_205 0 -1.8359328859465631e-05
GC_12_206 b_12 NI_12 NS_206 0 -1.7125560052692174e-06
GC_12_207 b_12 NI_12 NS_207 0 -4.6257679585013631e-04
GC_12_208 b_12 NI_12 NS_208 0 -2.2343191876900229e-04
GC_12_209 b_12 NI_12 NS_209 0 -9.6214933107039879e-07
GC_12_210 b_12 NI_12 NS_210 0 1.7060879721785364e-06
GC_12_211 b_12 NI_12 NS_211 0 5.5096224022562703e-05
GC_12_212 b_12 NI_12 NS_212 0 7.9463084264669222e-06
GC_12_213 b_12 NI_12 NS_213 0 -5.7752551927424562e-06
GC_12_214 b_12 NI_12 NS_214 0 -1.0983567740093290e-05
GC_12_215 b_12 NI_12 NS_215 0 -8.6041549836721342e-08
GC_12_216 b_12 NI_12 NS_216 0 1.4999175527107512e-06
GC_12_217 b_12 NI_12 NS_217 0 -7.6507448073493751e-07
GC_12_218 b_12 NI_12 NS_218 0 -8.2473616931111228e-07
GC_12_219 b_12 NI_12 NS_219 0 -1.4442635118354648e-04
GC_12_220 b_12 NI_12 NS_220 0 -7.1193339756234237e-06
GC_12_221 b_12 NI_12 NS_221 0 1.2540202002052658e-03
GC_12_222 b_12 NI_12 NS_222 0 -3.2026248872342691e-05
GC_12_223 b_12 NI_12 NS_223 0 8.1546736481860778e-04
GC_12_224 b_12 NI_12 NS_224 0 -5.7894156632457873e-04
GC_12_225 b_12 NI_12 NS_225 0 -2.7239275214320204e-04
GC_12_226 b_12 NI_12 NS_226 0 7.7376690266120138e-04
GC_12_227 b_12 NI_12 NS_227 0 -6.0919699001357297e-04
GC_12_228 b_12 NI_12 NS_228 0 1.2902447382293945e-04
GC_12_229 b_12 NI_12 NS_229 0 1.7009403280867003e-04
GC_12_230 b_12 NI_12 NS_230 0 -1.4359737393657075e-04
GC_12_231 b_12 NI_12 NS_231 0 -1.4322674767477923e-04
GC_12_232 b_12 NI_12 NS_232 0 -1.9327103589912936e-04
GC_12_233 b_12 NI_12 NS_233 0 -7.5152624367432040e-06
GC_12_234 b_12 NI_12 NS_234 0 1.8486941656585619e-05
GC_12_235 b_12 NI_12 NS_235 0 5.1042155099420377e-04
GC_12_236 b_12 NI_12 NS_236 0 -7.9716883597953967e-05
GC_12_237 b_12 NI_12 NS_237 0 1.4250158382220485e-05
GC_12_238 b_12 NI_12 NS_238 0 -4.2994163225600742e-05
GC_12_239 b_12 NI_12 NS_239 0 4.8058563424738699e-04
GC_12_240 b_12 NI_12 NS_240 0 -3.1871655525640452e-04
GC_12_241 b_12 NI_12 NS_241 0 -8.9583996100558454e-05
GC_12_242 b_12 NI_12 NS_242 0 -2.2334874758119544e-04
GC_12_243 b_12 NI_12 NS_243 0 1.6604558210091638e-06
GC_12_244 b_12 NI_12 NS_244 0 -2.8920547494820074e-05
GC_12_245 b_12 NI_12 NS_245 0 -4.7202523301515991e-05
GC_12_246 b_12 NI_12 NS_246 0 -1.4992322040419351e-04
GC_12_247 b_12 NI_12 NS_247 0 -3.0985337908212007e-03
GC_12_248 b_12 NI_12 NS_248 0 3.2699874768377995e-03
GC_12_249 b_12 NI_12 NS_249 0 6.7883969172459697e-06
GC_12_250 b_12 NI_12 NS_250 0 5.2403618431669862e-06
GC_12_251 b_12 NI_12 NS_251 0 2.8197714176977358e-03
GC_12_252 b_12 NI_12 NS_252 0 -1.1144627613033143e-03
GC_12_253 b_12 NI_12 NS_253 0 1.1482132040850822e-05
GC_12_254 b_12 NI_12 NS_254 0 5.4142568311679317e-06
GC_12_255 b_12 NI_12 NS_255 0 -4.5566564256111030e-05
GC_12_256 b_12 NI_12 NS_256 0 -2.6279788239282086e-04
GC_12_257 b_12 NI_12 NS_257 0 -3.3524201682488933e-05
GC_12_258 b_12 NI_12 NS_258 0 3.0850583774836745e-06
GC_12_259 b_12 NI_12 NS_259 0 2.8178598698298593e-05
GC_12_260 b_12 NI_12 NS_260 0 -3.9493520623938591e-06
GC_12_261 b_12 NI_12 NS_261 0 -1.1068944765603274e-05
GC_12_262 b_12 NI_12 NS_262 0 8.6936063229772718e-06
GC_12_263 b_12 NI_12 NS_263 0 2.9997972066185850e-04
GC_12_264 b_12 NI_12 NS_264 0 1.2609752805396168e-04
GC_12_265 b_12 NI_12 NS_265 0 2.7416821053949381e-03
GC_12_266 b_12 NI_12 NS_266 0 4.1168496062033942e-05
GC_12_267 b_12 NI_12 NS_267 0 -1.7998031526939632e-03
GC_12_268 b_12 NI_12 NS_268 0 -1.0956975879347574e-03
GC_12_269 b_12 NI_12 NS_269 0 1.4061287677789749e-03
GC_12_270 b_12 NI_12 NS_270 0 7.0213036245064895e-04
GC_12_271 b_12 NI_12 NS_271 0 4.4494701136611807e-05
GC_12_272 b_12 NI_12 NS_272 0 6.0761409488069615e-05
GC_12_273 b_12 NI_12 NS_273 0 4.0868527091089988e-04
GC_12_274 b_12 NI_12 NS_274 0 2.8035047528356198e-05
GC_12_275 b_12 NI_12 NS_275 0 6.1039431012392621e-04
GC_12_276 b_12 NI_12 NS_276 0 -1.3317933062945157e-03
GC_12_277 b_12 NI_12 NS_277 0 4.2358957623543685e-05
GC_12_278 b_12 NI_12 NS_278 0 1.2273835103602547e-04
GC_12_279 b_12 NI_12 NS_279 0 9.7907626279921979e-06
GC_12_280 b_12 NI_12 NS_280 0 7.0033702330230690e-04
GC_12_281 b_12 NI_12 NS_281 0 -8.1819293741059847e-05
GC_12_282 b_12 NI_12 NS_282 0 2.7092583160882384e-05
GC_12_283 b_12 NI_12 NS_283 0 -2.0444835456807914e-04
GC_12_284 b_12 NI_12 NS_284 0 2.8030879047198724e-04
GC_12_285 b_12 NI_12 NS_285 0 -4.0192522852989424e-05
GC_12_286 b_12 NI_12 NS_286 0 1.2817891194834529e-04
GC_12_287 b_12 NI_12 NS_287 0 -1.8759764286511772e-05
GC_12_288 b_12 NI_12 NS_288 0 -5.5203906824540243e-05
GC_12_289 b_12 NI_12 NS_289 0 -1.2490526480872274e-05
GC_12_290 b_12 NI_12 NS_290 0 6.3122935733288797e-05
GC_12_291 b_12 NI_12 NS_291 0 1.9078896444233153e-04
GC_12_292 b_12 NI_12 NS_292 0 4.4062811619574425e-04
GC_12_293 b_12 NI_12 NS_293 0 -9.5864328012914176e-06
GC_12_294 b_12 NI_12 NS_294 0 -2.3338414436469194e-06
GC_12_295 b_12 NI_12 NS_295 0 -9.9191686899032763e-05
GC_12_296 b_12 NI_12 NS_296 0 -3.7418946851503371e-05
GC_12_297 b_12 NI_12 NS_297 0 -1.0967008848027721e-06
GC_12_298 b_12 NI_12 NS_298 0 -6.6645484130595018e-07
GC_12_299 b_12 NI_12 NS_299 0 -4.7273373415018693e-05
GC_12_300 b_12 NI_12 NS_300 0 -8.4486613005345924e-05
GC_12_301 b_12 NI_12 NS_301 0 -3.2869429490164524e-06
GC_12_302 b_12 NI_12 NS_302 0 -5.2571843691307783e-06
GC_12_303 b_12 NI_12 NS_303 0 2.8977118799773766e-08
GC_12_304 b_12 NI_12 NS_304 0 -1.8341953382239372e-07
GC_12_305 b_12 NI_12 NS_305 0 -1.9804352499984247e-07
GC_12_306 b_12 NI_12 NS_306 0 -6.8285135772943587e-07
GC_12_307 b_12 NI_12 NS_307 0 -8.7484558690521395e-05
GC_12_308 b_12 NI_12 NS_308 0 -3.9080144668703048e-05
GC_12_309 b_12 NI_12 NS_309 0 -2.0376969194448673e-03
GC_12_310 b_12 NI_12 NS_310 0 -2.6979148551804755e-04
GC_12_311 b_12 NI_12 NS_311 0 9.8746942026836496e-04
GC_12_312 b_12 NI_12 NS_312 0 6.2089334503077171e-04
GC_12_313 b_12 NI_12 NS_313 0 -1.6023503573726525e-03
GC_12_314 b_12 NI_12 NS_314 0 -1.0182016742717745e-03
GC_12_315 b_12 NI_12 NS_315 0 -1.5221769099956354e-04
GC_12_316 b_12 NI_12 NS_316 0 -3.5021747089980748e-04
GC_12_317 b_12 NI_12 NS_317 0 2.7047197216471651e-04
GC_12_318 b_12 NI_12 NS_318 0 -1.3273472071456146e-04
GC_12_319 b_12 NI_12 NS_319 0 1.8394262161598366e-05
GC_12_320 b_12 NI_12 NS_320 0 -7.8835916883229968e-04
GC_12_321 b_12 NI_12 NS_321 0 1.1315950055285412e-06
GC_12_322 b_12 NI_12 NS_322 0 2.5322931791419846e-05
GC_12_323 b_12 NI_12 NS_323 0 1.9640154351980592e-04
GC_12_324 b_12 NI_12 NS_324 0 -3.7604674853667405e-04
GC_12_325 b_12 NI_12 NS_325 0 1.6413426706888130e-05
GC_12_326 b_12 NI_12 NS_326 0 -2.2490592156737270e-05
GC_12_327 b_12 NI_12 NS_327 0 4.6980028007794335e-04
GC_12_328 b_12 NI_12 NS_328 0 -2.8035645497090524e-04
GC_12_329 b_12 NI_12 NS_329 0 -5.2532684292244679e-05
GC_12_330 b_12 NI_12 NS_330 0 -1.2391619079189025e-04
GC_12_331 b_12 NI_12 NS_331 0 1.1188319458938586e-05
GC_12_332 b_12 NI_12 NS_332 0 -1.7939387653389714e-05
GC_12_333 b_12 NI_12 NS_333 0 -2.4806303414456570e-05
GC_12_334 b_12 NI_12 NS_334 0 -1.0140405251283147e-04
GC_12_335 b_12 NI_12 NS_335 0 -1.0091146194478656e-03
GC_12_336 b_12 NI_12 NS_336 0 2.6860199449809524e-03
GC_12_337 b_12 NI_12 NS_337 0 -1.3367844716032680e-06
GC_12_338 b_12 NI_12 NS_338 0 -8.5138660233521044e-07
GC_12_339 b_12 NI_12 NS_339 0 1.7787760506601106e-03
GC_12_340 b_12 NI_12 NS_340 0 -1.0063314776676548e-03
GC_12_341 b_12 NI_12 NS_341 0 3.9880543851292852e-06
GC_12_342 b_12 NI_12 NS_342 0 2.0130104597856281e-06
GC_12_343 b_12 NI_12 NS_343 0 -1.2995156888333847e-04
GC_12_344 b_12 NI_12 NS_344 0 -3.9594109249477731e-06
GC_12_345 b_12 NI_12 NS_345 0 -9.3783845159120568e-06
GC_12_346 b_12 NI_12 NS_346 0 3.0116554144618495e-06
GC_12_347 b_12 NI_12 NS_347 0 1.7798938505660059e-05
GC_12_348 b_12 NI_12 NS_348 0 2.4251323756866087e-07
GC_12_349 b_12 NI_12 NS_349 0 -4.5695707036083107e-06
GC_12_350 b_12 NI_12 NS_350 0 2.4362469572924428e-06
GC_12_351 b_12 NI_12 NS_351 0 1.2410760115777570e-04
GC_12_352 b_12 NI_12 NS_352 0 6.9885891917227736e-05
GC_12_353 b_12 NI_12 NS_353 0 6.2350542206847825e-02
GC_12_354 b_12 NI_12 NS_354 0 -7.6655238742362553e-05
GC_12_355 b_12 NI_12 NS_355 0 -6.3061911194363550e-03
GC_12_356 b_12 NI_12 NS_356 0 -2.5760123201772596e-03
GC_12_357 b_12 NI_12 NS_357 0 4.1561119705232673e-03
GC_12_358 b_12 NI_12 NS_358 0 2.6622431684536528e-03
GC_12_359 b_12 NI_12 NS_359 0 1.8528782085229758e-05
GC_12_360 b_12 NI_12 NS_360 0 1.7264092657374648e-05
GC_12_361 b_12 NI_12 NS_361 0 1.3250795595782735e-03
GC_12_362 b_12 NI_12 NS_362 0 1.5410622119305648e-03
GC_12_363 b_12 NI_12 NS_363 0 -3.0663438037846762e-04
GC_12_364 b_12 NI_12 NS_364 0 -3.0277794352990531e-04
GC_12_365 b_12 NI_12 NS_365 0 -6.5925268981015931e-05
GC_12_366 b_12 NI_12 NS_366 0 7.1505999997253109e-05
GC_12_367 b_12 NI_12 NS_367 0 -4.4716097059574814e-03
GC_12_368 b_12 NI_12 NS_368 0 9.1005488843021523e-04
GC_12_369 b_12 NI_12 NS_369 0 -8.4331119166457331e-05
GC_12_370 b_12 NI_12 NS_370 0 -5.7373344946614351e-05
GC_12_371 b_12 NI_12 NS_371 0 -5.0364603618903621e-04
GC_12_372 b_12 NI_12 NS_372 0 6.7167669751616750e-04
GC_12_373 b_12 NI_12 NS_373 0 3.8218817594644816e-04
GC_12_374 b_12 NI_12 NS_374 0 2.1974337075793978e-04
GC_12_375 b_12 NI_12 NS_375 0 -3.8368825840179244e-05
GC_12_376 b_12 NI_12 NS_376 0 -5.5206536578351493e-05
GC_12_377 b_12 NI_12 NS_377 0 -4.5984203314002805e-05
GC_12_378 b_12 NI_12 NS_378 0 8.1003859137751050e-05
GC_12_379 b_12 NI_12 NS_379 0 -2.2101035521148683e-03
GC_12_380 b_12 NI_12 NS_380 0 -4.9286261333404786e-03
GC_12_381 b_12 NI_12 NS_381 0 8.8201569393824121e-06
GC_12_382 b_12 NI_12 NS_382 0 3.1308145198061283e-05
GC_12_383 b_12 NI_12 NS_383 0 -1.0172721443567736e-03
GC_12_384 b_12 NI_12 NS_384 0 2.0857168392405989e-03
GC_12_385 b_12 NI_12 NS_385 0 -3.9419795713055606e-06
GC_12_386 b_12 NI_12 NS_386 0 9.8955693879682906e-06
GC_12_387 b_12 NI_12 NS_387 0 1.1473988216559635e-03
GC_12_388 b_12 NI_12 NS_388 0 -1.9937431007269933e-04
GC_12_389 b_12 NI_12 NS_389 0 -9.1484455381306974e-06
GC_12_390 b_12 NI_12 NS_390 0 -1.4434541503616389e-05
GC_12_391 b_12 NI_12 NS_391 0 2.8249065378592359e-06
GC_12_392 b_12 NI_12 NS_392 0 2.5727351489596320e-07
GC_12_393 b_12 NI_12 NS_393 0 1.9039410050006792e-06
GC_12_394 b_12 NI_12 NS_394 0 3.8167548275675512e-06
GC_12_395 b_12 NI_12 NS_395 0 1.3994629963121416e-04
GC_12_396 b_12 NI_12 NS_396 0 -6.3155412303413010e-05
GC_12_397 b_12 NI_12 NS_397 0 2.4173200764673894e-03
GC_12_398 b_12 NI_12 NS_398 0 -8.9963953402805662e-04
GC_12_399 b_12 NI_12 NS_399 0 3.9215896045025501e-03
GC_12_400 b_12 NI_12 NS_400 0 1.5934910656430613e-03
GC_12_401 b_12 NI_12 NS_401 0 -5.1951684061074411e-03
GC_12_402 b_12 NI_12 NS_402 0 -2.2950835618066809e-03
GC_12_403 b_12 NI_12 NS_403 0 -1.9306587163976343e-05
GC_12_404 b_12 NI_12 NS_404 0 -3.2372028033765044e-04
GC_12_405 b_12 NI_12 NS_405 0 1.2198672016797874e-03
GC_12_406 b_12 NI_12 NS_406 0 7.2025048449754600e-05
GC_12_407 b_12 NI_12 NS_407 0 -1.1882254250867341e-04
GC_12_408 b_12 NI_12 NS_408 0 -4.9216401053154884e-04
GC_12_409 b_12 NI_12 NS_409 0 -3.0545348102446187e-05
GC_12_410 b_12 NI_12 NS_410 0 -3.9662352823076623e-05
GC_12_411 b_12 NI_12 NS_411 0 -1.4006382872237819e-03
GC_12_412 b_12 NI_12 NS_412 0 4.2432315932599554e-04
GC_12_413 b_12 NI_12 NS_413 0 2.4952484390707738e-05
GC_12_414 b_12 NI_12 NS_414 0 -3.2409263637192278e-05
GC_12_415 b_12 NI_12 NS_415 0 2.3828704876562490e-05
GC_12_416 b_12 NI_12 NS_416 0 -3.6215976694950372e-04
GC_12_417 b_12 NI_12 NS_417 0 1.8587166361036208e-04
GC_12_418 b_12 NI_12 NS_418 0 -6.1147365075184956e-05
GC_12_419 b_12 NI_12 NS_419 0 -8.6207220029495928e-06
GC_12_420 b_12 NI_12 NS_420 0 -4.8737169574516055e-05
GC_12_421 b_12 NI_12 NS_421 0 -6.4513434790561082e-05
GC_12_422 b_12 NI_12 NS_422 0 -1.2458553948630960e-04
GC_12_423 b_12 NI_12 NS_423 0 1.8961261735367337e-03
GC_12_424 b_12 NI_12 NS_424 0 -4.9493402790130219e-04
GC_12_425 b_12 NI_12 NS_425 0 -3.6844538244122207e-05
GC_12_426 b_12 NI_12 NS_426 0 -3.0272954603568499e-05
GC_12_427 b_12 NI_12 NS_427 0 6.2331791862606841e-04
GC_12_428 b_12 NI_12 NS_428 0 -7.2798220536480932e-04
GC_12_429 b_12 NI_12 NS_429 0 -1.0089473556025659e-05
GC_12_430 b_12 NI_12 NS_430 0 1.2150397117948731e-05
GC_12_431 b_12 NI_12 NS_431 0 4.2947275634415622e-04
GC_12_432 b_12 NI_12 NS_432 0 4.8341743755956571e-04
GC_12_433 b_12 NI_12 NS_433 0 -6.9441858103714550e-07
GC_12_434 b_12 NI_12 NS_434 0 -1.4088778972271764e-05
GC_12_435 b_12 NI_12 NS_435 0 2.8826109087496175e-05
GC_12_436 b_12 NI_12 NS_436 0 4.8882504768930376e-07
GC_12_437 b_12 NI_12 NS_437 0 1.9709692660327817e-05
GC_12_438 b_12 NI_12 NS_438 0 -7.9146041111601873e-06
GC_12_439 b_12 NI_12 NS_439 0 -6.7909409960086796e-05
GC_12_440 b_12 NI_12 NS_440 0 2.3598926367086550e-04
GC_12_441 b_12 NI_12 NS_441 0 -4.2708164759708826e-04
GC_12_442 b_12 NI_12 NS_442 0 1.0643826866945264e-02
GC_12_443 b_12 NI_12 NS_443 0 -6.8704980320661874e-03
GC_12_444 b_12 NI_12 NS_444 0 -5.0120136606891918e-03
GC_12_445 b_12 NI_12 NS_445 0 -1.1447835455601900e-02
GC_12_446 b_12 NI_12 NS_446 0 1.0735562467621891e-03
GC_12_447 b_12 NI_12 NS_447 0 -7.3720617920908871e-06
GC_12_448 b_12 NI_12 NS_448 0 4.4728455443595965e-04
GC_12_449 b_12 NI_12 NS_449 0 1.2785105033435568e-03
GC_12_450 b_12 NI_12 NS_450 0 1.3899937933297640e-03
GC_12_451 b_12 NI_12 NS_451 0 3.2307851457270874e-03
GC_12_452 b_12 NI_12 NS_452 0 -1.4843900157400043e-03
GC_12_453 b_12 NI_12 NS_453 0 -1.3201530188005617e-06
GC_12_454 b_12 NI_12 NS_454 0 1.8361673199479217e-04
GC_12_455 b_12 NI_12 NS_455 0 3.0586200535160511e-03
GC_12_456 b_12 NI_12 NS_456 0 -1.0036044362568795e-03
GC_12_457 b_12 NI_12 NS_457 0 -3.6793167563789502e-05
GC_12_458 b_12 NI_12 NS_458 0 -8.9992844752383128e-06
GC_12_459 b_12 NI_12 NS_459 0 2.2235484117139482e-04
GC_12_460 b_12 NI_12 NS_460 0 2.0825856965312682e-04
GC_12_461 b_12 NI_12 NS_461 0 -9.1313663242178922e-05
GC_12_462 b_12 NI_12 NS_462 0 -1.7871927752417869e-07
GC_12_463 b_12 NI_12 NS_463 0 1.0552693721233872e-06
GC_12_464 b_12 NI_12 NS_464 0 -3.6284964867472331e-05
GC_12_465 b_12 NI_12 NS_465 0 -2.6579763599013045e-05
GC_12_466 b_12 NI_12 NS_466 0 4.9701355719089212e-05
GC_12_467 b_12 NI_12 NS_467 0 -5.4520826573199038e-04
GC_12_468 b_12 NI_12 NS_468 0 -6.7363334585057201e-04
GC_12_469 b_12 NI_12 NS_469 0 -1.5672381782325288e-06
GC_12_470 b_12 NI_12 NS_470 0 1.4085058367739669e-05
GC_12_471 b_12 NI_12 NS_471 0 -3.0121106132893771e-04
GC_12_472 b_12 NI_12 NS_472 0 5.2550430815185970e-04
GC_12_473 b_12 NI_12 NS_473 0 -1.4415676554340978e-06
GC_12_474 b_12 NI_12 NS_474 0 -7.4825903051447398e-07
GC_12_475 b_12 NI_12 NS_475 0 -5.8512335176419802e-06
GC_12_476 b_12 NI_12 NS_476 0 -1.2587912901515215e-04
GC_12_477 b_12 NI_12 NS_477 0 -7.1245037160220574e-09
GC_12_478 b_12 NI_12 NS_478 0 -1.6376168552425791e-06
GC_12_479 b_12 NI_12 NS_479 0 6.1888673415090894e-07
GC_12_480 b_12 NI_12 NS_480 0 8.9686813024106555e-08
GC_12_481 b_12 NI_12 NS_481 0 4.5856719700087051e-09
GC_12_482 b_12 NI_12 NS_482 0 -1.6803763439052693e-06
GC_12_483 b_12 NI_12 NS_483 0 -2.9751339538169018e-05
GC_12_484 b_12 NI_12 NS_484 0 -4.9532285572861893e-05
GC_12_485 b_12 NI_12 NS_485 0 -2.0974161974278516e-01
GC_12_486 b_12 NI_12 NS_486 0 8.5122560968368208e-03
GC_12_487 b_12 NI_12 NS_487 0 3.9389624399706058e-03
GC_12_488 b_12 NI_12 NS_488 0 6.3447891261458117e-03
GC_12_489 b_12 NI_12 NS_489 0 6.3735057916426393e-03
GC_12_490 b_12 NI_12 NS_490 0 -1.4728768484797523e-03
GC_12_491 b_12 NI_12 NS_491 0 1.0220457765955364e-03
GC_12_492 b_12 NI_12 NS_492 0 -2.5402354827195375e-04
GC_12_493 b_12 NI_12 NS_493 0 3.8323176271744311e-05
GC_12_494 b_12 NI_12 NS_494 0 1.4305840645968105e-03
GC_12_495 b_12 NI_12 NS_495 0 4.8532954886492292e-03
GC_12_496 b_12 NI_12 NS_496 0 2.0735074719675523e-03
GC_12_497 b_12 NI_12 NS_497 0 -2.1428855732649553e-04
GC_12_498 b_12 NI_12 NS_498 0 2.8146793344386250e-04
GC_12_499 b_12 NI_12 NS_499 0 1.3880798227345191e-03
GC_12_500 b_12 NI_12 NS_500 0 7.3954976629484626e-03
GC_12_501 b_12 NI_12 NS_501 0 -7.9388241417946729e-05
GC_12_502 b_12 NI_12 NS_502 0 8.1311494185085860e-05
GC_12_503 b_12 NI_12 NS_503 0 -4.2764070548124408e-04
GC_12_504 b_12 NI_12 NS_504 0 3.3126683248566762e-03
GC_12_505 b_12 NI_12 NS_505 0 5.1276143498414097e-04
GC_12_506 b_12 NI_12 NS_506 0 -2.0132379956791806e-04
GC_12_507 b_12 NI_12 NS_507 0 -1.1580927713229575e-04
GC_12_508 b_12 NI_12 NS_508 0 1.3690672201205554e-04
GC_12_509 b_12 NI_12 NS_509 0 1.9752176253350615e-05
GC_12_510 b_12 NI_12 NS_510 0 3.0510444002575873e-05
GC_12_511 b_12 NI_12 NS_511 0 -1.9135773487144819e-02
GC_12_512 b_12 NI_12 NS_512 0 -3.4522295129271610e-04
GC_12_513 b_12 NI_12 NS_513 0 2.9900381666650800e-05
GC_12_514 b_12 NI_12 NS_514 0 -2.0080412497363155e-05
GC_12_515 b_12 NI_12 NS_515 0 4.7909050580139589e-03
GC_12_516 b_12 NI_12 NS_516 0 4.8255635979699684e-03
GC_12_517 b_12 NI_12 NS_517 0 8.8003491761243698e-07
GC_12_518 b_12 NI_12 NS_518 0 3.8585949969754123e-05
GC_12_519 b_12 NI_12 NS_519 0 1.5599100431221676e-03
GC_12_520 b_12 NI_12 NS_520 0 -2.5655838691137512e-03
GC_12_521 b_12 NI_12 NS_521 0 -5.6200639145160372e-05
GC_12_522 b_12 NI_12 NS_522 0 -1.9485297041601074e-05
GC_12_523 b_12 NI_12 NS_523 0 1.8693252513548583e-05
GC_12_524 b_12 NI_12 NS_524 0 -1.3870211867820562e-05
GC_12_525 b_12 NI_12 NS_525 0 3.0673982222364725e-05
GC_12_526 b_12 NI_12 NS_526 0 6.2243233909538465e-06
GC_12_527 b_12 NI_12 NS_527 0 4.8466378628223055e-04
GC_12_528 b_12 NI_12 NS_528 0 -4.9870876752896058e-04
GD_12_1 b_12 NI_12 NA_1 0 -1.4221113416605051e-02
GD_12_2 b_12 NI_12 NA_2 0 -2.9557136715395861e-03
GD_12_3 b_12 NI_12 NA_3 0 -1.2056772305508588e-02
GD_12_4 b_12 NI_12 NA_4 0 -3.3553895468513822e-03
GD_12_5 b_12 NI_12 NA_5 0 3.8252618377357952e-03
GD_12_6 b_12 NI_12 NA_6 0 -3.3694698104132226e-03
GD_12_7 b_12 NI_12 NA_7 0 -4.8329132536127561e-03
GD_12_8 b_12 NI_12 NA_8 0 -2.1945666340195840e-04
GD_12_9 b_12 NI_12 NA_9 0 -6.4891693247787929e-02
GD_12_10 b_12 NI_12 NA_10 0 -8.6526583901853273e-03
GD_12_11 b_12 NI_12 NA_11 0 2.2570012410937008e-03
GD_12_12 b_12 NI_12 NA_12 0 2.6886836568734046e-01
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+00
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-02
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+00
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-02
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+00
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-02
*
* Impinging wave, port 4
RA_4 NA_4 0 3.5355339059327378e+00
FA_4 0 NA_4 VI_4 1.0
GA_4 0 NA_4 a_4 b_4 2.0000000000000000e-02
*
* Impinging wave, port 5
RA_5 NA_5 0 3.5355339059327378e+00
FA_5 0 NA_5 VI_5 1.0
GA_5 0 NA_5 a_5 b_5 2.0000000000000000e-02
*
* Impinging wave, port 6
RA_6 NA_6 0 3.5355339059327378e+00
FA_6 0 NA_6 VI_6 1.0
GA_6 0 NA_6 a_6 b_6 2.0000000000000000e-02
*
* Impinging wave, port 7
RA_7 NA_7 0 3.5355339059327378e+00
FA_7 0 NA_7 VI_7 1.0
GA_7 0 NA_7 a_7 b_7 2.0000000000000000e-02
*
* Impinging wave, port 8
RA_8 NA_8 0 3.5355339059327378e+00
FA_8 0 NA_8 VI_8 1.0
GA_8 0 NA_8 a_8 b_8 2.0000000000000000e-02
*
* Impinging wave, port 9
RA_9 NA_9 0 3.5355339059327378e+00
FA_9 0 NA_9 VI_9 1.0
GA_9 0 NA_9 a_9 b_9 2.0000000000000000e-02
*
* Impinging wave, port 10
RA_10 NA_10 0 3.5355339059327378e+00
FA_10 0 NA_10 VI_10 1.0
GA_10 0 NA_10 a_10 b_10 2.0000000000000000e-02
*
* Impinging wave, port 11
RA_11 NA_11 0 3.5355339059327378e+00
FA_11 0 NA_11 VI_11 1.0
GA_11 0 NA_11 a_11 b_11 2.0000000000000000e-02
*
* Impinging wave, port 12
RA_12 NA_12 0 3.5355339059327378e+00
FA_12 0 NA_12 VI_12 1.0
GA_12 0 NA_12 a_12 b_12 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-13
RS_1 NS_1 0 1.2063458770185771e+00
GS_1_1 0 NS_1 NA_1 0 1.6921379288850509e+00
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-13
RS_2 NS_2 0 2.0414994648771170e+01
GS_2_1 0 NS_2 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 3/4
CS_3 NS_3 0 9.9999999999999998e-13
CS_4 NS_4 0 9.9999999999999998e-13
RS_3 NS_3 0 2.2164632983638530e+01
RS_4 NS_4 0 2.2164632983638530e+01
GL_3 0 NS_3 NS_4 0 6.2432580119989492e-02
GL_4 0 NS_4 NS_3 0 -6.2432580119989492e-02
GS_3_1 0 NS_3 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 5/6
CS_5 NS_5 0 9.9999999999999998e-13
CS_6 NS_6 0 9.9999999999999998e-13
RS_5 NS_5 0 2.4208144339458560e+01
RS_6 NS_6 0 2.4208144339458560e+01
GL_5 0 NS_5 NS_6 0 8.7759448763363015e-02
GL_6 0 NS_6 NS_5 0 -8.7759448763363015e-02
GS_5_1 0 NS_5 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 7/8
CS_7 NS_7 0 9.9999999999999998e-13
CS_8 NS_8 0 9.9999999999999998e-13
RS_7 NS_7 0 1.3097029666184031e+02
RS_8 NS_8 0 1.3097029666184031e+02
GL_7 0 NS_7 NS_8 0 2.9672291989323329e-01
GL_8 0 NS_8 NS_7 0 -2.9672291989323329e-01
GS_7_1 0 NS_7 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 9/10
CS_9 NS_9 0 9.9999999999999998e-13
CS_10 NS_10 0 9.9999999999999998e-13
RS_9 NS_9 0 3.2672536376024027e+01
RS_10 NS_10 0 3.2672536376024027e+01
GL_9 0 NS_9 NS_10 0 1.2489866711430768e-01
GL_10 0 NS_10 NS_9 0 -1.2489866711430768e-01
GS_9_1 0 NS_9 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 11/12
CS_11 NS_11 0 9.9999999999999998e-13
CS_12 NS_12 0 9.9999999999999998e-13
RS_11 NS_11 0 3.6741731246022816e+01
RS_12 NS_12 0 3.6741731246022816e+01
GL_11 0 NS_11 NS_12 0 1.6399845549232167e-01
GL_12 0 NS_12 NS_11 0 -1.6399845549232167e-01
GS_11_1 0 NS_11 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 13/14
CS_13 NS_13 0 9.9999999999999998e-13
CS_14 NS_14 0 9.9999999999999998e-13
RS_13 NS_13 0 8.3646036557163740e+01
RS_14 NS_14 0 8.3646036557163740e+01
GL_13 0 NS_13 NS_14 0 1.6830719130342967e-01
GL_14 0 NS_14 NS_13 0 -1.6830719130342967e-01
GS_13_1 0 NS_13 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 15/16
CS_15 NS_15 0 9.9999999999999998e-13
CS_16 NS_16 0 9.9999999999999998e-13
RS_15 NS_15 0 4.0307732865054554e+01
RS_16 NS_16 0 4.0307732865054554e+01
GL_15 0 NS_15 NS_16 0 1.8890575271706389e-01
GL_16 0 NS_16 NS_15 0 -1.8890575271706389e-01
GS_15_1 0 NS_15 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 17/18
CS_17 NS_17 0 9.9999999999999998e-13
CS_18 NS_18 0 9.9999999999999998e-13
RS_17 NS_17 0 1.4268073111996583e+02
RS_18 NS_18 0 1.4268073111996583e+02
GL_17 0 NS_17 NS_18 0 1.9419078929943706e-01
GL_18 0 NS_18 NS_17 0 -1.9419078929943706e-01
GS_17_1 0 NS_17 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 19/20
CS_19 NS_19 0 9.9999999999999998e-13
CS_20 NS_20 0 9.9999999999999998e-13
RS_19 NS_19 0 7.1679198821979867e+01
RS_20 NS_20 0 7.1679198821979867e+01
GL_19 0 NS_19 NS_20 0 2.0702628270375376e-01
GL_20 0 NS_20 NS_19 0 -2.0702628270375376e-01
GS_19_1 0 NS_19 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 21/22
CS_21 NS_21 0 9.9999999999999998e-13
CS_22 NS_22 0 9.9999999999999998e-13
RS_21 NS_21 0 1.6005864146684806e+02
RS_22 NS_22 0 1.6005864146684809e+02
GL_21 0 NS_21 NS_22 0 2.5423900390253934e-01
GL_22 0 NS_22 NS_21 0 -2.5423900390253934e-01
GS_21_1 0 NS_21 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 23/24
CS_23 NS_23 0 9.9999999999999998e-13
CS_24 NS_24 0 9.9999999999999998e-13
RS_23 NS_23 0 1.9181463552142085e+02
RS_24 NS_24 0 1.9181463552142085e+02
GL_23 0 NS_23 NS_24 0 2.1188941693262670e-01
GL_24 0 NS_24 NS_23 0 -2.1188941693262670e-01
GS_23_1 0 NS_23 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 25/26
CS_25 NS_25 0 9.9999999999999998e-13
CS_26 NS_26 0 9.9999999999999998e-13
RS_25 NS_25 0 2.5689115313648813e+02
RS_26 NS_26 0 2.5689115313648813e+02
GL_25 0 NS_25 NS_26 0 2.1774212061821885e-01
GL_26 0 NS_26 NS_25 0 -2.1774212061821885e-01
GS_25_1 0 NS_25 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 27/28
CS_27 NS_27 0 9.9999999999999998e-13
CS_28 NS_28 0 9.9999999999999998e-13
RS_27 NS_27 0 6.2765149843829192e+01
RS_28 NS_28 0 6.2765149843829192e+01
GL_27 0 NS_27 NS_28 0 2.3246082537351351e-01
GL_28 0 NS_28 NS_27 0 -2.3246082537351351e-01
GS_27_1 0 NS_27 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 29/30
CS_29 NS_29 0 9.9999999999999998e-13
CS_30 NS_30 0 9.9999999999999998e-13
RS_29 NS_29 0 3.5419967361311882e+02
RS_30 NS_30 0 3.5419967361311882e+02
GL_29 0 NS_29 NS_30 0 2.2268031336810420e-01
GL_30 0 NS_30 NS_29 0 -2.2268031336810420e-01
GS_29_1 0 NS_29 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 31/32
CS_31 NS_31 0 9.9999999999999998e-13
CS_32 NS_32 0 9.9999999999999998e-13
RS_31 NS_31 0 9.0838548010669172e+01
RS_32 NS_32 0 9.0838548010669186e+01
GL_31 0 NS_31 NS_32 0 2.2647420085995260e-01
GL_32 0 NS_32 NS_31 0 -2.2647420085995260e-01
GS_31_1 0 NS_31 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 33/34
CS_33 NS_33 0 9.9999999999999998e-13
CS_34 NS_34 0 9.9999999999999998e-13
RS_33 NS_33 0 5.0298322136619066e+02
RS_34 NS_34 0 5.0298322136619078e+02
GL_33 0 NS_33 NS_34 0 2.4757175091537195e-01
GL_34 0 NS_34 NS_33 0 -2.4757175091537195e-01
GS_33_1 0 NS_33 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 35/36
CS_35 NS_35 0 9.9999999999999998e-13
CS_36 NS_36 0 9.9999999999999998e-13
RS_35 NS_35 0 1.1113846377285431e+02
RS_36 NS_36 0 1.1113846377285431e+02
GL_35 0 NS_35 NS_36 0 2.4529156966751164e-01
GL_36 0 NS_36 NS_35 0 -2.4529156966751164e-01
GS_35_1 0 NS_35 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 37/38
CS_37 NS_37 0 9.9999999999999998e-13
CS_38 NS_38 0 9.9999999999999998e-13
RS_37 NS_37 0 4.1132635267896995e+02
RS_38 NS_38 0 4.1132635267896990e+02
GL_37 0 NS_37 NS_38 0 2.4323159344727399e-01
GL_38 0 NS_38 NS_37 0 -2.4323159344727399e-01
GS_37_1 0 NS_37 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 39/40
CS_39 NS_39 0 9.9999999999999998e-13
CS_40 NS_40 0 9.9999999999999998e-13
RS_39 NS_39 0 6.1483243702508491e+02
RS_40 NS_40 0 6.1483243702508491e+02
GL_39 0 NS_39 NS_40 0 2.3313794138995145e-01
GL_40 0 NS_40 NS_39 0 -2.3313794138995145e-01
GS_39_1 0 NS_39 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 41/42
CS_41 NS_41 0 9.9999999999999998e-13
CS_42 NS_42 0 9.9999999999999998e-13
RS_41 NS_41 0 6.0708452252497170e+02
RS_42 NS_42 0 6.0708452252497170e+02
GL_41 0 NS_41 NS_42 0 2.3828547054015958e-01
GL_42 0 NS_42 NS_41 0 -2.3828547054015958e-01
GS_41_1 0 NS_41 NA_1 0 1.6921379288850509e+00
*
* Complex pair n. 43/44
CS_43 NS_43 0 9.9999999999999998e-13
CS_44 NS_44 0 9.9999999999999998e-13
RS_43 NS_43 0 1.9238303220034285e+02
RS_44 NS_44 0 1.9238303220034285e+02
GL_43 0 NS_43 NS_44 0 2.3639447764395666e-01
GL_44 0 NS_44 NS_43 0 -2.3639447764395666e-01
GS_43_1 0 NS_43 NA_1 0 1.6921379288850509e+00
*
* Real pole n. 45
CS_45 NS_45 0 9.9999999999999998e-13
RS_45 NS_45 0 1.2063458770185771e+00
GS_45_2 0 NS_45 NA_2 0 1.6921379288850509e+00
*
* Real pole n. 46
CS_46 NS_46 0 9.9999999999999998e-13
RS_46 NS_46 0 2.0414994648771170e+01
GS_46_2 0 NS_46 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 47/48
CS_47 NS_47 0 9.9999999999999998e-13
CS_48 NS_48 0 9.9999999999999998e-13
RS_47 NS_47 0 2.2164632983638530e+01
RS_48 NS_48 0 2.2164632983638530e+01
GL_47 0 NS_47 NS_48 0 6.2432580119989492e-02
GL_48 0 NS_48 NS_47 0 -6.2432580119989492e-02
GS_47_2 0 NS_47 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 49/50
CS_49 NS_49 0 9.9999999999999998e-13
CS_50 NS_50 0 9.9999999999999998e-13
RS_49 NS_49 0 2.4208144339458560e+01
RS_50 NS_50 0 2.4208144339458560e+01
GL_49 0 NS_49 NS_50 0 8.7759448763363015e-02
GL_50 0 NS_50 NS_49 0 -8.7759448763363015e-02
GS_49_2 0 NS_49 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 51/52
CS_51 NS_51 0 9.9999999999999998e-13
CS_52 NS_52 0 9.9999999999999998e-13
RS_51 NS_51 0 1.3097029666184031e+02
RS_52 NS_52 0 1.3097029666184031e+02
GL_51 0 NS_51 NS_52 0 2.9672291989323329e-01
GL_52 0 NS_52 NS_51 0 -2.9672291989323329e-01
GS_51_2 0 NS_51 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 53/54
CS_53 NS_53 0 9.9999999999999998e-13
CS_54 NS_54 0 9.9999999999999998e-13
RS_53 NS_53 0 3.2672536376024027e+01
RS_54 NS_54 0 3.2672536376024027e+01
GL_53 0 NS_53 NS_54 0 1.2489866711430768e-01
GL_54 0 NS_54 NS_53 0 -1.2489866711430768e-01
GS_53_2 0 NS_53 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 55/56
CS_55 NS_55 0 9.9999999999999998e-13
CS_56 NS_56 0 9.9999999999999998e-13
RS_55 NS_55 0 3.6741731246022816e+01
RS_56 NS_56 0 3.6741731246022816e+01
GL_55 0 NS_55 NS_56 0 1.6399845549232167e-01
GL_56 0 NS_56 NS_55 0 -1.6399845549232167e-01
GS_55_2 0 NS_55 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 57/58
CS_57 NS_57 0 9.9999999999999998e-13
CS_58 NS_58 0 9.9999999999999998e-13
RS_57 NS_57 0 8.3646036557163740e+01
RS_58 NS_58 0 8.3646036557163740e+01
GL_57 0 NS_57 NS_58 0 1.6830719130342967e-01
GL_58 0 NS_58 NS_57 0 -1.6830719130342967e-01
GS_57_2 0 NS_57 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 59/60
CS_59 NS_59 0 9.9999999999999998e-13
CS_60 NS_60 0 9.9999999999999998e-13
RS_59 NS_59 0 4.0307732865054554e+01
RS_60 NS_60 0 4.0307732865054554e+01
GL_59 0 NS_59 NS_60 0 1.8890575271706389e-01
GL_60 0 NS_60 NS_59 0 -1.8890575271706389e-01
GS_59_2 0 NS_59 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 61/62
CS_61 NS_61 0 9.9999999999999998e-13
CS_62 NS_62 0 9.9999999999999998e-13
RS_61 NS_61 0 1.4268073111996583e+02
RS_62 NS_62 0 1.4268073111996583e+02
GL_61 0 NS_61 NS_62 0 1.9419078929943706e-01
GL_62 0 NS_62 NS_61 0 -1.9419078929943706e-01
GS_61_2 0 NS_61 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 63/64
CS_63 NS_63 0 9.9999999999999998e-13
CS_64 NS_64 0 9.9999999999999998e-13
RS_63 NS_63 0 7.1679198821979867e+01
RS_64 NS_64 0 7.1679198821979867e+01
GL_63 0 NS_63 NS_64 0 2.0702628270375376e-01
GL_64 0 NS_64 NS_63 0 -2.0702628270375376e-01
GS_63_2 0 NS_63 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 65/66
CS_65 NS_65 0 9.9999999999999998e-13
CS_66 NS_66 0 9.9999999999999998e-13
RS_65 NS_65 0 1.6005864146684806e+02
RS_66 NS_66 0 1.6005864146684809e+02
GL_65 0 NS_65 NS_66 0 2.5423900390253934e-01
GL_66 0 NS_66 NS_65 0 -2.5423900390253934e-01
GS_65_2 0 NS_65 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 67/68
CS_67 NS_67 0 9.9999999999999998e-13
CS_68 NS_68 0 9.9999999999999998e-13
RS_67 NS_67 0 1.9181463552142085e+02
RS_68 NS_68 0 1.9181463552142085e+02
GL_67 0 NS_67 NS_68 0 2.1188941693262670e-01
GL_68 0 NS_68 NS_67 0 -2.1188941693262670e-01
GS_67_2 0 NS_67 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 69/70
CS_69 NS_69 0 9.9999999999999998e-13
CS_70 NS_70 0 9.9999999999999998e-13
RS_69 NS_69 0 2.5689115313648813e+02
RS_70 NS_70 0 2.5689115313648813e+02
GL_69 0 NS_69 NS_70 0 2.1774212061821885e-01
GL_70 0 NS_70 NS_69 0 -2.1774212061821885e-01
GS_69_2 0 NS_69 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 71/72
CS_71 NS_71 0 9.9999999999999998e-13
CS_72 NS_72 0 9.9999999999999998e-13
RS_71 NS_71 0 6.2765149843829192e+01
RS_72 NS_72 0 6.2765149843829192e+01
GL_71 0 NS_71 NS_72 0 2.3246082537351351e-01
GL_72 0 NS_72 NS_71 0 -2.3246082537351351e-01
GS_71_2 0 NS_71 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 73/74
CS_73 NS_73 0 9.9999999999999998e-13
CS_74 NS_74 0 9.9999999999999998e-13
RS_73 NS_73 0 3.5419967361311882e+02
RS_74 NS_74 0 3.5419967361311882e+02
GL_73 0 NS_73 NS_74 0 2.2268031336810420e-01
GL_74 0 NS_74 NS_73 0 -2.2268031336810420e-01
GS_73_2 0 NS_73 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 75/76
CS_75 NS_75 0 9.9999999999999998e-13
CS_76 NS_76 0 9.9999999999999998e-13
RS_75 NS_75 0 9.0838548010669172e+01
RS_76 NS_76 0 9.0838548010669186e+01
GL_75 0 NS_75 NS_76 0 2.2647420085995260e-01
GL_76 0 NS_76 NS_75 0 -2.2647420085995260e-01
GS_75_2 0 NS_75 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 77/78
CS_77 NS_77 0 9.9999999999999998e-13
CS_78 NS_78 0 9.9999999999999998e-13
RS_77 NS_77 0 5.0298322136619066e+02
RS_78 NS_78 0 5.0298322136619078e+02
GL_77 0 NS_77 NS_78 0 2.4757175091537195e-01
GL_78 0 NS_78 NS_77 0 -2.4757175091537195e-01
GS_77_2 0 NS_77 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 79/80
CS_79 NS_79 0 9.9999999999999998e-13
CS_80 NS_80 0 9.9999999999999998e-13
RS_79 NS_79 0 1.1113846377285431e+02
RS_80 NS_80 0 1.1113846377285431e+02
GL_79 0 NS_79 NS_80 0 2.4529156966751164e-01
GL_80 0 NS_80 NS_79 0 -2.4529156966751164e-01
GS_79_2 0 NS_79 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 81/82
CS_81 NS_81 0 9.9999999999999998e-13
CS_82 NS_82 0 9.9999999999999998e-13
RS_81 NS_81 0 4.1132635267896995e+02
RS_82 NS_82 0 4.1132635267896990e+02
GL_81 0 NS_81 NS_82 0 2.4323159344727399e-01
GL_82 0 NS_82 NS_81 0 -2.4323159344727399e-01
GS_81_2 0 NS_81 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 83/84
CS_83 NS_83 0 9.9999999999999998e-13
CS_84 NS_84 0 9.9999999999999998e-13
RS_83 NS_83 0 6.1483243702508491e+02
RS_84 NS_84 0 6.1483243702508491e+02
GL_83 0 NS_83 NS_84 0 2.3313794138995145e-01
GL_84 0 NS_84 NS_83 0 -2.3313794138995145e-01
GS_83_2 0 NS_83 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 85/86
CS_85 NS_85 0 9.9999999999999998e-13
CS_86 NS_86 0 9.9999999999999998e-13
RS_85 NS_85 0 6.0708452252497170e+02
RS_86 NS_86 0 6.0708452252497170e+02
GL_85 0 NS_85 NS_86 0 2.3828547054015958e-01
GL_86 0 NS_86 NS_85 0 -2.3828547054015958e-01
GS_85_2 0 NS_85 NA_2 0 1.6921379288850509e+00
*
* Complex pair n. 87/88
CS_87 NS_87 0 9.9999999999999998e-13
CS_88 NS_88 0 9.9999999999999998e-13
RS_87 NS_87 0 1.9238303220034285e+02
RS_88 NS_88 0 1.9238303220034285e+02
GL_87 0 NS_87 NS_88 0 2.3639447764395666e-01
GL_88 0 NS_88 NS_87 0 -2.3639447764395666e-01
GS_87_2 0 NS_87 NA_2 0 1.6921379288850509e+00
*
* Real pole n. 89
CS_89 NS_89 0 9.9999999999999998e-13
RS_89 NS_89 0 1.2063458770185771e+00
GS_89_3 0 NS_89 NA_3 0 1.6921379288850509e+00
*
* Real pole n. 90
CS_90 NS_90 0 9.9999999999999998e-13
RS_90 NS_90 0 2.0414994648771170e+01
GS_90_3 0 NS_90 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 91/92
CS_91 NS_91 0 9.9999999999999998e-13
CS_92 NS_92 0 9.9999999999999998e-13
RS_91 NS_91 0 2.2164632983638530e+01
RS_92 NS_92 0 2.2164632983638530e+01
GL_91 0 NS_91 NS_92 0 6.2432580119989492e-02
GL_92 0 NS_92 NS_91 0 -6.2432580119989492e-02
GS_91_3 0 NS_91 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 93/94
CS_93 NS_93 0 9.9999999999999998e-13
CS_94 NS_94 0 9.9999999999999998e-13
RS_93 NS_93 0 2.4208144339458560e+01
RS_94 NS_94 0 2.4208144339458560e+01
GL_93 0 NS_93 NS_94 0 8.7759448763363015e-02
GL_94 0 NS_94 NS_93 0 -8.7759448763363015e-02
GS_93_3 0 NS_93 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 95/96
CS_95 NS_95 0 9.9999999999999998e-13
CS_96 NS_96 0 9.9999999999999998e-13
RS_95 NS_95 0 1.3097029666184031e+02
RS_96 NS_96 0 1.3097029666184031e+02
GL_95 0 NS_95 NS_96 0 2.9672291989323329e-01
GL_96 0 NS_96 NS_95 0 -2.9672291989323329e-01
GS_95_3 0 NS_95 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 97/98
CS_97 NS_97 0 9.9999999999999998e-13
CS_98 NS_98 0 9.9999999999999998e-13
RS_97 NS_97 0 3.2672536376024027e+01
RS_98 NS_98 0 3.2672536376024027e+01
GL_97 0 NS_97 NS_98 0 1.2489866711430768e-01
GL_98 0 NS_98 NS_97 0 -1.2489866711430768e-01
GS_97_3 0 NS_97 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 99/100
CS_99 NS_99 0 9.9999999999999998e-13
CS_100 NS_100 0 9.9999999999999998e-13
RS_99 NS_99 0 3.6741731246022816e+01
RS_100 NS_100 0 3.6741731246022816e+01
GL_99 0 NS_99 NS_100 0 1.6399845549232167e-01
GL_100 0 NS_100 NS_99 0 -1.6399845549232167e-01
GS_99_3 0 NS_99 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 101/102
CS_101 NS_101 0 9.9999999999999998e-13
CS_102 NS_102 0 9.9999999999999998e-13
RS_101 NS_101 0 8.3646036557163740e+01
RS_102 NS_102 0 8.3646036557163740e+01
GL_101 0 NS_101 NS_102 0 1.6830719130342967e-01
GL_102 0 NS_102 NS_101 0 -1.6830719130342967e-01
GS_101_3 0 NS_101 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 103/104
CS_103 NS_103 0 9.9999999999999998e-13
CS_104 NS_104 0 9.9999999999999998e-13
RS_103 NS_103 0 4.0307732865054554e+01
RS_104 NS_104 0 4.0307732865054554e+01
GL_103 0 NS_103 NS_104 0 1.8890575271706389e-01
GL_104 0 NS_104 NS_103 0 -1.8890575271706389e-01
GS_103_3 0 NS_103 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 105/106
CS_105 NS_105 0 9.9999999999999998e-13
CS_106 NS_106 0 9.9999999999999998e-13
RS_105 NS_105 0 1.4268073111996583e+02
RS_106 NS_106 0 1.4268073111996583e+02
GL_105 0 NS_105 NS_106 0 1.9419078929943706e-01
GL_106 0 NS_106 NS_105 0 -1.9419078929943706e-01
GS_105_3 0 NS_105 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 107/108
CS_107 NS_107 0 9.9999999999999998e-13
CS_108 NS_108 0 9.9999999999999998e-13
RS_107 NS_107 0 7.1679198821979867e+01
RS_108 NS_108 0 7.1679198821979867e+01
GL_107 0 NS_107 NS_108 0 2.0702628270375376e-01
GL_108 0 NS_108 NS_107 0 -2.0702628270375376e-01
GS_107_3 0 NS_107 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 109/110
CS_109 NS_109 0 9.9999999999999998e-13
CS_110 NS_110 0 9.9999999999999998e-13
RS_109 NS_109 0 1.6005864146684806e+02
RS_110 NS_110 0 1.6005864146684809e+02
GL_109 0 NS_109 NS_110 0 2.5423900390253934e-01
GL_110 0 NS_110 NS_109 0 -2.5423900390253934e-01
GS_109_3 0 NS_109 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 111/112
CS_111 NS_111 0 9.9999999999999998e-13
CS_112 NS_112 0 9.9999999999999998e-13
RS_111 NS_111 0 1.9181463552142085e+02
RS_112 NS_112 0 1.9181463552142085e+02
GL_111 0 NS_111 NS_112 0 2.1188941693262670e-01
GL_112 0 NS_112 NS_111 0 -2.1188941693262670e-01
GS_111_3 0 NS_111 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 113/114
CS_113 NS_113 0 9.9999999999999998e-13
CS_114 NS_114 0 9.9999999999999998e-13
RS_113 NS_113 0 2.5689115313648813e+02
RS_114 NS_114 0 2.5689115313648813e+02
GL_113 0 NS_113 NS_114 0 2.1774212061821885e-01
GL_114 0 NS_114 NS_113 0 -2.1774212061821885e-01
GS_113_3 0 NS_113 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 115/116
CS_115 NS_115 0 9.9999999999999998e-13
CS_116 NS_116 0 9.9999999999999998e-13
RS_115 NS_115 0 6.2765149843829192e+01
RS_116 NS_116 0 6.2765149843829192e+01
GL_115 0 NS_115 NS_116 0 2.3246082537351351e-01
GL_116 0 NS_116 NS_115 0 -2.3246082537351351e-01
GS_115_3 0 NS_115 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 117/118
CS_117 NS_117 0 9.9999999999999998e-13
CS_118 NS_118 0 9.9999999999999998e-13
RS_117 NS_117 0 3.5419967361311882e+02
RS_118 NS_118 0 3.5419967361311882e+02
GL_117 0 NS_117 NS_118 0 2.2268031336810420e-01
GL_118 0 NS_118 NS_117 0 -2.2268031336810420e-01
GS_117_3 0 NS_117 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 119/120
CS_119 NS_119 0 9.9999999999999998e-13
CS_120 NS_120 0 9.9999999999999998e-13
RS_119 NS_119 0 9.0838548010669172e+01
RS_120 NS_120 0 9.0838548010669186e+01
GL_119 0 NS_119 NS_120 0 2.2647420085995260e-01
GL_120 0 NS_120 NS_119 0 -2.2647420085995260e-01
GS_119_3 0 NS_119 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 121/122
CS_121 NS_121 0 9.9999999999999998e-13
CS_122 NS_122 0 9.9999999999999998e-13
RS_121 NS_121 0 5.0298322136619066e+02
RS_122 NS_122 0 5.0298322136619078e+02
GL_121 0 NS_121 NS_122 0 2.4757175091537195e-01
GL_122 0 NS_122 NS_121 0 -2.4757175091537195e-01
GS_121_3 0 NS_121 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 123/124
CS_123 NS_123 0 9.9999999999999998e-13
CS_124 NS_124 0 9.9999999999999998e-13
RS_123 NS_123 0 1.1113846377285431e+02
RS_124 NS_124 0 1.1113846377285431e+02
GL_123 0 NS_123 NS_124 0 2.4529156966751164e-01
GL_124 0 NS_124 NS_123 0 -2.4529156966751164e-01
GS_123_3 0 NS_123 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 125/126
CS_125 NS_125 0 9.9999999999999998e-13
CS_126 NS_126 0 9.9999999999999998e-13
RS_125 NS_125 0 4.1132635267896995e+02
RS_126 NS_126 0 4.1132635267896990e+02
GL_125 0 NS_125 NS_126 0 2.4323159344727399e-01
GL_126 0 NS_126 NS_125 0 -2.4323159344727399e-01
GS_125_3 0 NS_125 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 127/128
CS_127 NS_127 0 9.9999999999999998e-13
CS_128 NS_128 0 9.9999999999999998e-13
RS_127 NS_127 0 6.1483243702508491e+02
RS_128 NS_128 0 6.1483243702508491e+02
GL_127 0 NS_127 NS_128 0 2.3313794138995145e-01
GL_128 0 NS_128 NS_127 0 -2.3313794138995145e-01
GS_127_3 0 NS_127 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 129/130
CS_129 NS_129 0 9.9999999999999998e-13
CS_130 NS_130 0 9.9999999999999998e-13
RS_129 NS_129 0 6.0708452252497170e+02
RS_130 NS_130 0 6.0708452252497170e+02
GL_129 0 NS_129 NS_130 0 2.3828547054015958e-01
GL_130 0 NS_130 NS_129 0 -2.3828547054015958e-01
GS_129_3 0 NS_129 NA_3 0 1.6921379288850509e+00
*
* Complex pair n. 131/132
CS_131 NS_131 0 9.9999999999999998e-13
CS_132 NS_132 0 9.9999999999999998e-13
RS_131 NS_131 0 1.9238303220034285e+02
RS_132 NS_132 0 1.9238303220034285e+02
GL_131 0 NS_131 NS_132 0 2.3639447764395666e-01
GL_132 0 NS_132 NS_131 0 -2.3639447764395666e-01
GS_131_3 0 NS_131 NA_3 0 1.6921379288850509e+00
*
* Real pole n. 133
CS_133 NS_133 0 9.9999999999999998e-13
RS_133 NS_133 0 1.2063458770185771e+00
GS_133_4 0 NS_133 NA_4 0 1.6921379288850509e+00
*
* Real pole n. 134
CS_134 NS_134 0 9.9999999999999998e-13
RS_134 NS_134 0 2.0414994648771170e+01
GS_134_4 0 NS_134 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 135/136
CS_135 NS_135 0 9.9999999999999998e-13
CS_136 NS_136 0 9.9999999999999998e-13
RS_135 NS_135 0 2.2164632983638530e+01
RS_136 NS_136 0 2.2164632983638530e+01
GL_135 0 NS_135 NS_136 0 6.2432580119989492e-02
GL_136 0 NS_136 NS_135 0 -6.2432580119989492e-02
GS_135_4 0 NS_135 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 137/138
CS_137 NS_137 0 9.9999999999999998e-13
CS_138 NS_138 0 9.9999999999999998e-13
RS_137 NS_137 0 2.4208144339458560e+01
RS_138 NS_138 0 2.4208144339458560e+01
GL_137 0 NS_137 NS_138 0 8.7759448763363015e-02
GL_138 0 NS_138 NS_137 0 -8.7759448763363015e-02
GS_137_4 0 NS_137 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 139/140
CS_139 NS_139 0 9.9999999999999998e-13
CS_140 NS_140 0 9.9999999999999998e-13
RS_139 NS_139 0 1.3097029666184031e+02
RS_140 NS_140 0 1.3097029666184031e+02
GL_139 0 NS_139 NS_140 0 2.9672291989323329e-01
GL_140 0 NS_140 NS_139 0 -2.9672291989323329e-01
GS_139_4 0 NS_139 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 141/142
CS_141 NS_141 0 9.9999999999999998e-13
CS_142 NS_142 0 9.9999999999999998e-13
RS_141 NS_141 0 3.2672536376024027e+01
RS_142 NS_142 0 3.2672536376024027e+01
GL_141 0 NS_141 NS_142 0 1.2489866711430768e-01
GL_142 0 NS_142 NS_141 0 -1.2489866711430768e-01
GS_141_4 0 NS_141 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 143/144
CS_143 NS_143 0 9.9999999999999998e-13
CS_144 NS_144 0 9.9999999999999998e-13
RS_143 NS_143 0 3.6741731246022816e+01
RS_144 NS_144 0 3.6741731246022816e+01
GL_143 0 NS_143 NS_144 0 1.6399845549232167e-01
GL_144 0 NS_144 NS_143 0 -1.6399845549232167e-01
GS_143_4 0 NS_143 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 145/146
CS_145 NS_145 0 9.9999999999999998e-13
CS_146 NS_146 0 9.9999999999999998e-13
RS_145 NS_145 0 8.3646036557163740e+01
RS_146 NS_146 0 8.3646036557163740e+01
GL_145 0 NS_145 NS_146 0 1.6830719130342967e-01
GL_146 0 NS_146 NS_145 0 -1.6830719130342967e-01
GS_145_4 0 NS_145 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 147/148
CS_147 NS_147 0 9.9999999999999998e-13
CS_148 NS_148 0 9.9999999999999998e-13
RS_147 NS_147 0 4.0307732865054554e+01
RS_148 NS_148 0 4.0307732865054554e+01
GL_147 0 NS_147 NS_148 0 1.8890575271706389e-01
GL_148 0 NS_148 NS_147 0 -1.8890575271706389e-01
GS_147_4 0 NS_147 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 149/150
CS_149 NS_149 0 9.9999999999999998e-13
CS_150 NS_150 0 9.9999999999999998e-13
RS_149 NS_149 0 1.4268073111996583e+02
RS_150 NS_150 0 1.4268073111996583e+02
GL_149 0 NS_149 NS_150 0 1.9419078929943706e-01
GL_150 0 NS_150 NS_149 0 -1.9419078929943706e-01
GS_149_4 0 NS_149 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 151/152
CS_151 NS_151 0 9.9999999999999998e-13
CS_152 NS_152 0 9.9999999999999998e-13
RS_151 NS_151 0 7.1679198821979867e+01
RS_152 NS_152 0 7.1679198821979867e+01
GL_151 0 NS_151 NS_152 0 2.0702628270375376e-01
GL_152 0 NS_152 NS_151 0 -2.0702628270375376e-01
GS_151_4 0 NS_151 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 153/154
CS_153 NS_153 0 9.9999999999999998e-13
CS_154 NS_154 0 9.9999999999999998e-13
RS_153 NS_153 0 1.6005864146684806e+02
RS_154 NS_154 0 1.6005864146684809e+02
GL_153 0 NS_153 NS_154 0 2.5423900390253934e-01
GL_154 0 NS_154 NS_153 0 -2.5423900390253934e-01
GS_153_4 0 NS_153 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 155/156
CS_155 NS_155 0 9.9999999999999998e-13
CS_156 NS_156 0 9.9999999999999998e-13
RS_155 NS_155 0 1.9181463552142085e+02
RS_156 NS_156 0 1.9181463552142085e+02
GL_155 0 NS_155 NS_156 0 2.1188941693262670e-01
GL_156 0 NS_156 NS_155 0 -2.1188941693262670e-01
GS_155_4 0 NS_155 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 157/158
CS_157 NS_157 0 9.9999999999999998e-13
CS_158 NS_158 0 9.9999999999999998e-13
RS_157 NS_157 0 2.5689115313648813e+02
RS_158 NS_158 0 2.5689115313648813e+02
GL_157 0 NS_157 NS_158 0 2.1774212061821885e-01
GL_158 0 NS_158 NS_157 0 -2.1774212061821885e-01
GS_157_4 0 NS_157 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 159/160
CS_159 NS_159 0 9.9999999999999998e-13
CS_160 NS_160 0 9.9999999999999998e-13
RS_159 NS_159 0 6.2765149843829192e+01
RS_160 NS_160 0 6.2765149843829192e+01
GL_159 0 NS_159 NS_160 0 2.3246082537351351e-01
GL_160 0 NS_160 NS_159 0 -2.3246082537351351e-01
GS_159_4 0 NS_159 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 161/162
CS_161 NS_161 0 9.9999999999999998e-13
CS_162 NS_162 0 9.9999999999999998e-13
RS_161 NS_161 0 3.5419967361311882e+02
RS_162 NS_162 0 3.5419967361311882e+02
GL_161 0 NS_161 NS_162 0 2.2268031336810420e-01
GL_162 0 NS_162 NS_161 0 -2.2268031336810420e-01
GS_161_4 0 NS_161 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 163/164
CS_163 NS_163 0 9.9999999999999998e-13
CS_164 NS_164 0 9.9999999999999998e-13
RS_163 NS_163 0 9.0838548010669172e+01
RS_164 NS_164 0 9.0838548010669186e+01
GL_163 0 NS_163 NS_164 0 2.2647420085995260e-01
GL_164 0 NS_164 NS_163 0 -2.2647420085995260e-01
GS_163_4 0 NS_163 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 165/166
CS_165 NS_165 0 9.9999999999999998e-13
CS_166 NS_166 0 9.9999999999999998e-13
RS_165 NS_165 0 5.0298322136619066e+02
RS_166 NS_166 0 5.0298322136619078e+02
GL_165 0 NS_165 NS_166 0 2.4757175091537195e-01
GL_166 0 NS_166 NS_165 0 -2.4757175091537195e-01
GS_165_4 0 NS_165 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 167/168
CS_167 NS_167 0 9.9999999999999998e-13
CS_168 NS_168 0 9.9999999999999998e-13
RS_167 NS_167 0 1.1113846377285431e+02
RS_168 NS_168 0 1.1113846377285431e+02
GL_167 0 NS_167 NS_168 0 2.4529156966751164e-01
GL_168 0 NS_168 NS_167 0 -2.4529156966751164e-01
GS_167_4 0 NS_167 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 169/170
CS_169 NS_169 0 9.9999999999999998e-13
CS_170 NS_170 0 9.9999999999999998e-13
RS_169 NS_169 0 4.1132635267896995e+02
RS_170 NS_170 0 4.1132635267896990e+02
GL_169 0 NS_169 NS_170 0 2.4323159344727399e-01
GL_170 0 NS_170 NS_169 0 -2.4323159344727399e-01
GS_169_4 0 NS_169 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 171/172
CS_171 NS_171 0 9.9999999999999998e-13
CS_172 NS_172 0 9.9999999999999998e-13
RS_171 NS_171 0 6.1483243702508491e+02
RS_172 NS_172 0 6.1483243702508491e+02
GL_171 0 NS_171 NS_172 0 2.3313794138995145e-01
GL_172 0 NS_172 NS_171 0 -2.3313794138995145e-01
GS_171_4 0 NS_171 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 173/174
CS_173 NS_173 0 9.9999999999999998e-13
CS_174 NS_174 0 9.9999999999999998e-13
RS_173 NS_173 0 6.0708452252497170e+02
RS_174 NS_174 0 6.0708452252497170e+02
GL_173 0 NS_173 NS_174 0 2.3828547054015958e-01
GL_174 0 NS_174 NS_173 0 -2.3828547054015958e-01
GS_173_4 0 NS_173 NA_4 0 1.6921379288850509e+00
*
* Complex pair n. 175/176
CS_175 NS_175 0 9.9999999999999998e-13
CS_176 NS_176 0 9.9999999999999998e-13
RS_175 NS_175 0 1.9238303220034285e+02
RS_176 NS_176 0 1.9238303220034285e+02
GL_175 0 NS_175 NS_176 0 2.3639447764395666e-01
GL_176 0 NS_176 NS_175 0 -2.3639447764395666e-01
GS_175_4 0 NS_175 NA_4 0 1.6921379288850509e+00
*
* Real pole n. 177
CS_177 NS_177 0 9.9999999999999998e-13
RS_177 NS_177 0 1.2063458770185771e+00
GS_177_5 0 NS_177 NA_5 0 1.6921379288850509e+00
*
* Real pole n. 178
CS_178 NS_178 0 9.9999999999999998e-13
RS_178 NS_178 0 2.0414994648771170e+01
GS_178_5 0 NS_178 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 179/180
CS_179 NS_179 0 9.9999999999999998e-13
CS_180 NS_180 0 9.9999999999999998e-13
RS_179 NS_179 0 2.2164632983638530e+01
RS_180 NS_180 0 2.2164632983638530e+01
GL_179 0 NS_179 NS_180 0 6.2432580119989492e-02
GL_180 0 NS_180 NS_179 0 -6.2432580119989492e-02
GS_179_5 0 NS_179 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 181/182
CS_181 NS_181 0 9.9999999999999998e-13
CS_182 NS_182 0 9.9999999999999998e-13
RS_181 NS_181 0 2.4208144339458560e+01
RS_182 NS_182 0 2.4208144339458560e+01
GL_181 0 NS_181 NS_182 0 8.7759448763363015e-02
GL_182 0 NS_182 NS_181 0 -8.7759448763363015e-02
GS_181_5 0 NS_181 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 183/184
CS_183 NS_183 0 9.9999999999999998e-13
CS_184 NS_184 0 9.9999999999999998e-13
RS_183 NS_183 0 1.3097029666184031e+02
RS_184 NS_184 0 1.3097029666184031e+02
GL_183 0 NS_183 NS_184 0 2.9672291989323329e-01
GL_184 0 NS_184 NS_183 0 -2.9672291989323329e-01
GS_183_5 0 NS_183 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 185/186
CS_185 NS_185 0 9.9999999999999998e-13
CS_186 NS_186 0 9.9999999999999998e-13
RS_185 NS_185 0 3.2672536376024027e+01
RS_186 NS_186 0 3.2672536376024027e+01
GL_185 0 NS_185 NS_186 0 1.2489866711430768e-01
GL_186 0 NS_186 NS_185 0 -1.2489866711430768e-01
GS_185_5 0 NS_185 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 187/188
CS_187 NS_187 0 9.9999999999999998e-13
CS_188 NS_188 0 9.9999999999999998e-13
RS_187 NS_187 0 3.6741731246022816e+01
RS_188 NS_188 0 3.6741731246022816e+01
GL_187 0 NS_187 NS_188 0 1.6399845549232167e-01
GL_188 0 NS_188 NS_187 0 -1.6399845549232167e-01
GS_187_5 0 NS_187 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 189/190
CS_189 NS_189 0 9.9999999999999998e-13
CS_190 NS_190 0 9.9999999999999998e-13
RS_189 NS_189 0 8.3646036557163740e+01
RS_190 NS_190 0 8.3646036557163740e+01
GL_189 0 NS_189 NS_190 0 1.6830719130342967e-01
GL_190 0 NS_190 NS_189 0 -1.6830719130342967e-01
GS_189_5 0 NS_189 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 191/192
CS_191 NS_191 0 9.9999999999999998e-13
CS_192 NS_192 0 9.9999999999999998e-13
RS_191 NS_191 0 4.0307732865054554e+01
RS_192 NS_192 0 4.0307732865054554e+01
GL_191 0 NS_191 NS_192 0 1.8890575271706389e-01
GL_192 0 NS_192 NS_191 0 -1.8890575271706389e-01
GS_191_5 0 NS_191 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 193/194
CS_193 NS_193 0 9.9999999999999998e-13
CS_194 NS_194 0 9.9999999999999998e-13
RS_193 NS_193 0 1.4268073111996583e+02
RS_194 NS_194 0 1.4268073111996583e+02
GL_193 0 NS_193 NS_194 0 1.9419078929943706e-01
GL_194 0 NS_194 NS_193 0 -1.9419078929943706e-01
GS_193_5 0 NS_193 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 195/196
CS_195 NS_195 0 9.9999999999999998e-13
CS_196 NS_196 0 9.9999999999999998e-13
RS_195 NS_195 0 7.1679198821979867e+01
RS_196 NS_196 0 7.1679198821979867e+01
GL_195 0 NS_195 NS_196 0 2.0702628270375376e-01
GL_196 0 NS_196 NS_195 0 -2.0702628270375376e-01
GS_195_5 0 NS_195 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 197/198
CS_197 NS_197 0 9.9999999999999998e-13
CS_198 NS_198 0 9.9999999999999998e-13
RS_197 NS_197 0 1.6005864146684806e+02
RS_198 NS_198 0 1.6005864146684809e+02
GL_197 0 NS_197 NS_198 0 2.5423900390253934e-01
GL_198 0 NS_198 NS_197 0 -2.5423900390253934e-01
GS_197_5 0 NS_197 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 199/200
CS_199 NS_199 0 9.9999999999999998e-13
CS_200 NS_200 0 9.9999999999999998e-13
RS_199 NS_199 0 1.9181463552142085e+02
RS_200 NS_200 0 1.9181463552142085e+02
GL_199 0 NS_199 NS_200 0 2.1188941693262670e-01
GL_200 0 NS_200 NS_199 0 -2.1188941693262670e-01
GS_199_5 0 NS_199 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 201/202
CS_201 NS_201 0 9.9999999999999998e-13
CS_202 NS_202 0 9.9999999999999998e-13
RS_201 NS_201 0 2.5689115313648813e+02
RS_202 NS_202 0 2.5689115313648813e+02
GL_201 0 NS_201 NS_202 0 2.1774212061821885e-01
GL_202 0 NS_202 NS_201 0 -2.1774212061821885e-01
GS_201_5 0 NS_201 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 203/204
CS_203 NS_203 0 9.9999999999999998e-13
CS_204 NS_204 0 9.9999999999999998e-13
RS_203 NS_203 0 6.2765149843829192e+01
RS_204 NS_204 0 6.2765149843829192e+01
GL_203 0 NS_203 NS_204 0 2.3246082537351351e-01
GL_204 0 NS_204 NS_203 0 -2.3246082537351351e-01
GS_203_5 0 NS_203 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 205/206
CS_205 NS_205 0 9.9999999999999998e-13
CS_206 NS_206 0 9.9999999999999998e-13
RS_205 NS_205 0 3.5419967361311882e+02
RS_206 NS_206 0 3.5419967361311882e+02
GL_205 0 NS_205 NS_206 0 2.2268031336810420e-01
GL_206 0 NS_206 NS_205 0 -2.2268031336810420e-01
GS_205_5 0 NS_205 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 207/208
CS_207 NS_207 0 9.9999999999999998e-13
CS_208 NS_208 0 9.9999999999999998e-13
RS_207 NS_207 0 9.0838548010669172e+01
RS_208 NS_208 0 9.0838548010669186e+01
GL_207 0 NS_207 NS_208 0 2.2647420085995260e-01
GL_208 0 NS_208 NS_207 0 -2.2647420085995260e-01
GS_207_5 0 NS_207 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 209/210
CS_209 NS_209 0 9.9999999999999998e-13
CS_210 NS_210 0 9.9999999999999998e-13
RS_209 NS_209 0 5.0298322136619066e+02
RS_210 NS_210 0 5.0298322136619078e+02
GL_209 0 NS_209 NS_210 0 2.4757175091537195e-01
GL_210 0 NS_210 NS_209 0 -2.4757175091537195e-01
GS_209_5 0 NS_209 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 211/212
CS_211 NS_211 0 9.9999999999999998e-13
CS_212 NS_212 0 9.9999999999999998e-13
RS_211 NS_211 0 1.1113846377285431e+02
RS_212 NS_212 0 1.1113846377285431e+02
GL_211 0 NS_211 NS_212 0 2.4529156966751164e-01
GL_212 0 NS_212 NS_211 0 -2.4529156966751164e-01
GS_211_5 0 NS_211 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 213/214
CS_213 NS_213 0 9.9999999999999998e-13
CS_214 NS_214 0 9.9999999999999998e-13
RS_213 NS_213 0 4.1132635267896995e+02
RS_214 NS_214 0 4.1132635267896990e+02
GL_213 0 NS_213 NS_214 0 2.4323159344727399e-01
GL_214 0 NS_214 NS_213 0 -2.4323159344727399e-01
GS_213_5 0 NS_213 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 215/216
CS_215 NS_215 0 9.9999999999999998e-13
CS_216 NS_216 0 9.9999999999999998e-13
RS_215 NS_215 0 6.1483243702508491e+02
RS_216 NS_216 0 6.1483243702508491e+02
GL_215 0 NS_215 NS_216 0 2.3313794138995145e-01
GL_216 0 NS_216 NS_215 0 -2.3313794138995145e-01
GS_215_5 0 NS_215 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 217/218
CS_217 NS_217 0 9.9999999999999998e-13
CS_218 NS_218 0 9.9999999999999998e-13
RS_217 NS_217 0 6.0708452252497170e+02
RS_218 NS_218 0 6.0708452252497170e+02
GL_217 0 NS_217 NS_218 0 2.3828547054015958e-01
GL_218 0 NS_218 NS_217 0 -2.3828547054015958e-01
GS_217_5 0 NS_217 NA_5 0 1.6921379288850509e+00
*
* Complex pair n. 219/220
CS_219 NS_219 0 9.9999999999999998e-13
CS_220 NS_220 0 9.9999999999999998e-13
RS_219 NS_219 0 1.9238303220034285e+02
RS_220 NS_220 0 1.9238303220034285e+02
GL_219 0 NS_219 NS_220 0 2.3639447764395666e-01
GL_220 0 NS_220 NS_219 0 -2.3639447764395666e-01
GS_219_5 0 NS_219 NA_5 0 1.6921379288850509e+00
*
* Real pole n. 221
CS_221 NS_221 0 9.9999999999999998e-13
RS_221 NS_221 0 1.2063458770185771e+00
GS_221_6 0 NS_221 NA_6 0 1.6921379288850509e+00
*
* Real pole n. 222
CS_222 NS_222 0 9.9999999999999998e-13
RS_222 NS_222 0 2.0414994648771170e+01
GS_222_6 0 NS_222 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 223/224
CS_223 NS_223 0 9.9999999999999998e-13
CS_224 NS_224 0 9.9999999999999998e-13
RS_223 NS_223 0 2.2164632983638530e+01
RS_224 NS_224 0 2.2164632983638530e+01
GL_223 0 NS_223 NS_224 0 6.2432580119989492e-02
GL_224 0 NS_224 NS_223 0 -6.2432580119989492e-02
GS_223_6 0 NS_223 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 225/226
CS_225 NS_225 0 9.9999999999999998e-13
CS_226 NS_226 0 9.9999999999999998e-13
RS_225 NS_225 0 2.4208144339458560e+01
RS_226 NS_226 0 2.4208144339458560e+01
GL_225 0 NS_225 NS_226 0 8.7759448763363015e-02
GL_226 0 NS_226 NS_225 0 -8.7759448763363015e-02
GS_225_6 0 NS_225 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 227/228
CS_227 NS_227 0 9.9999999999999998e-13
CS_228 NS_228 0 9.9999999999999998e-13
RS_227 NS_227 0 1.3097029666184031e+02
RS_228 NS_228 0 1.3097029666184031e+02
GL_227 0 NS_227 NS_228 0 2.9672291989323329e-01
GL_228 0 NS_228 NS_227 0 -2.9672291989323329e-01
GS_227_6 0 NS_227 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 229/230
CS_229 NS_229 0 9.9999999999999998e-13
CS_230 NS_230 0 9.9999999999999998e-13
RS_229 NS_229 0 3.2672536376024027e+01
RS_230 NS_230 0 3.2672536376024027e+01
GL_229 0 NS_229 NS_230 0 1.2489866711430768e-01
GL_230 0 NS_230 NS_229 0 -1.2489866711430768e-01
GS_229_6 0 NS_229 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 231/232
CS_231 NS_231 0 9.9999999999999998e-13
CS_232 NS_232 0 9.9999999999999998e-13
RS_231 NS_231 0 3.6741731246022816e+01
RS_232 NS_232 0 3.6741731246022816e+01
GL_231 0 NS_231 NS_232 0 1.6399845549232167e-01
GL_232 0 NS_232 NS_231 0 -1.6399845549232167e-01
GS_231_6 0 NS_231 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 233/234
CS_233 NS_233 0 9.9999999999999998e-13
CS_234 NS_234 0 9.9999999999999998e-13
RS_233 NS_233 0 8.3646036557163740e+01
RS_234 NS_234 0 8.3646036557163740e+01
GL_233 0 NS_233 NS_234 0 1.6830719130342967e-01
GL_234 0 NS_234 NS_233 0 -1.6830719130342967e-01
GS_233_6 0 NS_233 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 235/236
CS_235 NS_235 0 9.9999999999999998e-13
CS_236 NS_236 0 9.9999999999999998e-13
RS_235 NS_235 0 4.0307732865054554e+01
RS_236 NS_236 0 4.0307732865054554e+01
GL_235 0 NS_235 NS_236 0 1.8890575271706389e-01
GL_236 0 NS_236 NS_235 0 -1.8890575271706389e-01
GS_235_6 0 NS_235 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 237/238
CS_237 NS_237 0 9.9999999999999998e-13
CS_238 NS_238 0 9.9999999999999998e-13
RS_237 NS_237 0 1.4268073111996583e+02
RS_238 NS_238 0 1.4268073111996583e+02
GL_237 0 NS_237 NS_238 0 1.9419078929943706e-01
GL_238 0 NS_238 NS_237 0 -1.9419078929943706e-01
GS_237_6 0 NS_237 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 239/240
CS_239 NS_239 0 9.9999999999999998e-13
CS_240 NS_240 0 9.9999999999999998e-13
RS_239 NS_239 0 7.1679198821979867e+01
RS_240 NS_240 0 7.1679198821979867e+01
GL_239 0 NS_239 NS_240 0 2.0702628270375376e-01
GL_240 0 NS_240 NS_239 0 -2.0702628270375376e-01
GS_239_6 0 NS_239 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 241/242
CS_241 NS_241 0 9.9999999999999998e-13
CS_242 NS_242 0 9.9999999999999998e-13
RS_241 NS_241 0 1.6005864146684806e+02
RS_242 NS_242 0 1.6005864146684809e+02
GL_241 0 NS_241 NS_242 0 2.5423900390253934e-01
GL_242 0 NS_242 NS_241 0 -2.5423900390253934e-01
GS_241_6 0 NS_241 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 243/244
CS_243 NS_243 0 9.9999999999999998e-13
CS_244 NS_244 0 9.9999999999999998e-13
RS_243 NS_243 0 1.9181463552142085e+02
RS_244 NS_244 0 1.9181463552142085e+02
GL_243 0 NS_243 NS_244 0 2.1188941693262670e-01
GL_244 0 NS_244 NS_243 0 -2.1188941693262670e-01
GS_243_6 0 NS_243 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 245/246
CS_245 NS_245 0 9.9999999999999998e-13
CS_246 NS_246 0 9.9999999999999998e-13
RS_245 NS_245 0 2.5689115313648813e+02
RS_246 NS_246 0 2.5689115313648813e+02
GL_245 0 NS_245 NS_246 0 2.1774212061821885e-01
GL_246 0 NS_246 NS_245 0 -2.1774212061821885e-01
GS_245_6 0 NS_245 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 247/248
CS_247 NS_247 0 9.9999999999999998e-13
CS_248 NS_248 0 9.9999999999999998e-13
RS_247 NS_247 0 6.2765149843829192e+01
RS_248 NS_248 0 6.2765149843829192e+01
GL_247 0 NS_247 NS_248 0 2.3246082537351351e-01
GL_248 0 NS_248 NS_247 0 -2.3246082537351351e-01
GS_247_6 0 NS_247 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 249/250
CS_249 NS_249 0 9.9999999999999998e-13
CS_250 NS_250 0 9.9999999999999998e-13
RS_249 NS_249 0 3.5419967361311882e+02
RS_250 NS_250 0 3.5419967361311882e+02
GL_249 0 NS_249 NS_250 0 2.2268031336810420e-01
GL_250 0 NS_250 NS_249 0 -2.2268031336810420e-01
GS_249_6 0 NS_249 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 251/252
CS_251 NS_251 0 9.9999999999999998e-13
CS_252 NS_252 0 9.9999999999999998e-13
RS_251 NS_251 0 9.0838548010669172e+01
RS_252 NS_252 0 9.0838548010669186e+01
GL_251 0 NS_251 NS_252 0 2.2647420085995260e-01
GL_252 0 NS_252 NS_251 0 -2.2647420085995260e-01
GS_251_6 0 NS_251 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 253/254
CS_253 NS_253 0 9.9999999999999998e-13
CS_254 NS_254 0 9.9999999999999998e-13
RS_253 NS_253 0 5.0298322136619066e+02
RS_254 NS_254 0 5.0298322136619078e+02
GL_253 0 NS_253 NS_254 0 2.4757175091537195e-01
GL_254 0 NS_254 NS_253 0 -2.4757175091537195e-01
GS_253_6 0 NS_253 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 255/256
CS_255 NS_255 0 9.9999999999999998e-13
CS_256 NS_256 0 9.9999999999999998e-13
RS_255 NS_255 0 1.1113846377285431e+02
RS_256 NS_256 0 1.1113846377285431e+02
GL_255 0 NS_255 NS_256 0 2.4529156966751164e-01
GL_256 0 NS_256 NS_255 0 -2.4529156966751164e-01
GS_255_6 0 NS_255 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 257/258
CS_257 NS_257 0 9.9999999999999998e-13
CS_258 NS_258 0 9.9999999999999998e-13
RS_257 NS_257 0 4.1132635267896995e+02
RS_258 NS_258 0 4.1132635267896990e+02
GL_257 0 NS_257 NS_258 0 2.4323159344727399e-01
GL_258 0 NS_258 NS_257 0 -2.4323159344727399e-01
GS_257_6 0 NS_257 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 259/260
CS_259 NS_259 0 9.9999999999999998e-13
CS_260 NS_260 0 9.9999999999999998e-13
RS_259 NS_259 0 6.1483243702508491e+02
RS_260 NS_260 0 6.1483243702508491e+02
GL_259 0 NS_259 NS_260 0 2.3313794138995145e-01
GL_260 0 NS_260 NS_259 0 -2.3313794138995145e-01
GS_259_6 0 NS_259 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 261/262
CS_261 NS_261 0 9.9999999999999998e-13
CS_262 NS_262 0 9.9999999999999998e-13
RS_261 NS_261 0 6.0708452252497170e+02
RS_262 NS_262 0 6.0708452252497170e+02
GL_261 0 NS_261 NS_262 0 2.3828547054015958e-01
GL_262 0 NS_262 NS_261 0 -2.3828547054015958e-01
GS_261_6 0 NS_261 NA_6 0 1.6921379288850509e+00
*
* Complex pair n. 263/264
CS_263 NS_263 0 9.9999999999999998e-13
CS_264 NS_264 0 9.9999999999999998e-13
RS_263 NS_263 0 1.9238303220034285e+02
RS_264 NS_264 0 1.9238303220034285e+02
GL_263 0 NS_263 NS_264 0 2.3639447764395666e-01
GL_264 0 NS_264 NS_263 0 -2.3639447764395666e-01
GS_263_6 0 NS_263 NA_6 0 1.6921379288850509e+00
*
* Real pole n. 265
CS_265 NS_265 0 9.9999999999999998e-13
RS_265 NS_265 0 1.2063458770185771e+00
GS_265_7 0 NS_265 NA_7 0 1.6921379288850509e+00
*
* Real pole n. 266
CS_266 NS_266 0 9.9999999999999998e-13
RS_266 NS_266 0 2.0414994648771170e+01
GS_266_7 0 NS_266 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 267/268
CS_267 NS_267 0 9.9999999999999998e-13
CS_268 NS_268 0 9.9999999999999998e-13
RS_267 NS_267 0 2.2164632983638530e+01
RS_268 NS_268 0 2.2164632983638530e+01
GL_267 0 NS_267 NS_268 0 6.2432580119989492e-02
GL_268 0 NS_268 NS_267 0 -6.2432580119989492e-02
GS_267_7 0 NS_267 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 269/270
CS_269 NS_269 0 9.9999999999999998e-13
CS_270 NS_270 0 9.9999999999999998e-13
RS_269 NS_269 0 2.4208144339458560e+01
RS_270 NS_270 0 2.4208144339458560e+01
GL_269 0 NS_269 NS_270 0 8.7759448763363015e-02
GL_270 0 NS_270 NS_269 0 -8.7759448763363015e-02
GS_269_7 0 NS_269 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 271/272
CS_271 NS_271 0 9.9999999999999998e-13
CS_272 NS_272 0 9.9999999999999998e-13
RS_271 NS_271 0 1.3097029666184031e+02
RS_272 NS_272 0 1.3097029666184031e+02
GL_271 0 NS_271 NS_272 0 2.9672291989323329e-01
GL_272 0 NS_272 NS_271 0 -2.9672291989323329e-01
GS_271_7 0 NS_271 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 273/274
CS_273 NS_273 0 9.9999999999999998e-13
CS_274 NS_274 0 9.9999999999999998e-13
RS_273 NS_273 0 3.2672536376024027e+01
RS_274 NS_274 0 3.2672536376024027e+01
GL_273 0 NS_273 NS_274 0 1.2489866711430768e-01
GL_274 0 NS_274 NS_273 0 -1.2489866711430768e-01
GS_273_7 0 NS_273 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 275/276
CS_275 NS_275 0 9.9999999999999998e-13
CS_276 NS_276 0 9.9999999999999998e-13
RS_275 NS_275 0 3.6741731246022816e+01
RS_276 NS_276 0 3.6741731246022816e+01
GL_275 0 NS_275 NS_276 0 1.6399845549232167e-01
GL_276 0 NS_276 NS_275 0 -1.6399845549232167e-01
GS_275_7 0 NS_275 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 277/278
CS_277 NS_277 0 9.9999999999999998e-13
CS_278 NS_278 0 9.9999999999999998e-13
RS_277 NS_277 0 8.3646036557163740e+01
RS_278 NS_278 0 8.3646036557163740e+01
GL_277 0 NS_277 NS_278 0 1.6830719130342967e-01
GL_278 0 NS_278 NS_277 0 -1.6830719130342967e-01
GS_277_7 0 NS_277 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 279/280
CS_279 NS_279 0 9.9999999999999998e-13
CS_280 NS_280 0 9.9999999999999998e-13
RS_279 NS_279 0 4.0307732865054554e+01
RS_280 NS_280 0 4.0307732865054554e+01
GL_279 0 NS_279 NS_280 0 1.8890575271706389e-01
GL_280 0 NS_280 NS_279 0 -1.8890575271706389e-01
GS_279_7 0 NS_279 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 281/282
CS_281 NS_281 0 9.9999999999999998e-13
CS_282 NS_282 0 9.9999999999999998e-13
RS_281 NS_281 0 1.4268073111996583e+02
RS_282 NS_282 0 1.4268073111996583e+02
GL_281 0 NS_281 NS_282 0 1.9419078929943706e-01
GL_282 0 NS_282 NS_281 0 -1.9419078929943706e-01
GS_281_7 0 NS_281 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 283/284
CS_283 NS_283 0 9.9999999999999998e-13
CS_284 NS_284 0 9.9999999999999998e-13
RS_283 NS_283 0 7.1679198821979867e+01
RS_284 NS_284 0 7.1679198821979867e+01
GL_283 0 NS_283 NS_284 0 2.0702628270375376e-01
GL_284 0 NS_284 NS_283 0 -2.0702628270375376e-01
GS_283_7 0 NS_283 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 285/286
CS_285 NS_285 0 9.9999999999999998e-13
CS_286 NS_286 0 9.9999999999999998e-13
RS_285 NS_285 0 1.6005864146684806e+02
RS_286 NS_286 0 1.6005864146684809e+02
GL_285 0 NS_285 NS_286 0 2.5423900390253934e-01
GL_286 0 NS_286 NS_285 0 -2.5423900390253934e-01
GS_285_7 0 NS_285 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 287/288
CS_287 NS_287 0 9.9999999999999998e-13
CS_288 NS_288 0 9.9999999999999998e-13
RS_287 NS_287 0 1.9181463552142085e+02
RS_288 NS_288 0 1.9181463552142085e+02
GL_287 0 NS_287 NS_288 0 2.1188941693262670e-01
GL_288 0 NS_288 NS_287 0 -2.1188941693262670e-01
GS_287_7 0 NS_287 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 289/290
CS_289 NS_289 0 9.9999999999999998e-13
CS_290 NS_290 0 9.9999999999999998e-13
RS_289 NS_289 0 2.5689115313648813e+02
RS_290 NS_290 0 2.5689115313648813e+02
GL_289 0 NS_289 NS_290 0 2.1774212061821885e-01
GL_290 0 NS_290 NS_289 0 -2.1774212061821885e-01
GS_289_7 0 NS_289 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 291/292
CS_291 NS_291 0 9.9999999999999998e-13
CS_292 NS_292 0 9.9999999999999998e-13
RS_291 NS_291 0 6.2765149843829192e+01
RS_292 NS_292 0 6.2765149843829192e+01
GL_291 0 NS_291 NS_292 0 2.3246082537351351e-01
GL_292 0 NS_292 NS_291 0 -2.3246082537351351e-01
GS_291_7 0 NS_291 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 293/294
CS_293 NS_293 0 9.9999999999999998e-13
CS_294 NS_294 0 9.9999999999999998e-13
RS_293 NS_293 0 3.5419967361311882e+02
RS_294 NS_294 0 3.5419967361311882e+02
GL_293 0 NS_293 NS_294 0 2.2268031336810420e-01
GL_294 0 NS_294 NS_293 0 -2.2268031336810420e-01
GS_293_7 0 NS_293 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 295/296
CS_295 NS_295 0 9.9999999999999998e-13
CS_296 NS_296 0 9.9999999999999998e-13
RS_295 NS_295 0 9.0838548010669172e+01
RS_296 NS_296 0 9.0838548010669186e+01
GL_295 0 NS_295 NS_296 0 2.2647420085995260e-01
GL_296 0 NS_296 NS_295 0 -2.2647420085995260e-01
GS_295_7 0 NS_295 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 297/298
CS_297 NS_297 0 9.9999999999999998e-13
CS_298 NS_298 0 9.9999999999999998e-13
RS_297 NS_297 0 5.0298322136619066e+02
RS_298 NS_298 0 5.0298322136619078e+02
GL_297 0 NS_297 NS_298 0 2.4757175091537195e-01
GL_298 0 NS_298 NS_297 0 -2.4757175091537195e-01
GS_297_7 0 NS_297 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 299/300
CS_299 NS_299 0 9.9999999999999998e-13
CS_300 NS_300 0 9.9999999999999998e-13
RS_299 NS_299 0 1.1113846377285431e+02
RS_300 NS_300 0 1.1113846377285431e+02
GL_299 0 NS_299 NS_300 0 2.4529156966751164e-01
GL_300 0 NS_300 NS_299 0 -2.4529156966751164e-01
GS_299_7 0 NS_299 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 301/302
CS_301 NS_301 0 9.9999999999999998e-13
CS_302 NS_302 0 9.9999999999999998e-13
RS_301 NS_301 0 4.1132635267896995e+02
RS_302 NS_302 0 4.1132635267896990e+02
GL_301 0 NS_301 NS_302 0 2.4323159344727399e-01
GL_302 0 NS_302 NS_301 0 -2.4323159344727399e-01
GS_301_7 0 NS_301 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 303/304
CS_303 NS_303 0 9.9999999999999998e-13
CS_304 NS_304 0 9.9999999999999998e-13
RS_303 NS_303 0 6.1483243702508491e+02
RS_304 NS_304 0 6.1483243702508491e+02
GL_303 0 NS_303 NS_304 0 2.3313794138995145e-01
GL_304 0 NS_304 NS_303 0 -2.3313794138995145e-01
GS_303_7 0 NS_303 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 305/306
CS_305 NS_305 0 9.9999999999999998e-13
CS_306 NS_306 0 9.9999999999999998e-13
RS_305 NS_305 0 6.0708452252497170e+02
RS_306 NS_306 0 6.0708452252497170e+02
GL_305 0 NS_305 NS_306 0 2.3828547054015958e-01
GL_306 0 NS_306 NS_305 0 -2.3828547054015958e-01
GS_305_7 0 NS_305 NA_7 0 1.6921379288850509e+00
*
* Complex pair n. 307/308
CS_307 NS_307 0 9.9999999999999998e-13
CS_308 NS_308 0 9.9999999999999998e-13
RS_307 NS_307 0 1.9238303220034285e+02
RS_308 NS_308 0 1.9238303220034285e+02
GL_307 0 NS_307 NS_308 0 2.3639447764395666e-01
GL_308 0 NS_308 NS_307 0 -2.3639447764395666e-01
GS_307_7 0 NS_307 NA_7 0 1.6921379288850509e+00
*
* Real pole n. 309
CS_309 NS_309 0 9.9999999999999998e-13
RS_309 NS_309 0 1.2063458770185771e+00
GS_309_8 0 NS_309 NA_8 0 1.6921379288850509e+00
*
* Real pole n. 310
CS_310 NS_310 0 9.9999999999999998e-13
RS_310 NS_310 0 2.0414994648771170e+01
GS_310_8 0 NS_310 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 311/312
CS_311 NS_311 0 9.9999999999999998e-13
CS_312 NS_312 0 9.9999999999999998e-13
RS_311 NS_311 0 2.2164632983638530e+01
RS_312 NS_312 0 2.2164632983638530e+01
GL_311 0 NS_311 NS_312 0 6.2432580119989492e-02
GL_312 0 NS_312 NS_311 0 -6.2432580119989492e-02
GS_311_8 0 NS_311 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 313/314
CS_313 NS_313 0 9.9999999999999998e-13
CS_314 NS_314 0 9.9999999999999998e-13
RS_313 NS_313 0 2.4208144339458560e+01
RS_314 NS_314 0 2.4208144339458560e+01
GL_313 0 NS_313 NS_314 0 8.7759448763363015e-02
GL_314 0 NS_314 NS_313 0 -8.7759448763363015e-02
GS_313_8 0 NS_313 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 315/316
CS_315 NS_315 0 9.9999999999999998e-13
CS_316 NS_316 0 9.9999999999999998e-13
RS_315 NS_315 0 1.3097029666184031e+02
RS_316 NS_316 0 1.3097029666184031e+02
GL_315 0 NS_315 NS_316 0 2.9672291989323329e-01
GL_316 0 NS_316 NS_315 0 -2.9672291989323329e-01
GS_315_8 0 NS_315 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 317/318
CS_317 NS_317 0 9.9999999999999998e-13
CS_318 NS_318 0 9.9999999999999998e-13
RS_317 NS_317 0 3.2672536376024027e+01
RS_318 NS_318 0 3.2672536376024027e+01
GL_317 0 NS_317 NS_318 0 1.2489866711430768e-01
GL_318 0 NS_318 NS_317 0 -1.2489866711430768e-01
GS_317_8 0 NS_317 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 319/320
CS_319 NS_319 0 9.9999999999999998e-13
CS_320 NS_320 0 9.9999999999999998e-13
RS_319 NS_319 0 3.6741731246022816e+01
RS_320 NS_320 0 3.6741731246022816e+01
GL_319 0 NS_319 NS_320 0 1.6399845549232167e-01
GL_320 0 NS_320 NS_319 0 -1.6399845549232167e-01
GS_319_8 0 NS_319 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 321/322
CS_321 NS_321 0 9.9999999999999998e-13
CS_322 NS_322 0 9.9999999999999998e-13
RS_321 NS_321 0 8.3646036557163740e+01
RS_322 NS_322 0 8.3646036557163740e+01
GL_321 0 NS_321 NS_322 0 1.6830719130342967e-01
GL_322 0 NS_322 NS_321 0 -1.6830719130342967e-01
GS_321_8 0 NS_321 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 323/324
CS_323 NS_323 0 9.9999999999999998e-13
CS_324 NS_324 0 9.9999999999999998e-13
RS_323 NS_323 0 4.0307732865054554e+01
RS_324 NS_324 0 4.0307732865054554e+01
GL_323 0 NS_323 NS_324 0 1.8890575271706389e-01
GL_324 0 NS_324 NS_323 0 -1.8890575271706389e-01
GS_323_8 0 NS_323 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 325/326
CS_325 NS_325 0 9.9999999999999998e-13
CS_326 NS_326 0 9.9999999999999998e-13
RS_325 NS_325 0 1.4268073111996583e+02
RS_326 NS_326 0 1.4268073111996583e+02
GL_325 0 NS_325 NS_326 0 1.9419078929943706e-01
GL_326 0 NS_326 NS_325 0 -1.9419078929943706e-01
GS_325_8 0 NS_325 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 327/328
CS_327 NS_327 0 9.9999999999999998e-13
CS_328 NS_328 0 9.9999999999999998e-13
RS_327 NS_327 0 7.1679198821979867e+01
RS_328 NS_328 0 7.1679198821979867e+01
GL_327 0 NS_327 NS_328 0 2.0702628270375376e-01
GL_328 0 NS_328 NS_327 0 -2.0702628270375376e-01
GS_327_8 0 NS_327 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 329/330
CS_329 NS_329 0 9.9999999999999998e-13
CS_330 NS_330 0 9.9999999999999998e-13
RS_329 NS_329 0 1.6005864146684806e+02
RS_330 NS_330 0 1.6005864146684809e+02
GL_329 0 NS_329 NS_330 0 2.5423900390253934e-01
GL_330 0 NS_330 NS_329 0 -2.5423900390253934e-01
GS_329_8 0 NS_329 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 331/332
CS_331 NS_331 0 9.9999999999999998e-13
CS_332 NS_332 0 9.9999999999999998e-13
RS_331 NS_331 0 1.9181463552142085e+02
RS_332 NS_332 0 1.9181463552142085e+02
GL_331 0 NS_331 NS_332 0 2.1188941693262670e-01
GL_332 0 NS_332 NS_331 0 -2.1188941693262670e-01
GS_331_8 0 NS_331 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 333/334
CS_333 NS_333 0 9.9999999999999998e-13
CS_334 NS_334 0 9.9999999999999998e-13
RS_333 NS_333 0 2.5689115313648813e+02
RS_334 NS_334 0 2.5689115313648813e+02
GL_333 0 NS_333 NS_334 0 2.1774212061821885e-01
GL_334 0 NS_334 NS_333 0 -2.1774212061821885e-01
GS_333_8 0 NS_333 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 335/336
CS_335 NS_335 0 9.9999999999999998e-13
CS_336 NS_336 0 9.9999999999999998e-13
RS_335 NS_335 0 6.2765149843829192e+01
RS_336 NS_336 0 6.2765149843829192e+01
GL_335 0 NS_335 NS_336 0 2.3246082537351351e-01
GL_336 0 NS_336 NS_335 0 -2.3246082537351351e-01
GS_335_8 0 NS_335 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 337/338
CS_337 NS_337 0 9.9999999999999998e-13
CS_338 NS_338 0 9.9999999999999998e-13
RS_337 NS_337 0 3.5419967361311882e+02
RS_338 NS_338 0 3.5419967361311882e+02
GL_337 0 NS_337 NS_338 0 2.2268031336810420e-01
GL_338 0 NS_338 NS_337 0 -2.2268031336810420e-01
GS_337_8 0 NS_337 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 339/340
CS_339 NS_339 0 9.9999999999999998e-13
CS_340 NS_340 0 9.9999999999999998e-13
RS_339 NS_339 0 9.0838548010669172e+01
RS_340 NS_340 0 9.0838548010669186e+01
GL_339 0 NS_339 NS_340 0 2.2647420085995260e-01
GL_340 0 NS_340 NS_339 0 -2.2647420085995260e-01
GS_339_8 0 NS_339 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 341/342
CS_341 NS_341 0 9.9999999999999998e-13
CS_342 NS_342 0 9.9999999999999998e-13
RS_341 NS_341 0 5.0298322136619066e+02
RS_342 NS_342 0 5.0298322136619078e+02
GL_341 0 NS_341 NS_342 0 2.4757175091537195e-01
GL_342 0 NS_342 NS_341 0 -2.4757175091537195e-01
GS_341_8 0 NS_341 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 343/344
CS_343 NS_343 0 9.9999999999999998e-13
CS_344 NS_344 0 9.9999999999999998e-13
RS_343 NS_343 0 1.1113846377285431e+02
RS_344 NS_344 0 1.1113846377285431e+02
GL_343 0 NS_343 NS_344 0 2.4529156966751164e-01
GL_344 0 NS_344 NS_343 0 -2.4529156966751164e-01
GS_343_8 0 NS_343 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 345/346
CS_345 NS_345 0 9.9999999999999998e-13
CS_346 NS_346 0 9.9999999999999998e-13
RS_345 NS_345 0 4.1132635267896995e+02
RS_346 NS_346 0 4.1132635267896990e+02
GL_345 0 NS_345 NS_346 0 2.4323159344727399e-01
GL_346 0 NS_346 NS_345 0 -2.4323159344727399e-01
GS_345_8 0 NS_345 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 347/348
CS_347 NS_347 0 9.9999999999999998e-13
CS_348 NS_348 0 9.9999999999999998e-13
RS_347 NS_347 0 6.1483243702508491e+02
RS_348 NS_348 0 6.1483243702508491e+02
GL_347 0 NS_347 NS_348 0 2.3313794138995145e-01
GL_348 0 NS_348 NS_347 0 -2.3313794138995145e-01
GS_347_8 0 NS_347 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 349/350
CS_349 NS_349 0 9.9999999999999998e-13
CS_350 NS_350 0 9.9999999999999998e-13
RS_349 NS_349 0 6.0708452252497170e+02
RS_350 NS_350 0 6.0708452252497170e+02
GL_349 0 NS_349 NS_350 0 2.3828547054015958e-01
GL_350 0 NS_350 NS_349 0 -2.3828547054015958e-01
GS_349_8 0 NS_349 NA_8 0 1.6921379288850509e+00
*
* Complex pair n. 351/352
CS_351 NS_351 0 9.9999999999999998e-13
CS_352 NS_352 0 9.9999999999999998e-13
RS_351 NS_351 0 1.9238303220034285e+02
RS_352 NS_352 0 1.9238303220034285e+02
GL_351 0 NS_351 NS_352 0 2.3639447764395666e-01
GL_352 0 NS_352 NS_351 0 -2.3639447764395666e-01
GS_351_8 0 NS_351 NA_8 0 1.6921379288850509e+00
*
* Real pole n. 353
CS_353 NS_353 0 9.9999999999999998e-13
RS_353 NS_353 0 1.2063458770185771e+00
GS_353_9 0 NS_353 NA_9 0 1.6921379288850509e+00
*
* Real pole n. 354
CS_354 NS_354 0 9.9999999999999998e-13
RS_354 NS_354 0 2.0414994648771170e+01
GS_354_9 0 NS_354 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 355/356
CS_355 NS_355 0 9.9999999999999998e-13
CS_356 NS_356 0 9.9999999999999998e-13
RS_355 NS_355 0 2.2164632983638530e+01
RS_356 NS_356 0 2.2164632983638530e+01
GL_355 0 NS_355 NS_356 0 6.2432580119989492e-02
GL_356 0 NS_356 NS_355 0 -6.2432580119989492e-02
GS_355_9 0 NS_355 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 357/358
CS_357 NS_357 0 9.9999999999999998e-13
CS_358 NS_358 0 9.9999999999999998e-13
RS_357 NS_357 0 2.4208144339458560e+01
RS_358 NS_358 0 2.4208144339458560e+01
GL_357 0 NS_357 NS_358 0 8.7759448763363015e-02
GL_358 0 NS_358 NS_357 0 -8.7759448763363015e-02
GS_357_9 0 NS_357 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 359/360
CS_359 NS_359 0 9.9999999999999998e-13
CS_360 NS_360 0 9.9999999999999998e-13
RS_359 NS_359 0 1.3097029666184031e+02
RS_360 NS_360 0 1.3097029666184031e+02
GL_359 0 NS_359 NS_360 0 2.9672291989323329e-01
GL_360 0 NS_360 NS_359 0 -2.9672291989323329e-01
GS_359_9 0 NS_359 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 361/362
CS_361 NS_361 0 9.9999999999999998e-13
CS_362 NS_362 0 9.9999999999999998e-13
RS_361 NS_361 0 3.2672536376024027e+01
RS_362 NS_362 0 3.2672536376024027e+01
GL_361 0 NS_361 NS_362 0 1.2489866711430768e-01
GL_362 0 NS_362 NS_361 0 -1.2489866711430768e-01
GS_361_9 0 NS_361 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 363/364
CS_363 NS_363 0 9.9999999999999998e-13
CS_364 NS_364 0 9.9999999999999998e-13
RS_363 NS_363 0 3.6741731246022816e+01
RS_364 NS_364 0 3.6741731246022816e+01
GL_363 0 NS_363 NS_364 0 1.6399845549232167e-01
GL_364 0 NS_364 NS_363 0 -1.6399845549232167e-01
GS_363_9 0 NS_363 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 365/366
CS_365 NS_365 0 9.9999999999999998e-13
CS_366 NS_366 0 9.9999999999999998e-13
RS_365 NS_365 0 8.3646036557163740e+01
RS_366 NS_366 0 8.3646036557163740e+01
GL_365 0 NS_365 NS_366 0 1.6830719130342967e-01
GL_366 0 NS_366 NS_365 0 -1.6830719130342967e-01
GS_365_9 0 NS_365 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 367/368
CS_367 NS_367 0 9.9999999999999998e-13
CS_368 NS_368 0 9.9999999999999998e-13
RS_367 NS_367 0 4.0307732865054554e+01
RS_368 NS_368 0 4.0307732865054554e+01
GL_367 0 NS_367 NS_368 0 1.8890575271706389e-01
GL_368 0 NS_368 NS_367 0 -1.8890575271706389e-01
GS_367_9 0 NS_367 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 369/370
CS_369 NS_369 0 9.9999999999999998e-13
CS_370 NS_370 0 9.9999999999999998e-13
RS_369 NS_369 0 1.4268073111996583e+02
RS_370 NS_370 0 1.4268073111996583e+02
GL_369 0 NS_369 NS_370 0 1.9419078929943706e-01
GL_370 0 NS_370 NS_369 0 -1.9419078929943706e-01
GS_369_9 0 NS_369 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 371/372
CS_371 NS_371 0 9.9999999999999998e-13
CS_372 NS_372 0 9.9999999999999998e-13
RS_371 NS_371 0 7.1679198821979867e+01
RS_372 NS_372 0 7.1679198821979867e+01
GL_371 0 NS_371 NS_372 0 2.0702628270375376e-01
GL_372 0 NS_372 NS_371 0 -2.0702628270375376e-01
GS_371_9 0 NS_371 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 373/374
CS_373 NS_373 0 9.9999999999999998e-13
CS_374 NS_374 0 9.9999999999999998e-13
RS_373 NS_373 0 1.6005864146684806e+02
RS_374 NS_374 0 1.6005864146684809e+02
GL_373 0 NS_373 NS_374 0 2.5423900390253934e-01
GL_374 0 NS_374 NS_373 0 -2.5423900390253934e-01
GS_373_9 0 NS_373 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 375/376
CS_375 NS_375 0 9.9999999999999998e-13
CS_376 NS_376 0 9.9999999999999998e-13
RS_375 NS_375 0 1.9181463552142085e+02
RS_376 NS_376 0 1.9181463552142085e+02
GL_375 0 NS_375 NS_376 0 2.1188941693262670e-01
GL_376 0 NS_376 NS_375 0 -2.1188941693262670e-01
GS_375_9 0 NS_375 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 377/378
CS_377 NS_377 0 9.9999999999999998e-13
CS_378 NS_378 0 9.9999999999999998e-13
RS_377 NS_377 0 2.5689115313648813e+02
RS_378 NS_378 0 2.5689115313648813e+02
GL_377 0 NS_377 NS_378 0 2.1774212061821885e-01
GL_378 0 NS_378 NS_377 0 -2.1774212061821885e-01
GS_377_9 0 NS_377 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 379/380
CS_379 NS_379 0 9.9999999999999998e-13
CS_380 NS_380 0 9.9999999999999998e-13
RS_379 NS_379 0 6.2765149843829192e+01
RS_380 NS_380 0 6.2765149843829192e+01
GL_379 0 NS_379 NS_380 0 2.3246082537351351e-01
GL_380 0 NS_380 NS_379 0 -2.3246082537351351e-01
GS_379_9 0 NS_379 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 381/382
CS_381 NS_381 0 9.9999999999999998e-13
CS_382 NS_382 0 9.9999999999999998e-13
RS_381 NS_381 0 3.5419967361311882e+02
RS_382 NS_382 0 3.5419967361311882e+02
GL_381 0 NS_381 NS_382 0 2.2268031336810420e-01
GL_382 0 NS_382 NS_381 0 -2.2268031336810420e-01
GS_381_9 0 NS_381 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 383/384
CS_383 NS_383 0 9.9999999999999998e-13
CS_384 NS_384 0 9.9999999999999998e-13
RS_383 NS_383 0 9.0838548010669172e+01
RS_384 NS_384 0 9.0838548010669186e+01
GL_383 0 NS_383 NS_384 0 2.2647420085995260e-01
GL_384 0 NS_384 NS_383 0 -2.2647420085995260e-01
GS_383_9 0 NS_383 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 385/386
CS_385 NS_385 0 9.9999999999999998e-13
CS_386 NS_386 0 9.9999999999999998e-13
RS_385 NS_385 0 5.0298322136619066e+02
RS_386 NS_386 0 5.0298322136619078e+02
GL_385 0 NS_385 NS_386 0 2.4757175091537195e-01
GL_386 0 NS_386 NS_385 0 -2.4757175091537195e-01
GS_385_9 0 NS_385 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 387/388
CS_387 NS_387 0 9.9999999999999998e-13
CS_388 NS_388 0 9.9999999999999998e-13
RS_387 NS_387 0 1.1113846377285431e+02
RS_388 NS_388 0 1.1113846377285431e+02
GL_387 0 NS_387 NS_388 0 2.4529156966751164e-01
GL_388 0 NS_388 NS_387 0 -2.4529156966751164e-01
GS_387_9 0 NS_387 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 389/390
CS_389 NS_389 0 9.9999999999999998e-13
CS_390 NS_390 0 9.9999999999999998e-13
RS_389 NS_389 0 4.1132635267896995e+02
RS_390 NS_390 0 4.1132635267896990e+02
GL_389 0 NS_389 NS_390 0 2.4323159344727399e-01
GL_390 0 NS_390 NS_389 0 -2.4323159344727399e-01
GS_389_9 0 NS_389 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 391/392
CS_391 NS_391 0 9.9999999999999998e-13
CS_392 NS_392 0 9.9999999999999998e-13
RS_391 NS_391 0 6.1483243702508491e+02
RS_392 NS_392 0 6.1483243702508491e+02
GL_391 0 NS_391 NS_392 0 2.3313794138995145e-01
GL_392 0 NS_392 NS_391 0 -2.3313794138995145e-01
GS_391_9 0 NS_391 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 393/394
CS_393 NS_393 0 9.9999999999999998e-13
CS_394 NS_394 0 9.9999999999999998e-13
RS_393 NS_393 0 6.0708452252497170e+02
RS_394 NS_394 0 6.0708452252497170e+02
GL_393 0 NS_393 NS_394 0 2.3828547054015958e-01
GL_394 0 NS_394 NS_393 0 -2.3828547054015958e-01
GS_393_9 0 NS_393 NA_9 0 1.6921379288850509e+00
*
* Complex pair n. 395/396
CS_395 NS_395 0 9.9999999999999998e-13
CS_396 NS_396 0 9.9999999999999998e-13
RS_395 NS_395 0 1.9238303220034285e+02
RS_396 NS_396 0 1.9238303220034285e+02
GL_395 0 NS_395 NS_396 0 2.3639447764395666e-01
GL_396 0 NS_396 NS_395 0 -2.3639447764395666e-01
GS_395_9 0 NS_395 NA_9 0 1.6921379288850509e+00
*
* Real pole n. 397
CS_397 NS_397 0 9.9999999999999998e-13
RS_397 NS_397 0 1.2063458770185771e+00
GS_397_10 0 NS_397 NA_10 0 1.6921379288850509e+00
*
* Real pole n. 398
CS_398 NS_398 0 9.9999999999999998e-13
RS_398 NS_398 0 2.0414994648771170e+01
GS_398_10 0 NS_398 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 399/400
CS_399 NS_399 0 9.9999999999999998e-13
CS_400 NS_400 0 9.9999999999999998e-13
RS_399 NS_399 0 2.2164632983638530e+01
RS_400 NS_400 0 2.2164632983638530e+01
GL_399 0 NS_399 NS_400 0 6.2432580119989492e-02
GL_400 0 NS_400 NS_399 0 -6.2432580119989492e-02
GS_399_10 0 NS_399 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 401/402
CS_401 NS_401 0 9.9999999999999998e-13
CS_402 NS_402 0 9.9999999999999998e-13
RS_401 NS_401 0 2.4208144339458560e+01
RS_402 NS_402 0 2.4208144339458560e+01
GL_401 0 NS_401 NS_402 0 8.7759448763363015e-02
GL_402 0 NS_402 NS_401 0 -8.7759448763363015e-02
GS_401_10 0 NS_401 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 403/404
CS_403 NS_403 0 9.9999999999999998e-13
CS_404 NS_404 0 9.9999999999999998e-13
RS_403 NS_403 0 1.3097029666184031e+02
RS_404 NS_404 0 1.3097029666184031e+02
GL_403 0 NS_403 NS_404 0 2.9672291989323329e-01
GL_404 0 NS_404 NS_403 0 -2.9672291989323329e-01
GS_403_10 0 NS_403 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 405/406
CS_405 NS_405 0 9.9999999999999998e-13
CS_406 NS_406 0 9.9999999999999998e-13
RS_405 NS_405 0 3.2672536376024027e+01
RS_406 NS_406 0 3.2672536376024027e+01
GL_405 0 NS_405 NS_406 0 1.2489866711430768e-01
GL_406 0 NS_406 NS_405 0 -1.2489866711430768e-01
GS_405_10 0 NS_405 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 407/408
CS_407 NS_407 0 9.9999999999999998e-13
CS_408 NS_408 0 9.9999999999999998e-13
RS_407 NS_407 0 3.6741731246022816e+01
RS_408 NS_408 0 3.6741731246022816e+01
GL_407 0 NS_407 NS_408 0 1.6399845549232167e-01
GL_408 0 NS_408 NS_407 0 -1.6399845549232167e-01
GS_407_10 0 NS_407 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 409/410
CS_409 NS_409 0 9.9999999999999998e-13
CS_410 NS_410 0 9.9999999999999998e-13
RS_409 NS_409 0 8.3646036557163740e+01
RS_410 NS_410 0 8.3646036557163740e+01
GL_409 0 NS_409 NS_410 0 1.6830719130342967e-01
GL_410 0 NS_410 NS_409 0 -1.6830719130342967e-01
GS_409_10 0 NS_409 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 411/412
CS_411 NS_411 0 9.9999999999999998e-13
CS_412 NS_412 0 9.9999999999999998e-13
RS_411 NS_411 0 4.0307732865054554e+01
RS_412 NS_412 0 4.0307732865054554e+01
GL_411 0 NS_411 NS_412 0 1.8890575271706389e-01
GL_412 0 NS_412 NS_411 0 -1.8890575271706389e-01
GS_411_10 0 NS_411 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 413/414
CS_413 NS_413 0 9.9999999999999998e-13
CS_414 NS_414 0 9.9999999999999998e-13
RS_413 NS_413 0 1.4268073111996583e+02
RS_414 NS_414 0 1.4268073111996583e+02
GL_413 0 NS_413 NS_414 0 1.9419078929943706e-01
GL_414 0 NS_414 NS_413 0 -1.9419078929943706e-01
GS_413_10 0 NS_413 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 415/416
CS_415 NS_415 0 9.9999999999999998e-13
CS_416 NS_416 0 9.9999999999999998e-13
RS_415 NS_415 0 7.1679198821979867e+01
RS_416 NS_416 0 7.1679198821979867e+01
GL_415 0 NS_415 NS_416 0 2.0702628270375376e-01
GL_416 0 NS_416 NS_415 0 -2.0702628270375376e-01
GS_415_10 0 NS_415 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 417/418
CS_417 NS_417 0 9.9999999999999998e-13
CS_418 NS_418 0 9.9999999999999998e-13
RS_417 NS_417 0 1.6005864146684806e+02
RS_418 NS_418 0 1.6005864146684809e+02
GL_417 0 NS_417 NS_418 0 2.5423900390253934e-01
GL_418 0 NS_418 NS_417 0 -2.5423900390253934e-01
GS_417_10 0 NS_417 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 419/420
CS_419 NS_419 0 9.9999999999999998e-13
CS_420 NS_420 0 9.9999999999999998e-13
RS_419 NS_419 0 1.9181463552142085e+02
RS_420 NS_420 0 1.9181463552142085e+02
GL_419 0 NS_419 NS_420 0 2.1188941693262670e-01
GL_420 0 NS_420 NS_419 0 -2.1188941693262670e-01
GS_419_10 0 NS_419 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 421/422
CS_421 NS_421 0 9.9999999999999998e-13
CS_422 NS_422 0 9.9999999999999998e-13
RS_421 NS_421 0 2.5689115313648813e+02
RS_422 NS_422 0 2.5689115313648813e+02
GL_421 0 NS_421 NS_422 0 2.1774212061821885e-01
GL_422 0 NS_422 NS_421 0 -2.1774212061821885e-01
GS_421_10 0 NS_421 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 423/424
CS_423 NS_423 0 9.9999999999999998e-13
CS_424 NS_424 0 9.9999999999999998e-13
RS_423 NS_423 0 6.2765149843829192e+01
RS_424 NS_424 0 6.2765149843829192e+01
GL_423 0 NS_423 NS_424 0 2.3246082537351351e-01
GL_424 0 NS_424 NS_423 0 -2.3246082537351351e-01
GS_423_10 0 NS_423 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 425/426
CS_425 NS_425 0 9.9999999999999998e-13
CS_426 NS_426 0 9.9999999999999998e-13
RS_425 NS_425 0 3.5419967361311882e+02
RS_426 NS_426 0 3.5419967361311882e+02
GL_425 0 NS_425 NS_426 0 2.2268031336810420e-01
GL_426 0 NS_426 NS_425 0 -2.2268031336810420e-01
GS_425_10 0 NS_425 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 427/428
CS_427 NS_427 0 9.9999999999999998e-13
CS_428 NS_428 0 9.9999999999999998e-13
RS_427 NS_427 0 9.0838548010669172e+01
RS_428 NS_428 0 9.0838548010669186e+01
GL_427 0 NS_427 NS_428 0 2.2647420085995260e-01
GL_428 0 NS_428 NS_427 0 -2.2647420085995260e-01
GS_427_10 0 NS_427 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 429/430
CS_429 NS_429 0 9.9999999999999998e-13
CS_430 NS_430 0 9.9999999999999998e-13
RS_429 NS_429 0 5.0298322136619066e+02
RS_430 NS_430 0 5.0298322136619078e+02
GL_429 0 NS_429 NS_430 0 2.4757175091537195e-01
GL_430 0 NS_430 NS_429 0 -2.4757175091537195e-01
GS_429_10 0 NS_429 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 431/432
CS_431 NS_431 0 9.9999999999999998e-13
CS_432 NS_432 0 9.9999999999999998e-13
RS_431 NS_431 0 1.1113846377285431e+02
RS_432 NS_432 0 1.1113846377285431e+02
GL_431 0 NS_431 NS_432 0 2.4529156966751164e-01
GL_432 0 NS_432 NS_431 0 -2.4529156966751164e-01
GS_431_10 0 NS_431 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 433/434
CS_433 NS_433 0 9.9999999999999998e-13
CS_434 NS_434 0 9.9999999999999998e-13
RS_433 NS_433 0 4.1132635267896995e+02
RS_434 NS_434 0 4.1132635267896990e+02
GL_433 0 NS_433 NS_434 0 2.4323159344727399e-01
GL_434 0 NS_434 NS_433 0 -2.4323159344727399e-01
GS_433_10 0 NS_433 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 435/436
CS_435 NS_435 0 9.9999999999999998e-13
CS_436 NS_436 0 9.9999999999999998e-13
RS_435 NS_435 0 6.1483243702508491e+02
RS_436 NS_436 0 6.1483243702508491e+02
GL_435 0 NS_435 NS_436 0 2.3313794138995145e-01
GL_436 0 NS_436 NS_435 0 -2.3313794138995145e-01
GS_435_10 0 NS_435 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 437/438
CS_437 NS_437 0 9.9999999999999998e-13
CS_438 NS_438 0 9.9999999999999998e-13
RS_437 NS_437 0 6.0708452252497170e+02
RS_438 NS_438 0 6.0708452252497170e+02
GL_437 0 NS_437 NS_438 0 2.3828547054015958e-01
GL_438 0 NS_438 NS_437 0 -2.3828547054015958e-01
GS_437_10 0 NS_437 NA_10 0 1.6921379288850509e+00
*
* Complex pair n. 439/440
CS_439 NS_439 0 9.9999999999999998e-13
CS_440 NS_440 0 9.9999999999999998e-13
RS_439 NS_439 0 1.9238303220034285e+02
RS_440 NS_440 0 1.9238303220034285e+02
GL_439 0 NS_439 NS_440 0 2.3639447764395666e-01
GL_440 0 NS_440 NS_439 0 -2.3639447764395666e-01
GS_439_10 0 NS_439 NA_10 0 1.6921379288850509e+00
*
* Real pole n. 441
CS_441 NS_441 0 9.9999999999999998e-13
RS_441 NS_441 0 1.2063458770185771e+00
GS_441_11 0 NS_441 NA_11 0 1.6921379288850509e+00
*
* Real pole n. 442
CS_442 NS_442 0 9.9999999999999998e-13
RS_442 NS_442 0 2.0414994648771170e+01
GS_442_11 0 NS_442 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 443/444
CS_443 NS_443 0 9.9999999999999998e-13
CS_444 NS_444 0 9.9999999999999998e-13
RS_443 NS_443 0 2.2164632983638530e+01
RS_444 NS_444 0 2.2164632983638530e+01
GL_443 0 NS_443 NS_444 0 6.2432580119989492e-02
GL_444 0 NS_444 NS_443 0 -6.2432580119989492e-02
GS_443_11 0 NS_443 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 445/446
CS_445 NS_445 0 9.9999999999999998e-13
CS_446 NS_446 0 9.9999999999999998e-13
RS_445 NS_445 0 2.4208144339458560e+01
RS_446 NS_446 0 2.4208144339458560e+01
GL_445 0 NS_445 NS_446 0 8.7759448763363015e-02
GL_446 0 NS_446 NS_445 0 -8.7759448763363015e-02
GS_445_11 0 NS_445 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 447/448
CS_447 NS_447 0 9.9999999999999998e-13
CS_448 NS_448 0 9.9999999999999998e-13
RS_447 NS_447 0 1.3097029666184031e+02
RS_448 NS_448 0 1.3097029666184031e+02
GL_447 0 NS_447 NS_448 0 2.9672291989323329e-01
GL_448 0 NS_448 NS_447 0 -2.9672291989323329e-01
GS_447_11 0 NS_447 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 449/450
CS_449 NS_449 0 9.9999999999999998e-13
CS_450 NS_450 0 9.9999999999999998e-13
RS_449 NS_449 0 3.2672536376024027e+01
RS_450 NS_450 0 3.2672536376024027e+01
GL_449 0 NS_449 NS_450 0 1.2489866711430768e-01
GL_450 0 NS_450 NS_449 0 -1.2489866711430768e-01
GS_449_11 0 NS_449 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 451/452
CS_451 NS_451 0 9.9999999999999998e-13
CS_452 NS_452 0 9.9999999999999998e-13
RS_451 NS_451 0 3.6741731246022816e+01
RS_452 NS_452 0 3.6741731246022816e+01
GL_451 0 NS_451 NS_452 0 1.6399845549232167e-01
GL_452 0 NS_452 NS_451 0 -1.6399845549232167e-01
GS_451_11 0 NS_451 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 453/454
CS_453 NS_453 0 9.9999999999999998e-13
CS_454 NS_454 0 9.9999999999999998e-13
RS_453 NS_453 0 8.3646036557163740e+01
RS_454 NS_454 0 8.3646036557163740e+01
GL_453 0 NS_453 NS_454 0 1.6830719130342967e-01
GL_454 0 NS_454 NS_453 0 -1.6830719130342967e-01
GS_453_11 0 NS_453 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 455/456
CS_455 NS_455 0 9.9999999999999998e-13
CS_456 NS_456 0 9.9999999999999998e-13
RS_455 NS_455 0 4.0307732865054554e+01
RS_456 NS_456 0 4.0307732865054554e+01
GL_455 0 NS_455 NS_456 0 1.8890575271706389e-01
GL_456 0 NS_456 NS_455 0 -1.8890575271706389e-01
GS_455_11 0 NS_455 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 457/458
CS_457 NS_457 0 9.9999999999999998e-13
CS_458 NS_458 0 9.9999999999999998e-13
RS_457 NS_457 0 1.4268073111996583e+02
RS_458 NS_458 0 1.4268073111996583e+02
GL_457 0 NS_457 NS_458 0 1.9419078929943706e-01
GL_458 0 NS_458 NS_457 0 -1.9419078929943706e-01
GS_457_11 0 NS_457 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 459/460
CS_459 NS_459 0 9.9999999999999998e-13
CS_460 NS_460 0 9.9999999999999998e-13
RS_459 NS_459 0 7.1679198821979867e+01
RS_460 NS_460 0 7.1679198821979867e+01
GL_459 0 NS_459 NS_460 0 2.0702628270375376e-01
GL_460 0 NS_460 NS_459 0 -2.0702628270375376e-01
GS_459_11 0 NS_459 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 461/462
CS_461 NS_461 0 9.9999999999999998e-13
CS_462 NS_462 0 9.9999999999999998e-13
RS_461 NS_461 0 1.6005864146684806e+02
RS_462 NS_462 0 1.6005864146684809e+02
GL_461 0 NS_461 NS_462 0 2.5423900390253934e-01
GL_462 0 NS_462 NS_461 0 -2.5423900390253934e-01
GS_461_11 0 NS_461 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 463/464
CS_463 NS_463 0 9.9999999999999998e-13
CS_464 NS_464 0 9.9999999999999998e-13
RS_463 NS_463 0 1.9181463552142085e+02
RS_464 NS_464 0 1.9181463552142085e+02
GL_463 0 NS_463 NS_464 0 2.1188941693262670e-01
GL_464 0 NS_464 NS_463 0 -2.1188941693262670e-01
GS_463_11 0 NS_463 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 465/466
CS_465 NS_465 0 9.9999999999999998e-13
CS_466 NS_466 0 9.9999999999999998e-13
RS_465 NS_465 0 2.5689115313648813e+02
RS_466 NS_466 0 2.5689115313648813e+02
GL_465 0 NS_465 NS_466 0 2.1774212061821885e-01
GL_466 0 NS_466 NS_465 0 -2.1774212061821885e-01
GS_465_11 0 NS_465 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 467/468
CS_467 NS_467 0 9.9999999999999998e-13
CS_468 NS_468 0 9.9999999999999998e-13
RS_467 NS_467 0 6.2765149843829192e+01
RS_468 NS_468 0 6.2765149843829192e+01
GL_467 0 NS_467 NS_468 0 2.3246082537351351e-01
GL_468 0 NS_468 NS_467 0 -2.3246082537351351e-01
GS_467_11 0 NS_467 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 469/470
CS_469 NS_469 0 9.9999999999999998e-13
CS_470 NS_470 0 9.9999999999999998e-13
RS_469 NS_469 0 3.5419967361311882e+02
RS_470 NS_470 0 3.5419967361311882e+02
GL_469 0 NS_469 NS_470 0 2.2268031336810420e-01
GL_470 0 NS_470 NS_469 0 -2.2268031336810420e-01
GS_469_11 0 NS_469 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 471/472
CS_471 NS_471 0 9.9999999999999998e-13
CS_472 NS_472 0 9.9999999999999998e-13
RS_471 NS_471 0 9.0838548010669172e+01
RS_472 NS_472 0 9.0838548010669186e+01
GL_471 0 NS_471 NS_472 0 2.2647420085995260e-01
GL_472 0 NS_472 NS_471 0 -2.2647420085995260e-01
GS_471_11 0 NS_471 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 473/474
CS_473 NS_473 0 9.9999999999999998e-13
CS_474 NS_474 0 9.9999999999999998e-13
RS_473 NS_473 0 5.0298322136619066e+02
RS_474 NS_474 0 5.0298322136619078e+02
GL_473 0 NS_473 NS_474 0 2.4757175091537195e-01
GL_474 0 NS_474 NS_473 0 -2.4757175091537195e-01
GS_473_11 0 NS_473 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 475/476
CS_475 NS_475 0 9.9999999999999998e-13
CS_476 NS_476 0 9.9999999999999998e-13
RS_475 NS_475 0 1.1113846377285431e+02
RS_476 NS_476 0 1.1113846377285431e+02
GL_475 0 NS_475 NS_476 0 2.4529156966751164e-01
GL_476 0 NS_476 NS_475 0 -2.4529156966751164e-01
GS_475_11 0 NS_475 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 477/478
CS_477 NS_477 0 9.9999999999999998e-13
CS_478 NS_478 0 9.9999999999999998e-13
RS_477 NS_477 0 4.1132635267896995e+02
RS_478 NS_478 0 4.1132635267896990e+02
GL_477 0 NS_477 NS_478 0 2.4323159344727399e-01
GL_478 0 NS_478 NS_477 0 -2.4323159344727399e-01
GS_477_11 0 NS_477 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 479/480
CS_479 NS_479 0 9.9999999999999998e-13
CS_480 NS_480 0 9.9999999999999998e-13
RS_479 NS_479 0 6.1483243702508491e+02
RS_480 NS_480 0 6.1483243702508491e+02
GL_479 0 NS_479 NS_480 0 2.3313794138995145e-01
GL_480 0 NS_480 NS_479 0 -2.3313794138995145e-01
GS_479_11 0 NS_479 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 481/482
CS_481 NS_481 0 9.9999999999999998e-13
CS_482 NS_482 0 9.9999999999999998e-13
RS_481 NS_481 0 6.0708452252497170e+02
RS_482 NS_482 0 6.0708452252497170e+02
GL_481 0 NS_481 NS_482 0 2.3828547054015958e-01
GL_482 0 NS_482 NS_481 0 -2.3828547054015958e-01
GS_481_11 0 NS_481 NA_11 0 1.6921379288850509e+00
*
* Complex pair n. 483/484
CS_483 NS_483 0 9.9999999999999998e-13
CS_484 NS_484 0 9.9999999999999998e-13
RS_483 NS_483 0 1.9238303220034285e+02
RS_484 NS_484 0 1.9238303220034285e+02
GL_483 0 NS_483 NS_484 0 2.3639447764395666e-01
GL_484 0 NS_484 NS_483 0 -2.3639447764395666e-01
GS_483_11 0 NS_483 NA_11 0 1.6921379288850509e+00
*
* Real pole n. 485
CS_485 NS_485 0 9.9999999999999998e-13
RS_485 NS_485 0 1.2063458770185771e+00
GS_485_12 0 NS_485 NA_12 0 1.6921379288850509e+00
*
* Real pole n. 486
CS_486 NS_486 0 9.9999999999999998e-13
RS_486 NS_486 0 2.0414994648771170e+01
GS_486_12 0 NS_486 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 487/488
CS_487 NS_487 0 9.9999999999999998e-13
CS_488 NS_488 0 9.9999999999999998e-13
RS_487 NS_487 0 2.2164632983638530e+01
RS_488 NS_488 0 2.2164632983638530e+01
GL_487 0 NS_487 NS_488 0 6.2432580119989492e-02
GL_488 0 NS_488 NS_487 0 -6.2432580119989492e-02
GS_487_12 0 NS_487 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 489/490
CS_489 NS_489 0 9.9999999999999998e-13
CS_490 NS_490 0 9.9999999999999998e-13
RS_489 NS_489 0 2.4208144339458560e+01
RS_490 NS_490 0 2.4208144339458560e+01
GL_489 0 NS_489 NS_490 0 8.7759448763363015e-02
GL_490 0 NS_490 NS_489 0 -8.7759448763363015e-02
GS_489_12 0 NS_489 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 491/492
CS_491 NS_491 0 9.9999999999999998e-13
CS_492 NS_492 0 9.9999999999999998e-13
RS_491 NS_491 0 1.3097029666184031e+02
RS_492 NS_492 0 1.3097029666184031e+02
GL_491 0 NS_491 NS_492 0 2.9672291989323329e-01
GL_492 0 NS_492 NS_491 0 -2.9672291989323329e-01
GS_491_12 0 NS_491 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 493/494
CS_493 NS_493 0 9.9999999999999998e-13
CS_494 NS_494 0 9.9999999999999998e-13
RS_493 NS_493 0 3.2672536376024027e+01
RS_494 NS_494 0 3.2672536376024027e+01
GL_493 0 NS_493 NS_494 0 1.2489866711430768e-01
GL_494 0 NS_494 NS_493 0 -1.2489866711430768e-01
GS_493_12 0 NS_493 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 495/496
CS_495 NS_495 0 9.9999999999999998e-13
CS_496 NS_496 0 9.9999999999999998e-13
RS_495 NS_495 0 3.6741731246022816e+01
RS_496 NS_496 0 3.6741731246022816e+01
GL_495 0 NS_495 NS_496 0 1.6399845549232167e-01
GL_496 0 NS_496 NS_495 0 -1.6399845549232167e-01
GS_495_12 0 NS_495 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 497/498
CS_497 NS_497 0 9.9999999999999998e-13
CS_498 NS_498 0 9.9999999999999998e-13
RS_497 NS_497 0 8.3646036557163740e+01
RS_498 NS_498 0 8.3646036557163740e+01
GL_497 0 NS_497 NS_498 0 1.6830719130342967e-01
GL_498 0 NS_498 NS_497 0 -1.6830719130342967e-01
GS_497_12 0 NS_497 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 499/500
CS_499 NS_499 0 9.9999999999999998e-13
CS_500 NS_500 0 9.9999999999999998e-13
RS_499 NS_499 0 4.0307732865054554e+01
RS_500 NS_500 0 4.0307732865054554e+01
GL_499 0 NS_499 NS_500 0 1.8890575271706389e-01
GL_500 0 NS_500 NS_499 0 -1.8890575271706389e-01
GS_499_12 0 NS_499 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 501/502
CS_501 NS_501 0 9.9999999999999998e-13
CS_502 NS_502 0 9.9999999999999998e-13
RS_501 NS_501 0 1.4268073111996583e+02
RS_502 NS_502 0 1.4268073111996583e+02
GL_501 0 NS_501 NS_502 0 1.9419078929943706e-01
GL_502 0 NS_502 NS_501 0 -1.9419078929943706e-01
GS_501_12 0 NS_501 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 503/504
CS_503 NS_503 0 9.9999999999999998e-13
CS_504 NS_504 0 9.9999999999999998e-13
RS_503 NS_503 0 7.1679198821979867e+01
RS_504 NS_504 0 7.1679198821979867e+01
GL_503 0 NS_503 NS_504 0 2.0702628270375376e-01
GL_504 0 NS_504 NS_503 0 -2.0702628270375376e-01
GS_503_12 0 NS_503 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 505/506
CS_505 NS_505 0 9.9999999999999998e-13
CS_506 NS_506 0 9.9999999999999998e-13
RS_505 NS_505 0 1.6005864146684806e+02
RS_506 NS_506 0 1.6005864146684809e+02
GL_505 0 NS_505 NS_506 0 2.5423900390253934e-01
GL_506 0 NS_506 NS_505 0 -2.5423900390253934e-01
GS_505_12 0 NS_505 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 507/508
CS_507 NS_507 0 9.9999999999999998e-13
CS_508 NS_508 0 9.9999999999999998e-13
RS_507 NS_507 0 1.9181463552142085e+02
RS_508 NS_508 0 1.9181463552142085e+02
GL_507 0 NS_507 NS_508 0 2.1188941693262670e-01
GL_508 0 NS_508 NS_507 0 -2.1188941693262670e-01
GS_507_12 0 NS_507 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 509/510
CS_509 NS_509 0 9.9999999999999998e-13
CS_510 NS_510 0 9.9999999999999998e-13
RS_509 NS_509 0 2.5689115313648813e+02
RS_510 NS_510 0 2.5689115313648813e+02
GL_509 0 NS_509 NS_510 0 2.1774212061821885e-01
GL_510 0 NS_510 NS_509 0 -2.1774212061821885e-01
GS_509_12 0 NS_509 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 511/512
CS_511 NS_511 0 9.9999999999999998e-13
CS_512 NS_512 0 9.9999999999999998e-13
RS_511 NS_511 0 6.2765149843829192e+01
RS_512 NS_512 0 6.2765149843829192e+01
GL_511 0 NS_511 NS_512 0 2.3246082537351351e-01
GL_512 0 NS_512 NS_511 0 -2.3246082537351351e-01
GS_511_12 0 NS_511 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 513/514
CS_513 NS_513 0 9.9999999999999998e-13
CS_514 NS_514 0 9.9999999999999998e-13
RS_513 NS_513 0 3.5419967361311882e+02
RS_514 NS_514 0 3.5419967361311882e+02
GL_513 0 NS_513 NS_514 0 2.2268031336810420e-01
GL_514 0 NS_514 NS_513 0 -2.2268031336810420e-01
GS_513_12 0 NS_513 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 515/516
CS_515 NS_515 0 9.9999999999999998e-13
CS_516 NS_516 0 9.9999999999999998e-13
RS_515 NS_515 0 9.0838548010669172e+01
RS_516 NS_516 0 9.0838548010669186e+01
GL_515 0 NS_515 NS_516 0 2.2647420085995260e-01
GL_516 0 NS_516 NS_515 0 -2.2647420085995260e-01
GS_515_12 0 NS_515 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 517/518
CS_517 NS_517 0 9.9999999999999998e-13
CS_518 NS_518 0 9.9999999999999998e-13
RS_517 NS_517 0 5.0298322136619066e+02
RS_518 NS_518 0 5.0298322136619078e+02
GL_517 0 NS_517 NS_518 0 2.4757175091537195e-01
GL_518 0 NS_518 NS_517 0 -2.4757175091537195e-01
GS_517_12 0 NS_517 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 519/520
CS_519 NS_519 0 9.9999999999999998e-13
CS_520 NS_520 0 9.9999999999999998e-13
RS_519 NS_519 0 1.1113846377285431e+02
RS_520 NS_520 0 1.1113846377285431e+02
GL_519 0 NS_519 NS_520 0 2.4529156966751164e-01
GL_520 0 NS_520 NS_519 0 -2.4529156966751164e-01
GS_519_12 0 NS_519 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 521/522
CS_521 NS_521 0 9.9999999999999998e-13
CS_522 NS_522 0 9.9999999999999998e-13
RS_521 NS_521 0 4.1132635267896995e+02
RS_522 NS_522 0 4.1132635267896990e+02
GL_521 0 NS_521 NS_522 0 2.4323159344727399e-01
GL_522 0 NS_522 NS_521 0 -2.4323159344727399e-01
GS_521_12 0 NS_521 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 523/524
CS_523 NS_523 0 9.9999999999999998e-13
CS_524 NS_524 0 9.9999999999999998e-13
RS_523 NS_523 0 6.1483243702508491e+02
RS_524 NS_524 0 6.1483243702508491e+02
GL_523 0 NS_523 NS_524 0 2.3313794138995145e-01
GL_524 0 NS_524 NS_523 0 -2.3313794138995145e-01
GS_523_12 0 NS_523 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 525/526
CS_525 NS_525 0 9.9999999999999998e-13
CS_526 NS_526 0 9.9999999999999998e-13
RS_525 NS_525 0 6.0708452252497170e+02
RS_526 NS_526 0 6.0708452252497170e+02
GL_525 0 NS_525 NS_526 0 2.3828547054015958e-01
GL_526 0 NS_526 NS_525 0 -2.3828547054015958e-01
GS_525_12 0 NS_525 NA_12 0 1.6921379288850509e+00
*
* Complex pair n. 527/528
CS_527 NS_527 0 9.9999999999999998e-13
CS_528 NS_528 0 9.9999999999999998e-13
RS_527 NS_527 0 1.9238303220034285e+02
RS_528 NS_528 0 1.9238303220034285e+02
GL_527 0 NS_527 NS_528 0 2.3639447764395666e-01
GL_528 0 NS_528 NS_527 0 -2.3639447764395666e-01
GS_527_12 0 NS_527 NA_12 0 1.6921379288850509e+00
*
******************************


.ends
*******************
* End of subcircuit
*******************
